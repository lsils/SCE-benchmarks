module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n113 , n114 , n115 , n116 , n117 , n118 , n120 , n121 , n122 , n123 , n124 , n126 , n127 , n128 , n129 , n131 , n132 , n133 , n135 , n137 , n138 , n139 , n141 , n143 , n144 , n145 , n147 , n148 , n149 , n151 , n152 , n153 , n154 , n155 , n157 , n158 , n159 , n160 , n161 , n162 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 ;
  buffer buf_n131( .i (x15), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n135( .i (x16), .o (n135) );
  buffer buf_n141( .i (x18), .o (n141) );
  assign n268 = n135 | n141 ;
  buffer buf_n269( .i (n268), .o (n269) );
  assign n276 = n133 & ~n269 ;
  buffer buf_n137( .i (x17), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n143( .i (x19), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  assign n277 = n139 & n145 ;
  assign n278 = n135 & ~n141 ;
  buffer buf_n279( .i (n278), .o (n279) );
  assign n286 = ( n139 & n145 ) | ( n139 & n279 ) | ( n145 & n279 ) ;
  assign n287 = ( n276 & ~n277 ) | ( n276 & n286 ) | ( ~n277 & n286 ) ;
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n147( .i (x20), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  assign n294 = n137 | n143 ;
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = n149 | n295 ;
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n126( .i (x14), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n270( .i (n269), .o (n270) );
  assign n298 = n129 & ~n270 ;
  assign n299 = ( n149 & ~n279 ) | ( n149 & n295 ) | ( ~n279 & n295 ) ;
  buffer buf_n300( .i (n299), .o (n300) );
  assign n301 = ( n297 & n298 ) | ( n297 & ~n300 ) | ( n298 & ~n300 ) ;
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n120( .i (x13), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n271( .i (n270), .o (n271) );
  assign n307 = n124 & ~n271 ;
  buffer buf_n151( .i (x21), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  assign n308 = ( n155 & ~n281 ) | ( n155 & n297 ) | ( ~n281 & n297 ) ;
  assign n309 = n148 | n152 ;
  assign n310 = n295 | n309 ;
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  assign n313 = ( n307 & ~n308 ) | ( n307 & n312 ) | ( ~n308 & n312 ) ;
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n113( .i (x12), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n272( .i (n271), .o (n272) );
  assign n318 = n118 & ~n272 ;
  buffer buf_n157( .i (x22), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  assign n319 = n161 | n311 ;
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n282( .i (n281), .o (n282) );
  assign n321 = ( n162 & ~n282 ) | ( n162 & n312 ) | ( ~n282 & n312 ) ;
  assign n322 = ( n318 & n320 ) | ( n318 & ~n321 ) | ( n320 & ~n321 ) ;
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n105( .i (x11), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n273( .i (n272), .o (n273) );
  assign n326 = n111 & ~n273 ;
  buffer buf_n164( .i (x23), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n283( .i (n282), .o (n283) );
  assign n327 = ( n170 & ~n283 ) | ( n170 & n320 ) | ( ~n283 & n320 ) ;
  assign n328 = n158 | n165 ;
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  assign n332 = n312 | n331 ;
  buffer buf_n333( .i (n332), .o (n333) );
  assign n334 = ( n326 & ~n327 ) | ( n326 & n333 ) | ( ~n327 & n333 ) ;
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n96( .i (x10), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n274( .i (n273), .o (n274) );
  assign n337 = n103 & ~n274 ;
  buffer buf_n172( .i (x24), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n284( .i (n283), .o (n284) );
  assign n338 = ( n179 & ~n284 ) | ( n179 & n333 ) | ( ~n284 & n333 ) ;
  assign n339 = n175 | n329 ;
  assign n340 = n311 | n339 ;
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  assign n344 = ( n337 & ~n338 ) | ( n337 & n343 ) | ( ~n338 & n343 ) ;
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n87( .i (x9), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  assign n346 = n94 & ~n274 ;
  buffer buf_n181( .i (x25), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  assign n347 = n188 | n342 ;
  assign n348 = ( n188 & ~n284 ) | ( n188 & n342 ) | ( ~n284 & n342 ) ;
  assign n349 = ( n346 & n347 ) | ( n346 & ~n348 ) | ( n347 & ~n348 ) ;
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n77( .i (x8), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n275( .i (n274), .o (n275) );
  assign n351 = n85 & ~n275 ;
  buffer buf_n190( .i (x26), .o (n190) );
  assign n352 = n181 | n190 ;
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  assign n360 = n343 | n359 ;
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  assign n361 = ~n197 & n284 ;
  buffer buf_n362( .i (n283), .o (n362) );
  assign n363 = ( n188 & n197 ) | ( n188 & ~n362 ) | ( n197 & ~n362 ) ;
  assign n364 = ( n343 & ~n361 ) | ( n343 & n363 ) | ( ~n361 & n363 ) ;
  assign n365 = ( n351 & n360 ) | ( n351 & ~n364 ) | ( n360 & ~n364 ) ;
  buffer buf_n67( .i (x7), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  assign n366 = n75 & ~n275 ;
  buffer buf_n199( .i (x27), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  assign n367 = n203 | n355 ;
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  assign n371 = n343 | n370 ;
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  assign n372 = ~n206 & n362 ;
  assign n373 = ( n206 & n358 ) | ( n206 & ~n362 ) | ( n358 & ~n362 ) ;
  buffer buf_n374( .i (n342), .o (n374) );
  assign n375 = ( ~n372 & n373 ) | ( ~n372 & n374 ) | ( n373 & n374 ) ;
  assign n376 = ( n366 & n371 ) | ( n366 & ~n375 ) | ( n371 & ~n375 ) ;
  buffer buf_n58( .i (x6), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  assign n377 = n65 & ~n274 ;
  buffer buf_n208( .i (x28), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  assign n378 = n200 | n209 ;
  assign n379 = n353 | n378 ;
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  assign n384 = n341 | n382 ;
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n386 = ~n214 & n283 ;
  buffer buf_n387( .i (n282), .o (n387) );
  assign n388 = ( n214 & n368 ) | ( n214 & ~n387 ) | ( n368 & ~n387 ) ;
  buffer buf_n389( .i (n341), .o (n389) );
  assign n390 = ( ~n386 & n388 ) | ( ~n386 & n389 ) | ( n388 & n389 ) ;
  assign n391 = ( n377 & n385 ) | ( n377 & ~n390 ) | ( n385 & ~n390 ) ;
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n48( .i (x5), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  assign n393 = n56 & ~n275 ;
  buffer buf_n216( .i (x29), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n383( .i (n382), .o (n383) );
  assign n394 = n223 | n383 ;
  assign n395 = n374 | n394 ;
  assign n396 = ~n223 & n362 ;
  buffer buf_n397( .i (n387), .o (n397) );
  assign n398 = ( n223 & n383 ) | ( n223 & ~n397 ) | ( n383 & ~n397 ) ;
  assign n399 = ( n374 & ~n396 ) | ( n374 & n398 ) | ( ~n396 & n398 ) ;
  assign n400 = ( n393 & n395 ) | ( n393 & ~n399 ) | ( n395 & ~n399 ) ;
  buffer buf_n225( .i (x30), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  assign n401 = n222 & ~n231 ;
  assign n402 = n397 & n401 ;
  buffer buf_n39( .i (x4), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n403( .i (n273), .o (n403) );
  assign n404 = n46 & ~n403 ;
  assign n405 = n402 | n404 ;
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n232( .i (n231), .o (n232) );
  assign n406 = ~n231 & n382 ;
  assign n407 = ( ~n232 & n389 ) | ( ~n232 & n406 ) | ( n389 & n406 ) ;
  assign n408 = ( n221 & ~n230 ) | ( n221 & n282 ) | ( ~n230 & n282 ) ;
  assign n409 = n382 | n408 ;
  assign n410 = n389 | n409 ;
  assign n411 = ( n285 & n407 ) | ( n285 & ~n410 ) | ( n407 & ~n410 ) ;
  assign n412 = n405 | n411 ;
  buffer buf_n30( .i (x3), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  assign n413 = n37 & ~n403 ;
  buffer buf_n234( .i (x31), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n414( .i (n281), .o (n414) );
  assign n415 = ~n239 & n414 ;
  buffer buf_n416( .i (n415), .o (n416) );
  assign n418 = n217 | n226 ;
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  assign n424 = n416 & n423 ;
  assign n425 = n413 | n424 ;
  buffer buf_n240( .i (n239), .o (n240) );
  assign n426 = n240 & n387 ;
  assign n427 = ~n423 & n426 ;
  assign n428 = n385 | n427 ;
  buffer buf_n417( .i (n416), .o (n417) );
  assign n429 = n383 & ~n416 ;
  assign n430 = ( n374 & ~n417 ) | ( n374 & n429 ) | ( ~n417 & n429 ) ;
  assign n431 = ( n425 & n428 ) | ( n425 & ~n430 ) | ( n428 & ~n430 ) ;
  buffer buf_n21( .i (x2), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  assign n432 = n28 & ~n403 ;
  buffer buf_n242( .i (x32), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  assign n433 = ~n247 & n414 ;
  buffer buf_n434( .i (n433), .o (n434) );
  assign n436 = n239 | n421 ;
  buffer buf_n437( .i (n436), .o (n437) );
  assign n438 = n434 & n437 ;
  assign n439 = n432 | n438 ;
  buffer buf_n248( .i (n247), .o (n248) );
  assign n440 = n248 & n387 ;
  assign n441 = ~n437 & n440 ;
  assign n442 = n385 | n441 ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n443 = n383 & ~n434 ;
  buffer buf_n444( .i (n389), .o (n444) );
  assign n445 = ( ~n435 & n443 ) | ( ~n435 & n444 ) | ( n443 & n444 ) ;
  assign n446 = ( n439 & n442 ) | ( n439 & ~n445 ) | ( n442 & ~n445 ) ;
  buffer buf_n12( .i (x1), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  assign n447 = n19 & ~n403 ;
  buffer buf_n250( .i (x33), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  assign n448 = n236 | n244 ;
  assign n449 = n419 | n448 ;
  assign n450 = n380 | n449 ;
  buffer buf_n451( .i (n450), .o (n451) );
  assign n452 = n341 | n451 ;
  assign n453 = ( n257 & ~n397 ) | ( n257 & n452 ) | ( ~n397 & n452 ) ;
  assign n454 = n175 | n253 ;
  assign n455 = n330 | n454 ;
  assign n456 = n312 | n455 ;
  assign n457 = n451 | n456 ;
  buffer buf_n458( .i (n457), .o (n458) );
  assign n459 = ( n447 & ~n453 ) | ( n447 & n458 ) | ( ~n453 & n458 ) ;
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  assign n461 = n10 & ~n275 ;
  buffer buf_n259( .i (x34), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  assign n462 = n267 | n458 ;
  assign n463 = ( n267 & ~n285 ) | ( n267 & n458 ) | ( ~n285 & n458 ) ;
  assign n464 = ( n461 & n462 ) | ( n461 & ~n463 ) | ( n462 & ~n463 ) ;
  assign y0 = ~n293 ;
  assign y1 = ~n306 ;
  assign y2 = ~n317 ;
  assign y3 = ~n325 ;
  assign y4 = ~n336 ;
  assign y5 = ~n345 ;
  assign y6 = ~n350 ;
  assign y7 = ~n365 ;
  assign y8 = ~n376 ;
  assign y9 = ~n392 ;
  assign y10 = ~n400 ;
  assign y11 = ~n412 ;
  assign y12 = ~n431 ;
  assign y13 = ~n446 ;
  assign y14 = ~n460 ;
  assign y15 = ~n464 ;
endmodule
