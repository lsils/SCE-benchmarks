module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( a_44_ , a_5_ , a_38_ , a_43_ , a_20_ , a_27_ , a_8_ , a_40_ , a_47_ , a_11_ , a_0_ , a_6_ , a_16_ , a_9_ , a_31_ , a_4_ , a_30_ , a_35_ , a_26_ , a_19_ , a_7_ , a_13_ , a_45_ , a_34_ , a_42_ , a_14_ , a_41_ , a_17_ , a_37_ , a_18_ , a_29_ , a_21_ , a_32_ , a_22_ , a_36_ , a_3_ , a_28_ , a_46_ , a_25_ , a_10_ , a_12_ , a_33_ , a_24_ , a_1_ , a_15_ , a_2_ , a_39_ , a_23_ , b_47_ , b_43_ , b_40_ , b_11_ , b_7_ , b_5_ , b_32_ , b_17_ , b_29_ , b_25_ , b_12_ , b_16_ , b_1_ , b_42_ , b_0_ , b_28_ , b_9_ , b_36_ , b_2_ , b_20_ , b_41_ , b_33_ , b_31_ , b_34_ , b_13_ , b_21_ , b_35_ , b_39_ , b_27_ , b_46_ , b_4_ , b_14_ , b_37_ , b_22_ , b_6_ , b_38_ , b_18_ , b_15_ , b_30_ , b_8_ , b_26_ , b_24_ , b_19_ , b_23_ , b_10_ , b_3_ , b_45_ , b_44_ );
  input a_44_ , a_5_ , a_38_ , a_43_ , a_20_ , a_27_ , a_8_ , a_40_ , a_47_ , a_11_ , a_0_ , a_6_ , a_16_ , a_9_ , a_31_ , a_4_ , a_30_ , a_35_ , a_26_ , a_19_ , a_7_ , a_13_ , a_45_ , a_34_ , a_42_ , a_14_ , a_41_ , a_17_ , a_37_ , a_18_ , a_29_ , a_21_ , a_32_ , a_22_ , a_36_ , a_3_ , a_28_ , a_46_ , a_25_ , a_10_ , a_12_ , a_33_ , a_24_ , a_1_ , a_15_ , a_2_ , a_39_ , a_23_ ;
  output b_47_ , b_43_ , b_40_ , b_11_ , b_7_ , b_5_ , b_32_ , b_17_ , b_29_ , b_25_ , b_12_ , b_16_ , b_1_ , b_42_ , b_0_ , b_28_ , b_9_ , b_36_ , b_2_ , b_20_ , b_41_ , b_33_ , b_31_ , b_34_ , b_13_ , b_21_ , b_35_ , b_39_ , b_27_ , b_46_ , b_4_ , b_14_ , b_37_ , b_22_ , b_6_ , b_38_ , b_18_ , b_15_ , b_30_ , b_8_ , b_26_ , b_24_ , b_19_ , b_23_ , b_10_ , b_3_ , b_45_ , b_44_ ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 ;
  buffer buf_n102( .i (a_33_), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n71( .i (a_35_), .o (n71) );
  buffer buf_n78( .i (a_34_), .o (n78) );
  assign n113 = n71 & n78 ;
  assign n114 = n103 & n113 ;
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n69( .i (a_30_), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n67( .i (a_31_), .o (n67) );
  buffer buf_n90( .i (a_32_), .o (n90) );
  assign n116 = n67 | n90 ;
  assign n117 = n70 | n116 ;
  buffer buf_n118( .i (n117), .o (n118) );
  assign n119 = n115 & n118 ;
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  assign n122 = n71 | n78 ;
  assign n123 = n103 | n122 ;
  buffer buf_n124( .i (n123), .o (n124) );
  assign n125 = n67 & n90 ;
  assign n126 = n70 & n125 ;
  buffer buf_n127( .i (n126), .o (n127) );
  assign n128 = n124 & n127 ;
  buffer buf_n129( .i (n128), .o (n129) );
  assign n130 = ( n71 & n78 ) | ( n71 & n102 ) | ( n78 & n102 ) ;
  buffer buf_n131( .i (n130), .o (n131) );
  assign n132 = ( n67 & n69 ) | ( n67 & n90 ) | ( n69 & n90 ) ;
  buffer buf_n133( .i (n132), .o (n133) );
  assign n134 = n131 & n133 ;
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  assign n137 = n129 & n136 ;
  assign n138 = n121 & n137 ;
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n54( .i (a_27_), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n87( .i (a_29_), .o (n87) );
  buffer buf_n96( .i (a_28_), .o (n96) );
  assign n140 = n87 & n96 ;
  assign n141 = n55 & n140 ;
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n104( .i (a_24_), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n72( .i (a_26_), .o (n72) );
  buffer buf_n98( .i (a_25_), .o (n98) );
  assign n143 = n72 | n98 ;
  assign n144 = n105 | n143 ;
  buffer buf_n145( .i (n144), .o (n145) );
  assign n146 = n142 | n145 ;
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  assign n149 = ( n54 & n87 ) | ( n54 & n96 ) | ( n87 & n96 ) ;
  buffer buf_n150( .i (n149), .o (n150) );
  assign n151 = ( n72 & n98 ) | ( n72 & n104 ) | ( n98 & n104 ) ;
  buffer buf_n152( .i (n151), .o (n152) );
  assign n153 = n150 | n152 ;
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  assign n156 = n87 | n96 ;
  assign n157 = n55 | n156 ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n159 = n72 & n98 ;
  assign n160 = n105 & n159 ;
  buffer buf_n161( .i (n160), .o (n161) );
  assign n162 = n158 | n161 ;
  buffer buf_n163( .i (n162), .o (n163) );
  assign n164 = n155 | n163 ;
  assign n165 = n148 | n164 ;
  buffer buf_n166( .i (n165), .o (n166) );
  assign n167 = n139 & n166 ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = n115 | n118 ;
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  assign n172 = n124 | n127 ;
  buffer buf_n173( .i (n172), .o (n173) );
  assign n174 = n131 | n133 ;
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  assign n177 = n173 & n176 ;
  assign n178 = n171 & n177 ;
  buffer buf_n179( .i (n178), .o (n179) );
  assign n180 = n142 & n145 ;
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  assign n183 = n150 & n152 ;
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  assign n186 = n158 & n161 ;
  buffer buf_n187( .i (n186), .o (n187) );
  assign n188 = n185 | n187 ;
  assign n189 = n182 | n188 ;
  buffer buf_n190( .i (n189), .o (n190) );
  assign n191 = n179 & n190 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = n168 & n192 ;
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  assign n196 = ( n120 & n129 ) | ( n120 & n136 ) | ( n129 & n136 ) ;
  buffer buf_n197( .i (n196), .o (n197) );
  assign n198 = ( n147 & n155 ) | ( n147 & n163 ) | ( n155 & n163 ) ;
  buffer buf_n199( .i (n198), .o (n199) );
  assign n200 = n197 & n199 ;
  buffer buf_n201( .i (n200), .o (n201) );
  assign n202 = ( n170 & n173 ) | ( n170 & n176 ) | ( n173 & n176 ) ;
  buffer buf_n203( .i (n202), .o (n203) );
  assign n204 = ( n181 & n185 ) | ( n181 & n187 ) | ( n185 & n187 ) ;
  buffer buf_n205( .i (n204), .o (n205) );
  assign n206 = n203 & n205 ;
  buffer buf_n207( .i (n206), .o (n207) );
  assign n208 = n201 & n207 ;
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  assign n211 = n129 | n136 ;
  assign n212 = n121 | n211 ;
  buffer buf_n213( .i (n212), .o (n213) );
  assign n214 = n155 & n163 ;
  assign n215 = n148 & n214 ;
  buffer buf_n216( .i (n215), .o (n216) );
  assign n217 = n213 & n216 ;
  buffer buf_n218( .i (n217), .o (n218) );
  assign n219 = n173 | n176 ;
  assign n220 = n171 | n219 ;
  buffer buf_n221( .i (n220), .o (n221) );
  assign n222 = n185 & n187 ;
  assign n223 = n182 & n222 ;
  buffer buf_n224( .i (n223), .o (n224) );
  assign n225 = n221 & n224 ;
  buffer buf_n226( .i (n225), .o (n226) );
  assign n227 = n218 & n226 ;
  buffer buf_n228( .i (n227), .o (n228) );
  assign n229 = n210 & n228 ;
  assign n230 = n195 & n229 ;
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n110( .i (a_39_), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n57( .i (a_40_), .o (n57) );
  buffer buf_n82( .i (a_41_), .o (n82) );
  assign n232 = n57 & n82 ;
  assign n233 = n111 & n232 ;
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n92( .i (a_36_), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n51( .i (a_38_), .o (n51) );
  buffer buf_n84( .i (a_37_), .o (n84) );
  assign n235 = n51 | n84 ;
  assign n236 = n93 | n235 ;
  buffer buf_n237( .i (n236), .o (n237) );
  assign n238 = n234 & n237 ;
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  assign n241 = n57 | n82 ;
  assign n242 = n111 | n241 ;
  buffer buf_n243( .i (n242), .o (n243) );
  assign n244 = n51 & n84 ;
  assign n245 = n93 & n244 ;
  buffer buf_n246( .i (n245), .o (n246) );
  assign n247 = n243 & n246 ;
  buffer buf_n248( .i (n247), .o (n248) );
  assign n249 = ( n57 & n82 ) | ( n57 & n110 ) | ( n82 & n110 ) ;
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = ( n51 & n84 ) | ( n51 & n92 ) | ( n84 & n92 ) ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n253 = n250 & n252 ;
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  assign n256 = n248 | n255 ;
  assign n257 = n240 | n256 ;
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n49( .i (a_44_), .o (n49) );
  buffer buf_n52( .i (a_43_), .o (n52) );
  buffer buf_n79( .i (a_42_), .o (n79) );
  assign n259 = ( n49 & n52 ) | ( n49 & n79 ) | ( n52 & n79 ) ;
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n58( .i (a_47_), .o (n58) );
  buffer buf_n76( .i (a_45_), .o (n76) );
  buffer buf_n97( .i (a_46_), .o (n97) );
  assign n261 = ( n58 & n76 ) | ( n58 & n97 ) | ( n76 & n97 ) ;
  buffer buf_n262( .i (n261), .o (n262) );
  assign n263 = n260 | n262 ;
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n80( .i (n79), .o (n80) );
  assign n266 = n49 & n52 ;
  assign n267 = n80 & n266 ;
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n77( .i (n76), .o (n77) );
  assign n269 = n58 | n97 ;
  assign n270 = n77 | n269 ;
  buffer buf_n271( .i (n270), .o (n271) );
  assign n272 = n268 | n271 ;
  buffer buf_n273( .i (n272), .o (n273) );
  assign n274 = n265 & n273 ;
  assign n275 = n58 & n97 ;
  assign n276 = n77 & n275 ;
  buffer buf_n277( .i (n276), .o (n277) );
  assign n278 = n49 | n52 ;
  assign n279 = n80 | n278 ;
  buffer buf_n280( .i (n279), .o (n280) );
  assign n281 = n277 | n280 ;
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  assign n284 = n274 & n283 ;
  buffer buf_n285( .i (n284), .o (n285) );
  assign n286 = n258 | n285 ;
  buffer buf_n287( .i (n286), .o (n287) );
  assign n288 = n234 | n237 ;
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  assign n291 = n243 | n246 ;
  buffer buf_n292( .i (n291), .o (n292) );
  assign n293 = n250 | n252 ;
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = n292 | n295 ;
  assign n297 = n290 | n296 ;
  buffer buf_n298( .i (n297), .o (n298) );
  assign n299 = n260 & n262 ;
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  assign n302 = n268 & n271 ;
  buffer buf_n303( .i (n302), .o (n303) );
  assign n304 = n301 & n303 ;
  assign n305 = n277 & n280 ;
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  assign n308 = n304 & n307 ;
  buffer buf_n309( .i (n308), .o (n309) );
  assign n310 = n298 | n309 ;
  buffer buf_n311( .i (n310), .o (n311) );
  assign n312 = n287 | n311 ;
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  assign n315 = n248 & n255 ;
  assign n316 = n240 & n315 ;
  buffer buf_n317( .i (n316), .o (n317) );
  assign n318 = n265 | n273 ;
  assign n319 = n283 | n318 ;
  buffer buf_n320( .i (n319), .o (n320) );
  assign n321 = n317 | n320 ;
  buffer buf_n322( .i (n321), .o (n322) );
  assign n323 = n292 & n295 ;
  assign n324 = n290 & n323 ;
  buffer buf_n325( .i (n324), .o (n325) );
  assign n326 = n301 | n303 ;
  assign n327 = n307 | n326 ;
  buffer buf_n328( .i (n327), .o (n328) );
  assign n329 = n325 | n328 ;
  buffer buf_n330( .i (n329), .o (n330) );
  assign n331 = n322 | n330 ;
  buffer buf_n332( .i (n331), .o (n332) );
  assign n333 = ( n239 & n248 ) | ( n239 & n255 ) | ( n248 & n255 ) ;
  buffer buf_n334( .i (n333), .o (n334) );
  assign n335 = ( n265 & n273 ) | ( n265 & n282 ) | ( n273 & n282 ) ;
  buffer buf_n336( .i (n335), .o (n336) );
  assign n337 = n334 | n336 ;
  buffer buf_n338( .i (n337), .o (n338) );
  assign n339 = ( n289 & n292 ) | ( n289 & n295 ) | ( n292 & n295 ) ;
  buffer buf_n340( .i (n339), .o (n340) );
  assign n341 = ( n301 & n303 ) | ( n301 & n306 ) | ( n303 & n306 ) ;
  buffer buf_n342( .i (n341), .o (n342) );
  assign n343 = n340 | n342 ;
  buffer buf_n344( .i (n343), .o (n344) );
  assign n345 = n338 | n344 ;
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  assign n348 = n332 | n347 ;
  assign n349 = n314 | n348 ;
  buffer buf_n350( .i (n349), .o (n350) );
  assign n351 = n231 & n350 ;
  buffer buf_n352( .i (n351), .o (n352) );
  assign n353 = n139 | n166 ;
  buffer buf_n354( .i (n353), .o (n354) );
  assign n355 = n179 | n190 ;
  buffer buf_n356( .i (n355), .o (n356) );
  assign n357 = n354 & n356 ;
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  assign n360 = n213 | n216 ;
  buffer buf_n361( .i (n360), .o (n361) );
  assign n362 = n221 | n224 ;
  buffer buf_n363( .i (n362), .o (n363) );
  assign n364 = n361 & n363 ;
  buffer buf_n365( .i (n364), .o (n365) );
  assign n366 = n197 | n199 ;
  buffer buf_n367( .i (n366), .o (n367) );
  assign n368 = n203 | n205 ;
  buffer buf_n369( .i (n368), .o (n369) );
  assign n370 = n367 & n369 ;
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  assign n373 = n365 & n372 ;
  assign n374 = n359 & n373 ;
  buffer buf_n375( .i (n374), .o (n375) );
  assign n376 = n258 & n285 ;
  buffer buf_n377( .i (n376), .o (n377) );
  assign n378 = n298 & n309 ;
  buffer buf_n379( .i (n378), .o (n379) );
  assign n380 = n377 | n379 ;
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  assign n383 = n317 & n320 ;
  buffer buf_n384( .i (n383), .o (n384) );
  assign n385 = n325 & n328 ;
  buffer buf_n386( .i (n385), .o (n386) );
  assign n387 = n384 | n386 ;
  buffer buf_n388( .i (n387), .o (n388) );
  assign n389 = n334 & n336 ;
  buffer buf_n390( .i (n389), .o (n390) );
  assign n391 = n340 & n342 ;
  buffer buf_n392( .i (n391), .o (n392) );
  assign n393 = n390 | n392 ;
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  assign n396 = n388 | n395 ;
  assign n397 = n382 | n396 ;
  buffer buf_n398( .i (n397), .o (n398) );
  assign n399 = n375 & n398 ;
  buffer buf_n400( .i (n399), .o (n400) );
  assign n401 = n352 & n400 ;
  buffer buf_n402( .i (n401), .o (n402) );
  assign n403 = n168 | n192 ;
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  assign n406 = n201 | n207 ;
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  assign n409 = n218 | n226 ;
  buffer buf_n410( .i (n409), .o (n410) );
  assign n411 = n408 & n410 ;
  assign n412 = n405 & n411 ;
  buffer buf_n413( .i (n412), .o (n413) );
  assign n414 = n287 & n311 ;
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  assign n417 = n322 & n330 ;
  buffer buf_n418( .i (n417), .o (n418) );
  assign n419 = n338 & n344 ;
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  assign n422 = n418 | n421 ;
  assign n423 = n416 | n422 ;
  buffer buf_n424( .i (n423), .o (n424) );
  assign n425 = n413 & n424 ;
  buffer buf_n426( .i (n425), .o (n426) );
  assign n427 = n354 | n356 ;
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  assign n430 = n361 | n363 ;
  buffer buf_n431( .i (n430), .o (n431) );
  assign n432 = n367 | n369 ;
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  assign n435 = n431 & n434 ;
  assign n436 = n429 & n435 ;
  buffer buf_n437( .i (n436), .o (n437) );
  assign n438 = n377 & n379 ;
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  assign n441 = n384 & n386 ;
  buffer buf_n442( .i (n441), .o (n442) );
  assign n443 = n390 & n392 ;
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  assign n446 = n442 | n445 ;
  assign n447 = n440 | n446 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = n437 & n448 ;
  buffer buf_n450( .i (n449), .o (n450) );
  assign n451 = n426 & n450 ;
  buffer buf_n452( .i (n451), .o (n452) );
  assign n453 = n402 & n452 ;
  buffer buf_n454( .i (n453), .o (n454) );
  assign n455 = ( n194 & n210 ) | ( n194 & n228 ) | ( n210 & n228 ) ;
  buffer buf_n456( .i (n455), .o (n456) );
  assign n457 = ( n313 & n332 ) | ( n313 & n347 ) | ( n332 & n347 ) ;
  buffer buf_n458( .i (n457), .o (n458) );
  assign n459 = n456 & n458 ;
  buffer buf_n460( .i (n459), .o (n460) );
  assign n461 = ( n358 & n365 ) | ( n358 & n372 ) | ( n365 & n372 ) ;
  buffer buf_n462( .i (n461), .o (n462) );
  assign n463 = ( n381 & n388 ) | ( n381 & n395 ) | ( n388 & n395 ) ;
  buffer buf_n464( .i (n463), .o (n464) );
  assign n465 = n462 & n464 ;
  buffer buf_n466( .i (n465), .o (n466) );
  assign n467 = n460 & n466 ;
  buffer buf_n468( .i (n467), .o (n468) );
  assign n469 = ( n404 & n408 ) | ( n404 & n410 ) | ( n408 & n410 ) ;
  buffer buf_n470( .i (n469), .o (n470) );
  assign n471 = ( n415 & n418 ) | ( n415 & n421 ) | ( n418 & n421 ) ;
  buffer buf_n472( .i (n471), .o (n472) );
  assign n473 = n470 & n472 ;
  buffer buf_n474( .i (n473), .o (n474) );
  assign n475 = ( n428 & n431 ) | ( n428 & n434 ) | ( n431 & n434 ) ;
  buffer buf_n476( .i (n475), .o (n476) );
  assign n477 = ( n439 & n442 ) | ( n439 & n445 ) | ( n442 & n445 ) ;
  buffer buf_n478( .i (n477), .o (n478) );
  assign n479 = n476 & n478 ;
  buffer buf_n480( .i (n479), .o (n480) );
  assign n481 = n474 & n480 ;
  buffer buf_n482( .i (n481), .o (n482) );
  assign n483 = n468 & n482 ;
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  assign n486 = n454 & n485 ;
  assign n487 = n210 | n228 ;
  assign n488 = n195 | n487 ;
  buffer buf_n489( .i (n488), .o (n489) );
  assign n490 = n332 & n347 ;
  assign n491 = n314 & n490 ;
  buffer buf_n492( .i (n491), .o (n492) );
  assign n493 = n489 & n492 ;
  buffer buf_n494( .i (n493), .o (n494) );
  assign n495 = n365 | n372 ;
  assign n496 = n359 | n495 ;
  buffer buf_n497( .i (n496), .o (n497) );
  assign n498 = n388 & n395 ;
  assign n499 = n382 & n498 ;
  buffer buf_n500( .i (n499), .o (n500) );
  assign n501 = n497 & n500 ;
  buffer buf_n502( .i (n501), .o (n502) );
  assign n503 = n494 & n502 ;
  buffer buf_n504( .i (n503), .o (n504) );
  assign n505 = n408 | n410 ;
  assign n506 = n405 | n505 ;
  buffer buf_n507( .i (n506), .o (n507) );
  assign n508 = n418 & n421 ;
  assign n509 = n416 & n508 ;
  buffer buf_n510( .i (n509), .o (n510) );
  assign n511 = n507 & n510 ;
  buffer buf_n512( .i (n511), .o (n512) );
  assign n513 = n431 | n434 ;
  assign n514 = n429 | n513 ;
  buffer buf_n515( .i (n514), .o (n515) );
  assign n516 = n442 & n445 ;
  assign n517 = n440 & n516 ;
  buffer buf_n518( .i (n517), .o (n518) );
  assign n519 = n515 & n518 ;
  buffer buf_n520( .i (n519), .o (n520) );
  assign n521 = n512 & n520 ;
  buffer buf_n522( .i (n521), .o (n522) );
  assign n523 = n504 & n522 ;
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  assign n526 = n486 & n525 ;
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n65( .i (a_9_), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n59( .i (a_11_), .o (n59) );
  buffer buf_n99( .i (a_10_), .o (n99) );
  assign n528 = n59 & n99 ;
  assign n529 = n66 & n528 ;
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n62( .i (a_6_), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n56( .i (a_8_), .o (n56) );
  buffer buf_n74( .i (a_7_), .o (n74) );
  assign n531 = n56 | n74 ;
  assign n532 = n63 | n531 ;
  buffer buf_n533( .i (n532), .o (n533) );
  assign n534 = n530 & n533 ;
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  assign n537 = n59 | n99 ;
  assign n538 = n66 | n537 ;
  buffer buf_n539( .i (n538), .o (n539) );
  assign n540 = n56 & n74 ;
  assign n541 = n63 & n540 ;
  buffer buf_n542( .i (n541), .o (n542) );
  assign n543 = n539 & n542 ;
  buffer buf_n544( .i (n543), .o (n544) );
  assign n545 = ( n59 & n65 ) | ( n59 & n99 ) | ( n65 & n99 ) ;
  buffer buf_n546( .i (n545), .o (n546) );
  assign n547 = ( n56 & n62 ) | ( n56 & n74 ) | ( n62 & n74 ) ;
  buffer buf_n548( .i (n547), .o (n548) );
  assign n549 = n546 & n548 ;
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  assign n552 = n544 & n551 ;
  assign n553 = n536 & n552 ;
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n94( .i (a_3_), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n50( .i (a_5_), .o (n50) );
  buffer buf_n68( .i (a_4_), .o (n68) );
  assign n555 = n50 & n68 ;
  assign n556 = n95 & n555 ;
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n60( .i (a_0_), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n106( .i (a_1_), .o (n106) );
  buffer buf_n109( .i (a_2_), .o (n109) );
  assign n558 = n106 | n109 ;
  assign n559 = n61 | n558 ;
  buffer buf_n560( .i (n559), .o (n560) );
  assign n561 = n557 | n560 ;
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  assign n564 = n50 | n68 ;
  assign n565 = n95 | n564 ;
  buffer buf_n566( .i (n565), .o (n566) );
  assign n567 = n106 & n109 ;
  assign n568 = n61 & n567 ;
  buffer buf_n569( .i (n568), .o (n569) );
  assign n570 = n566 | n569 ;
  buffer buf_n571( .i (n570), .o (n571) );
  assign n572 = ( n50 & n68 ) | ( n50 & n94 ) | ( n68 & n94 ) ;
  buffer buf_n573( .i (n572), .o (n573) );
  assign n574 = ( n60 & n106 ) | ( n60 & n109 ) | ( n106 & n109 ) ;
  buffer buf_n575( .i (n574), .o (n575) );
  assign n576 = n573 | n575 ;
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  assign n579 = n571 | n578 ;
  assign n580 = n563 | n579 ;
  buffer buf_n581( .i (n580), .o (n581) );
  assign n582 = n554 & n581 ;
  buffer buf_n583( .i (n582), .o (n583) );
  assign n584 = n530 | n533 ;
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  assign n587 = n539 | n542 ;
  buffer buf_n588( .i (n587), .o (n588) );
  assign n589 = n546 | n548 ;
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  assign n592 = n588 & n591 ;
  assign n593 = n586 & n592 ;
  buffer buf_n594( .i (n593), .o (n594) );
  assign n595 = n557 & n560 ;
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  assign n598 = n566 & n569 ;
  buffer buf_n599( .i (n598), .o (n599) );
  assign n600 = n573 & n575 ;
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  assign n603 = n599 | n602 ;
  assign n604 = n597 | n603 ;
  buffer buf_n605( .i (n604), .o (n605) );
  assign n606 = n594 & n605 ;
  buffer buf_n607( .i (n606), .o (n607) );
  assign n608 = n583 & n607 ;
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  assign n611 = n544 | n551 ;
  assign n612 = n536 | n611 ;
  buffer buf_n613( .i (n612), .o (n613) );
  assign n614 = n571 & n578 ;
  assign n615 = n563 & n614 ;
  buffer buf_n616( .i (n615), .o (n616) );
  assign n617 = n613 & n616 ;
  buffer buf_n618( .i (n617), .o (n618) );
  assign n619 = n588 | n591 ;
  assign n620 = n586 | n619 ;
  buffer buf_n621( .i (n620), .o (n621) );
  assign n622 = n599 & n602 ;
  assign n623 = n597 & n622 ;
  buffer buf_n624( .i (n623), .o (n624) );
  assign n625 = n621 & n624 ;
  buffer buf_n626( .i (n625), .o (n626) );
  assign n627 = n618 & n626 ;
  buffer buf_n628( .i (n627), .o (n628) );
  assign n629 = ( n535 & n544 ) | ( n535 & n551 ) | ( n544 & n551 ) ;
  buffer buf_n630( .i (n629), .o (n630) );
  assign n631 = ( n562 & n571 ) | ( n562 & n578 ) | ( n571 & n578 ) ;
  buffer buf_n632( .i (n631), .o (n632) );
  assign n633 = n630 & n632 ;
  buffer buf_n634( .i (n633), .o (n634) );
  assign n635 = ( n585 & n588 ) | ( n585 & n591 ) | ( n588 & n591 ) ;
  buffer buf_n636( .i (n635), .o (n636) );
  assign n637 = ( n596 & n599 ) | ( n596 & n602 ) | ( n599 & n602 ) ;
  buffer buf_n638( .i (n637), .o (n638) );
  assign n639 = n636 & n638 ;
  buffer buf_n640( .i (n639), .o (n640) );
  assign n641 = n634 & n640 ;
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  assign n644 = n628 & n643 ;
  assign n645 = n610 & n644 ;
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n88( .i (a_21_), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n91( .i (a_22_), .o (n91) );
  buffer buf_n112( .i (a_23_), .o (n112) );
  assign n647 = n91 & n112 ;
  assign n648 = n89 & n647 ;
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n85( .i (a_18_), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n53( .i (a_20_), .o (n53) );
  buffer buf_n73( .i (a_19_), .o (n73) );
  assign n650 = n53 | n73 ;
  assign n651 = n86 | n650 ;
  buffer buf_n652( .i (n651), .o (n652) );
  assign n653 = n649 | n652 ;
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  assign n656 = n91 | n112 ;
  assign n657 = n89 | n656 ;
  buffer buf_n658( .i (n657), .o (n658) );
  assign n659 = n53 & n73 ;
  assign n660 = n86 & n659 ;
  buffer buf_n661( .i (n660), .o (n661) );
  assign n662 = n658 | n661 ;
  buffer buf_n663( .i (n662), .o (n663) );
  assign n664 = ( n88 & n91 ) | ( n88 & n112 ) | ( n91 & n112 ) ;
  buffer buf_n665( .i (n664), .o (n665) );
  assign n666 = ( n53 & n73 ) | ( n53 & n85 ) | ( n73 & n85 ) ;
  buffer buf_n667( .i (n666), .o (n667) );
  assign n668 = n665 | n667 ;
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  assign n671 = n663 & n670 ;
  assign n672 = n655 & n671 ;
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n107( .i (a_15_), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n64( .i (a_16_), .o (n64) );
  buffer buf_n83( .i (a_17_), .o (n83) );
  assign n674 = n64 & n83 ;
  assign n675 = n108 & n674 ;
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n100( .i (a_12_), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n75( .i (a_13_), .o (n75) );
  buffer buf_n81( .i (a_14_), .o (n81) );
  assign n677 = n75 | n81 ;
  assign n678 = n101 | n677 ;
  buffer buf_n679( .i (n678), .o (n679) );
  assign n680 = n676 & n679 ;
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  assign n683 = n64 | n83 ;
  assign n684 = n108 | n683 ;
  buffer buf_n685( .i (n684), .o (n685) );
  assign n686 = n75 & n81 ;
  assign n687 = n101 & n686 ;
  buffer buf_n688( .i (n687), .o (n688) );
  assign n689 = n685 & n688 ;
  buffer buf_n690( .i (n689), .o (n690) );
  assign n691 = ( n64 & n83 ) | ( n64 & n107 ) | ( n83 & n107 ) ;
  buffer buf_n692( .i (n691), .o (n692) );
  assign n693 = ( n75 & n81 ) | ( n75 & n100 ) | ( n81 & n100 ) ;
  buffer buf_n694( .i (n693), .o (n694) );
  assign n695 = n692 & n694 ;
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  assign n698 = n690 | n697 ;
  assign n699 = n682 | n698 ;
  buffer buf_n700( .i (n699), .o (n700) );
  assign n701 = n673 | n700 ;
  buffer buf_n702( .i (n701), .o (n702) );
  assign n703 = n649 & n652 ;
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  assign n706 = n658 & n661 ;
  buffer buf_n707( .i (n706), .o (n707) );
  assign n708 = n665 & n667 ;
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  assign n711 = n707 & n710 ;
  assign n712 = n705 & n711 ;
  buffer buf_n713( .i (n712), .o (n713) );
  assign n714 = n685 | n688 ;
  buffer buf_n715( .i (n714), .o (n715) );
  assign n716 = n692 | n694 ;
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  assign n719 = n715 | n718 ;
  assign n720 = n676 | n679 ;
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  assign n723 = n719 | n722 ;
  buffer buf_n724( .i (n723), .o (n724) );
  assign n725 = n713 | n724 ;
  buffer buf_n726( .i (n725), .o (n726) );
  assign n727 = n702 | n726 ;
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  assign n730 = n663 | n670 ;
  assign n731 = n655 | n730 ;
  buffer buf_n732( .i (n731), .o (n732) );
  assign n733 = n690 & n697 ;
  assign n734 = n682 & n733 ;
  buffer buf_n735( .i (n734), .o (n735) );
  assign n736 = n732 | n735 ;
  buffer buf_n737( .i (n736), .o (n737) );
  assign n738 = n707 | n710 ;
  assign n739 = n705 | n738 ;
  buffer buf_n740( .i (n739), .o (n740) );
  assign n741 = n715 & n718 ;
  assign n742 = n722 & n741 ;
  buffer buf_n743( .i (n742), .o (n743) );
  assign n744 = n740 | n743 ;
  buffer buf_n745( .i (n744), .o (n745) );
  assign n746 = n737 | n745 ;
  buffer buf_n747( .i (n746), .o (n747) );
  assign n748 = ( n654 & n663 ) | ( n654 & n670 ) | ( n663 & n670 ) ;
  buffer buf_n749( .i (n748), .o (n749) );
  assign n750 = ( n681 & n690 ) | ( n681 & n697 ) | ( n690 & n697 ) ;
  buffer buf_n751( .i (n750), .o (n751) );
  assign n752 = n749 | n751 ;
  buffer buf_n753( .i (n752), .o (n753) );
  assign n754 = ( n704 & n707 ) | ( n704 & n710 ) | ( n707 & n710 ) ;
  buffer buf_n755( .i (n754), .o (n755) );
  assign n756 = ( n715 & n718 ) | ( n715 & n721 ) | ( n718 & n721 ) ;
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = n755 | n757 ;
  buffer buf_n759( .i (n758), .o (n759) );
  assign n760 = n753 | n759 ;
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  assign n763 = n747 | n762 ;
  assign n764 = n729 | n763 ;
  buffer buf_n765( .i (n764), .o (n765) );
  assign n766 = n646 | n765 ;
  buffer buf_n767( .i (n766), .o (n767) );
  assign n768 = n554 | n581 ;
  buffer buf_n769( .i (n768), .o (n769) );
  assign n770 = n594 | n605 ;
  buffer buf_n771( .i (n770), .o (n771) );
  assign n772 = n769 & n771 ;
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  assign n775 = n630 | n632 ;
  buffer buf_n776( .i (n775), .o (n776) );
  assign n777 = n636 | n638 ;
  buffer buf_n778( .i (n777), .o (n778) );
  assign n779 = n776 & n778 ;
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  assign n782 = n613 | n616 ;
  buffer buf_n783( .i (n782), .o (n783) );
  assign n784 = n621 | n624 ;
  buffer buf_n785( .i (n784), .o (n785) );
  assign n786 = n783 & n785 ;
  buffer buf_n787( .i (n786), .o (n787) );
  assign n788 = n781 & n787 ;
  assign n789 = n774 & n788 ;
  buffer buf_n790( .i (n789), .o (n790) );
  assign n791 = n673 & n700 ;
  buffer buf_n792( .i (n791), .o (n792) );
  assign n793 = n713 & n724 ;
  buffer buf_n794( .i (n793), .o (n794) );
  assign n795 = n792 | n794 ;
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  assign n798 = n732 & n735 ;
  buffer buf_n799( .i (n798), .o (n799) );
  assign n800 = n740 & n743 ;
  buffer buf_n801( .i (n800), .o (n801) );
  assign n802 = n799 | n801 ;
  buffer buf_n803( .i (n802), .o (n803) );
  assign n804 = n749 & n751 ;
  buffer buf_n805( .i (n804), .o (n805) );
  assign n806 = n755 & n757 ;
  buffer buf_n807( .i (n806), .o (n807) );
  assign n808 = n805 | n807 ;
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  assign n811 = n803 | n810 ;
  assign n812 = n797 | n811 ;
  buffer buf_n813( .i (n812), .o (n813) );
  assign n814 = n790 | n813 ;
  buffer buf_n815( .i (n814), .o (n815) );
  assign n816 = n767 | n815 ;
  buffer buf_n817( .i (n816), .o (n817) );
  assign n818 = n618 | n626 ;
  buffer buf_n819( .i (n818), .o (n819) );
  assign n820 = n634 | n640 ;
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  assign n823 = n819 & n822 ;
  assign n824 = n583 | n607 ;
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  assign n827 = n823 & n826 ;
  buffer buf_n828( .i (n827), .o (n828) );
  assign n829 = n702 & n726 ;
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  assign n832 = n737 & n745 ;
  buffer buf_n833( .i (n832), .o (n833) );
  assign n834 = n753 & n759 ;
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  assign n837 = n833 | n836 ;
  assign n838 = n831 | n837 ;
  buffer buf_n839( .i (n838), .o (n839) );
  assign n840 = n828 | n839 ;
  buffer buf_n841( .i (n840), .o (n841) );
  assign n842 = n769 | n771 ;
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  assign n845 = n776 | n778 ;
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  assign n848 = n783 | n785 ;
  buffer buf_n849( .i (n848), .o (n849) );
  assign n850 = n847 & n849 ;
  assign n851 = n844 & n850 ;
  buffer buf_n852( .i (n851), .o (n852) );
  assign n853 = n792 & n794 ;
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  assign n856 = n799 & n801 ;
  buffer buf_n857( .i (n856), .o (n857) );
  assign n858 = n805 & n807 ;
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  assign n861 = n857 | n860 ;
  assign n862 = n855 | n861 ;
  buffer buf_n863( .i (n862), .o (n863) );
  assign n864 = n852 | n863 ;
  buffer buf_n865( .i (n864), .o (n865) );
  assign n866 = n841 | n865 ;
  buffer buf_n867( .i (n866), .o (n867) );
  assign n868 = n817 | n867 ;
  buffer buf_n869( .i (n868), .o (n869) );
  assign n870 = ( n609 & n628 ) | ( n609 & n643 ) | ( n628 & n643 ) ;
  buffer buf_n871( .i (n870), .o (n871) );
  assign n872 = ( n728 & n747 ) | ( n728 & n762 ) | ( n747 & n762 ) ;
  buffer buf_n873( .i (n872), .o (n873) );
  assign n874 = n871 | n873 ;
  buffer buf_n875( .i (n874), .o (n875) );
  assign n876 = ( n773 & n781 ) | ( n773 & n787 ) | ( n781 & n787 ) ;
  buffer buf_n877( .i (n876), .o (n877) );
  assign n878 = ( n796 & n803 ) | ( n796 & n810 ) | ( n803 & n810 ) ;
  buffer buf_n879( .i (n878), .o (n879) );
  assign n880 = n877 | n879 ;
  buffer buf_n881( .i (n880), .o (n881) );
  assign n882 = n875 | n881 ;
  buffer buf_n883( .i (n882), .o (n883) );
  assign n884 = ( n819 & n822 ) | ( n819 & n825 ) | ( n822 & n825 ) ;
  buffer buf_n885( .i (n884), .o (n885) );
  assign n886 = ( n830 & n833 ) | ( n830 & n836 ) | ( n833 & n836 ) ;
  buffer buf_n887( .i (n886), .o (n887) );
  assign n888 = n885 | n887 ;
  buffer buf_n889( .i (n888), .o (n889) );
  assign n890 = ( n843 & n847 ) | ( n843 & n849 ) | ( n847 & n849 ) ;
  buffer buf_n891( .i (n890), .o (n891) );
  assign n892 = ( n854 & n857 ) | ( n854 & n860 ) | ( n857 & n860 ) ;
  buffer buf_n893( .i (n892), .o (n893) );
  assign n894 = n891 | n893 ;
  buffer buf_n895( .i (n894), .o (n895) );
  assign n896 = n889 | n895 ;
  buffer buf_n897( .i (n896), .o (n897) );
  assign n898 = n883 | n897 ;
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  assign n901 = n869 | n900 ;
  assign n902 = n628 | n643 ;
  assign n903 = n610 | n902 ;
  buffer buf_n904( .i (n903), .o (n904) );
  assign n905 = n747 & n762 ;
  assign n906 = n729 & n905 ;
  buffer buf_n907( .i (n906), .o (n907) );
  assign n908 = n904 | n907 ;
  buffer buf_n909( .i (n908), .o (n909) );
  assign n910 = n781 | n787 ;
  assign n911 = n774 | n910 ;
  buffer buf_n912( .i (n911), .o (n912) );
  assign n913 = n803 & n810 ;
  assign n914 = n797 & n913 ;
  buffer buf_n915( .i (n914), .o (n915) );
  assign n916 = n912 | n915 ;
  buffer buf_n917( .i (n916), .o (n917) );
  assign n918 = n909 | n917 ;
  buffer buf_n919( .i (n918), .o (n919) );
  assign n920 = n819 | n822 ;
  assign n921 = n826 | n920 ;
  buffer buf_n922( .i (n921), .o (n922) );
  assign n923 = n833 & n836 ;
  assign n924 = n831 & n923 ;
  buffer buf_n925( .i (n924), .o (n925) );
  assign n926 = n922 | n925 ;
  buffer buf_n927( .i (n926), .o (n927) );
  assign n928 = n847 | n849 ;
  assign n929 = n844 | n928 ;
  buffer buf_n930( .i (n929), .o (n930) );
  assign n931 = n857 & n860 ;
  assign n932 = n855 & n931 ;
  buffer buf_n933( .i (n932), .o (n933) );
  assign n934 = n930 | n933 ;
  buffer buf_n935( .i (n934), .o (n935) );
  assign n936 = n927 | n935 ;
  buffer buf_n937( .i (n936), .o (n937) );
  assign n938 = n919 | n937 ;
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  assign n941 = n901 | n940 ;
  buffer buf_n942( .i (n941), .o (n942) );
  assign n943 = n527 | n942 ;
  buffer buf_n944( .i (n943), .o (n944) );
  assign n945 = n231 | n350 ;
  buffer buf_n946( .i (n945), .o (n946) );
  assign n947 = n375 | n398 ;
  buffer buf_n948( .i (n947), .o (n948) );
  assign n949 = n946 & n948 ;
  buffer buf_n950( .i (n949), .o (n950) );
  assign n951 = n413 | n424 ;
  buffer buf_n952( .i (n951), .o (n952) );
  assign n953 = n437 | n448 ;
  buffer buf_n954( .i (n953), .o (n954) );
  assign n955 = n952 & n954 ;
  buffer buf_n956( .i (n955), .o (n956) );
  assign n957 = n950 & n956 ;
  buffer buf_n958( .i (n957), .o (n958) );
  assign n959 = n456 | n458 ;
  buffer buf_n960( .i (n959), .o (n960) );
  assign n961 = n462 | n464 ;
  buffer buf_n962( .i (n961), .o (n962) );
  assign n963 = n960 & n962 ;
  buffer buf_n964( .i (n963), .o (n964) );
  assign n965 = n470 | n472 ;
  buffer buf_n966( .i (n965), .o (n966) );
  assign n967 = n476 | n478 ;
  buffer buf_n968( .i (n967), .o (n968) );
  assign n969 = n966 & n968 ;
  buffer buf_n970( .i (n969), .o (n970) );
  assign n971 = n964 & n970 ;
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  assign n974 = n958 & n973 ;
  assign n975 = n489 | n492 ;
  buffer buf_n976( .i (n975), .o (n976) );
  assign n977 = n497 | n500 ;
  buffer buf_n978( .i (n977), .o (n978) );
  assign n979 = n976 & n978 ;
  buffer buf_n980( .i (n979), .o (n980) );
  assign n981 = n507 | n510 ;
  buffer buf_n982( .i (n981), .o (n982) );
  assign n983 = n515 | n518 ;
  buffer buf_n984( .i (n983), .o (n984) );
  assign n985 = n982 & n984 ;
  buffer buf_n986( .i (n985), .o (n986) );
  assign n987 = n980 & n986 ;
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  assign n990 = n974 & n989 ;
  buffer buf_n991( .i (n990), .o (n991) );
  assign n992 = n646 & n765 ;
  buffer buf_n993( .i (n992), .o (n993) );
  assign n994 = n790 & n813 ;
  buffer buf_n995( .i (n994), .o (n995) );
  assign n996 = n993 | n995 ;
  buffer buf_n997( .i (n996), .o (n997) );
  assign n998 = n828 & n839 ;
  buffer buf_n999( .i (n998), .o (n999) );
  assign n1000 = n852 & n863 ;
  buffer buf_n1001( .i (n1000), .o (n1001) );
  assign n1002 = n999 | n1001 ;
  buffer buf_n1003( .i (n1002), .o (n1003) );
  assign n1004 = n997 | n1003 ;
  buffer buf_n1005( .i (n1004), .o (n1005) );
  assign n1006 = n871 & n873 ;
  buffer buf_n1007( .i (n1006), .o (n1007) );
  assign n1008 = n877 & n879 ;
  buffer buf_n1009( .i (n1008), .o (n1009) );
  assign n1010 = n1007 | n1009 ;
  buffer buf_n1011( .i (n1010), .o (n1011) );
  assign n1012 = n885 & n887 ;
  buffer buf_n1013( .i (n1012), .o (n1013) );
  assign n1014 = n891 & n893 ;
  buffer buf_n1015( .i (n1014), .o (n1015) );
  assign n1016 = n1013 | n1015 ;
  buffer buf_n1017( .i (n1016), .o (n1017) );
  assign n1018 = n1011 | n1017 ;
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  assign n1021 = n1005 | n1020 ;
  assign n1022 = n904 & n907 ;
  buffer buf_n1023( .i (n1022), .o (n1023) );
  assign n1024 = n912 & n915 ;
  buffer buf_n1025( .i (n1024), .o (n1025) );
  assign n1026 = n1023 | n1025 ;
  buffer buf_n1027( .i (n1026), .o (n1027) );
  assign n1028 = n922 & n925 ;
  buffer buf_n1029( .i (n1028), .o (n1029) );
  assign n1030 = n930 & n933 ;
  buffer buf_n1031( .i (n1030), .o (n1031) );
  assign n1032 = n1029 | n1031 ;
  buffer buf_n1033( .i (n1032), .o (n1033) );
  assign n1034 = n1027 | n1033 ;
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  assign n1037 = n1021 | n1036 ;
  buffer buf_n1038( .i (n1037), .o (n1038) );
  assign n1039 = n991 | n1038 ;
  buffer buf_n1040( .i (n1039), .o (n1040) );
  assign n1041 = n944 | n1040 ;
  buffer buf_n1042( .i (n1041), .o (n1042) );
  assign n1043 = n352 | n400 ;
  buffer buf_n1044( .i (n1043), .o (n1044) );
  assign n1045 = n426 | n450 ;
  buffer buf_n1046( .i (n1045), .o (n1046) );
  assign n1047 = n1044 & n1046 ;
  buffer buf_n1048( .i (n1047), .o (n1048) );
  assign n1049 = n460 | n466 ;
  buffer buf_n1050( .i (n1049), .o (n1050) );
  assign n1051 = n474 | n480 ;
  buffer buf_n1052( .i (n1051), .o (n1052) );
  assign n1053 = n1050 & n1052 ;
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  assign n1056 = n1048 & n1055 ;
  assign n1057 = n494 | n502 ;
  buffer buf_n1058( .i (n1057), .o (n1058) );
  assign n1059 = n512 | n520 ;
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1061 = n1058 & n1060 ;
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  assign n1064 = n1056 & n1063 ;
  buffer buf_n1065( .i (n1064), .o (n1065) );
  assign n1066 = n767 & n815 ;
  buffer buf_n1067( .i (n1066), .o (n1067) );
  assign n1068 = n841 & n865 ;
  buffer buf_n1069( .i (n1068), .o (n1069) );
  assign n1070 = n1067 | n1069 ;
  buffer buf_n1071( .i (n1070), .o (n1071) );
  assign n1072 = n875 & n881 ;
  buffer buf_n1073( .i (n1072), .o (n1073) );
  assign n1074 = n889 & n895 ;
  buffer buf_n1075( .i (n1074), .o (n1075) );
  assign n1076 = n1073 | n1075 ;
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  assign n1079 = n1071 | n1078 ;
  assign n1080 = n909 & n917 ;
  buffer buf_n1081( .i (n1080), .o (n1081) );
  assign n1082 = n927 & n935 ;
  buffer buf_n1083( .i (n1082), .o (n1083) );
  assign n1084 = n1081 | n1083 ;
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  assign n1087 = n1079 | n1086 ;
  buffer buf_n1088( .i (n1087), .o (n1088) );
  assign n1089 = n1065 | n1088 ;
  buffer buf_n1090( .i (n1089), .o (n1090) );
  assign n1091 = n946 | n948 ;
  buffer buf_n1092( .i (n1091), .o (n1092) );
  assign n1093 = n952 | n954 ;
  buffer buf_n1094( .i (n1093), .o (n1094) );
  assign n1095 = n1092 & n1094 ;
  buffer buf_n1096( .i (n1095), .o (n1096) );
  assign n1097 = n960 | n962 ;
  buffer buf_n1098( .i (n1097), .o (n1098) );
  assign n1099 = n966 | n968 ;
  buffer buf_n1100( .i (n1099), .o (n1100) );
  assign n1101 = n1098 & n1100 ;
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  assign n1104 = n1096 & n1103 ;
  assign n1105 = n976 | n978 ;
  buffer buf_n1106( .i (n1105), .o (n1106) );
  assign n1107 = n982 | n984 ;
  buffer buf_n1108( .i (n1107), .o (n1108) );
  assign n1109 = n1106 & n1108 ;
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  assign n1112 = n1104 & n1111 ;
  buffer buf_n1113( .i (n1112), .o (n1113) );
  assign n1114 = n993 & n995 ;
  buffer buf_n1115( .i (n1114), .o (n1115) );
  assign n1116 = n999 & n1001 ;
  buffer buf_n1117( .i (n1116), .o (n1117) );
  assign n1118 = n1115 | n1117 ;
  buffer buf_n1119( .i (n1118), .o (n1119) );
  assign n1120 = n1007 & n1009 ;
  buffer buf_n1121( .i (n1120), .o (n1121) );
  assign n1122 = n1013 & n1015 ;
  buffer buf_n1123( .i (n1122), .o (n1123) );
  assign n1124 = n1121 | n1123 ;
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  assign n1127 = n1119 | n1126 ;
  assign n1128 = n1023 & n1025 ;
  buffer buf_n1129( .i (n1128), .o (n1129) );
  assign n1130 = n1029 & n1031 ;
  buffer buf_n1131( .i (n1130), .o (n1131) );
  assign n1132 = n1129 | n1131 ;
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  assign n1135 = n1127 | n1134 ;
  buffer buf_n1136( .i (n1135), .o (n1136) );
  assign n1137 = n1113 | n1136 ;
  buffer buf_n1138( .i (n1137), .o (n1138) );
  assign n1139 = n1090 | n1138 ;
  buffer buf_n1140( .i (n1139), .o (n1140) );
  assign n1141 = n1042 | n1140 ;
  buffer buf_n1142( .i (n1141), .o (n1142) );
  assign n1143 = n402 | n452 ;
  buffer buf_n1144( .i (n1143), .o (n1144) );
  assign n1145 = n468 | n482 ;
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  assign n1148 = n1144 & n1147 ;
  assign n1149 = n504 | n522 ;
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  assign n1152 = n1148 & n1151 ;
  buffer buf_n1153( .i (n1152), .o (n1153) );
  assign n1154 = n817 & n867 ;
  buffer buf_n1155( .i (n1154), .o (n1155) );
  assign n1156 = n883 & n897 ;
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  assign n1159 = n1155 | n1158 ;
  assign n1160 = n919 & n937 ;
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  assign n1163 = n1159 | n1162 ;
  buffer buf_n1164( .i (n1163), .o (n1164) );
  assign n1165 = n1153 | n1164 ;
  buffer buf_n1166( .i (n1165), .o (n1166) );
  assign n1167 = n950 | n956 ;
  buffer buf_n1168( .i (n1167), .o (n1168) );
  assign n1169 = n964 | n970 ;
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  assign n1172 = n1168 & n1171 ;
  assign n1173 = n980 | n986 ;
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  assign n1176 = n1172 & n1175 ;
  buffer buf_n1177( .i (n1176), .o (n1177) );
  assign n1178 = n997 & n1003 ;
  buffer buf_n1179( .i (n1178), .o (n1179) );
  assign n1180 = n1011 & n1017 ;
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  assign n1183 = n1179 | n1182 ;
  assign n1184 = n1027 & n1033 ;
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  assign n1187 = n1183 | n1186 ;
  buffer buf_n1188( .i (n1187), .o (n1188) );
  assign n1189 = n1177 | n1188 ;
  buffer buf_n1190( .i (n1189), .o (n1190) );
  assign n1191 = n1166 | n1190 ;
  buffer buf_n1192( .i (n1191), .o (n1192) );
  assign n1193 = n1044 | n1046 ;
  buffer buf_n1194( .i (n1193), .o (n1194) );
  assign n1195 = n1050 | n1052 ;
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  assign n1198 = n1194 & n1197 ;
  assign n1199 = n1058 | n1060 ;
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  assign n1202 = n1198 & n1201 ;
  buffer buf_n1203( .i (n1202), .o (n1203) );
  assign n1204 = n1067 & n1069 ;
  buffer buf_n1205( .i (n1204), .o (n1205) );
  assign n1206 = n1073 & n1075 ;
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  assign n1209 = n1205 | n1208 ;
  assign n1210 = n1081 & n1083 ;
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  assign n1213 = n1209 | n1212 ;
  buffer buf_n1214( .i (n1213), .o (n1214) );
  assign n1215 = n1203 | n1214 ;
  buffer buf_n1216( .i (n1215), .o (n1216) );
  assign n1217 = n1092 | n1094 ;
  buffer buf_n1218( .i (n1217), .o (n1218) );
  assign n1219 = n1098 | n1100 ;
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  assign n1222 = n1218 & n1221 ;
  assign n1223 = n1106 | n1108 ;
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  assign n1226 = n1222 & n1225 ;
  buffer buf_n1227( .i (n1226), .o (n1227) );
  assign n1228 = n1115 & n1117 ;
  buffer buf_n1229( .i (n1228), .o (n1229) );
  assign n1230 = n1121 & n1123 ;
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  assign n1233 = n1229 | n1232 ;
  assign n1234 = n1129 & n1131 ;
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  assign n1237 = n1233 | n1236 ;
  buffer buf_n1238( .i (n1237), .o (n1238) );
  assign n1239 = n1227 | n1238 ;
  buffer buf_n1240( .i (n1239), .o (n1240) );
  assign n1241 = n1216 | n1240 ;
  buffer buf_n1242( .i (n1241), .o (n1242) );
  assign n1243 = n1192 | n1242 ;
  buffer buf_n1244( .i (n1243), .o (n1244) );
  assign n1245 = n1142 | n1244 ;
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n1247( .i (n1246), .o (n1247) );
  assign n1248 = ( n454 & n485 ) | ( n454 & n524 ) | ( n485 & n524 ) ;
  buffer buf_n1249( .i (n1248), .o (n1249) );
  assign n1250 = ( n869 & n900 ) | ( n869 & n939 ) | ( n900 & n939 ) ;
  buffer buf_n1251( .i (n1250), .o (n1251) );
  assign n1252 = n1249 | n1251 ;
  buffer buf_n1253( .i (n1252), .o (n1253) );
  assign n1254 = ( n958 & n973 ) | ( n958 & n988 ) | ( n973 & n988 ) ;
  buffer buf_n1255( .i (n1254), .o (n1255) );
  assign n1256 = ( n1005 & n1020 ) | ( n1005 & n1035 ) | ( n1020 & n1035 ) ;
  buffer buf_n1257( .i (n1256), .o (n1257) );
  assign n1258 = n1255 | n1257 ;
  buffer buf_n1259( .i (n1258), .o (n1259) );
  assign n1260 = n1253 | n1259 ;
  buffer buf_n1261( .i (n1260), .o (n1261) );
  assign n1262 = ( n1048 & n1055 ) | ( n1048 & n1062 ) | ( n1055 & n1062 ) ;
  buffer buf_n1263( .i (n1262), .o (n1263) );
  assign n1264 = ( n1071 & n1078 ) | ( n1071 & n1085 ) | ( n1078 & n1085 ) ;
  buffer buf_n1265( .i (n1264), .o (n1265) );
  assign n1266 = n1263 | n1265 ;
  buffer buf_n1267( .i (n1266), .o (n1267) );
  assign n1268 = ( n1096 & n1103 ) | ( n1096 & n1110 ) | ( n1103 & n1110 ) ;
  buffer buf_n1269( .i (n1268), .o (n1269) );
  assign n1270 = ( n1119 & n1126 ) | ( n1119 & n1133 ) | ( n1126 & n1133 ) ;
  buffer buf_n1271( .i (n1270), .o (n1271) );
  assign n1272 = n1269 | n1271 ;
  buffer buf_n1273( .i (n1272), .o (n1273) );
  assign n1274 = n1267 | n1273 ;
  buffer buf_n1275( .i (n1274), .o (n1275) );
  assign n1276 = n1261 | n1275 ;
  buffer buf_n1277( .i (n1276), .o (n1277) );
  assign n1278 = ( n1144 & n1147 ) | ( n1144 & n1150 ) | ( n1147 & n1150 ) ;
  buffer buf_n1279( .i (n1278), .o (n1279) );
  assign n1280 = ( n1155 & n1158 ) | ( n1155 & n1161 ) | ( n1158 & n1161 ) ;
  buffer buf_n1281( .i (n1280), .o (n1281) );
  assign n1282 = n1279 | n1281 ;
  buffer buf_n1283( .i (n1282), .o (n1283) );
  assign n1284 = ( n1168 & n1171 ) | ( n1168 & n1174 ) | ( n1171 & n1174 ) ;
  buffer buf_n1285( .i (n1284), .o (n1285) );
  assign n1286 = ( n1179 & n1182 ) | ( n1179 & n1185 ) | ( n1182 & n1185 ) ;
  buffer buf_n1287( .i (n1286), .o (n1287) );
  assign n1288 = n1285 | n1287 ;
  buffer buf_n1289( .i (n1288), .o (n1289) );
  assign n1290 = n1283 | n1289 ;
  buffer buf_n1291( .i (n1290), .o (n1291) );
  assign n1292 = ( n1194 & n1197 ) | ( n1194 & n1200 ) | ( n1197 & n1200 ) ;
  buffer buf_n1293( .i (n1292), .o (n1293) );
  assign n1294 = ( n1205 & n1208 ) | ( n1205 & n1211 ) | ( n1208 & n1211 ) ;
  buffer buf_n1295( .i (n1294), .o (n1295) );
  assign n1296 = n1293 | n1295 ;
  buffer buf_n1297( .i (n1296), .o (n1297) );
  assign n1298 = ( n1218 & n1221 ) | ( n1218 & n1224 ) | ( n1221 & n1224 ) ;
  buffer buf_n1299( .i (n1298), .o (n1299) );
  assign n1300 = ( n1229 & n1232 ) | ( n1229 & n1235 ) | ( n1232 & n1235 ) ;
  buffer buf_n1301( .i (n1300), .o (n1301) );
  assign n1302 = n1299 | n1301 ;
  buffer buf_n1303( .i (n1302), .o (n1303) );
  assign n1304 = n1297 | n1303 ;
  buffer buf_n1305( .i (n1304), .o (n1305) );
  assign n1306 = n1291 | n1305 ;
  buffer buf_n1307( .i (n1306), .o (n1307) );
  assign n1308 = n1277 | n1307 ;
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  assign n1311 = n454 | n485 ;
  assign n1312 = n525 | n1311 ;
  buffer buf_n1313( .i (n1312), .o (n1313) );
  assign n1314 = n869 & n900 ;
  assign n1315 = n940 & n1314 ;
  buffer buf_n1316( .i (n1315), .o (n1316) );
  assign n1317 = n1313 | n1316 ;
  buffer buf_n1318( .i (n1317), .o (n1318) );
  assign n1319 = n958 | n973 ;
  assign n1320 = n989 | n1319 ;
  buffer buf_n1321( .i (n1320), .o (n1321) );
  assign n1322 = n1005 & n1020 ;
  assign n1323 = n1036 & n1322 ;
  buffer buf_n1324( .i (n1323), .o (n1324) );
  assign n1325 = n1321 | n1324 ;
  buffer buf_n1326( .i (n1325), .o (n1326) );
  assign n1327 = n1318 | n1326 ;
  buffer buf_n1328( .i (n1327), .o (n1328) );
  assign n1329 = n1048 | n1055 ;
  assign n1330 = n1063 | n1329 ;
  buffer buf_n1331( .i (n1330), .o (n1331) );
  assign n1332 = n1071 & n1078 ;
  assign n1333 = n1086 & n1332 ;
  buffer buf_n1334( .i (n1333), .o (n1334) );
  assign n1335 = n1331 | n1334 ;
  buffer buf_n1336( .i (n1335), .o (n1336) );
  assign n1337 = n1096 | n1103 ;
  assign n1338 = n1111 | n1337 ;
  buffer buf_n1339( .i (n1338), .o (n1339) );
  assign n1340 = n1119 & n1126 ;
  assign n1341 = n1134 & n1340 ;
  buffer buf_n1342( .i (n1341), .o (n1342) );
  assign n1343 = n1339 | n1342 ;
  buffer buf_n1344( .i (n1343), .o (n1344) );
  assign n1345 = n1336 | n1344 ;
  buffer buf_n1346( .i (n1345), .o (n1346) );
  assign n1347 = n1328 | n1346 ;
  buffer buf_n1348( .i (n1347), .o (n1348) );
  assign n1349 = n1144 | n1147 ;
  assign n1350 = n1151 | n1349 ;
  buffer buf_n1351( .i (n1350), .o (n1351) );
  assign n1352 = n1155 & n1158 ;
  assign n1353 = n1162 & n1352 ;
  buffer buf_n1354( .i (n1353), .o (n1354) );
  assign n1355 = n1351 | n1354 ;
  buffer buf_n1356( .i (n1355), .o (n1356) );
  assign n1357 = n1168 | n1171 ;
  assign n1358 = n1175 | n1357 ;
  buffer buf_n1359( .i (n1358), .o (n1359) );
  assign n1360 = n1179 & n1182 ;
  assign n1361 = n1186 & n1360 ;
  buffer buf_n1362( .i (n1361), .o (n1362) );
  assign n1363 = n1359 | n1362 ;
  buffer buf_n1364( .i (n1363), .o (n1364) );
  assign n1365 = n1356 | n1364 ;
  buffer buf_n1366( .i (n1365), .o (n1366) );
  assign n1367 = n1194 | n1197 ;
  assign n1368 = n1201 | n1367 ;
  buffer buf_n1369( .i (n1368), .o (n1369) );
  assign n1370 = n1205 & n1208 ;
  assign n1371 = n1212 & n1370 ;
  buffer buf_n1372( .i (n1371), .o (n1372) );
  assign n1373 = n1369 | n1372 ;
  buffer buf_n1374( .i (n1373), .o (n1374) );
  assign n1375 = n1218 | n1221 ;
  assign n1376 = n1225 | n1375 ;
  buffer buf_n1377( .i (n1376), .o (n1377) );
  assign n1378 = n1229 & n1232 ;
  assign n1379 = n1236 & n1378 ;
  buffer buf_n1380( .i (n1379), .o (n1380) );
  assign n1381 = n1377 | n1380 ;
  buffer buf_n1382( .i (n1381), .o (n1382) );
  assign n1383 = n1374 | n1382 ;
  buffer buf_n1384( .i (n1383), .o (n1384) );
  assign n1385 = n1366 | n1384 ;
  buffer buf_n1386( .i (n1385), .o (n1386) );
  assign n1387 = n1348 | n1386 ;
  buffer buf_n1388( .i (n1387), .o (n1388) );
  assign n1389 = n1310 | n1388 ;
  assign n1390 = n1247 | n1389 ;
  assign n1391 = n1142 & n1244 ;
  buffer buf_n1392( .i (n1391), .o (n1392) );
  assign n1394 = n1277 & n1307 ;
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  assign n1397 = n1348 & n1386 ;
  buffer buf_n1398( .i (n1397), .o (n1398) );
  assign n1399 = ( n1392 & n1396 ) | ( n1392 & n1398 ) | ( n1396 & n1398 ) ;
  assign n1400 = n1042 & n1140 ;
  buffer buf_n1401( .i (n1400), .o (n1401) );
  assign n1402 = n1192 & n1242 ;
  buffer buf_n1403( .i (n1402), .o (n1403) );
  assign n1404 = n1401 | n1403 ;
  buffer buf_n1405( .i (n1404), .o (n1405) );
  assign n1407 = n1261 & n1275 ;
  buffer buf_n1408( .i (n1407), .o (n1408) );
  assign n1409 = n1291 & n1305 ;
  buffer buf_n1410( .i (n1409), .o (n1410) );
  assign n1411 = n1408 | n1410 ;
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  assign n1414 = n1328 & n1346 ;
  buffer buf_n1415( .i (n1414), .o (n1415) );
  assign n1416 = n1366 & n1384 ;
  buffer buf_n1417( .i (n1416), .o (n1417) );
  assign n1418 = n1415 | n1417 ;
  buffer buf_n1419( .i (n1418), .o (n1419) );
  assign n1420 = ( n1405 & n1413 ) | ( n1405 & n1419 ) | ( n1413 & n1419 ) ;
  assign n1421 = n527 & n942 ;
  buffer buf_n1422( .i (n1421), .o (n1422) );
  assign n1423 = n991 & n1038 ;
  buffer buf_n1424( .i (n1423), .o (n1424) );
  assign n1425 = n1422 & n1424 ;
  buffer buf_n1426( .i (n1425), .o (n1426) );
  assign n1427 = n1065 & n1088 ;
  buffer buf_n1428( .i (n1427), .o (n1428) );
  assign n1429 = n1113 & n1136 ;
  buffer buf_n1430( .i (n1429), .o (n1430) );
  assign n1431 = n1428 & n1430 ;
  buffer buf_n1432( .i (n1431), .o (n1432) );
  assign n1433 = n1426 | n1432 ;
  buffer buf_n1434( .i (n1433), .o (n1434) );
  assign n1435 = n1153 & n1164 ;
  buffer buf_n1436( .i (n1435), .o (n1436) );
  assign n1437 = n1177 & n1188 ;
  buffer buf_n1438( .i (n1437), .o (n1438) );
  assign n1439 = n1436 & n1438 ;
  buffer buf_n1440( .i (n1439), .o (n1440) );
  assign n1441 = n1203 & n1214 ;
  buffer buf_n1442( .i (n1441), .o (n1442) );
  assign n1443 = n1227 & n1238 ;
  buffer buf_n1444( .i (n1443), .o (n1444) );
  assign n1445 = n1442 & n1444 ;
  buffer buf_n1446( .i (n1445), .o (n1446) );
  assign n1447 = n1440 | n1446 ;
  buffer buf_n1448( .i (n1447), .o (n1448) );
  assign n1449 = n1434 | n1448 ;
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  assign n1452 = n1249 & n1251 ;
  buffer buf_n1453( .i (n1452), .o (n1453) );
  assign n1454 = n1255 & n1257 ;
  buffer buf_n1455( .i (n1454), .o (n1455) );
  assign n1456 = n1453 & n1455 ;
  buffer buf_n1457( .i (n1456), .o (n1457) );
  assign n1458 = n1263 & n1265 ;
  buffer buf_n1459( .i (n1458), .o (n1459) );
  assign n1460 = n1269 & n1271 ;
  buffer buf_n1461( .i (n1460), .o (n1461) );
  assign n1462 = n1459 & n1461 ;
  buffer buf_n1463( .i (n1462), .o (n1463) );
  assign n1464 = n1457 | n1463 ;
  buffer buf_n1465( .i (n1464), .o (n1465) );
  assign n1466 = n1279 & n1281 ;
  buffer buf_n1467( .i (n1466), .o (n1467) );
  assign n1468 = n1285 & n1287 ;
  buffer buf_n1469( .i (n1468), .o (n1469) );
  assign n1470 = n1467 & n1469 ;
  buffer buf_n1471( .i (n1470), .o (n1471) );
  assign n1472 = n1293 & n1295 ;
  buffer buf_n1473( .i (n1472), .o (n1473) );
  assign n1474 = n1299 & n1301 ;
  buffer buf_n1475( .i (n1474), .o (n1475) );
  assign n1476 = n1473 & n1475 ;
  buffer buf_n1477( .i (n1476), .o (n1477) );
  assign n1478 = n1471 | n1477 ;
  buffer buf_n1479( .i (n1478), .o (n1479) );
  assign n1480 = n1465 | n1479 ;
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  assign n1483 = n1313 & n1316 ;
  buffer buf_n1484( .i (n1483), .o (n1484) );
  assign n1485 = n1321 & n1324 ;
  buffer buf_n1486( .i (n1485), .o (n1486) );
  assign n1487 = n1484 & n1486 ;
  buffer buf_n1488( .i (n1487), .o (n1488) );
  assign n1489 = n1331 & n1334 ;
  buffer buf_n1490( .i (n1489), .o (n1490) );
  assign n1491 = n1339 & n1342 ;
  buffer buf_n1492( .i (n1491), .o (n1492) );
  assign n1493 = n1490 & n1492 ;
  buffer buf_n1494( .i (n1493), .o (n1494) );
  assign n1495 = n1488 | n1494 ;
  buffer buf_n1496( .i (n1495), .o (n1496) );
  assign n1497 = n1351 & n1354 ;
  buffer buf_n1498( .i (n1497), .o (n1498) );
  assign n1499 = n1359 & n1362 ;
  buffer buf_n1500( .i (n1499), .o (n1500) );
  assign n1501 = n1498 & n1500 ;
  buffer buf_n1502( .i (n1501), .o (n1502) );
  assign n1503 = n1369 & n1372 ;
  buffer buf_n1504( .i (n1503), .o (n1504) );
  assign n1505 = n1377 & n1380 ;
  buffer buf_n1506( .i (n1505), .o (n1506) );
  assign n1507 = n1504 & n1506 ;
  buffer buf_n1508( .i (n1507), .o (n1508) );
  assign n1509 = n1502 | n1508 ;
  buffer buf_n1510( .i (n1509), .o (n1510) );
  assign n1511 = n1496 | n1510 ;
  buffer buf_n1512( .i (n1511), .o (n1512) );
  assign n1513 = n1482 | n1512 ;
  assign n1514 = n1451 | n1513 ;
  assign n1515 = n1434 & n1448 ;
  buffer buf_n1516( .i (n1515), .o (n1516) );
  assign n1518 = n1465 & n1479 ;
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  assign n1521 = n1496 & n1510 ;
  buffer buf_n1522( .i (n1521), .o (n1522) );
  assign n1523 = ( n1516 & n1520 ) | ( n1516 & n1522 ) | ( n1520 & n1522 ) ;
  assign n1524 = n1426 & n1432 ;
  buffer buf_n1525( .i (n1524), .o (n1525) );
  assign n1526 = n1440 & n1446 ;
  buffer buf_n1527( .i (n1526), .o (n1527) );
  assign n1528 = n1525 | n1527 ;
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  assign n1531 = n1457 & n1463 ;
  buffer buf_n1532( .i (n1531), .o (n1532) );
  assign n1533 = n1471 & n1477 ;
  buffer buf_n1534( .i (n1533), .o (n1534) );
  assign n1535 = n1532 | n1534 ;
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  assign n1538 = n1488 & n1494 ;
  buffer buf_n1539( .i (n1538), .o (n1539) );
  assign n1540 = n1502 & n1508 ;
  buffer buf_n1541( .i (n1540), .o (n1541) );
  assign n1542 = n1539 | n1541 ;
  buffer buf_n1543( .i (n1542), .o (n1543) );
  assign n1544 = n1537 | n1543 ;
  assign n1545 = n1530 | n1544 ;
  assign n1546 = n944 & n1040 ;
  buffer buf_n1547( .i (n1546), .o (n1547) );
  assign n1548 = n1090 & n1138 ;
  buffer buf_n1549( .i (n1548), .o (n1549) );
  assign n1550 = n1547 | n1549 ;
  buffer buf_n1551( .i (n1550), .o (n1551) );
  assign n1552 = n1166 & n1190 ;
  buffer buf_n1553( .i (n1552), .o (n1553) );
  assign n1554 = n1216 & n1240 ;
  buffer buf_n1555( .i (n1554), .o (n1555) );
  assign n1556 = n1553 | n1555 ;
  buffer buf_n1557( .i (n1556), .o (n1557) );
  assign n1558 = n1551 & n1557 ;
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  assign n1561 = n1253 & n1259 ;
  buffer buf_n1562( .i (n1561), .o (n1562) );
  assign n1563 = n1267 & n1273 ;
  buffer buf_n1564( .i (n1563), .o (n1564) );
  assign n1565 = n1562 | n1564 ;
  buffer buf_n1566( .i (n1565), .o (n1566) );
  assign n1567 = n1283 & n1289 ;
  buffer buf_n1568( .i (n1567), .o (n1568) );
  assign n1569 = n1297 & n1303 ;
  buffer buf_n1570( .i (n1569), .o (n1570) );
  assign n1571 = n1568 | n1570 ;
  buffer buf_n1572( .i (n1571), .o (n1572) );
  assign n1573 = n1566 & n1572 ;
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  assign n1576 = n1318 & n1326 ;
  buffer buf_n1577( .i (n1576), .o (n1577) );
  assign n1578 = n1336 & n1344 ;
  buffer buf_n1579( .i (n1578), .o (n1579) );
  assign n1580 = n1577 | n1579 ;
  buffer buf_n1581( .i (n1580), .o (n1581) );
  assign n1582 = n1356 & n1364 ;
  buffer buf_n1583( .i (n1582), .o (n1583) );
  assign n1584 = n1374 & n1382 ;
  buffer buf_n1585( .i (n1584), .o (n1585) );
  assign n1586 = n1583 | n1585 ;
  buffer buf_n1587( .i (n1586), .o (n1587) );
  assign n1588 = n1581 & n1587 ;
  buffer buf_n1589( .i (n1588), .o (n1589) );
  assign n1590 = n1575 | n1589 ;
  assign n1591 = n1560 | n1590 ;
  assign n1592 = n1422 | n1424 ;
  buffer buf_n1593( .i (n1592), .o (n1593) );
  assign n1594 = n1428 | n1430 ;
  buffer buf_n1595( .i (n1594), .o (n1595) );
  assign n1596 = n1593 & n1595 ;
  buffer buf_n1597( .i (n1596), .o (n1597) );
  assign n1598 = n1436 | n1438 ;
  buffer buf_n1599( .i (n1598), .o (n1599) );
  assign n1600 = n1442 | n1444 ;
  buffer buf_n1601( .i (n1600), .o (n1601) );
  assign n1602 = n1599 & n1601 ;
  buffer buf_n1603( .i (n1602), .o (n1603) );
  assign n1604 = n1597 | n1603 ;
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  assign n1607 = n1453 | n1455 ;
  buffer buf_n1608( .i (n1607), .o (n1608) );
  assign n1609 = n1459 | n1461 ;
  buffer buf_n1610( .i (n1609), .o (n1610) );
  assign n1611 = n1608 & n1610 ;
  buffer buf_n1612( .i (n1611), .o (n1612) );
  assign n1613 = n1467 | n1469 ;
  buffer buf_n1614( .i (n1613), .o (n1614) );
  assign n1615 = n1473 | n1475 ;
  buffer buf_n1616( .i (n1615), .o (n1616) );
  assign n1617 = n1614 & n1616 ;
  buffer buf_n1618( .i (n1617), .o (n1618) );
  assign n1619 = n1612 | n1618 ;
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n1621( .i (n1620), .o (n1621) );
  assign n1622 = n1484 | n1486 ;
  buffer buf_n1623( .i (n1622), .o (n1623) );
  assign n1624 = n1490 | n1492 ;
  buffer buf_n1625( .i (n1624), .o (n1625) );
  assign n1626 = n1623 & n1625 ;
  buffer buf_n1627( .i (n1626), .o (n1627) );
  assign n1628 = n1498 | n1500 ;
  buffer buf_n1629( .i (n1628), .o (n1629) );
  assign n1630 = n1504 | n1506 ;
  buffer buf_n1631( .i (n1630), .o (n1631) );
  assign n1632 = n1629 & n1631 ;
  buffer buf_n1633( .i (n1632), .o (n1633) );
  assign n1634 = n1627 | n1633 ;
  buffer buf_n1635( .i (n1634), .o (n1635) );
  assign n1636 = n1621 | n1635 ;
  assign n1637 = n1606 | n1636 ;
  assign n1638 = n1547 & n1549 ;
  buffer buf_n1639( .i (n1638), .o (n1639) );
  assign n1640 = n1553 & n1555 ;
  buffer buf_n1641( .i (n1640), .o (n1641) );
  assign n1642 = n1639 | n1641 ;
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  assign n1645 = n1562 & n1564 ;
  buffer buf_n1646( .i (n1645), .o (n1646) );
  assign n1647 = n1568 & n1570 ;
  buffer buf_n1648( .i (n1647), .o (n1648) );
  assign n1649 = n1646 | n1648 ;
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  assign n1652 = n1577 & n1579 ;
  buffer buf_n1653( .i (n1652), .o (n1653) );
  assign n1654 = n1583 & n1585 ;
  buffer buf_n1655( .i (n1654), .o (n1655) );
  assign n1656 = n1653 | n1655 ;
  buffer buf_n1657( .i (n1656), .o (n1657) );
  assign n1658 = n1651 | n1657 ;
  assign n1659 = n1644 | n1658 ;
  assign n1660 = n1639 & n1641 ;
  buffer buf_n1661( .i (n1660), .o (n1661) );
  assign n1663 = n1646 & n1648 ;
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  assign n1666 = n1653 & n1655 ;
  buffer buf_n1667( .i (n1666), .o (n1667) );
  assign n1668 = ( n1661 & n1665 ) | ( n1661 & n1667 ) | ( n1665 & n1667 ) ;
  assign n1669 = n1597 & n1603 ;
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  assign n1672 = n1612 & n1618 ;
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  assign n1675 = n1627 & n1633 ;
  buffer buf_n1676( .i (n1675), .o (n1676) );
  assign n1677 = n1674 & n1676 ;
  assign n1678 = n1671 & n1677 ;
  assign n1679 = ( n1605 & n1621 ) | ( n1605 & n1635 ) | ( n1621 & n1635 ) ;
  assign n1680 = n1525 & n1527 ;
  buffer buf_n1681( .i (n1680), .o (n1681) );
  assign n1683 = n1532 & n1534 ;
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  assign n1686 = n1539 & n1541 ;
  buffer buf_n1687( .i (n1686), .o (n1687) );
  assign n1688 = ( n1681 & n1685 ) | ( n1681 & n1687 ) | ( n1685 & n1687 ) ;
  buffer buf_n1393( .i (n1392), .o (n1393) );
  assign n1689 = n1396 & n1398 ;
  assign n1690 = n1393 & n1689 ;
  buffer buf_n1682( .i (n1681), .o (n1682) );
  assign n1691 = n1685 & n1687 ;
  assign n1692 = n1682 & n1691 ;
  assign n1693 = ( n1643 & n1651 ) | ( n1643 & n1657 ) | ( n1651 & n1657 ) ;
  assign n1694 = n1482 & n1512 ;
  assign n1695 = n1451 & n1694 ;
  assign n1696 = n1401 & n1403 ;
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  assign n1699 = n1408 & n1410 ;
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  assign n1702 = n1415 & n1417 ;
  buffer buf_n1703( .i (n1702), .o (n1703) );
  assign n1704 = n1701 & n1703 ;
  assign n1705 = n1698 & n1704 ;
  assign n1706 = n1685 | n1687 ;
  assign n1707 = n1682 | n1706 ;
  assign n1708 = n1593 | n1595 ;
  buffer buf_n1709( .i (n1708), .o (n1709) );
  assign n1710 = n1599 | n1601 ;
  buffer buf_n1711( .i (n1710), .o (n1711) );
  assign n1712 = n1709 & n1711 ;
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  assign n1715 = n1608 | n1610 ;
  buffer buf_n1716( .i (n1715), .o (n1716) );
  assign n1717 = n1614 | n1616 ;
  buffer buf_n1718( .i (n1717), .o (n1718) );
  assign n1719 = n1716 & n1718 ;
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  assign n1722 = n1623 | n1625 ;
  buffer buf_n1723( .i (n1722), .o (n1723) );
  assign n1724 = n1629 | n1631 ;
  buffer buf_n1725( .i (n1724), .o (n1725) );
  assign n1726 = n1723 & n1725 ;
  buffer buf_n1727( .i (n1726), .o (n1727) );
  assign n1728 = n1721 | n1727 ;
  assign n1729 = n1714 | n1728 ;
  buffer buf_n1406( .i (n1405), .o (n1406) );
  assign n1730 = n1413 | n1419 ;
  assign n1731 = n1406 | n1730 ;
  assign n1732 = n1551 | n1557 ;
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  assign n1735 = n1566 | n1572 ;
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  assign n1738 = n1581 | n1587 ;
  buffer buf_n1739( .i (n1738), .o (n1739) );
  assign n1740 = n1737 & n1739 ;
  assign n1741 = n1734 & n1740 ;
  assign n1742 = ( n1559 & n1575 ) | ( n1559 & n1589 ) | ( n1575 & n1589 ) ;
  assign n1743 = ( n1733 & n1737 ) | ( n1733 & n1739 ) | ( n1737 & n1739 ) ;
  assign n1744 = ( n1670 & n1674 ) | ( n1670 & n1676 ) | ( n1674 & n1676 ) ;
  assign n1745 = n1709 | n1711 ;
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  assign n1748 = n1716 | n1718 ;
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  assign n1751 = n1723 | n1725 ;
  buffer buf_n1752( .i (n1751), .o (n1752) );
  assign n1753 = n1750 & n1752 ;
  assign n1754 = n1747 & n1753 ;
  assign n1755 = n1737 | n1739 ;
  assign n1756 = n1734 | n1755 ;
  assign n1757 = n1413 & n1419 ;
  assign n1758 = n1406 & n1757 ;
  assign n1759 = n1651 & n1657 ;
  assign n1760 = n1644 & n1759 ;
  assign n1761 = ( n1246 & n1310 ) | ( n1246 & n1388 ) | ( n1310 & n1388 ) ;
  assign n1762 = ( n1529 & n1537 ) | ( n1529 & n1543 ) | ( n1537 & n1543 ) ;
  assign n1763 = n1674 | n1676 ;
  assign n1764 = n1671 | n1763 ;
  assign n1765 = ( n1697 & n1701 ) | ( n1697 & n1703 ) | ( n1701 & n1703 ) ;
  assign n1766 = ( n1746 & n1750 ) | ( n1746 & n1752 ) | ( n1750 & n1752 ) ;
  buffer buf_n1517( .i (n1516), .o (n1517) );
  assign n1767 = n1520 & n1522 ;
  assign n1768 = n1517 & n1767 ;
  assign n1769 = n1701 | n1703 ;
  assign n1770 = n1698 | n1769 ;
  assign n1771 = n1721 & n1727 ;
  assign n1772 = n1714 & n1771 ;
  assign n1773 = n1621 & n1635 ;
  assign n1774 = n1606 & n1773 ;
  assign n1775 = n1575 & n1589 ;
  assign n1776 = n1560 & n1775 ;
  assign n1777 = n1520 | n1522 ;
  assign n1778 = n1517 | n1777 ;
  buffer buf_n1662( .i (n1661), .o (n1662) );
  assign n1779 = n1665 | n1667 ;
  assign n1780 = n1662 | n1779 ;
  assign n1781 = n1665 & n1667 ;
  assign n1782 = n1662 & n1781 ;
  assign n1783 = ( n1713 & n1721 ) | ( n1713 & n1727 ) | ( n1721 & n1727 ) ;
  assign n1784 = n1750 | n1752 ;
  assign n1785 = n1747 | n1784 ;
  assign n1786 = ( n1450 & n1482 ) | ( n1450 & n1512 ) | ( n1482 & n1512 ) ;
  assign n1787 = n1537 & n1543 ;
  assign n1788 = n1530 & n1787 ;
  assign n1789 = n1310 & n1388 ;
  assign n1790 = n1247 & n1789 ;
  assign n1791 = n1396 | n1398 ;
  assign n1792 = n1393 | n1791 ;
  assign b_47_ = n1390 ;
  assign b_43_ = n1399 ;
  assign b_40_ = n1420 ;
  assign b_11_ = n1514 ;
  assign b_7_ = n1523 ;
  assign b_5_ = n1545 ;
  assign b_32_ = n1591 ;
  assign b_17_ = n1637 ;
  assign b_29_ = n1659 ;
  assign b_25_ = n1668 ;
  assign b_12_ = n1678 ;
  assign b_16_ = n1679 ;
  assign b_1_ = n1688 ;
  assign b_42_ = n1690 ;
  assign b_0_ = n1692 ;
  assign b_28_ = n1693 ;
  assign b_9_ = n1695 ;
  assign b_36_ = n1705 ;
  assign b_2_ = n1707 ;
  assign b_20_ = n1729 ;
  assign b_41_ = n1731 ;
  assign b_33_ = n1741 ;
  assign b_31_ = n1742 ;
  assign b_34_ = n1743 ;
  assign b_13_ = n1744 ;
  assign b_21_ = n1754 ;
  assign b_35_ = n1756 ;
  assign b_39_ = n1758 ;
  assign b_27_ = n1760 ;
  assign b_46_ = n1761 ;
  assign b_4_ = n1762 ;
  assign b_14_ = n1764 ;
  assign b_37_ = n1765 ;
  assign b_22_ = n1766 ;
  assign b_6_ = n1768 ;
  assign b_38_ = n1770 ;
  assign b_18_ = n1772 ;
  assign b_15_ = n1774 ;
  assign b_30_ = n1776 ;
  assign b_8_ = n1778 ;
  assign b_26_ = n1780 ;
  assign b_24_ = n1782 ;
  assign b_19_ = n1783 ;
  assign b_23_ = n1785 ;
  assign b_10_ = n1786 ;
  assign b_3_ = n1788 ;
  assign b_45_ = n1790 ;
  assign b_44_ = n1792 ;
endmodule
