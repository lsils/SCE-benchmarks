module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( N1 , N100 , N103 , N106 , N109 , N110 , N111 , N112 , N113 , N114 , N115 , N118 , N12 , N121 , N124 , N127 , N130 , N133 , N134 , N135 , N138 , N141 , N144 , N147 , N15 , N150 , N151 , N152 , N153 , N154 , N155 , N156 , N157 , N158 , N159 , N160 , N161 , N162 , N163 , N164 , N165 , N166 , N167 , N168 , N169 , N170 , N171 , N172 , N173 , N174 , N175 , N176 , N177 , N178 , N179 , N18 , N180 , N181 , N182 , N183 , N184 , N185 , N186 , N187 , N188 , N189 , N190 , N191 , N192 , N193 , N194 , N195 , N196 , N197 , N198 , N199 , N200 , N201 , N202 , N203 , N204 , N205 , N206 , N207 , N208 , N209 , N210 , N211 , N212 , N213 , N214 , N215 , N216 , N217 , N218 , N219 , N220 , N221 , N222 , N223 , N224 , N225 , N226 , N227 , N228 , N229 , N23 , N230 , N231 , N232 , N233 , N234 , N235 , N236 , N237 , N238 , N239 , N240 , N241_I , N242 , N245 , N248 , N251 , N254 , N257 , N26 , N260 , N263 , N267 , N271 , N274 , N277 , N280 , N283 , N286 , N289 , N29 , N293 , N296 , N299 , N303 , N307 , N310 , N313 , N316 , N319 , N32 , N322 , N325 , N328 , N331 , N334 , N337 , N340 , N343 , N346 , N349 , N35 , N352 , N355 , N358 , N361 , N364 , N367 , N38 , N382 , N41 , N44 , N47 , N5 , N50 , N53 , N54 , N55 , N56 , N57 , N58 , N59 , N60 , N61 , N62 , N63 , N64 , N65 , N66 , N69 , N70 , N73 , N74 , N75 , N76 , N77 , N78 , N79 , N80 , N81 , N82 , N83 , N84 , N85 , N86 , N87 , N88 , N89 , N9 , N94 , N97 , N10025 , N10101 , N10102 , N10103 , N10104 , N10109 , N10110 , N10111 , N10112 , N10350 , N10351 , N10352 , N10353 , N10574 , N10575 , N10576 , N10628 , N10632 , N10641 , N10704 , N10706 , N10711 , N10712 , N10713 , N10714 , N10715 , N10716 , N10717 , N10718 , N10729 , N10759 , N10760 , N10761 , N10762 , N10763 , N10827 , N10837 , N10838 , N10839 , N10840 , N10868 , N10869 , N10870 , N10871 , N10905 , N10906 , N10907 , N10908 , N1110 , N1111 , N1112 , N1113 , N1114 , N11333 , N11334 , N11340 , N11342 , N1489 , N1490 , N1781 , N241_O , N387 , N388 , N478 , N482 , N484 , N486 , N489 , N492 , N501 , N505 , N507 , N509 , N511 , N513 , N515 , N517 , N519 , N535 , N537 , N539 , N541 , N543 , N545 , N547 , N549 , N551 , N553 , N556 , N559 , N561 , N563 , N565 , N567 , N569 , N571 , N573 , N582 , N643 , N707 , N813 , N881 , N882 , N883 , N884 , N885 , N889 , N945 );
  input N1 , N100 , N103 , N106 , N109 , N110 , N111 , N112 , N113 , N114 , N115 , N118 , N12 , N121 , N124 , N127 , N130 , N133 , N134 , N135 , N138 , N141 , N144 , N147 , N15 , N150 , N151 , N152 , N153 , N154 , N155 , N156 , N157 , N158 , N159 , N160 , N161 , N162 , N163 , N164 , N165 , N166 , N167 , N168 , N169 , N170 , N171 , N172 , N173 , N174 , N175 , N176 , N177 , N178 , N179 , N18 , N180 , N181 , N182 , N183 , N184 , N185 , N186 , N187 , N188 , N189 , N190 , N191 , N192 , N193 , N194 , N195 , N196 , N197 , N198 , N199 , N200 , N201 , N202 , N203 , N204 , N205 , N206 , N207 , N208 , N209 , N210 , N211 , N212 , N213 , N214 , N215 , N216 , N217 , N218 , N219 , N220 , N221 , N222 , N223 , N224 , N225 , N226 , N227 , N228 , N229 , N23 , N230 , N231 , N232 , N233 , N234 , N235 , N236 , N237 , N238 , N239 , N240 , N241_I , N242 , N245 , N248 , N251 , N254 , N257 , N26 , N260 , N263 , N267 , N271 , N274 , N277 , N280 , N283 , N286 , N289 , N29 , N293 , N296 , N299 , N303 , N307 , N310 , N313 , N316 , N319 , N32 , N322 , N325 , N328 , N331 , N334 , N337 , N340 , N343 , N346 , N349 , N35 , N352 , N355 , N358 , N361 , N364 , N367 , N38 , N382 , N41 , N44 , N47 , N5 , N50 , N53 , N54 , N55 , N56 , N57 , N58 , N59 , N60 , N61 , N62 , N63 , N64 , N65 , N66 , N69 , N70 , N73 , N74 , N75 , N76 , N77 , N78 , N79 , N80 , N81 , N82 , N83 , N84 , N85 , N86 , N87 , N88 , N89 , N9 , N94 , N97 ;
  output N10025 , N10101 , N10102 , N10103 , N10104 , N10109 , N10110 , N10111 , N10112 , N10350 , N10351 , N10352 , N10353 , N10574 , N10575 , N10576 , N10628 , N10632 , N10641 , N10704 , N10706 , N10711 , N10712 , N10713 , N10714 , N10715 , N10716 , N10717 , N10718 , N10729 , N10759 , N10760 , N10761 , N10762 , N10763 , N10827 , N10837 , N10838 , N10839 , N10840 , N10868 , N10869 , N10870 , N10871 , N10905 , N10906 , N10907 , N10908 , N1110 , N1111 , N1112 , N1113 , N1114 , N11333 , N11334 , N11340 , N11342 , N1489 , N1490 , N1781 , N241_O , N387 , N388 , N478 , N482 , N484 , N486 , N489 , N492 , N501 , N505 , N507 , N509 , N511 , N513 , N515 , N517 , N519 , N535 , N537 , N539 , N541 , N543 , N545 , N547 , N549 , N551 , N553 , N556 , N559 , N561 , N563 , N565 , N567 , N569 , N571 , N573 , N582 , N643 , N707 , N813 , N881 , N882 , N883 , N884 , N885 , N889 , N945 ;
  wire n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 ;
  assign n208 = ~N18 & N41 ;
  buffer buf_n209( .i (n208), .o (n209) );
  assign n210 = ~N310 & n209 ;
  buffer buf_n211( .i (n210), .o (n211) );
  assign n216 = N18 | N41 ;
  assign n217 = N310 & ~n216 ;
  buffer buf_n218( .i (n217), .o (n218) );
  assign n224 = n211 | n218 ;
  buffer buf_n225( .i (n224), .o (n225) );
  assign n228 = N367 & ~n225 ;
  buffer buf_n229( .i (n228), .o (n229) );
  assign n230 = ~N367 & n225 ;
  buffer buf_n231( .i (n230), .o (n231) );
  assign n232 = ~n229 & ~n231 ;
  assign n233 = N267 & N382 ;
  buffer buf_n234( .i (n233), .o (n234) );
  assign n291 = ~N38 & n234 ;
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  assign n347 = N263 & n234 ;
  assign n348 = N38 & ~n347 ;
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  assign n402 = N263 & N382 ;
  buffer buf_n403( .i (n402), .o (n403) );
  assign n404 = N38 & n403 ;
  buffer buf_n405( .i (n404), .o (n405) );
  assign n409 = N38 | n403 ;
  buffer buf_n410( .i (n409), .o (n410) );
  assign n413 = ~n405 & n410 ;
  buffer buf_n414( .i (n413), .o (n414) );
  assign n415 = N12 & N9 ;
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  assign n421 = N18 & ~N213 ;
  buffer buf_n422( .i (n421), .o (n422) );
  assign n425 = n418 | n422 ;
  buffer buf_n426( .i (n425), .o (n426) );
  assign n427 = N260 | n426 ;
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  assign n430 = N18 & ~N214 ;
  buffer buf_n431( .i (n430), .o (n431) );
  assign n434 = n418 | n431 ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n436 = N257 | n435 ;
  buffer buf_n437( .i (n436), .o (n437) );
  assign n447 = N260 & n426 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = n437 | n448 ;
  assign n450 = n429 & n449 ;
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  assign n487 = N18 & ~N215 ;
  buffer buf_n488( .i (n487), .o (n488) );
  assign n491 = n418 | n488 ;
  buffer buf_n492( .i (n491), .o (n492) );
  assign n493 = N106 | n492 ;
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  assign n500 = N106 & n492 ;
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  assign n506 = N18 & ~N216 ;
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n510( .i (n417), .o (n510) );
  assign n511 = n507 | n510 ;
  buffer buf_n512( .i (n511), .o (n512) );
  assign n513 = N254 & n512 ;
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  assign n517 = N18 & ~N209 ;
  buffer buf_n518( .i (n517), .o (n518) );
  assign n519 = n510 | n518 ;
  buffer buf_n520( .i (n519), .o (n520) );
  assign n521 = N251 | n520 ;
  buffer buf_n522( .i (n521), .o (n522) );
  assign n567 = N254 | n512 ;
  buffer buf_n568( .i (n567), .o (n568) );
  assign n569 = n522 & n568 ;
  buffer buf_n570( .i (n569), .o (n570) );
  assign n571 = n516 | n570 ;
  buffer buf_n572( .i (n571), .o (n572) );
  assign n606 = n505 | n572 ;
  assign n607 = n499 & n606 ;
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  assign n640 = N257 & n435 ;
  buffer buf_n641( .i (n640), .o (n641) );
  assign n650 = n437 & ~n641 ;
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  assign n690 = n428 & ~n448 ;
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  assign n731 = n684 & n724 ;
  buffer buf_n732( .i (n731), .o (n732) );
  assign n734 = ~n638 & n732 ;
  assign n735 = n486 & ~n734 ;
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n419( .i (n418), .o (n419) );
  assign n736 = ~N153 & N18 ;
  buffer buf_n737( .i (n736), .o (n737) );
  assign n740 = n419 | n737 ;
  buffer buf_n741( .i (n740), .o (n741) );
  assign n742 = N303 & n741 ;
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  assign n777 = N303 | n741 ;
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  assign n811 = ~N154 & N18 ;
  buffer buf_n812( .i (n811), .o (n812) );
  assign n815 = n419 | n812 ;
  buffer buf_n816( .i (n815), .o (n816) );
  assign n817 = N299 & n816 ;
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  assign n824 = N299 | n816 ;
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  assign n829 = ~N155 & N18 ;
  buffer buf_n830( .i (n829), .o (n830) );
  assign n833 = n510 | n830 ;
  buffer buf_n834( .i (n833), .o (n834) );
  assign n835 = N296 & n834 ;
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  assign n839 = N296 | n834 ;
  buffer buf_n840( .i (n839), .o (n840) );
  assign n844 = ~N156 & N18 ;
  buffer buf_n845( .i (n844), .o (n845) );
  assign n848 = n510 | n845 ;
  buffer buf_n849( .i (n848), .o (n849) );
  assign n850 = N293 | n849 ;
  buffer buf_n851( .i (n850), .o (n851) );
  assign n883 = n840 & n851 ;
  buffer buf_n884( .i (n883), .o (n884) );
  assign n886 = n838 | n884 ;
  buffer buf_n887( .i (n886), .o (n887) );
  assign n915 = n828 & n887 ;
  buffer buf_n916( .i (n915), .o (n916) );
  assign n917 = n823 | n916 ;
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n885( .i (n884), .o (n885) );
  assign n941 = N293 & n849 ;
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  assign n973 = n837 | n943 ;
  buffer buf_n974( .i (n973), .o (n974) );
  assign n975 = n885 & ~n974 ;
  buffer buf_n976( .i (n975), .o (n976) );
  assign n1002 = ~n818 & n825 ;
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  assign n1034 = n976 & n1005 ;
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  assign n1037 = n918 & ~n1036 ;
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  assign n1060 = ~N157 & N18 ;
  buffer buf_n1061( .i (n417), .o (n1061) );
  assign n1062 = n1060 | n1061 ;
  buffer buf_n1063( .i (n1062), .o (n1063) );
  assign n1064 = N289 & n1063 ;
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  assign n1078 = N289 | n1063 ;
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  assign n1089 = N135 & ~N18 ;
  buffer buf_n1090( .i (n1089), .o (n1090) );
  assign n1091 = N158 & N18 ;
  assign n1092 = n1090 | n1091 ;
  buffer buf_n1093( .i (n1092), .o (n1093) );
  assign n1094 = N286 & ~n1093 ;
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  assign n1103 = ~N286 & n1093 ;
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  assign n1111 = N144 & ~N18 ;
  buffer buf_n1112( .i (n1111), .o (n1112) );
  assign n1113 = N159 & N18 ;
  assign n1114 = n1112 | n1113 ;
  buffer buf_n1115( .i (n1114), .o (n1115) );
  assign n1116 = ~N283 & n1115 ;
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  assign n1123 = N283 & ~n1115 ;
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  assign n1129 = N138 & ~N18 ;
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n1131 = N160 & N18 ;
  assign n1132 = n1130 | n1131 ;
  buffer buf_n1133( .i (n1132), .o (n1133) );
  assign n1134 = ~N280 & n1133 ;
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  assign n1138 = N147 & ~N18 ;
  buffer buf_n1139( .i (n1138), .o (n1139) );
  assign n1140 = N151 & N18 ;
  assign n1141 = n1139 | n1140 ;
  buffer buf_n1142( .i (n1141), .o (n1142) );
  assign n1143 = ~N277 & n1142 ;
  buffer buf_n1144( .i (n1143), .o (n1144) );
  assign n1180 = N280 & ~n1133 ;
  buffer buf_n1181( .i (n1180), .o (n1181) );
  assign n1182 = n1144 & ~n1181 ;
  buffer buf_n1183( .i (n1182), .o (n1183) );
  assign n1184 = n1137 | n1183 ;
  buffer buf_n1185( .i (n1184), .o (n1185) );
  assign n1212 = ~n1128 & n1185 ;
  assign n1213 = n1122 | n1212 ;
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  assign n1239 = n1110 | n1215 ;
  assign n1240 = ~n1102 & n1239 ;
  buffer buf_n1241( .i (n1240), .o (n1241) );
  assign n1263 = n1088 & ~n1241 ;
  buffer buf_n1264( .i (n1263), .o (n1264) );
  assign n1281 = N277 & ~n1142 ;
  buffer buf_n1282( .i (n1281), .o (n1282) );
  assign n1283 = n1144 | n1282 ;
  buffer buf_n1284( .i (n1283), .o (n1284) );
  assign n1316 = n1135 | n1181 ;
  buffer buf_n1317( .i (n1316), .o (n1317) );
  assign n1353 = n1284 | n1317 ;
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  assign n1380 = n1095 | n1104 ;
  buffer buf_n1381( .i (n1380), .o (n1381) );
  assign n1411 = n1117 | n1124 ;
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  assign n1443 = n1381 | n1414 ;
  buffer buf_n1444( .i (n1443), .o (n1444) );
  assign n1445 = n1356 | n1444 ;
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  assign n1453 = n1264 & n1451 ;
  assign n1454 = n1077 | n1453 ;
  buffer buf_n1455( .i (n1454), .o (n1455) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  assign n1470 = N18 & N219 ;
  assign n1471 = ~N18 & N66 ;
  buffer buf_n1472( .i (n1471), .o (n1472) );
  assign n1473 = n1470 | n1472 ;
  buffer buf_n1474( .i (n1473), .o (n1474) );
  assign n1475 = ~N364 & n1474 ;
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n1488( .i (n1487), .o (n1488) );
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  assign n1504 = N364 & ~n1474 ;
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n1522( .i (n1521), .o (n1522) );
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  assign n1532 = N18 & N220 ;
  assign n1533 = ~N18 & N50 ;
  buffer buf_n1534( .i (n1533), .o (n1534) );
  assign n1535 = n1532 | n1534 ;
  buffer buf_n1536( .i (n1535), .o (n1536) );
  assign n1537 = N361 & ~n1536 ;
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1543( .i (n1542), .o (n1543) );
  assign n1545 = ~N361 & n1536 ;
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  assign n1552 = N18 & N221 ;
  assign n1553 = ~N18 & N32 ;
  buffer buf_n1554( .i (n1553), .o (n1554) );
  assign n1555 = n1552 | n1554 ;
  buffer buf_n1556( .i (n1555), .o (n1556) );
  assign n1557 = N358 & ~n1556 ;
  buffer buf_n1558( .i (n1557), .o (n1558) );
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  assign n1561 = ~N358 & n1556 ;
  buffer buf_n1562( .i (n1561), .o (n1562) );
  assign n1564 = N18 & N222 ;
  assign n1565 = ~N18 & N35 ;
  buffer buf_n1566( .i (n1565), .o (n1566) );
  assign n1567 = n1564 | n1566 ;
  buffer buf_n1568( .i (n1567), .o (n1568) );
  assign n1569 = ~N355 & n1568 ;
  buffer buf_n1570( .i (n1569), .o (n1570) );
  assign n1594 = n1562 | n1570 ;
  buffer buf_n1595( .i (n1594), .o (n1595) );
  assign n1596 = ~n1560 & n1595 ;
  buffer buf_n1597( .i (n1596), .o (n1597) );
  assign n1618 = n1550 | n1597 ;
  assign n1619 = ~n1543 & n1618 ;
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  assign n1637 = n1558 | n1562 ;
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  assign n1663 = N355 & ~n1568 ;
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  assign n1689 = n1572 | n1666 ;
  buffer buf_n1690( .i (n1689), .o (n1690) );
  assign n1713 = n1640 | n1690 ;
  buffer buf_n1714( .i (n1713), .o (n1714) );
  assign n1732 = n1544 | n1714 ;
  assign n1733 = ~n1620 & n1732 ;
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n1633( .i (n1632), .o (n1633) );
  buffer buf_n1634( .i (n1633), .o (n1634) );
  buffer buf_n1635( .i (n1634), .o (n1635) );
  buffer buf_n1636( .i (n1635), .o (n1636) );
  assign n1750 = N18 & N217 ;
  assign n1751 = N118 & ~N18 ;
  buffer buf_n1752( .i (n1751), .o (n1752) );
  assign n1753 = n1750 | n1752 ;
  buffer buf_n1754( .i (n1753), .o (n1754) );
  assign n1755 = ~N340 & n1754 ;
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  assign n1780 = N18 & N226 ;
  assign n1781 = ~N18 & N97 ;
  buffer buf_n1782( .i (n1781), .o (n1782) );
  assign n1783 = n1780 | n1782 ;
  buffer buf_n1784( .i (n1783), .o (n1784) );
  assign n1785 = N343 & ~n1784 ;
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  assign n1789 = n1758 | n1788 ;
  buffer buf_n1790( .i (n1789), .o (n1790) );
  assign n1791 = N340 & ~n1754 ;
  buffer buf_n1792( .i (n1791), .o (n1792) );
  assign n1812 = ~N343 & n1784 ;
  buffer buf_n1813( .i (n1812), .o (n1813) );
  assign n1815 = n1792 | n1813 ;
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  buffer buf_n1818( .i (n1817), .o (n1818) );
  assign n1819 = n1790 | n1818 ;
  buffer buf_n1820( .i (n1819), .o (n1820) );
  assign n1821 = N18 & N224 ;
  assign n1822 = N121 & ~N18 ;
  buffer buf_n1823( .i (n1822), .o (n1823) );
  assign n1824 = n1821 | n1823 ;
  buffer buf_n1825( .i (n1824), .o (n1825) );
  assign n1826 = N349 & ~n1825 ;
  buffer buf_n1827( .i (n1826), .o (n1827) );
  assign n1836 = ~N349 & n1825 ;
  buffer buf_n1837( .i (n1836), .o (n1837) );
  assign n1847 = n1827 | n1837 ;
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  assign n1869 = N18 & N225 ;
  assign n1870 = ~N18 & N94 ;
  buffer buf_n1871( .i (n1870), .o (n1871) );
  assign n1872 = n1869 | n1871 ;
  buffer buf_n1873( .i (n1872), .o (n1873) );
  assign n1874 = N346 & ~n1873 ;
  buffer buf_n1875( .i (n1874), .o (n1875) );
  assign n1880 = ~N346 & n1873 ;
  buffer buf_n1881( .i (n1880), .o (n1881) );
  assign n1888 = n1875 | n1881 ;
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  buffer buf_n1891( .i (n1890), .o (n1891) );
  assign n1914 = n1850 | n1891 ;
  buffer buf_n1915( .i (n1914), .o (n1915) );
  assign n1916 = n1820 | n1915 ;
  buffer buf_n1917( .i (n1916), .o (n1917) );
  assign n1929 = N18 & N223 ;
  assign n1930 = ~N18 & N47 ;
  buffer buf_n1931( .i (n1930), .o (n1931) );
  assign n1932 = n1929 | n1931 ;
  buffer buf_n1933( .i (n1932), .o (n1933) );
  assign n1934 = ~N352 & n1933 ;
  buffer buf_n1935( .i (n1934), .o (n1935) );
  assign n1948 = N352 & ~n1933 ;
  buffer buf_n1949( .i (n1948), .o (n1949) );
  assign n1961 = n1935 | n1949 ;
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n1967( .i (n1966), .o (n1967) );
  buffer buf_n1968( .i (n1967), .o (n1968) );
  assign n1972 = n1917 | n1968 ;
  buffer buf_n1973( .i (n1972), .o (n1973) );
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  assign n1983 = N18 & N231 ;
  assign n1984 = N100 & ~N18 ;
  buffer buf_n1985( .i (n1984), .o (n1985) );
  assign n1986 = n1983 | n1985 ;
  buffer buf_n1987( .i (n1986), .o (n1987) );
  assign n1988 = N334 & ~n1987 ;
  buffer buf_n1989( .i (n1988), .o (n1989) );
  buffer buf_n1990( .i (n1989), .o (n1990) );
  buffer buf_n1991( .i (n1990), .o (n1991) );
  buffer buf_n1992( .i (n1991), .o (n1992) );
  buffer buf_n1993( .i (n1992), .o (n1993) );
  buffer buf_n1994( .i (n1993), .o (n1994) );
  buffer buf_n1995( .i (n1994), .o (n1995) );
  buffer buf_n1996( .i (n1995), .o (n1996) );
  assign n1997 = ~N334 & n1987 ;
  buffer buf_n1998( .i (n1997), .o (n1998) );
  buffer buf_n1999( .i (n1998), .o (n1999) );
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n2001( .i (n2000), .o (n2001) );
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n2003), .o (n2004) );
  assign n2005 = N18 & N232 ;
  assign n2006 = N124 & ~N18 ;
  buffer buf_n2007( .i (n2006), .o (n2007) );
  assign n2008 = n2005 | n2007 ;
  buffer buf_n2009( .i (n2008), .o (n2009) );
  assign n2010 = N331 & ~n2009 ;
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n2012( .i (n2011), .o (n2012) );
  buffer buf_n2013( .i (n2012), .o (n2013) );
  buffer buf_n2014( .i (n2013), .o (n2014) );
  buffer buf_n2015( .i (n2014), .o (n2015) );
  assign n2016 = ~N331 & n2009 ;
  buffer buf_n2017( .i (n2016), .o (n2017) );
  buffer buf_n2018( .i (n2017), .o (n2018) );
  buffer buf_n2019( .i (n2018), .o (n2019) );
  buffer buf_n2020( .i (n2019), .o (n2020) );
  assign n2021 = N18 & N233 ;
  assign n2022 = N127 & ~N18 ;
  buffer buf_n2023( .i (n2022), .o (n2023) );
  assign n2024 = n2021 | n2023 ;
  buffer buf_n2025( .i (n2024), .o (n2025) );
  assign n2026 = N328 & ~n2025 ;
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2028( .i (n2027), .o (n2028) );
  assign n2029 = ~N328 & n2025 ;
  buffer buf_n2030( .i (n2029), .o (n2030) );
  assign n2032 = N18 & N234 ;
  assign n2033 = N130 & ~N18 ;
  buffer buf_n2034( .i (n2033), .o (n2034) );
  assign n2035 = n2032 | n2034 ;
  buffer buf_n2036( .i (n2035), .o (n2036) );
  assign n2037 = ~N325 & n2036 ;
  buffer buf_n2038( .i (n2037), .o (n2038) );
  assign n2057 = n2030 | n2038 ;
  assign n2058 = ~n2028 & n2057 ;
  buffer buf_n2059( .i (n2058), .o (n2059) );
  assign n2076 = n2020 | n2059 ;
  assign n2077 = ~n2015 & n2076 ;
  buffer buf_n2078( .i (n2077), .o (n2078) );
  assign n2090 = n2004 | n2078 ;
  assign n2091 = ~n1996 & n2090 ;
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n2099( .i (n2098), .o (n2099) );
  buffer buf_n2100( .i (n2099), .o (n2100) );
  assign n2101 = N18 & N235 ;
  assign n2102 = N103 & ~N18 ;
  buffer buf_n2103( .i (n2102), .o (n2103) );
  assign n2104 = n2101 | n2103 ;
  buffer buf_n2105( .i (n2104), .o (n2105) );
  assign n2106 = ~N322 & n2105 ;
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n2111( .i (n2110), .o (n2111) );
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  assign n2120 = N322 & ~n2105 ;
  buffer buf_n2121( .i (n2120), .o (n2121) );
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  buffer buf_n2129( .i (n2128), .o (n2129) );
  buffer buf_n2130( .i (n2129), .o (n2130) );
  assign n2133 = N18 & N236 ;
  assign n2134 = ~N18 & N23 ;
  buffer buf_n2135( .i (n2134), .o (n2135) );
  assign n2136 = n2133 | n2135 ;
  buffer buf_n2137( .i (n2136), .o (n2137) );
  assign n2138 = N319 & ~n2137 ;
  buffer buf_n2139( .i (n2138), .o (n2139) );
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n2143( .i (n2142), .o (n2143) );
  buffer buf_n2144( .i (n2143), .o (n2144) );
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  assign n2149 = ~N319 & n2137 ;
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  buffer buf_n2152( .i (n2151), .o (n2152) );
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n2155( .i (n2154), .o (n2155) );
  assign n2156 = N18 & N237 ;
  assign n2157 = ~N18 & N26 ;
  buffer buf_n2158( .i (n2157), .o (n2158) );
  assign n2159 = n2156 | n2158 ;
  buffer buf_n2160( .i (n2159), .o (n2160) );
  assign n2161 = N316 & ~n2160 ;
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n2163( .i (n2162), .o (n2163) );
  buffer buf_n2164( .i (n2163), .o (n2164) );
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  assign n2166 = N18 & N238 ;
  assign n2167 = ~N18 & N29 ;
  buffer buf_n2168( .i (n2167), .o (n2168) );
  assign n2169 = n2166 | n2168 ;
  buffer buf_n2170( .i (n2169), .o (n2170) );
  assign n2171 = N313 & ~n2170 ;
  buffer buf_n2172( .i (n2171), .o (n2172) );
  assign n2176 = n213 & ~n2172 ;
  buffer buf_n2177( .i (n2176), .o (n2177) );
  assign n2178 = ~N316 & n2160 ;
  buffer buf_n2179( .i (n2178), .o (n2179) );
  assign n2180 = ~N313 & n2170 ;
  buffer buf_n2181( .i (n2180), .o (n2181) );
  assign n2184 = n2179 | n2181 ;
  buffer buf_n2185( .i (n2184), .o (n2185) );
  assign n2186 = n2177 | n2185 ;
  assign n2187 = ~n2165 & n2186 ;
  buffer buf_n2188( .i (n2187), .o (n2188) );
  assign n2192 = n2155 | n2188 ;
  buffer buf_n2193( .i (n2192), .o (n2193) );
  assign n2195 = ~n2146 & n2193 ;
  buffer buf_n2196( .i (n2195), .o (n2196) );
  assign n2197 = ~n2130 & n2196 ;
  assign n2198 = n2117 | n2197 ;
  buffer buf_n2199( .i (n2198), .o (n2199) );
  assign n2200 = N367 | n2199 ;
  buffer buf_n2201( .i (n2200), .o (n2201) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  buffer buf_n2119( .i (n2118), .o (n2119) );
  buffer buf_n2131( .i (n2130), .o (n2131) );
  buffer buf_n2132( .i (n2131), .o (n2132) );
  assign n2202 = n2162 | n2179 ;
  buffer buf_n2203( .i (n2202), .o (n2203) );
  buffer buf_n2204( .i (n2203), .o (n2204) );
  buffer buf_n2205( .i (n2204), .o (n2205) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  assign n2207 = n2172 | n2181 ;
  buffer buf_n2208( .i (n2207), .o (n2208) );
  assign n2211 = n227 | n2208 ;
  buffer buf_n2212( .i (n2211), .o (n2212) );
  assign n2213 = n2205 | n2212 ;
  buffer buf_n2214( .i (n2213), .o (n2214) );
  assign n2215 = n2139 | n2150 ;
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  assign n2225 = n2214 | n2220 ;
  buffer buf_n2226( .i (n2225), .o (n2226) );
  buffer buf_n2227( .i (n2226), .o (n2227) );
  assign n2228 = ~n2196 & n2227 ;
  buffer buf_n2229( .i (n2228), .o (n2229) );
  assign n2230 = n2132 | n2229 ;
  assign n2231 = ~n2119 & n2230 ;
  buffer buf_n2232( .i (n2231), .o (n2232) );
  assign n2233 = n2201 & ~n2232 ;
  buffer buf_n2234( .i (n2233), .o (n2234) );
  assign n2236 = n2027 | n2030 ;
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  assign n2256 = N325 & ~n2036 ;
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  assign n2274 = n2039 | n2258 ;
  buffer buf_n2275( .i (n2274), .o (n2275) );
  assign n2290 = n2238 | n2275 ;
  buffer buf_n2291( .i (n2290), .o (n2291) );
  assign n2292 = n2011 | n2017 ;
  buffer buf_n2293( .i (n2292), .o (n2293) );
  buffer buf_n2294( .i (n2293), .o (n2294) );
  assign n2313 = n1989 | n1998 ;
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  assign n2332 = n2294 | n2315 ;
  buffer buf_n2333( .i (n2332), .o (n2333) );
  assign n2334 = n2291 | n2333 ;
  buffer buf_n2335( .i (n2334), .o (n2335) );
  buffer buf_n2336( .i (n2335), .o (n2336) );
  buffer buf_n2337( .i (n2336), .o (n2337) );
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  buffer buf_n2340( .i (n2339), .o (n2340) );
  buffer buf_n2341( .i (n2340), .o (n2341) );
  buffer buf_n2342( .i (n2341), .o (n2342) );
  buffer buf_n2343( .i (n2342), .o (n2343) );
  buffer buf_n2344( .i (n2343), .o (n2344) );
  assign n2345 = n2234 & ~n2344 ;
  assign n2346 = n2100 | n2345 ;
  buffer buf_n2347( .i (n2346), .o (n2347) );
  assign n2350 = ~n1982 & n2347 ;
  buffer buf_n2351( .i (n2350), .o (n2351) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  buffer buf_n1954( .i (n1953), .o (n1954) );
  buffer buf_n1955( .i (n1954), .o (n1955) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  buffer buf_n1960( .i (n1959), .o (n1960) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  buffer buf_n1846( .i (n1845), .o (n1846) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  buffer buf_n1879( .i (n1878), .o (n1879) );
  buffer buf_n1814( .i (n1813), .o (n1814) );
  assign n2352 = n1757 | n1814 ;
  assign n2353 = ~n1788 & n2352 ;
  buffer buf_n2354( .i (n2353), .o (n2354) );
  assign n2375 = ~n1879 & n2354 ;
  buffer buf_n2376( .i (n2375), .o (n2376) );
  assign n2377 = n1887 | n2376 ;
  buffer buf_n2378( .i (n2377), .o (n2378) );
  assign n2391 = ~n1835 & n2378 ;
  assign n2392 = n1846 | n2391 ;
  buffer buf_n2393( .i (n2392), .o (n2393) );
  assign n2394 = ~n1960 & n2393 ;
  assign n2395 = n1947 | n2394 ;
  buffer buf_n2396( .i (n2395), .o (n2396) );
  buffer buf_n2397( .i (n2396), .o (n2397) );
  buffer buf_n2398( .i (n2397), .o (n2398) );
  buffer buf_n2399( .i (n2398), .o (n2399) );
  buffer buf_n2400( .i (n2399), .o (n2400) );
  buffer buf_n2401( .i (n2400), .o (n2401) );
  buffer buf_n2402( .i (n2401), .o (n2402) );
  buffer buf_n2403( .i (n2402), .o (n2403) );
  assign n2404 = n2351 | n2403 ;
  buffer buf_n2405( .i (n2404), .o (n2405) );
  assign n2409 = n1636 | n2405 ;
  assign n2410 = ~n1749 & n2409 ;
  buffer buf_n2411( .i (n2410), .o (n2411) );
  assign n2412 = ~n1531 & n2411 ;
  assign n2413 = n1503 | n2412 ;
  buffer buf_n2414( .i (n2413), .o (n2414) );
  assign n2419 = n1280 & ~n2414 ;
  assign n2420 = n1469 | n2419 ;
  buffer buf_n2421( .i (n2420), .o (n2421) );
  assign n2427 = n940 & n2421 ;
  assign n2428 = n1059 | n2427 ;
  buffer buf_n2429( .i (n2428), .o (n2429) );
  assign n2430 = n810 & n2429 ;
  assign n2431 = n776 | n2430 ;
  buffer buf_n2432( .i (n2431), .o (n2432) );
  assign n2439 = n494 & ~n501 ;
  buffer buf_n2440( .i (n2439), .o (n2440) );
  buffer buf_n2441( .i (n2440), .o (n2441) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  assign n2478 = N251 & n520 ;
  buffer buf_n2479( .i (n2478), .o (n2479) );
  assign n2480 = n522 & ~n2479 ;
  buffer buf_n2481( .i (n2480), .o (n2481) );
  assign n2522 = ~n514 & n568 ;
  buffer buf_n2523( .i (n2522), .o (n2523) );
  assign n2568 = n2481 & n2523 ;
  buffer buf_n2569( .i (n2568), .o (n2569) );
  assign n2602 = n2442 & n2569 ;
  buffer buf_n2603( .i (n2602), .o (n2603) );
  buffer buf_n2604( .i (n2603), .o (n2604) );
  buffer buf_n2605( .i (n2604), .o (n2605) );
  buffer buf_n2606( .i (n2605), .o (n2606) );
  buffer buf_n2607( .i (n2606), .o (n2607) );
  buffer buf_n2608( .i (n2607), .o (n2608) );
  buffer buf_n2609( .i (n2608), .o (n2609) );
  buffer buf_n2610( .i (n2609), .o (n2610) );
  buffer buf_n2611( .i (n2610), .o (n2611) );
  buffer buf_n2612( .i (n2611), .o (n2612) );
  buffer buf_n2613( .i (n2612), .o (n2613) );
  buffer buf_n2614( .i (n2613), .o (n2614) );
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  buffer buf_n2617( .i (n2616), .o (n2617) );
  buffer buf_n2618( .i (n2617), .o (n2618) );
  buffer buf_n2619( .i (n2618), .o (n2619) );
  buffer buf_n2620( .i (n2619), .o (n2620) );
  buffer buf_n2621( .i (n2620), .o (n2621) );
  buffer buf_n2622( .i (n2621), .o (n2622) );
  buffer buf_n2623( .i (n2622), .o (n2623) );
  buffer buf_n2624( .i (n2623), .o (n2624) );
  buffer buf_n2625( .i (n2624), .o (n2625) );
  buffer buf_n2626( .i (n2625), .o (n2626) );
  buffer buf_n2627( .i (n2626), .o (n2627) );
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  buffer buf_n2631( .i (n2630), .o (n2631) );
  buffer buf_n2632( .i (n2631), .o (n2632) );
  buffer buf_n2633( .i (n2632), .o (n2633) );
  assign n2634 = ~n2432 & n2633 ;
  buffer buf_n2635( .i (n2634), .o (n2635) );
  assign n2636 = n733 & n2635 ;
  assign n2637 = n735 & ~n2636 ;
  buffer buf_n2638( .i (n2637), .o (n2638) );
  buffer buf_n2639( .i (n2638), .o (n2639) );
  buffer buf_n2640( .i (n2639), .o (n2640) );
  buffer buf_n2641( .i (n2640), .o (n2641) );
  buffer buf_n2642( .i (n2641), .o (n2642) );
  buffer buf_n2643( .i (n2642), .o (n2643) );
  buffer buf_n2644( .i (n2643), .o (n2644) );
  buffer buf_n2645( .i (n2644), .o (n2645) );
  assign n2646 = n414 | n2645 ;
  buffer buf_n2647( .i (n2646), .o (n2647) );
  assign n2648 = ~n401 & n2647 ;
  assign n2649 = n346 | n2648 ;
  inverter inv_n2650( .i (n2649), .o (n2650) );
  assign n2651 = N245 & N271 ;
  buffer buf_n2652( .i (n2651), .o (n2652) );
  assign n2653 = ~N38 & N382 ;
  assign n2654 = ~n2652 & n2653 ;
  buffer buf_n2655( .i (n2654), .o (n2655) );
  buffer buf_n2656( .i (n2655), .o (n2656) );
  buffer buf_n2657( .i (n2656), .o (n2657) );
  buffer buf_n2658( .i (n2657), .o (n2658) );
  buffer buf_n2659( .i (n2658), .o (n2659) );
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2660), .o (n2661) );
  buffer buf_n2662( .i (n2661), .o (n2662) );
  buffer buf_n2663( .i (n2662), .o (n2663) );
  buffer buf_n2664( .i (n2663), .o (n2664) );
  buffer buf_n2665( .i (n2664), .o (n2665) );
  buffer buf_n2666( .i (n2665), .o (n2666) );
  buffer buf_n2667( .i (n2666), .o (n2667) );
  buffer buf_n2668( .i (n2667), .o (n2668) );
  buffer buf_n2669( .i (n2668), .o (n2669) );
  buffer buf_n2670( .i (n2669), .o (n2670) );
  buffer buf_n2671( .i (n2670), .o (n2671) );
  buffer buf_n2672( .i (n2671), .o (n2672) );
  buffer buf_n2673( .i (n2672), .o (n2673) );
  assign n2674 = ~N18 & N53 ;
  assign n2675 = N18 & ~N325 ;
  assign n2676 = n2674 | n2675 ;
  buffer buf_n2677( .i (n2676), .o (n2677) );
  buffer buf_n2678( .i (n2677), .o (n2678) );
  assign n2679 = N18 & N203 ;
  assign n2680 = n2034 | n2679 ;
  buffer buf_n2681( .i (n2680), .o (n2681) );
  assign n2682 = n2678 | n2681 ;
  buffer buf_n2683( .i (n2682), .o (n2683) );
  buffer buf_n2684( .i (n2683), .o (n2684) );
  buffer buf_n2685( .i (n2684), .o (n2685) );
  buffer buf_n2686( .i (n2685), .o (n2686) );
  buffer buf_n2687( .i (n2686), .o (n2687) );
  assign n2688 = ~N18 & N73 ;
  assign n2689 = N18 & ~N322 ;
  assign n2690 = n2688 | n2689 ;
  buffer buf_n2691( .i (n2690), .o (n2691) );
  buffer buf_n2692( .i (n2691), .o (n2692) );
  assign n2693 = N18 & N204 ;
  assign n2694 = n2103 | n2693 ;
  buffer buf_n2695( .i (n2694), .o (n2695) );
  assign n2696 = n2692 & n2695 ;
  buffer buf_n2697( .i (n2696), .o (n2697) );
  buffer buf_n2698( .i (n2697), .o (n2698) );
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n2700( .i (n2699), .o (n2700) );
  assign n2701 = ~N18 & N74 ;
  assign n2702 = N18 & ~N313 ;
  assign n2703 = n2701 | n2702 ;
  buffer buf_n2704( .i (n2703), .o (n2704) );
  assign n2705 = N18 & N207 ;
  assign n2706 = n2168 | n2705 ;
  buffer buf_n2707( .i (n2706), .o (n2707) );
  assign n2708 = n2704 & n2707 ;
  assign n2709 = N70 | N89 ;
  assign n2710 = n209 & n2709 ;
  assign n2711 = N18 | N70 ;
  buffer buf_n2712( .i (n2711), .o (n2712) );
  assign n2713 = N89 & n2712 ;
  assign n2714 = n2710 | n2713 ;
  buffer buf_n2715( .i (n2714), .o (n2715) );
  assign n2716 = n2708 | n2715 ;
  assign n2717 = ~N18 & N76 ;
  assign n2718 = N18 & ~N316 ;
  assign n2719 = n2717 | n2718 ;
  buffer buf_n2720( .i (n2719), .o (n2720) );
  assign n2721 = N18 & N206 ;
  assign n2722 = n2158 | n2721 ;
  buffer buf_n2723( .i (n2722), .o (n2723) );
  assign n2724 = n2720 | n2723 ;
  assign n2725 = n2704 | n2707 ;
  assign n2726 = n2724 & n2725 ;
  assign n2727 = n2716 & n2726 ;
  assign n2728 = n2720 & n2723 ;
  assign n2729 = ~N18 & N75 ;
  assign n2730 = N18 & ~N319 ;
  assign n2731 = n2729 | n2730 ;
  buffer buf_n2732( .i (n2731), .o (n2732) );
  assign n2735 = N18 & N205 ;
  assign n2736 = n2135 | n2735 ;
  buffer buf_n2737( .i (n2736), .o (n2737) );
  assign n2738 = n2732 & n2737 ;
  assign n2739 = n2728 | n2738 ;
  buffer buf_n2740( .i (n2739), .o (n2740) );
  assign n2741 = n2727 | n2740 ;
  assign n2742 = n2692 | n2695 ;
  assign n2743 = n2732 | n2737 ;
  assign n2744 = n2742 & n2743 ;
  buffer buf_n2745( .i (n2744), .o (n2745) );
  buffer buf_n2746( .i (n2745), .o (n2746) );
  assign n2747 = n2741 & n2746 ;
  assign n2748 = n2700 | n2747 ;
  assign n2749 = n2687 & n2748 ;
  assign n2750 = ~N18 & N54 ;
  assign n2751 = N18 & ~N328 ;
  assign n2752 = n2750 | n2751 ;
  buffer buf_n2753( .i (n2752), .o (n2753) );
  assign n2756 = N18 & N202 ;
  assign n2757 = n2023 | n2756 ;
  buffer buf_n2758( .i (n2757), .o (n2758) );
  assign n2759 = n2753 & n2758 ;
  assign n2760 = n2678 & n2681 ;
  assign n2761 = n2759 | n2760 ;
  buffer buf_n2762( .i (n2761), .o (n2762) );
  buffer buf_n2763( .i (n2762), .o (n2763) );
  buffer buf_n2764( .i (n2763), .o (n2764) );
  buffer buf_n2765( .i (n2764), .o (n2765) );
  buffer buf_n2766( .i (n2765), .o (n2766) );
  assign n2767 = n2749 | n2766 ;
  assign n2768 = ~N18 & N56 ;
  assign n2769 = N18 & ~N334 ;
  assign n2770 = n2768 | n2769 ;
  buffer buf_n2771( .i (n2770), .o (n2771) );
  buffer buf_n2772( .i (n2771), .o (n2772) );
  assign n2773 = N18 & N200 ;
  assign n2774 = n1985 | n2773 ;
  buffer buf_n2775( .i (n2774), .o (n2775) );
  assign n2776 = n2772 | n2775 ;
  buffer buf_n2777( .i (n2776), .o (n2777) );
  assign n2778 = ~N18 & N55 ;
  assign n2779 = N18 & ~N331 ;
  assign n2780 = n2778 | n2779 ;
  buffer buf_n2781( .i (n2780), .o (n2781) );
  buffer buf_n2782( .i (n2781), .o (n2782) );
  assign n2783 = N18 & N201 ;
  assign n2784 = n2007 | n2783 ;
  buffer buf_n2785( .i (n2784), .o (n2785) );
  assign n2786 = n2782 & n2785 ;
  buffer buf_n2787( .i (n2786), .o (n2787) );
  assign n2788 = n2777 & ~n2787 ;
  assign n2789 = n2753 | n2758 ;
  assign n2790 = n2782 | n2785 ;
  assign n2791 = n2789 & n2790 ;
  buffer buf_n2792( .i (n2791), .o (n2792) );
  assign n2793 = n2788 & n2792 ;
  buffer buf_n2794( .i (n2793), .o (n2794) );
  buffer buf_n2795( .i (n2794), .o (n2795) );
  buffer buf_n2796( .i (n2795), .o (n2796) );
  buffer buf_n2797( .i (n2796), .o (n2797) );
  assign n2798 = n2767 & n2797 ;
  assign n2799 = n2777 & n2787 ;
  assign n2800 = n2772 & n2775 ;
  assign n2801 = ~N18 & N77 ;
  assign n2802 = N18 & ~N340 ;
  assign n2803 = n2801 | n2802 ;
  buffer buf_n2804( .i (n2803), .o (n2804) );
  assign n2805 = N18 & N187 ;
  assign n2806 = n1752 | n2805 ;
  buffer buf_n2807( .i (n2806), .o (n2807) );
  assign n2808 = n2804 & n2807 ;
  assign n2809 = n2800 | n2808 ;
  buffer buf_n2810( .i (n2809), .o (n2810) );
  assign n2811 = n2799 | n2810 ;
  buffer buf_n2812( .i (n2811), .o (n2812) );
  buffer buf_n2813( .i (n2812), .o (n2813) );
  buffer buf_n2814( .i (n2813), .o (n2814) );
  buffer buf_n2815( .i (n2814), .o (n2815) );
  buffer buf_n2816( .i (n2815), .o (n2816) );
  assign n2817 = n2798 | n2816 ;
  assign n2818 = ~N18 & N81 ;
  assign n2819 = N18 & ~N349 ;
  assign n2820 = n2818 | n2819 ;
  buffer buf_n2821( .i (n2820), .o (n2821) );
  buffer buf_n2822( .i (n2821), .o (n2822) );
  assign n2823 = N18 & N194 ;
  assign n2824 = n1823 | n2823 ;
  buffer buf_n2825( .i (n2824), .o (n2825) );
  assign n2826 = n2822 & n2825 ;
  assign n2827 = ~N18 & N80 ;
  assign n2828 = N18 & ~N352 ;
  assign n2829 = n2827 | n2828 ;
  buffer buf_n2830( .i (n2829), .o (n2830) );
  buffer buf_n2831( .i (n2830), .o (n2831) );
  assign n2832 = N18 & N193 ;
  assign n2833 = n1931 | n2832 ;
  buffer buf_n2834( .i (n2833), .o (n2834) );
  assign n2835 = n2831 & n2834 ;
  assign n2836 = n2826 | n2835 ;
  buffer buf_n2837( .i (n2836), .o (n2837) );
  buffer buf_n2838( .i (n2837), .o (n2838) );
  assign n2839 = ~N18 & N59 ;
  assign n2840 = N18 & ~N346 ;
  assign n2841 = n2839 | n2840 ;
  buffer buf_n2842( .i (n2841), .o (n2842) );
  assign n2843 = N18 & N195 ;
  assign n2844 = n1871 | n2843 ;
  buffer buf_n2845( .i (n2844), .o (n2845) );
  assign n2846 = n2842 | n2845 ;
  buffer buf_n2847( .i (n2846), .o (n2847) );
  buffer buf_n2848( .i (n2847), .o (n2848) );
  assign n2849 = n2822 | n2825 ;
  buffer buf_n2850( .i (n2849), .o (n2850) );
  assign n2851 = n2831 | n2834 ;
  buffer buf_n2852( .i (n2851), .o (n2852) );
  assign n2854 = n2850 & n2852 ;
  assign n2855 = n2848 & n2854 ;
  assign n2856 = ~n2838 & n2855 ;
  buffer buf_n2857( .i (n2856), .o (n2857) );
  assign n2858 = ~N18 & N78 ;
  assign n2859 = N18 & ~N343 ;
  assign n2860 = n2858 | n2859 ;
  buffer buf_n2861( .i (n2860), .o (n2861) );
  assign n2862 = N18 & N196 ;
  assign n2863 = n1782 | n2862 ;
  buffer buf_n2864( .i (n2863), .o (n2864) );
  assign n2865 = n2861 & n2864 ;
  assign n2866 = n2842 & n2845 ;
  assign n2867 = n2865 | n2866 ;
  buffer buf_n2868( .i (n2867), .o (n2868) );
  assign n2872 = n2804 | n2807 ;
  assign n2873 = n2861 | n2864 ;
  assign n2874 = n2872 & n2873 ;
  buffer buf_n2875( .i (n2874), .o (n2875) );
  assign n2876 = ~n2868 & n2875 ;
  buffer buf_n2877( .i (n2876), .o (n2877) );
  buffer buf_n2878( .i (n2877), .o (n2878) );
  assign n2879 = n2857 & n2878 ;
  buffer buf_n2880( .i (n2879), .o (n2880) );
  buffer buf_n2881( .i (n2880), .o (n2881) );
  buffer buf_n2882( .i (n2881), .o (n2882) );
  assign n2883 = n2817 & n2882 ;
  buffer buf_n2869( .i (n2868), .o (n2869) );
  buffer buf_n2870( .i (n2869), .o (n2870) );
  buffer buf_n2871( .i (n2870), .o (n2871) );
  assign n2884 = n2857 & n2871 ;
  buffer buf_n2853( .i (n2852), .o (n2853) );
  assign n2885 = n2837 & n2853 ;
  buffer buf_n2886( .i (n2885), .o (n2886) );
  buffer buf_n2887( .i (n2886), .o (n2887) );
  buffer buf_n2888( .i (n2887), .o (n2888) );
  assign n2889 = n2884 | n2888 ;
  buffer buf_n2890( .i (n2889), .o (n2890) );
  buffer buf_n2891( .i (n2890), .o (n2891) );
  buffer buf_n2892( .i (n2891), .o (n2892) );
  assign n2893 = n2883 | n2892 ;
  assign n2894 = ~N18 & N62 ;
  assign n2895 = N18 & ~N364 ;
  assign n2896 = n2894 | n2895 ;
  buffer buf_n2897( .i (n2896), .o (n2897) );
  buffer buf_n2898( .i (n2897), .o (n2898) );
  assign n2899 = N18 & N189 ;
  assign n2900 = n1472 | n2899 ;
  buffer buf_n2901( .i (n2900), .o (n2901) );
  assign n2902 = n2898 | n2901 ;
  buffer buf_n2903( .i (n2902), .o (n2903) );
  assign n2904 = ~N18 & N61 ;
  assign n2905 = N18 & ~N361 ;
  assign n2906 = n2904 | n2905 ;
  buffer buf_n2907( .i (n2906), .o (n2907) );
  buffer buf_n2908( .i (n2907), .o (n2908) );
  assign n2909 = N18 & N190 ;
  assign n2910 = n1534 | n2909 ;
  buffer buf_n2911( .i (n2910), .o (n2911) );
  assign n2912 = n2908 & n2911 ;
  buffer buf_n2913( .i (n2912), .o (n2913) );
  assign n2914 = n2903 & ~n2913 ;
  assign n2915 = n2898 & n2901 ;
  buffer buf_n2916( .i (n2915), .o (n2916) );
  assign n2918 = n2908 | n2911 ;
  buffer buf_n2919( .i (n2918), .o (n2919) );
  assign n2920 = ~n2916 & n2919 ;
  assign n2921 = n2914 & n2920 ;
  buffer buf_n2922( .i (n2921), .o (n2922) );
  assign n2923 = ~N18 & N60 ;
  assign n2924 = N18 & ~N358 ;
  assign n2925 = n2923 | n2924 ;
  buffer buf_n2926( .i (n2925), .o (n2926) );
  assign n2927 = N18 & N191 ;
  assign n2928 = n1554 | n2927 ;
  buffer buf_n2929( .i (n2928), .o (n2929) );
  assign n2930 = n2926 & n2929 ;
  assign n2931 = ~N18 & N79 ;
  assign n2932 = N18 & ~N355 ;
  assign n2933 = n2931 | n2932 ;
  buffer buf_n2934( .i (n2933), .o (n2934) );
  assign n2935 = N18 & N192 ;
  assign n2936 = n1566 | n2935 ;
  buffer buf_n2937( .i (n2936), .o (n2937) );
  assign n2938 = n2934 & n2937 ;
  assign n2939 = n2930 | n2938 ;
  buffer buf_n2940( .i (n2939), .o (n2940) );
  assign n2941 = n2926 | n2929 ;
  buffer buf_n2942( .i (n2941), .o (n2942) );
  assign n2944 = n2934 | n2937 ;
  buffer buf_n2945( .i (n2944), .o (n2945) );
  assign n2946 = n2942 & n2945 ;
  assign n2947 = ~n2940 & n2946 ;
  buffer buf_n2948( .i (n2947), .o (n2948) );
  assign n2949 = n2922 & n2948 ;
  buffer buf_n2950( .i (n2949), .o (n2950) );
  buffer buf_n2951( .i (n2950), .o (n2951) );
  buffer buf_n2952( .i (n2951), .o (n2952) );
  buffer buf_n2953( .i (n2952), .o (n2953) );
  buffer buf_n2954( .i (n2953), .o (n2954) );
  buffer buf_n2955( .i (n2954), .o (n2955) );
  assign n2956 = n2893 & n2955 ;
  buffer buf_n2943( .i (n2942), .o (n2943) );
  assign n2957 = n2940 & n2943 ;
  buffer buf_n2958( .i (n2957), .o (n2958) );
  assign n2959 = n2922 & n2958 ;
  buffer buf_n2917( .i (n2916), .o (n2917) );
  assign n2960 = n2903 & n2913 ;
  assign n2961 = n2917 | n2960 ;
  buffer buf_n2962( .i (n2961), .o (n2962) );
  buffer buf_n2963( .i (n2962), .o (n2963) );
  assign n2964 = n2959 | n2963 ;
  buffer buf_n2965( .i (n2964), .o (n2965) );
  buffer buf_n2966( .i (n2965), .o (n2966) );
  buffer buf_n2967( .i (n2966), .o (n2967) );
  buffer buf_n2968( .i (n2967), .o (n2968) );
  buffer buf_n2969( .i (n2968), .o (n2969) );
  buffer buf_n2970( .i (n2969), .o (n2970) );
  assign n2971 = n2956 | n2970 ;
  buffer buf_n2972( .i (n2971), .o (n2972) );
  assign n2973 = ~N18 & N64 ;
  assign n2974 = N18 & ~N289 ;
  assign n2975 = n2973 | n2974 ;
  buffer buf_n2976( .i (n2975), .o (n2976) );
  assign n2977 = ~N177 & N18 ;
  assign n2978 = n1061 | n2977 ;
  buffer buf_n2979( .i (n2978), .o (n2979) );
  assign n2980 = n2976 & ~n2979 ;
  assign n2981 = ~N18 & N85 ;
  assign n2982 = N18 & ~N286 ;
  assign n2983 = n2981 | n2982 ;
  buffer buf_n2984( .i (n2983), .o (n2984) );
  assign n2985 = N178 & N18 ;
  assign n2986 = n1090 | n2985 ;
  buffer buf_n2987( .i (n2986), .o (n2987) );
  assign n2988 = n2984 & n2987 ;
  assign n2989 = n2980 | n2988 ;
  buffer buf_n2990( .i (n2989), .o (n2990) );
  assign n2991 = ~n2976 & n2979 ;
  buffer buf_n2992( .i (n2991), .o (n2992) );
  assign n2994 = n2984 | n2987 ;
  buffer buf_n2995( .i (n2994), .o (n2995) );
  assign n2996 = ~n2992 & n2995 ;
  assign n2997 = ~n2990 & n2996 ;
  buffer buf_n2998( .i (n2997), .o (n2998) );
  assign n2999 = ~N18 & N84 ;
  assign n3000 = N18 & ~N283 ;
  assign n3001 = n2999 | n3000 ;
  buffer buf_n3002( .i (n3001), .o (n3002) );
  assign n3005 = N179 & N18 ;
  assign n3006 = n1112 | n3005 ;
  buffer buf_n3007( .i (n3006), .o (n3007) );
  assign n3008 = n3002 & n3007 ;
  assign n3009 = ~N18 & N83 ;
  assign n3010 = N18 & ~N280 ;
  assign n3011 = n3009 | n3010 ;
  buffer buf_n3012( .i (n3011), .o (n3012) );
  assign n3015 = N18 & N180 ;
  assign n3016 = n1130 | n3015 ;
  buffer buf_n3017( .i (n3016), .o (n3017) );
  assign n3018 = n3012 & n3017 ;
  assign n3019 = n3008 | n3018 ;
  buffer buf_n3020( .i (n3019), .o (n3020) );
  assign n3021 = n3002 | n3007 ;
  buffer buf_n3022( .i (n3021), .o (n3022) );
  assign n3024 = n3012 | n3017 ;
  buffer buf_n3025( .i (n3024), .o (n3025) );
  assign n3026 = n3022 & n3025 ;
  assign n3027 = ~n3020 & n3026 ;
  buffer buf_n3028( .i (n3027), .o (n3028) );
  buffer buf_n3029( .i (n3028), .o (n3029) );
  buffer buf_n3030( .i (n3029), .o (n3030) );
  assign n3031 = n2998 & n3030 ;
  buffer buf_n3032( .i (n3031), .o (n3032) );
  assign n3033 = ~N18 & N65 ;
  assign n3034 = N18 & ~N277 ;
  assign n3035 = n3033 | n3034 ;
  buffer buf_n3036( .i (n3035), .o (n3036) );
  buffer buf_n3037( .i (n3036), .o (n3037) );
  assign n3038 = N171 & N18 ;
  assign n3039 = n1139 | n3038 ;
  buffer buf_n3040( .i (n3039), .o (n3040) );
  assign n3041 = n3037 & n3040 ;
  buffer buf_n3042( .i (n3041), .o (n3042) );
  assign n3050 = n3037 | n3040 ;
  buffer buf_n3051( .i (n3050), .o (n3051) );
  assign n3052 = ~n3042 & n3051 ;
  buffer buf_n3053( .i (n3052), .o (n3053) );
  buffer buf_n3054( .i (n3053), .o (n3054) );
  buffer buf_n3055( .i (n3054), .o (n3055) );
  buffer buf_n3056( .i (n3055), .o (n3056) );
  buffer buf_n3057( .i (n3056), .o (n3057) );
  buffer buf_n3058( .i (n3057), .o (n3058) );
  assign n3059 = n3032 & n3058 ;
  buffer buf_n3060( .i (n3059), .o (n3060) );
  buffer buf_n3061( .i (n3060), .o (n3061) );
  buffer buf_n3062( .i (n3061), .o (n3062) );
  buffer buf_n3063( .i (n3062), .o (n3063) );
  buffer buf_n3064( .i (n3063), .o (n3064) );
  assign n3065 = n2972 & n3064 ;
  buffer buf_n3043( .i (n3042), .o (n3043) );
  buffer buf_n3044( .i (n3043), .o (n3044) );
  buffer buf_n3045( .i (n3044), .o (n3045) );
  buffer buf_n3046( .i (n3045), .o (n3046) );
  buffer buf_n3047( .i (n3046), .o (n3047) );
  buffer buf_n3048( .i (n3047), .o (n3048) );
  buffer buf_n3049( .i (n3048), .o (n3049) );
  assign n3066 = n3032 & n3049 ;
  buffer buf_n3023( .i (n3022), .o (n3023) );
  assign n3067 = n3020 & n3023 ;
  buffer buf_n3068( .i (n3067), .o (n3068) );
  buffer buf_n3069( .i (n3068), .o (n3069) );
  buffer buf_n3070( .i (n3069), .o (n3070) );
  assign n3071 = n2998 & n3070 ;
  buffer buf_n2993( .i (n2992), .o (n2993) );
  assign n3072 = n2990 & ~n2993 ;
  buffer buf_n3073( .i (n3072), .o (n3073) );
  buffer buf_n3074( .i (n3073), .o (n3074) );
  assign n3075 = n3071 | n3074 ;
  buffer buf_n3076( .i (n3075), .o (n3076) );
  assign n3077 = n3066 | n3076 ;
  buffer buf_n3078( .i (n3077), .o (n3078) );
  buffer buf_n3079( .i (n3078), .o (n3079) );
  buffer buf_n3080( .i (n3079), .o (n3080) );
  buffer buf_n3081( .i (n3080), .o (n3081) );
  buffer buf_n3082( .i (n3081), .o (n3082) );
  assign n3083 = n3065 | n3082 ;
  assign n3084 = N109 & ~N18 ;
  assign n3085 = N18 & ~N299 ;
  assign n3086 = n3084 | n3085 ;
  buffer buf_n3087( .i (n3086), .o (n3087) );
  assign n3088 = ~N174 & N18 ;
  buffer buf_n3089( .i (n3088), .o (n3089) );
  assign n3092 = n1061 | n3089 ;
  buffer buf_n3093( .i (n3092), .o (n3093) );
  assign n3094 = n3087 & ~n3093 ;
  assign n3095 = N110 & ~N18 ;
  assign n3096 = N18 & ~N303 ;
  assign n3097 = n3095 | n3096 ;
  buffer buf_n3098( .i (n3097), .o (n3098) );
  assign n3099 = ~N173 & N18 ;
  buffer buf_n3100( .i (n3099), .o (n3100) );
  assign n3103 = n1061 | n3100 ;
  buffer buf_n3104( .i (n3103), .o (n3104) );
  assign n3105 = n3098 & ~n3104 ;
  assign n3106 = n3094 | n3105 ;
  buffer buf_n3107( .i (n3106), .o (n3107) );
  assign n3108 = ~n3087 & n3093 ;
  buffer buf_n3109( .i (n3108), .o (n3109) );
  assign n3110 = ~n3098 & n3104 ;
  buffer buf_n3111( .i (n3110), .o (n3111) );
  assign n3113 = n3109 | n3111 ;
  assign n3114 = n3107 | n3113 ;
  buffer buf_n3115( .i (n3114), .o (n3115) );
  assign n3116 = ~N18 & N86 ;
  assign n3117 = N18 & ~N296 ;
  assign n3118 = n3116 | n3117 ;
  buffer buf_n3119( .i (n3118), .o (n3119) );
  buffer buf_n3120( .i (n3119), .o (n3120) );
  buffer buf_n3121( .i (n3120), .o (n3121) );
  buffer buf_n3122( .i (n3121), .o (n3122) );
  assign n3123 = ~N175 & N18 ;
  buffer buf_n3124( .i (n3123), .o (n3124) );
  buffer buf_n3127( .i (n417), .o (n3127) );
  assign n3128 = n3124 | n3127 ;
  buffer buf_n3129( .i (n3128), .o (n3129) );
  assign n3130 = n3122 & ~n3129 ;
  assign n3131 = ~N18 & N63 ;
  assign n3132 = N18 & ~N293 ;
  assign n3133 = n3131 | n3132 ;
  buffer buf_n3134( .i (n3133), .o (n3134) );
  buffer buf_n3135( .i (n3134), .o (n3135) );
  buffer buf_n3136( .i (n3135), .o (n3136) );
  buffer buf_n3137( .i (n3136), .o (n3137) );
  assign n3138 = ~N176 & N18 ;
  buffer buf_n3139( .i (n3138), .o (n3139) );
  assign n3142 = n3127 | n3139 ;
  buffer buf_n3143( .i (n3142), .o (n3143) );
  assign n3144 = n3137 & ~n3143 ;
  assign n3145 = n3130 | n3144 ;
  buffer buf_n3146( .i (n3145), .o (n3146) );
  assign n3147 = ~n3122 & n3129 ;
  buffer buf_n3148( .i (n3147), .o (n3148) );
  assign n3150 = ~n3137 & n3143 ;
  buffer buf_n3151( .i (n3150), .o (n3151) );
  assign n3152 = n3148 | n3151 ;
  assign n3153 = n3146 | n3152 ;
  buffer buf_n3154( .i (n3153), .o (n3154) );
  assign n3155 = n3115 | n3154 ;
  buffer buf_n3156( .i (n3155), .o (n3156) );
  buffer buf_n3157( .i (n3156), .o (n3157) );
  buffer buf_n3158( .i (n3157), .o (n3158) );
  buffer buf_n3159( .i (n3158), .o (n3159) );
  buffer buf_n3160( .i (n3159), .o (n3160) );
  buffer buf_n3161( .i (n3160), .o (n3161) );
  buffer buf_n3162( .i (n3161), .o (n3162) );
  buffer buf_n3163( .i (n3162), .o (n3163) );
  buffer buf_n3164( .i (n3163), .o (n3164) );
  assign n3165 = n3083 & ~n3164 ;
  buffer buf_n3149( .i (n3148), .o (n3149) );
  assign n3166 = n3146 & ~n3149 ;
  buffer buf_n3167( .i (n3166), .o (n3167) );
  assign n3168 = ~n3115 & n3167 ;
  buffer buf_n3112( .i (n3111), .o (n3112) );
  assign n3169 = n3107 & ~n3112 ;
  buffer buf_n3170( .i (n3169), .o (n3170) );
  buffer buf_n3171( .i (n3170), .o (n3171) );
  assign n3172 = n3168 | n3171 ;
  buffer buf_n3173( .i (n3172), .o (n3173) );
  buffer buf_n3174( .i (n3173), .o (n3174) );
  buffer buf_n3175( .i (n3174), .o (n3175) );
  buffer buf_n3176( .i (n3175), .o (n3176) );
  buffer buf_n3177( .i (n3176), .o (n3177) );
  buffer buf_n3178( .i (n3177), .o (n3178) );
  buffer buf_n3179( .i (n3178), .o (n3179) );
  buffer buf_n3180( .i (n3179), .o (n3180) );
  buffer buf_n3181( .i (n3180), .o (n3181) );
  assign n3182 = n3165 | n3181 ;
  assign n3183 = ~N18 & N87 ;
  assign n3184 = ~N106 & N18 ;
  assign n3185 = n3183 | n3184 ;
  buffer buf_n3186( .i (n3185), .o (n3186) );
  assign n3187 = ~N168 & N18 ;
  buffer buf_n3188( .i (n3187), .o (n3188) );
  assign n3191 = n3127 | n3188 ;
  buffer buf_n3192( .i (n3191), .o (n3192) );
  assign n3193 = ~n3186 & n3192 ;
  buffer buf_n3194( .i (n3193), .o (n3194) );
  buffer buf_n3195( .i (n3194), .o (n3195) );
  buffer buf_n3196( .i (n3195), .o (n3196) );
  assign n3197 = ~N18 & N88 ;
  assign n3198 = N18 & ~N260 ;
  assign n3199 = n3197 | n3198 ;
  buffer buf_n3200( .i (n3199), .o (n3200) );
  assign n3201 = ~N166 & N18 ;
  buffer buf_n3202( .i (n3201), .o (n3202) );
  assign n3205 = n3127 | n3202 ;
  buffer buf_n3206( .i (n3205), .o (n3206) );
  assign n3207 = ~n3200 & n3206 ;
  buffer buf_n3208( .i (n3207), .o (n3208) );
  assign n3210 = n3200 & ~n3206 ;
  buffer buf_n3211( .i (n3210), .o (n3211) );
  assign n3212 = n3208 | n3211 ;
  assign n3213 = N112 & ~N18 ;
  assign n3214 = N18 & ~N257 ;
  assign n3215 = n3213 | n3214 ;
  buffer buf_n3216( .i (n3215), .o (n3216) );
  assign n3217 = ~N167 & N18 ;
  buffer buf_n3218( .i (n3217), .o (n3218) );
  buffer buf_n3221( .i (n416), .o (n3221) );
  buffer buf_n3222( .i (n3221), .o (n3222) );
  assign n3223 = n3218 | n3222 ;
  buffer buf_n3224( .i (n3223), .o (n3224) );
  assign n3225 = n3216 & ~n3224 ;
  buffer buf_n3226( .i (n3225), .o (n3226) );
  assign n3227 = ~n3216 & n3224 ;
  buffer buf_n3228( .i (n3227), .o (n3228) );
  assign n3229 = n3226 | n3228 ;
  assign n3230 = n3212 | n3229 ;
  assign n3231 = n3196 | n3230 ;
  buffer buf_n3232( .i (n3231), .o (n3232) );
  buffer buf_n420( .i (n419), .o (n420) );
  assign n3233 = N113 & ~N18 ;
  assign n3234 = N18 & ~N251 ;
  assign n3235 = n3233 | n3234 ;
  buffer buf_n3236( .i (n3235), .o (n3236) );
  assign n3237 = ~n420 & n3236 ;
  assign n3238 = N111 & ~N18 ;
  assign n3239 = N18 & ~N254 ;
  assign n3240 = n3238 | n3239 ;
  buffer buf_n3241( .i (n3240), .o (n3241) );
  assign n3242 = ~N169 & N18 ;
  buffer buf_n3243( .i (n3242), .o (n3243) );
  assign n3246 = n3222 | n3243 ;
  buffer buf_n3247( .i (n3246), .o (n3247) );
  assign n3248 = n3241 & ~n3247 ;
  assign n3249 = n3237 | n3248 ;
  buffer buf_n3250( .i (n3249), .o (n3250) );
  buffer buf_n3251( .i (n3250), .o (n3251) );
  assign n3252 = n420 & ~n3236 ;
  buffer buf_n3253( .i (n3252), .o (n3253) );
  buffer buf_n3254( .i (n3253), .o (n3254) );
  assign n3255 = n3186 & ~n3192 ;
  buffer buf_n3256( .i (n3255), .o (n3256) );
  assign n3259 = ~n3241 & n3247 ;
  buffer buf_n3260( .i (n3259), .o (n3260) );
  assign n3262 = n3256 | n3260 ;
  assign n3263 = n3254 | n3262 ;
  assign n3264 = n3251 | n3263 ;
  buffer buf_n3265( .i (n3264), .o (n3265) );
  assign n3266 = n3232 | n3265 ;
  buffer buf_n3267( .i (n3266), .o (n3267) );
  buffer buf_n3268( .i (n3267), .o (n3268) );
  buffer buf_n3269( .i (n3268), .o (n3269) );
  buffer buf_n3270( .i (n3269), .o (n3270) );
  buffer buf_n3271( .i (n3270), .o (n3271) );
  buffer buf_n3272( .i (n3271), .o (n3272) );
  buffer buf_n3273( .i (n3272), .o (n3273) );
  buffer buf_n3274( .i (n3273), .o (n3274) );
  buffer buf_n3275( .i (n3274), .o (n3275) );
  buffer buf_n3276( .i (n3275), .o (n3276) );
  assign n3277 = n3182 & ~n3276 ;
  buffer buf_n3257( .i (n3256), .o (n3257) );
  buffer buf_n3258( .i (n3257), .o (n3258) );
  buffer buf_n3261( .i (n3260), .o (n3261) );
  assign n3278 = n3250 & ~n3261 ;
  assign n3279 = n3258 | n3278 ;
  buffer buf_n3280( .i (n3279), .o (n3280) );
  assign n3281 = ~n3232 & n3280 ;
  assign n3282 = N245 | N271 ;
  buffer buf_n3283( .i (n3282), .o (n3283) );
  assign n3284 = N382 & ~n3283 ;
  assign n3285 = N38 & ~n3284 ;
  buffer buf_n3286( .i (n3285), .o (n3286) );
  buffer buf_n3287( .i (n3286), .o (n3287) );
  buffer buf_n3209( .i (n3208), .o (n3209) );
  assign n3288 = n3211 | n3226 ;
  assign n3289 = ~n3209 & n3288 ;
  assign n3290 = n3287 | n3289 ;
  buffer buf_n3291( .i (n3290), .o (n3291) );
  buffer buf_n3292( .i (n3291), .o (n3292) );
  assign n3293 = n3281 | n3292 ;
  buffer buf_n3294( .i (n3293), .o (n3294) );
  buffer buf_n3295( .i (n3294), .o (n3295) );
  buffer buf_n3296( .i (n3295), .o (n3296) );
  buffer buf_n3297( .i (n3296), .o (n3297) );
  buffer buf_n3298( .i (n3297), .o (n3298) );
  buffer buf_n3299( .i (n3298), .o (n3299) );
  buffer buf_n3300( .i (n3299), .o (n3300) );
  buffer buf_n3301( .i (n3300), .o (n3301) );
  buffer buf_n3302( .i (n3301), .o (n3302) );
  buffer buf_n3303( .i (n3302), .o (n3303) );
  assign n3304 = n3277 | n3303 ;
  assign n3305 = ~n2673 & n3304 ;
  buffer buf_n3306( .i (n3305), .o (n3306) );
  assign n3307 = n2107 | n2121 ;
  buffer buf_n3308( .i (n3307), .o (n3308) );
  buffer buf_n3309( .i (n3308), .o (n3309) );
  buffer buf_n3310( .i (n3309), .o (n3310) );
  buffer buf_n3311( .i (n3310), .o (n3311) );
  buffer buf_n3312( .i (n3311), .o (n3312) );
  buffer buf_n3313( .i (n3312), .o (n3313) );
  buffer buf_n3314( .i (n3313), .o (n3314) );
  buffer buf_n3315( .i (n3314), .o (n3315) );
  buffer buf_n3316( .i (n3315), .o (n3316) );
  buffer buf_n3317( .i (n3316), .o (n3317) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2194( .i (n2193), .o (n2194) );
  assign n3318 = N367 & ~n2214 ;
  buffer buf_n3319( .i (n3318), .o (n3319) );
  assign n3320 = n2194 | n3319 ;
  assign n3321 = ~n2148 & n3320 ;
  buffer buf_n3322( .i (n3321), .o (n3322) );
  assign n3323 = ~n3317 & n3322 ;
  assign n3324 = n3317 & ~n3322 ;
  assign n3325 = ~n3323 & ~n3324 ;
  buffer buf_n2221( .i (n2220), .o (n2221) );
  buffer buf_n2222( .i (n2221), .o (n2222) );
  buffer buf_n2223( .i (n2222), .o (n2223) );
  buffer buf_n2224( .i (n2223), .o (n2224) );
  buffer buf_n2189( .i (n2188), .o (n2189) );
  buffer buf_n2190( .i (n2189), .o (n2190) );
  buffer buf_n2191( .i (n2190), .o (n2191) );
  assign n3326 = n2191 | n3319 ;
  buffer buf_n3327( .i (n3326), .o (n3327) );
  assign n3328 = n2224 & n3327 ;
  assign n3329 = n2224 | n3327 ;
  assign n3330 = n3328 | ~n3329 ;
  buffer buf_n2206( .i (n2205), .o (n2206) );
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n2175( .i (n2174), .o (n2175) );
  assign n3331 = n213 | n2181 ;
  buffer buf_n3332( .i (n3331), .o (n3332) );
  assign n3333 = n229 | n3332 ;
  assign n3334 = ~n2175 & n3333 ;
  buffer buf_n3335( .i (n3334), .o (n3335) );
  assign n3336 = n2206 & n3335 ;
  assign n3337 = n2206 | n3335 ;
  assign n3338 = n3336 | ~n3337 ;
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  assign n3339 = n215 | n229 ;
  buffer buf_n3340( .i (n3339), .o (n3340) );
  assign n3341 = n2210 | n3340 ;
  assign n3342 = n2210 & n3340 ;
  assign n3343 = ~n3341 | n3342 ;
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n2321( .i (n2320), .o (n2321) );
  buffer buf_n2322( .i (n2321), .o (n2322) );
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2325( .i (n2324), .o (n2325) );
  buffer buf_n2326( .i (n2325), .o (n2326) );
  buffer buf_n2327( .i (n2326), .o (n2327) );
  buffer buf_n2328( .i (n2327), .o (n2328) );
  buffer buf_n2329( .i (n2328), .o (n2329) );
  buffer buf_n2330( .i (n2329), .o (n2330) );
  buffer buf_n2331( .i (n2330), .o (n2331) );
  buffer buf_n2079( .i (n2078), .o (n2079) );
  buffer buf_n2080( .i (n2079), .o (n2080) );
  buffer buf_n2081( .i (n2080), .o (n2081) );
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2089( .i (n2088), .o (n2089) );
  buffer buf_n2295( .i (n2294), .o (n2295) );
  buffer buf_n2296( .i (n2295), .o (n2296) );
  assign n3344 = n2291 | n2296 ;
  buffer buf_n3345( .i (n3344), .o (n3345) );
  buffer buf_n3346( .i (n3345), .o (n3346) );
  buffer buf_n3347( .i (n3346), .o (n3347) );
  buffer buf_n3348( .i (n3347), .o (n3348) );
  buffer buf_n3349( .i (n3348), .o (n3349) );
  buffer buf_n3350( .i (n3349), .o (n3350) );
  buffer buf_n3351( .i (n3350), .o (n3351) );
  buffer buf_n3352( .i (n3351), .o (n3352) );
  buffer buf_n3353( .i (n3352), .o (n3353) );
  buffer buf_n3354( .i (n3353), .o (n3354) );
  assign n3355 = n2234 & ~n3354 ;
  assign n3356 = n2089 | n3355 ;
  buffer buf_n3357( .i (n3356), .o (n3357) );
  assign n3358 = n2331 | n3357 ;
  assign n3359 = n2331 & n3357 ;
  assign n3360 = ~n3358 | n3359 ;
  buffer buf_n2297( .i (n2296), .o (n2297) );
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  buffer buf_n2307( .i (n2306), .o (n2307) );
  buffer buf_n2308( .i (n2307), .o (n2308) );
  buffer buf_n2309( .i (n2308), .o (n2309) );
  buffer buf_n2310( .i (n2309), .o (n2310) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  buffer buf_n2064( .i (n2063), .o (n2064) );
  buffer buf_n2065( .i (n2064), .o (n2065) );
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n2073( .i (n2072), .o (n2073) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n2075( .i (n2074), .o (n2075) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  buffer buf_n2250( .i (n2249), .o (n2250) );
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  buffer buf_n2265( .i (n2264), .o (n2265) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  buffer buf_n2269( .i (n2268), .o (n2269) );
  buffer buf_n2270( .i (n2269), .o (n2270) );
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2273( .i (n2272), .o (n2273) );
  assign n3361 = n2234 & ~n2273 ;
  buffer buf_n3362( .i (n3361), .o (n3362) );
  assign n3363 = ~n2253 & n3362 ;
  assign n3364 = n2075 | n3363 ;
  buffer buf_n3365( .i (n3364), .o (n3365) );
  assign n3366 = n2312 | n3365 ;
  assign n3367 = n2312 & n3365 ;
  assign n3368 = ~n3366 | n3367 ;
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  buffer buf_n2055( .i (n2054), .o (n2055) );
  buffer buf_n2056( .i (n2055), .o (n2056) );
  assign n3369 = n2056 | n3362 ;
  buffer buf_n3370( .i (n3369), .o (n3370) );
  assign n3371 = n2255 | n3370 ;
  assign n3372 = n2255 & n3370 ;
  assign n3373 = ~n3371 | n3372 ;
  buffer buf_n2235( .i (n2234), .o (n2235) );
  buffer buf_n2276( .i (n2275), .o (n2276) );
  buffer buf_n2277( .i (n2276), .o (n2277) );
  buffer buf_n2278( .i (n2277), .o (n2278) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  buffer buf_n2280( .i (n2279), .o (n2280) );
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n2289( .i (n2288), .o (n2289) );
  assign n3374 = n2235 & n2289 ;
  assign n3375 = n2235 | n2289 ;
  assign n3376 = n3374 | ~n3375 ;
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  assign n3377 = n739 & ~n816 ;
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  assign n3378 = ~n741 & n814 ;
  assign n3379 = n3377 | n3378 ;
  buffer buf_n3380( .i (n3379), .o (n3380) );
  buffer buf_n3381( .i (n3380), .o (n3381) );
  buffer buf_n3382( .i (n3381), .o (n3382) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  assign n3383 = n832 & ~n849 ;
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  assign n3384 = ~n834 & n847 ;
  assign n3385 = n3383 | n3384 ;
  buffer buf_n3386( .i (n3385), .o (n3386) );
  assign n3387 = N141 & ~N18 ;
  buffer buf_n3388( .i (n3387), .o (n3388) );
  assign n3389 = N161 & N18 ;
  assign n3390 = n3388 | n3389 ;
  buffer buf_n3391( .i (n3390), .o (n3391) );
  assign n3392 = n1142 | n3391 ;
  assign n3393 = n1142 & n3391 ;
  assign n3394 = n3392 & ~n3393 ;
  buffer buf_n3395( .i (n3394), .o (n3395) );
  buffer buf_n3396( .i (n3395), .o (n3396) );
  buffer buf_n3397( .i (n3396), .o (n3397) );
  assign n3398 = n3386 | n3397 ;
  assign n3399 = n3386 & n3397 ;
  assign n3400 = n3398 & ~n3399 ;
  buffer buf_n3401( .i (n3400), .o (n3401) );
  assign n3402 = n3382 & ~n3401 ;
  assign n3403 = ~n3382 & n3401 ;
  assign n3404 = n3402 | n3403 ;
  buffer buf_n3405( .i (n3404), .o (n3405) );
  assign n3406 = n1063 & ~n1093 ;
  assign n3407 = ~n1063 & n1093 ;
  assign n3408 = n3406 | n3407 ;
  buffer buf_n3409( .i (n3408), .o (n3409) );
  assign n3410 = n1115 & n1133 ;
  assign n3411 = n1115 | n1133 ;
  assign n3412 = ~n3410 & n3411 ;
  buffer buf_n3413( .i (n3412), .o (n3413) );
  buffer buf_n3414( .i (n3413), .o (n3414) );
  buffer buf_n3415( .i (n3414), .o (n3415) );
  assign n3416 = n3409 & n3415 ;
  assign n3417 = n3409 | n3415 ;
  assign n3418 = ~n3416 & n3417 ;
  buffer buf_n3419( .i (n3418), .o (n3419) );
  buffer buf_n3420( .i (n3419), .o (n3420) );
  buffer buf_n3421( .i (n3420), .o (n3421) );
  buffer buf_n3422( .i (n3421), .o (n3422) );
  assign n3423 = ~n3405 & n3422 ;
  buffer buf_n3424( .i (n3423), .o (n3424) );
  assign n3425 = n518 & ~n3222 ;
  buffer buf_n3426( .i (n3425), .o (n3426) );
  buffer buf_n3427( .i (n3426), .o (n3427) );
  buffer buf_n3428( .i (n3427), .o (n3428) );
  buffer buf_n3429( .i (n3428), .o (n3429) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  assign n3430 = n424 & ~n435 ;
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  assign n3431 = ~n426 & n433 ;
  assign n3432 = n3430 | n3431 ;
  buffer buf_n3433( .i (n3432), .o (n3433) );
  assign n3434 = n3429 | n3433 ;
  assign n3435 = n3429 & n3433 ;
  assign n3436 = n3434 & ~n3435 ;
  buffer buf_n3437( .i (n3436), .o (n3437) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  assign n3438 = n490 & ~n512 ;
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  assign n3439 = ~n492 & n509 ;
  assign n3440 = n3438 | n3439 ;
  buffer buf_n3441( .i (n3440), .o (n3441) );
  assign n3442 = N18 & ~n419 ;
  buffer buf_n3443( .i (n3442), .o (n3443) );
  assign n3444 = N211 | N212 ;
  assign n3445 = N211 & N212 ;
  assign n3446 = n3444 & ~n3445 ;
  assign n3447 = n3443 & n3446 ;
  buffer buf_n3448( .i (n3447), .o (n3448) );
  assign n3449 = ~n3441 & n3448 ;
  assign n3450 = n3441 & ~n3448 ;
  assign n3451 = n3449 | n3450 ;
  buffer buf_n3452( .i (n3451), .o (n3452) );
  assign n3453 = n3437 | n3452 ;
  assign n3454 = n3437 & n3452 ;
  assign n3455 = n3453 & ~n3454 ;
  buffer buf_n3456( .i (n3455), .o (n3456) );
  buffer buf_n3457( .i (n3456), .o (n3457) );
  assign n3458 = n3405 & ~n3422 ;
  assign n3459 = n3457 | n3458 ;
  assign n3460 = n3424 | n3459 ;
  assign n3461 = N18 & N229 ;
  assign n3462 = n209 | n3461 ;
  buffer buf_n3463( .i (n3462), .o (n3463) );
  assign n3464 = ~n2009 & n3463 ;
  assign n3465 = n2009 & ~n3463 ;
  assign n3466 = n3464 | n3465 ;
  buffer buf_n3467( .i (n3466), .o (n3467) );
  assign n3468 = n1987 & ~n2137 ;
  assign n3469 = ~n1987 & n2137 ;
  assign n3470 = n3468 | n3469 ;
  buffer buf_n3471( .i (n3470), .o (n3471) );
  assign n3472 = ~n3467 & n3471 ;
  assign n3473 = n3467 & ~n3471 ;
  assign n3474 = n3472 | n3473 ;
  buffer buf_n3475( .i (n3474), .o (n3475) );
  buffer buf_n3476( .i (n3475), .o (n3476) );
  buffer buf_n3477( .i (n3476), .o (n3477) );
  buffer buf_n3478( .i (n3477), .o (n3478) );
  assign n3479 = ~n2105 & n2160 ;
  assign n3480 = n2105 & ~n2160 ;
  assign n3481 = n3479 | n3480 ;
  buffer buf_n3482( .i (n3481), .o (n3482) );
  buffer buf_n3483( .i (n3482), .o (n3483) );
  buffer buf_n3484( .i (n3483), .o (n3484) );
  buffer buf_n3485( .i (n3484), .o (n3485) );
  assign n3486 = n2025 & ~n2036 ;
  assign n3487 = ~n2025 & n2036 ;
  assign n3488 = n3486 | n3487 ;
  buffer buf_n3489( .i (n3488), .o (n3489) );
  assign n3490 = N18 & N239 ;
  assign n3491 = ~N18 & N44 ;
  buffer buf_n3492( .i (n3491), .o (n3492) );
  assign n3493 = n3490 | n3492 ;
  buffer buf_n3494( .i (n3493), .o (n3494) );
  assign n3495 = n2170 | n3494 ;
  assign n3496 = n2170 & n3494 ;
  assign n3497 = n3495 & ~n3496 ;
  buffer buf_n3498( .i (n3497), .o (n3498) );
  assign n3499 = n3489 & ~n3498 ;
  assign n3500 = ~n3489 & n3498 ;
  assign n3501 = n3499 | n3500 ;
  buffer buf_n3502( .i (n3501), .o (n3502) );
  assign n3503 = n3485 | n3502 ;
  assign n3504 = n3485 & n3502 ;
  assign n3505 = n3503 & ~n3504 ;
  buffer buf_n3506( .i (n3505), .o (n3506) );
  assign n3507 = ~n3478 & n3506 ;
  assign n3508 = n3478 & ~n3506 ;
  assign n3509 = n3507 | n3508 ;
  assign n3510 = ~n1825 & n1933 ;
  assign n3511 = n1825 & ~n1933 ;
  assign n3512 = n3510 | n3511 ;
  buffer buf_n3513( .i (n3512), .o (n3513) );
  assign n3514 = n1784 & n1873 ;
  assign n3515 = n1784 | n1873 ;
  assign n3516 = ~n3514 & n3515 ;
  buffer buf_n3517( .i (n3516), .o (n3517) );
  assign n3518 = n3513 & ~n3517 ;
  assign n3519 = ~n3513 & n3517 ;
  assign n3520 = n3518 | n3519 ;
  buffer buf_n3521( .i (n3520), .o (n3521) );
  buffer buf_n3522( .i (n3521), .o (n3522) );
  buffer buf_n3523( .i (n3522), .o (n3523) );
  buffer buf_n3524( .i (n3523), .o (n3524) );
  assign n3525 = N18 & N227 ;
  assign n3526 = N115 & ~N18 ;
  buffer buf_n3527( .i (n3526), .o (n3527) );
  assign n3528 = n3525 | n3527 ;
  buffer buf_n3529( .i (n3528), .o (n3529) );
  assign n3530 = n1754 | n3529 ;
  assign n3531 = n1754 & n3529 ;
  assign n3532 = n3530 & ~n3531 ;
  buffer buf_n3533( .i (n3532), .o (n3533) );
  buffer buf_n3534( .i (n3533), .o (n3534) );
  buffer buf_n3535( .i (n3534), .o (n3535) );
  buffer buf_n3536( .i (n3535), .o (n3536) );
  assign n3537 = n1474 & ~n1536 ;
  assign n3538 = ~n1474 & n1536 ;
  assign n3539 = n3537 | n3538 ;
  buffer buf_n3540( .i (n3539), .o (n3540) );
  assign n3541 = n1556 & n1568 ;
  assign n3542 = n1556 | n1568 ;
  assign n3543 = ~n3541 & n3542 ;
  buffer buf_n3544( .i (n3543), .o (n3544) );
  assign n3545 = n3540 | n3544 ;
  assign n3546 = n3540 & n3544 ;
  assign n3547 = n3545 & ~n3546 ;
  buffer buf_n3548( .i (n3547), .o (n3548) );
  assign n3549 = ~n3536 & n3548 ;
  assign n3550 = n3536 & ~n3548 ;
  assign n3551 = n3549 | n3550 ;
  buffer buf_n3552( .i (n3551), .o (n3552) );
  assign n3553 = n3524 & ~n3552 ;
  assign n3554 = ~n3524 & n3552 ;
  assign n3555 = n3553 | n3554 ;
  assign n3556 = n3509 & n3555 ;
  buffer buf_n3557( .i (n3556), .o (n3557) );
  buffer buf_n3558( .i (n3557), .o (n3558) );
  assign n3559 = ~n3460 & n3558 ;
  buffer buf_n3560( .i (n3559), .o (n3560) );
  inverter inv_n5030( .i (n3560), .o (n5030) );
  assign n3561 = N114 & ~N18 ;
  assign n3562 = N18 & ~N248 ;
  assign n3563 = n3561 | n3562 ;
  buffer buf_n3564( .i (n3563), .o (n3564) );
  assign n3565 = n3236 & n3564 ;
  assign n3566 = n3236 | n3564 ;
  assign n3567 = ~n3565 & n3566 ;
  buffer buf_n3568( .i (n3567), .o (n3568) );
  assign n3569 = n3200 & ~n3216 ;
  assign n3570 = ~n3200 & n3216 ;
  assign n3571 = n3569 | n3570 ;
  buffer buf_n3572( .i (n3571), .o (n3572) );
  assign n3573 = ~n3568 & n3572 ;
  assign n3574 = n3568 & ~n3572 ;
  assign n3575 = n3573 | n3574 ;
  buffer buf_n3576( .i (n3575), .o (n3576) );
  assign n3577 = n3186 & n3241 ;
  assign n3578 = n3186 | n3241 ;
  assign n3579 = ~n3577 & n3578 ;
  buffer buf_n3580( .i (n3579), .o (n3580) );
  assign n3581 = N263 & ~N267 ;
  assign n3582 = ~N263 & N267 ;
  assign n3583 = n3581 | n3582 ;
  assign n3584 = N18 & n3583 ;
  assign n3585 = N18 | n2652 ;
  assign n3586 = n3283 & ~n3585 ;
  assign n3587 = n3584 | n3586 ;
  buffer buf_n3588( .i (n3587), .o (n3588) );
  assign n3589 = ~n3580 & n3588 ;
  assign n3590 = n3580 & ~n3588 ;
  assign n3591 = n3589 | n3590 ;
  buffer buf_n3592( .i (n3591), .o (n3592) );
  assign n3593 = ~n3576 & n3592 ;
  assign n3594 = n3576 & ~n3592 ;
  assign n3595 = n3593 | n3594 ;
  assign n3596 = N18 & N310 ;
  assign n3597 = n2712 & ~n3596 ;
  buffer buf_n3598( .i (n3597), .o (n3598) );
  assign n3599 = ~N18 & N69 ;
  assign n3600 = N18 & ~N307 ;
  assign n3601 = n3599 | n3600 ;
  buffer buf_n3602( .i (n3601), .o (n3602) );
  assign n3603 = n3598 & n3602 ;
  assign n3604 = n3598 | n3602 ;
  assign n3605 = ~n3603 & n3604 ;
  buffer buf_n3606( .i (n3605), .o (n3606) );
  assign n3607 = n2704 & n2720 ;
  assign n3608 = n2704 | n2720 ;
  assign n3609 = ~n3607 & n3608 ;
  buffer buf_n3610( .i (n3609), .o (n3610) );
  assign n3611 = n3606 & ~n3610 ;
  assign n3612 = ~n3606 & n3610 ;
  assign n3613 = n3611 | n3612 ;
  buffer buf_n3614( .i (n3613), .o (n3614) );
  buffer buf_n3615( .i (n3614), .o (n3615) );
  buffer buf_n3616( .i (n3615), .o (n3616) );
  buffer buf_n2754( .i (n2753), .o (n2754) );
  buffer buf_n2755( .i (n2754), .o (n2755) );
  assign n3617 = n2771 & ~n2781 ;
  assign n3618 = ~n2771 & n2781 ;
  assign n3619 = n3617 | n3618 ;
  buffer buf_n3620( .i (n3619), .o (n3620) );
  assign n3621 = n2755 & ~n3620 ;
  assign n3622 = ~n2755 & n3620 ;
  assign n3623 = n3621 | n3622 ;
  buffer buf_n3624( .i (n3623), .o (n3624) );
  buffer buf_n2733( .i (n2732), .o (n2733) );
  buffer buf_n2734( .i (n2733), .o (n2734) );
  assign n3625 = n2677 & n2691 ;
  assign n3626 = n2677 | n2691 ;
  assign n3627 = ~n3625 & n3626 ;
  buffer buf_n3628( .i (n3627), .o (n3628) );
  assign n3629 = n2734 & n3628 ;
  assign n3630 = n2734 | n3628 ;
  assign n3631 = ~n3629 & n3630 ;
  buffer buf_n3632( .i (n3631), .o (n3632) );
  assign n3633 = ~n3624 & n3632 ;
  assign n3634 = n3624 & ~n3632 ;
  assign n3635 = n3633 | n3634 ;
  buffer buf_n3636( .i (n3635), .o (n3636) );
  assign n3637 = ~n3616 & n3636 ;
  assign n3638 = n3616 & ~n3636 ;
  assign n3639 = n3637 | n3638 ;
  assign n3640 = n3595 & n3639 ;
  assign n3641 = n2821 & n2830 ;
  assign n3642 = n2821 | n2830 ;
  assign n3643 = ~n3641 & n3642 ;
  buffer buf_n3644( .i (n3643), .o (n3644) );
  assign n3645 = n2897 & ~n2907 ;
  assign n3646 = ~n2897 & n2907 ;
  assign n3647 = n3645 | n3646 ;
  buffer buf_n3648( .i (n3647), .o (n3648) );
  assign n3649 = n3644 | n3648 ;
  assign n3650 = n3644 & n3648 ;
  assign n3651 = n3649 & ~n3650 ;
  buffer buf_n3652( .i (n3651), .o (n3652) );
  assign n3653 = n2842 & n2861 ;
  assign n3654 = n2842 | n2861 ;
  assign n3655 = ~n3653 & n3654 ;
  buffer buf_n3656( .i (n3655), .o (n3656) );
  buffer buf_n3657( .i (n3656), .o (n3657) );
  buffer buf_n3658( .i (n3657), .o (n3658) );
  assign n3659 = ~n3652 & n3658 ;
  assign n3660 = n3652 & ~n3658 ;
  assign n3661 = n3659 | n3660 ;
  buffer buf_n3662( .i (n3661), .o (n3662) );
  assign n3663 = n2926 & n2934 ;
  assign n3664 = n2926 | n2934 ;
  assign n3665 = ~n3663 & n3664 ;
  buffer buf_n3666( .i (n3665), .o (n3666) );
  assign n3667 = ~N18 & N58 ;
  assign n3668 = N18 & ~N337 ;
  assign n3669 = n3667 | n3668 ;
  buffer buf_n3670( .i (n3669), .o (n3670) );
  assign n3671 = n2804 & n3670 ;
  assign n3672 = n2804 | n3670 ;
  assign n3673 = ~n3671 & n3672 ;
  buffer buf_n3674( .i (n3673), .o (n3674) );
  assign n3675 = n3666 | n3674 ;
  assign n3676 = n3666 & n3674 ;
  assign n3677 = n3675 & ~n3676 ;
  buffer buf_n3678( .i (n3677), .o (n3678) );
  buffer buf_n3679( .i (n3678), .o (n3679) );
  buffer buf_n3680( .i (n3679), .o (n3680) );
  assign n3681 = n3662 & ~n3680 ;
  assign n3682 = ~n3662 & n3680 ;
  assign n3683 = n3681 | n3682 ;
  assign n3684 = n2976 & n2984 ;
  assign n3685 = n2976 | n2984 ;
  assign n3686 = ~n3684 & n3685 ;
  buffer buf_n3687( .i (n3686), .o (n3687) );
  assign n3688 = ~n3087 & n3098 ;
  assign n3689 = n3087 & ~n3098 ;
  assign n3690 = n3688 | n3689 ;
  buffer buf_n3691( .i (n3690), .o (n3691) );
  assign n3692 = ~n3687 & n3691 ;
  assign n3693 = n3687 & ~n3691 ;
  assign n3694 = n3692 | n3693 ;
  buffer buf_n3695( .i (n3694), .o (n3695) );
  buffer buf_n3003( .i (n3002), .o (n3003) );
  buffer buf_n3004( .i (n3003), .o (n3004) );
  assign n3696 = ~N18 & N82 ;
  assign n3697 = N18 & ~N274 ;
  assign n3698 = n3696 | n3697 ;
  buffer buf_n3699( .i (n3698), .o (n3699) );
  assign n3700 = n3036 & ~n3699 ;
  assign n3701 = ~n3036 & n3699 ;
  assign n3702 = n3700 | n3701 ;
  buffer buf_n3703( .i (n3702), .o (n3703) );
  assign n3704 = n3004 | n3703 ;
  assign n3705 = n3004 & n3703 ;
  assign n3706 = n3704 & ~n3705 ;
  buffer buf_n3707( .i (n3706), .o (n3707) );
  buffer buf_n3013( .i (n3012), .o (n3013) );
  buffer buf_n3014( .i (n3013), .o (n3014) );
  assign n3708 = n3119 & ~n3134 ;
  assign n3709 = ~n3119 & n3134 ;
  assign n3710 = n3708 | n3709 ;
  buffer buf_n3711( .i (n3710), .o (n3711) );
  assign n3712 = n3014 & n3711 ;
  assign n3713 = n3014 | n3711 ;
  assign n3714 = ~n3712 & n3713 ;
  buffer buf_n3715( .i (n3714), .o (n3715) );
  assign n3716 = n3707 & n3715 ;
  assign n3717 = n3707 | n3715 ;
  assign n3718 = ~n3716 & n3717 ;
  buffer buf_n3719( .i (n3718), .o (n3719) );
  assign n3720 = n3695 & n3719 ;
  assign n3721 = n3695 | n3719 ;
  assign n3722 = ~n3720 & n3721 ;
  assign n3723 = n3683 & n3722 ;
  assign n3724 = n3640 & n3723 ;
  buffer buf_n3725( .i (n3724), .o (n3725) );
  inverter inv_n5031( .i (n3725), .o (n5031) );
  assign n3729 = ~N170 & n3443 ;
  buffer buf_n3730( .i (n3729), .o (n3730) );
  buffer buf_n3203( .i (n3202), .o (n3203) );
  buffer buf_n3204( .i (n3203), .o (n3204) );
  assign n3731 = n3204 & ~n3224 ;
  buffer buf_n3219( .i (n3218), .o (n3219) );
  buffer buf_n3220( .i (n3219), .o (n3220) );
  assign n3732 = ~n3206 & n3220 ;
  assign n3733 = n3731 | n3732 ;
  buffer buf_n3734( .i (n3733), .o (n3734) );
  assign n3735 = ~n3730 & n3734 ;
  assign n3736 = n3730 & ~n3734 ;
  assign n3737 = n3735 | n3736 ;
  buffer buf_n3738( .i (n3737), .o (n3738) );
  buffer buf_n3189( .i (n3188), .o (n3189) );
  buffer buf_n3190( .i (n3189), .o (n3190) );
  assign n3739 = n3190 & ~n3247 ;
  buffer buf_n3244( .i (n3243), .o (n3244) );
  buffer buf_n3245( .i (n3244), .o (n3245) );
  assign n3740 = ~n3192 & n3245 ;
  assign n3741 = n3739 | n3740 ;
  buffer buf_n3742( .i (n3741), .o (n3742) );
  assign n3743 = ~N164 & N165 ;
  assign n3744 = N164 & ~N165 ;
  assign n3745 = n3743 | n3744 ;
  assign n3746 = n3443 & n3745 ;
  buffer buf_n3747( .i (n3746), .o (n3747) );
  assign n3748 = n3742 | n3747 ;
  assign n3749 = n3742 & n3747 ;
  assign n3750 = n3748 & ~n3749 ;
  buffer buf_n3751( .i (n3750), .o (n3751) );
  assign n3752 = n3738 | n3751 ;
  assign n3753 = n3738 & n3751 ;
  assign n3754 = n3752 & ~n3753 ;
  buffer buf_n3755( .i (n3754), .o (n3755) );
  assign n3756 = n2845 & n2864 ;
  assign n3757 = n2845 | n2864 ;
  assign n3758 = ~n3756 & n3757 ;
  buffer buf_n3759( .i (n3758), .o (n3759) );
  buffer buf_n3760( .i (n3759), .o (n3760) );
  buffer buf_n3761( .i (n3760), .o (n3761) );
  buffer buf_n3762( .i (n3761), .o (n3762) );
  assign n3763 = n2901 & ~n2911 ;
  assign n3764 = ~n2901 & n2911 ;
  assign n3765 = n3763 | n3764 ;
  buffer buf_n3766( .i (n3765), .o (n3766) );
  assign n3767 = n2929 & n2937 ;
  assign n3768 = n2929 | n2937 ;
  assign n3769 = ~n3767 & n3768 ;
  buffer buf_n3770( .i (n3769), .o (n3770) );
  assign n3771 = ~n3766 & n3770 ;
  assign n3772 = n3766 & ~n3770 ;
  assign n3773 = n3771 | n3772 ;
  buffer buf_n3774( .i (n3773), .o (n3774) );
  assign n3775 = n3762 & n3774 ;
  assign n3776 = n3762 | n3774 ;
  assign n3777 = ~n3775 & n3776 ;
  buffer buf_n3778( .i (n3777), .o (n3778) );
  assign n3779 = n2825 & n2834 ;
  assign n3780 = n2825 | n2834 ;
  assign n3781 = ~n3779 & n3780 ;
  buffer buf_n3782( .i (n3781), .o (n3782) );
  assign n3783 = N18 & N197 ;
  assign n3784 = n3527 | n3783 ;
  buffer buf_n3785( .i (n3784), .o (n3785) );
  assign n3786 = n2807 | n3785 ;
  assign n3787 = n2807 & n3785 ;
  assign n3788 = n3786 & ~n3787 ;
  buffer buf_n3789( .i (n3788), .o (n3789) );
  assign n3790 = ~n3782 & n3789 ;
  assign n3791 = n3782 & ~n3789 ;
  assign n3792 = n3790 | n3791 ;
  buffer buf_n3793( .i (n3792), .o (n3793) );
  buffer buf_n3794( .i (n3793), .o (n3794) );
  buffer buf_n3795( .i (n3794), .o (n3795) );
  buffer buf_n3796( .i (n3795), .o (n3796) );
  assign n3797 = n3778 | n3796 ;
  assign n3798 = n3778 & n3796 ;
  assign n3799 = n3797 & ~n3798 ;
  assign n3800 = ~n3755 & n3799 ;
  buffer buf_n3801( .i (n3800), .o (n3801) );
  buffer buf_n3802( .i (n3801), .o (n3802) );
  assign n3803 = N18 & N181 ;
  assign n3804 = n3388 | n3803 ;
  buffer buf_n3805( .i (n3804), .o (n3805) );
  assign n3806 = n3040 & ~n3805 ;
  assign n3807 = ~n3040 & n3805 ;
  assign n3808 = n3806 | n3807 ;
  buffer buf_n3809( .i (n3808), .o (n3809) );
  buffer buf_n3810( .i (n3809), .o (n3810) );
  buffer buf_n3811( .i (n3810), .o (n3811) );
  buffer buf_n3812( .i (n3811), .o (n3812) );
  buffer buf_n3813( .i (n3812), .o (n3813) );
  buffer buf_n3814( .i (n3813), .o (n3814) );
  buffer buf_n3101( .i (n3100), .o (n3101) );
  buffer buf_n3102( .i (n3101), .o (n3102) );
  assign n3815 = ~n3093 & n3102 ;
  buffer buf_n3090( .i (n3089), .o (n3090) );
  buffer buf_n3091( .i (n3090), .o (n3091) );
  assign n3816 = n3091 & ~n3104 ;
  assign n3817 = n3815 | n3816 ;
  buffer buf_n3818( .i (n3817), .o (n3818) );
  buffer buf_n3125( .i (n3124), .o (n3125) );
  buffer buf_n3126( .i (n3125), .o (n3126) );
  assign n3819 = n3126 & ~n3143 ;
  buffer buf_n3140( .i (n3139), .o (n3140) );
  buffer buf_n3141( .i (n3140), .o (n3141) );
  assign n3820 = ~n3129 & n3141 ;
  assign n3821 = n3819 | n3820 ;
  buffer buf_n3822( .i (n3821), .o (n3822) );
  assign n3823 = n3818 | n3822 ;
  assign n3824 = n3818 & n3822 ;
  assign n3825 = n3823 & ~n3824 ;
  buffer buf_n3826( .i (n3825), .o (n3826) );
  assign n3827 = ~n3814 & n3826 ;
  assign n3828 = n3814 & ~n3826 ;
  assign n3829 = n3827 | n3828 ;
  buffer buf_n3830( .i (n3829), .o (n3830) );
  assign n3831 = n2979 & n2987 ;
  assign n3832 = n2979 | n2987 ;
  assign n3833 = ~n3831 & n3832 ;
  buffer buf_n3834( .i (n3833), .o (n3834) );
  assign n3835 = n3007 & n3017 ;
  assign n3836 = n3007 | n3017 ;
  assign n3837 = ~n3835 & n3836 ;
  buffer buf_n3838( .i (n3837), .o (n3838) );
  buffer buf_n3839( .i (n3838), .o (n3839) );
  buffer buf_n3840( .i (n3839), .o (n3840) );
  assign n3841 = ~n3834 & n3840 ;
  assign n3842 = n3834 & ~n3840 ;
  assign n3843 = n3841 | n3842 ;
  buffer buf_n3844( .i (n3843), .o (n3844) );
  buffer buf_n3845( .i (n3844), .o (n3845) );
  buffer buf_n3846( .i (n3845), .o (n3846) );
  buffer buf_n3847( .i (n3846), .o (n3847) );
  assign n3848 = ~n3830 & n3847 ;
  assign n3849 = n3830 & ~n3847 ;
  assign n3850 = n3848 | n3849 ;
  assign n3851 = N18 & N208 ;
  assign n3852 = n3492 | n3851 ;
  buffer buf_n3853( .i (n3852), .o (n3853) );
  assign n3854 = N18 & N198 ;
  assign n3855 = n209 | n3854 ;
  buffer buf_n3856( .i (n3855), .o (n3856) );
  assign n3857 = n3853 | n3856 ;
  assign n3858 = n3853 & n3856 ;
  assign n3859 = n3857 & ~n3858 ;
  buffer buf_n3860( .i (n3859), .o (n3860) );
  buffer buf_n3861( .i (n3860), .o (n3861) );
  buffer buf_n3862( .i (n3861), .o (n3862) );
  buffer buf_n3863( .i (n3862), .o (n3863) );
  assign n3864 = n2707 & n2723 ;
  assign n3865 = n2707 | n2723 ;
  assign n3866 = ~n3864 & n3865 ;
  buffer buf_n3867( .i (n3866), .o (n3867) );
  assign n3868 = n2695 & ~n2737 ;
  assign n3869 = ~n2695 & n2737 ;
  assign n3870 = n3868 | n3869 ;
  buffer buf_n3871( .i (n3870), .o (n3871) );
  assign n3872 = n3867 | n3871 ;
  assign n3873 = n3867 & n3871 ;
  assign n3874 = n3872 & ~n3873 ;
  buffer buf_n3875( .i (n3874), .o (n3875) );
  assign n3876 = n3863 | n3875 ;
  assign n3877 = n3863 & n3875 ;
  assign n3878 = n3876 & ~n3877 ;
  buffer buf_n3879( .i (n3878), .o (n3879) );
  assign n3880 = n2775 & ~n2785 ;
  assign n3881 = ~n2775 & n2785 ;
  assign n3882 = n3880 | n3881 ;
  buffer buf_n3883( .i (n3882), .o (n3883) );
  assign n3884 = n2681 & n2758 ;
  assign n3885 = n2681 | n2758 ;
  assign n3886 = ~n3884 & n3885 ;
  buffer buf_n3887( .i (n3886), .o (n3887) );
  assign n3888 = n3883 | n3887 ;
  assign n3889 = n3883 & n3887 ;
  assign n3890 = n3888 & ~n3889 ;
  buffer buf_n3891( .i (n3890), .o (n3891) );
  buffer buf_n3892( .i (n3891), .o (n3892) );
  buffer buf_n3893( .i (n3892), .o (n3893) );
  buffer buf_n3894( .i (n3893), .o (n3894) );
  assign n3895 = n3879 & n3894 ;
  assign n3896 = n3879 | n3894 ;
  assign n3897 = ~n3895 & n3896 ;
  buffer buf_n3898( .i (n3897), .o (n3898) );
  buffer buf_n3899( .i (n3898), .o (n3899) );
  assign n3900 = ~n3850 & n3899 ;
  assign n3901 = n3802 & n3900 ;
  buffer buf_n3902( .i (n3901), .o (n3902) );
  inverter inv_n5032( .i (n3902), .o (n5032) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n2416( .i (n2415), .o (n2416) );
  buffer buf_n2417( .i (n2416), .o (n2417) );
  buffer buf_n2418( .i (n2417), .o (n2418) );
  assign n3903 = ~n1315 & n2418 ;
  buffer buf_n3904( .i (n3903), .o (n3904) );
  assign n3905 = n1315 & ~n2418 ;
  buffer buf_n3906( .i (n3905), .o (n3906) );
  assign n3907 = ~n3904 & ~n3906 ;
  buffer buf_n2433( .i (n2432), .o (n2433) );
  buffer buf_n2434( .i (n2433), .o (n2434) );
  buffer buf_n2435( .i (n2434), .o (n2435) );
  buffer buf_n2436( .i (n2435), .o (n2436) );
  buffer buf_n2437( .i (n2436), .o (n2437) );
  buffer buf_n2438( .i (n2437), .o (n2438) );
  buffer buf_n2482( .i (n2481), .o (n2482) );
  buffer buf_n2483( .i (n2482), .o (n2483) );
  buffer buf_n2484( .i (n2483), .o (n2484) );
  buffer buf_n2485( .i (n2484), .o (n2485) );
  buffer buf_n2486( .i (n2485), .o (n2486) );
  buffer buf_n2487( .i (n2486), .o (n2487) );
  buffer buf_n2488( .i (n2487), .o (n2488) );
  buffer buf_n2489( .i (n2488), .o (n2489) );
  buffer buf_n2490( .i (n2489), .o (n2490) );
  buffer buf_n2491( .i (n2490), .o (n2491) );
  buffer buf_n2492( .i (n2491), .o (n2492) );
  buffer buf_n2493( .i (n2492), .o (n2493) );
  buffer buf_n2494( .i (n2493), .o (n2494) );
  buffer buf_n2495( .i (n2494), .o (n2495) );
  buffer buf_n2496( .i (n2495), .o (n2496) );
  buffer buf_n2497( .i (n2496), .o (n2497) );
  buffer buf_n2498( .i (n2497), .o (n2498) );
  buffer buf_n2499( .i (n2498), .o (n2499) );
  buffer buf_n2500( .i (n2499), .o (n2500) );
  buffer buf_n2501( .i (n2500), .o (n2501) );
  buffer buf_n2502( .i (n2501), .o (n2502) );
  buffer buf_n2503( .i (n2502), .o (n2503) );
  buffer buf_n2504( .i (n2503), .o (n2504) );
  buffer buf_n2505( .i (n2504), .o (n2505) );
  buffer buf_n2506( .i (n2505), .o (n2506) );
  buffer buf_n2507( .i (n2506), .o (n2507) );
  buffer buf_n2508( .i (n2507), .o (n2508) );
  buffer buf_n2509( .i (n2508), .o (n2509) );
  buffer buf_n2510( .i (n2509), .o (n2510) );
  buffer buf_n2511( .i (n2510), .o (n2511) );
  buffer buf_n2512( .i (n2511), .o (n2512) );
  buffer buf_n2513( .i (n2512), .o (n2513) );
  buffer buf_n2514( .i (n2513), .o (n2514) );
  buffer buf_n2515( .i (n2514), .o (n2515) );
  buffer buf_n2516( .i (n2515), .o (n2516) );
  buffer buf_n2517( .i (n2516), .o (n2517) );
  buffer buf_n2518( .i (n2517), .o (n2518) );
  buffer buf_n2519( .i (n2518), .o (n2519) );
  buffer buf_n2520( .i (n2519), .o (n2520) );
  buffer buf_n2521( .i (n2520), .o (n2521) );
  assign n3908 = ~n2438 & n2521 ;
  buffer buf_n3909( .i (n3908), .o (n3909) );
  assign n3910 = n2438 & ~n2521 ;
  buffer buf_n3911( .i (n3910), .o (n3911) );
  assign n3912 = ~n3909 & ~n3911 ;
  assign n3913 = ~n1065 & n1079 ;
  buffer buf_n3914( .i (n3913), .o (n3914) );
  buffer buf_n3915( .i (n3914), .o (n3915) );
  buffer buf_n3916( .i (n3915), .o (n3916) );
  buffer buf_n3917( .i (n3916), .o (n3917) );
  buffer buf_n3918( .i (n3917), .o (n3918) );
  buffer buf_n3919( .i (n3918), .o (n3919) );
  buffer buf_n3920( .i (n3919), .o (n3920) );
  buffer buf_n3921( .i (n3920), .o (n3921) );
  buffer buf_n3922( .i (n3921), .o (n3922) );
  buffer buf_n3923( .i (n3922), .o (n3923) );
  buffer buf_n3924( .i (n3923), .o (n3924) );
  buffer buf_n3925( .i (n3924), .o (n3925) );
  buffer buf_n3926( .i (n3925), .o (n3926) );
  buffer buf_n3927( .i (n3926), .o (n3927) );
  buffer buf_n3928( .i (n3927), .o (n3928) );
  buffer buf_n3929( .i (n3928), .o (n3929) );
  buffer buf_n3930( .i (n3929), .o (n3930) );
  buffer buf_n3931( .i (n3930), .o (n3931) );
  buffer buf_n3932( .i (n3931), .o (n3932) );
  buffer buf_n3933( .i (n3932), .o (n3933) );
  buffer buf_n3934( .i (n3933), .o (n3934) );
  buffer buf_n3935( .i (n3934), .o (n3935) );
  buffer buf_n3936( .i (n3935), .o (n3936) );
  buffer buf_n3937( .i (n3936), .o (n3937) );
  buffer buf_n3938( .i (n3937), .o (n3938) );
  buffer buf_n3939( .i (n3938), .o (n3939) );
  buffer buf_n3940( .i (n3939), .o (n3940) );
  buffer buf_n3941( .i (n3940), .o (n3941) );
  buffer buf_n3942( .i (n3941), .o (n3942) );
  buffer buf_n3943( .i (n3942), .o (n3943) );
  buffer buf_n3944( .i (n3943), .o (n3944) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n1247( .i (n1246), .o (n1247) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  assign n3945 = n1354 | n1414 ;
  buffer buf_n3946( .i (n3945), .o (n3946) );
  buffer buf_n3947( .i (n3946), .o (n3947) );
  buffer buf_n3948( .i (n3947), .o (n3948) );
  buffer buf_n3949( .i (n3948), .o (n3949) );
  buffer buf_n3950( .i (n3949), .o (n3950) );
  buffer buf_n3951( .i (n3950), .o (n3951) );
  buffer buf_n3952( .i (n3951), .o (n3952) );
  buffer buf_n3953( .i (n3952), .o (n3953) );
  buffer buf_n3954( .i (n3953), .o (n3954) );
  buffer buf_n3955( .i (n3954), .o (n3955) );
  buffer buf_n3956( .i (n3955), .o (n3956) );
  buffer buf_n3957( .i (n3956), .o (n3957) );
  buffer buf_n3958( .i (n3957), .o (n3958) );
  buffer buf_n3959( .i (n3958), .o (n3959) );
  buffer buf_n3960( .i (n3959), .o (n3960) );
  buffer buf_n3961( .i (n3960), .o (n3961) );
  buffer buf_n3962( .i (n3961), .o (n3962) );
  buffer buf_n3963( .i (n3962), .o (n3963) );
  buffer buf_n3964( .i (n3963), .o (n3964) );
  buffer buf_n3965( .i (n3964), .o (n3965) );
  buffer buf_n3966( .i (n3965), .o (n3966) );
  buffer buf_n3967( .i (n3966), .o (n3967) );
  buffer buf_n3968( .i (n3967), .o (n3968) );
  buffer buf_n3969( .i (n3968), .o (n3969) );
  assign n3970 = n2414 & ~n3969 ;
  buffer buf_n3971( .i (n3970), .o (n3971) );
  assign n3972 = ~n1408 & n3971 ;
  assign n3973 = n1262 | n3972 ;
  buffer buf_n3974( .i (n3973), .o (n3974) );
  assign n3975 = n3944 & ~n3974 ;
  assign n3976 = ~n3944 & n3974 ;
  assign n3977 = n3975 | n3976 ;
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  assign n3978 = n1238 | n3971 ;
  buffer buf_n3979( .i (n3978), .o (n3979) );
  assign n3980 = n1410 | n3979 ;
  assign n3981 = n1410 & n3979 ;
  assign n3982 = ~n3980 | n3981 ;
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  assign n3983 = ~n1379 & n2414 ;
  assign n3984 = n1211 | n3983 ;
  buffer buf_n3985( .i (n3984), .o (n3985) );
  assign n3986 = n1442 & n3985 ;
  assign n3987 = n1442 | n3985 ;
  assign n3988 = n3986 | ~n3987 ;
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  assign n3989 = n1179 | n3904 ;
  buffer buf_n3990( .i (n3989), .o (n3990) );
  assign n3991 = n1352 | n3990 ;
  assign n3992 = n1352 & n3990 ;
  assign n3993 = ~n3991 | n3992 ;
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  assign n3994 = n609 | n649 ;
  assign n3995 = n446 & n3994 ;
  buffer buf_n3996( .i (n3995), .o (n3996) );
  buffer buf_n3997( .i (n3996), .o (n3997) );
  buffer buf_n3998( .i (n3997), .o (n3998) );
  buffer buf_n3999( .i (n3998), .o (n3999) );
  buffer buf_n4000( .i (n3999), .o (n4000) );
  buffer buf_n4001( .i (n4000), .o (n4001) );
  buffer buf_n4002( .i (n4001), .o (n4002) );
  buffer buf_n4003( .i (n4002), .o (n4003) );
  buffer buf_n4004( .i (n4003), .o (n4004) );
  buffer buf_n4005( .i (n4004), .o (n4005) );
  buffer buf_n4006( .i (n4005), .o (n4006) );
  buffer buf_n4007( .i (n4006), .o (n4007) );
  buffer buf_n4008( .i (n4007), .o (n4008) );
  buffer buf_n4009( .i (n4008), .o (n4009) );
  buffer buf_n4010( .i (n4009), .o (n4010) );
  buffer buf_n4011( .i (n4010), .o (n4011) );
  buffer buf_n4012( .i (n4011), .o (n4012) );
  buffer buf_n4013( .i (n4012), .o (n4013) );
  buffer buf_n4014( .i (n4013), .o (n4014) );
  buffer buf_n4015( .i (n4014), .o (n4015) );
  buffer buf_n4016( .i (n4015), .o (n4016) );
  buffer buf_n4017( .i (n4016), .o (n4017) );
  buffer buf_n4018( .i (n4017), .o (n4018) );
  buffer buf_n4019( .i (n4018), .o (n4019) );
  buffer buf_n4020( .i (n4019), .o (n4020) );
  buffer buf_n4021( .i (n4020), .o (n4021) );
  buffer buf_n4022( .i (n4021), .o (n4022) );
  buffer buf_n4023( .i (n4022), .o (n4023) );
  buffer buf_n4024( .i (n4023), .o (n4024) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  assign n4025 = n687 & n2635 ;
  assign n4026 = n4024 & ~n4025 ;
  buffer buf_n4027( .i (n4026), .o (n4027) );
  assign n4028 = n730 & n4027 ;
  assign n4029 = n730 | n4027 ;
  assign n4030 = n4028 | ~n4029 ;
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n639( .i (n638), .o (n639) );
  assign n4031 = n639 & ~n2635 ;
  buffer buf_n4032( .i (n4031), .o (n4032) );
  assign n4033 = n689 | n4032 ;
  assign n4034 = n689 & n4032 ;
  assign n4035 = ~n4033 | n4034 ;
  buffer buf_n2443( .i (n2442), .o (n2443) );
  buffer buf_n2444( .i (n2443), .o (n2444) );
  buffer buf_n2445( .i (n2444), .o (n2445) );
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n2448( .i (n2447), .o (n2448) );
  buffer buf_n2449( .i (n2448), .o (n2449) );
  buffer buf_n2450( .i (n2449), .o (n2450) );
  buffer buf_n2451( .i (n2450), .o (n2451) );
  buffer buf_n2452( .i (n2451), .o (n2452) );
  buffer buf_n2453( .i (n2452), .o (n2453) );
  buffer buf_n2454( .i (n2453), .o (n2454) );
  buffer buf_n2455( .i (n2454), .o (n2455) );
  buffer buf_n2456( .i (n2455), .o (n2456) );
  buffer buf_n2457( .i (n2456), .o (n2457) );
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n2460( .i (n2459), .o (n2460) );
  buffer buf_n2461( .i (n2460), .o (n2461) );
  buffer buf_n2462( .i (n2461), .o (n2462) );
  buffer buf_n2463( .i (n2462), .o (n2463) );
  buffer buf_n2464( .i (n2463), .o (n2464) );
  buffer buf_n2465( .i (n2464), .o (n2465) );
  buffer buf_n2466( .i (n2465), .o (n2466) );
  buffer buf_n2467( .i (n2466), .o (n2467) );
  buffer buf_n2468( .i (n2467), .o (n2468) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  buffer buf_n2470( .i (n2469), .o (n2470) );
  buffer buf_n2471( .i (n2470), .o (n2471) );
  buffer buf_n2472( .i (n2471), .o (n2472) );
  buffer buf_n2473( .i (n2472), .o (n2473) );
  buffer buf_n2474( .i (n2473), .o (n2474) );
  buffer buf_n2475( .i (n2474), .o (n2475) );
  buffer buf_n2476( .i (n2475), .o (n2476) );
  buffer buf_n2477( .i (n2476), .o (n2477) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n2570( .i (n2569), .o (n2570) );
  buffer buf_n2571( .i (n2570), .o (n2571) );
  buffer buf_n2572( .i (n2571), .o (n2572) );
  buffer buf_n2573( .i (n2572), .o (n2573) );
  buffer buf_n2574( .i (n2573), .o (n2574) );
  buffer buf_n2575( .i (n2574), .o (n2575) );
  buffer buf_n2576( .i (n2575), .o (n2576) );
  buffer buf_n2577( .i (n2576), .o (n2577) );
  buffer buf_n2578( .i (n2577), .o (n2578) );
  buffer buf_n2579( .i (n2578), .o (n2579) );
  buffer buf_n2580( .i (n2579), .o (n2580) );
  buffer buf_n2581( .i (n2580), .o (n2581) );
  buffer buf_n2582( .i (n2581), .o (n2582) );
  buffer buf_n2583( .i (n2582), .o (n2583) );
  buffer buf_n2584( .i (n2583), .o (n2584) );
  buffer buf_n2585( .i (n2584), .o (n2585) );
  buffer buf_n2586( .i (n2585), .o (n2586) );
  buffer buf_n2587( .i (n2586), .o (n2587) );
  buffer buf_n2588( .i (n2587), .o (n2588) );
  buffer buf_n2589( .i (n2588), .o (n2589) );
  buffer buf_n2590( .i (n2589), .o (n2590) );
  buffer buf_n2591( .i (n2590), .o (n2591) );
  buffer buf_n2592( .i (n2591), .o (n2592) );
  buffer buf_n2593( .i (n2592), .o (n2593) );
  buffer buf_n2594( .i (n2593), .o (n2594) );
  buffer buf_n2595( .i (n2594), .o (n2595) );
  buffer buf_n2596( .i (n2595), .o (n2596) );
  buffer buf_n2597( .i (n2596), .o (n2597) );
  buffer buf_n2598( .i (n2597), .o (n2598) );
  buffer buf_n2599( .i (n2598), .o (n2599) );
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  assign n4036 = ~n2432 & n2601 ;
  assign n4037 = n605 & ~n4036 ;
  buffer buf_n4038( .i (n4037), .o (n4038) );
  assign n4039 = n2477 | n4038 ;
  assign n4040 = n2477 & n4038 ;
  assign n4041 = ~n4039 | n4040 ;
  buffer buf_n2524( .i (n2523), .o (n2524) );
  buffer buf_n2525( .i (n2524), .o (n2525) );
  buffer buf_n2526( .i (n2525), .o (n2526) );
  buffer buf_n2527( .i (n2526), .o (n2527) );
  buffer buf_n2528( .i (n2527), .o (n2528) );
  buffer buf_n2529( .i (n2528), .o (n2529) );
  buffer buf_n2530( .i (n2529), .o (n2530) );
  buffer buf_n2531( .i (n2530), .o (n2531) );
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n2532), .o (n2533) );
  buffer buf_n2534( .i (n2533), .o (n2534) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  buffer buf_n2536( .i (n2535), .o (n2536) );
  buffer buf_n2537( .i (n2536), .o (n2537) );
  buffer buf_n2538( .i (n2537), .o (n2538) );
  buffer buf_n2539( .i (n2538), .o (n2539) );
  buffer buf_n2540( .i (n2539), .o (n2540) );
  buffer buf_n2541( .i (n2540), .o (n2541) );
  buffer buf_n2542( .i (n2541), .o (n2542) );
  buffer buf_n2543( .i (n2542), .o (n2543) );
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  buffer buf_n2551( .i (n2550), .o (n2551) );
  buffer buf_n2552( .i (n2551), .o (n2552) );
  buffer buf_n2553( .i (n2552), .o (n2553) );
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2555( .i (n2554), .o (n2555) );
  buffer buf_n2556( .i (n2555), .o (n2556) );
  buffer buf_n2557( .i (n2556), .o (n2557) );
  buffer buf_n2558( .i (n2557), .o (n2558) );
  buffer buf_n2559( .i (n2558), .o (n2559) );
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  buffer buf_n2563( .i (n2562), .o (n2563) );
  buffer buf_n2564( .i (n2563), .o (n2564) );
  buffer buf_n2565( .i (n2564), .o (n2565) );
  buffer buf_n2566( .i (n2565), .o (n2566) );
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  assign n4042 = n566 & ~n3909 ;
  buffer buf_n4043( .i (n4042), .o (n4043) );
  assign n4044 = ~n2567 & n4043 ;
  assign n4045 = n2567 & ~n4043 ;
  assign n4046 = ~n4044 & ~n4045 ;
  assign n4047 = N150 & N184 ;
  assign n4048 = N228 & N240 ;
  assign n4049 = n4047 & n4048 ;
  buffer buf_n4050( .i (n4049), .o (n4050) );
  assign n4051 = N152 & N210 ;
  assign n4052 = N218 & N230 ;
  assign n4053 = n4051 & n4052 ;
  buffer buf_n4054( .i (n4053), .o (n4054) );
  assign n4055 = n4050 & n4054 ;
  assign n4056 = N182 & N183 ;
  assign n4057 = N185 & N186 ;
  assign n4058 = n4056 & n4057 ;
  buffer buf_n4059( .i (n4058), .o (n4059) );
  assign n4060 = N162 & N172 ;
  assign n4061 = N188 & N199 ;
  assign n4062 = n4060 & n4061 ;
  buffer buf_n4063( .i (n4062), .o (n4063) );
  assign n4064 = n4059 & n4063 ;
  assign n4065 = n4055 & n4064 ;
  assign n4066 = n3560 & n4065 ;
  buffer buf_n3726( .i (n3725), .o (n3726) );
  buffer buf_n3727( .i (n3726), .o (n3727) );
  buffer buf_n3728( .i (n3727), .o (n3728) );
  assign n4067 = n3728 & n3902 ;
  assign n4068 = ~n4066 | ~n4067 ;
  assign n4069 = ~n743 & n778 ;
  buffer buf_n4070( .i (n4069), .o (n4070) );
  buffer buf_n4071( .i (n4070), .o (n4071) );
  buffer buf_n4072( .i (n4071), .o (n4072) );
  buffer buf_n4073( .i (n4072), .o (n4073) );
  buffer buf_n4074( .i (n4073), .o (n4074) );
  buffer buf_n4075( .i (n4074), .o (n4075) );
  buffer buf_n4076( .i (n4075), .o (n4076) );
  buffer buf_n4077( .i (n4076), .o (n4077) );
  buffer buf_n4078( .i (n4077), .o (n4078) );
  buffer buf_n4079( .i (n4078), .o (n4079) );
  buffer buf_n4080( .i (n4079), .o (n4080) );
  buffer buf_n4081( .i (n4080), .o (n4081) );
  buffer buf_n4082( .i (n4081), .o (n4082) );
  buffer buf_n4083( .i (n4082), .o (n4083) );
  buffer buf_n4084( .i (n4083), .o (n4084) );
  buffer buf_n4085( .i (n4084), .o (n4085) );
  buffer buf_n4086( .i (n4085), .o (n4086) );
  buffer buf_n4087( .i (n4086), .o (n4087) );
  buffer buf_n4088( .i (n4087), .o (n4088) );
  buffer buf_n4089( .i (n4088), .o (n4089) );
  buffer buf_n4090( .i (n4089), .o (n4090) );
  buffer buf_n4091( .i (n4090), .o (n4091) );
  buffer buf_n4092( .i (n4091), .o (n4092) );
  buffer buf_n4093( .i (n4092), .o (n4093) );
  buffer buf_n4094( .i (n4093), .o (n4094) );
  buffer buf_n4095( .i (n4094), .o (n4095) );
  buffer buf_n4096( .i (n4095), .o (n4096) );
  buffer buf_n4097( .i (n4096), .o (n4097) );
  buffer buf_n4098( .i (n4097), .o (n4098) );
  buffer buf_n4099( .i (n4098), .o (n4099) );
  buffer buf_n4100( .i (n4099), .o (n4100) );
  assign n4101 = n2429 | n4100 ;
  assign n4102 = n2429 & n4100 ;
  assign n4103 = ~n4101 | n4102 ;
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  assign n4104 = n1001 & ~n2421 ;
  assign n4105 = n914 & ~n4104 ;
  buffer buf_n4106( .i (n4105), .o (n4106) );
  assign n4107 = n1033 & n4106 ;
  assign n4108 = n1033 | n4106 ;
  assign n4109 = n4107 | ~n4108 ;
  assign n4110 = ~n836 & n840 ;
  buffer buf_n4111( .i (n4110), .o (n4111) );
  buffer buf_n4112( .i (n4111), .o (n4112) );
  buffer buf_n4113( .i (n4112), .o (n4113) );
  buffer buf_n4114( .i (n4113), .o (n4114) );
  buffer buf_n4115( .i (n4114), .o (n4115) );
  buffer buf_n4116( .i (n4115), .o (n4116) );
  buffer buf_n4117( .i (n4116), .o (n4117) );
  buffer buf_n4118( .i (n4117), .o (n4118) );
  buffer buf_n4119( .i (n4118), .o (n4119) );
  buffer buf_n4120( .i (n4119), .o (n4120) );
  buffer buf_n4121( .i (n4120), .o (n4121) );
  buffer buf_n4122( .i (n4121), .o (n4122) );
  buffer buf_n4123( .i (n4122), .o (n4123) );
  buffer buf_n4124( .i (n4123), .o (n4124) );
  buffer buf_n4125( .i (n4124), .o (n4125) );
  buffer buf_n4126( .i (n4125), .o (n4126) );
  buffer buf_n4127( .i (n4126), .o (n4127) );
  buffer buf_n4128( .i (n4127), .o (n4128) );
  buffer buf_n4129( .i (n4128), .o (n4129) );
  buffer buf_n4130( .i (n4129), .o (n4130) );
  buffer buf_n4131( .i (n4130), .o (n4131) );
  buffer buf_n4132( .i (n4131), .o (n4132) );
  buffer buf_n4133( .i (n4132), .o (n4133) );
  buffer buf_n4134( .i (n4133), .o (n4134) );
  buffer buf_n4135( .i (n4134), .o (n4135) );
  buffer buf_n4136( .i (n4135), .o (n4136) );
  buffer buf_n4137( .i (n4136), .o (n4137) );
  buffer buf_n4138( .i (n4137), .o (n4138) );
  buffer buf_n4139( .i (n4138), .o (n4139) );
  buffer buf_n4140( .i (n4139), .o (n4140) );
  buffer buf_n4141( .i (n4140), .o (n4141) );
  buffer buf_n4142( .i (n4141), .o (n4142) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  assign n4143 = n972 | n2421 ;
  assign n4144 = n882 & n4143 ;
  buffer buf_n4145( .i (n4144), .o (n4145) );
  assign n4146 = n4142 & ~n4145 ;
  assign n4147 = ~n4142 & n4145 ;
  assign n4148 = ~n4146 & ~n4147 ;
  buffer buf_n2422( .i (n2421), .o (n2422) );
  buffer buf_n2423( .i (n2422), .o (n2423) );
  buffer buf_n2424( .i (n2423), .o (n2424) );
  buffer buf_n2425( .i (n2424), .o (n2425) );
  buffer buf_n2426( .i (n2425), .o (n2426) );
  assign n4149 = n853 & ~n944 ;
  buffer buf_n4150( .i (n4149), .o (n4150) );
  buffer buf_n4151( .i (n4150), .o (n4151) );
  buffer buf_n4152( .i (n4151), .o (n4152) );
  buffer buf_n4153( .i (n4152), .o (n4153) );
  buffer buf_n4154( .i (n4153), .o (n4154) );
  buffer buf_n4155( .i (n4154), .o (n4155) );
  buffer buf_n4156( .i (n4155), .o (n4156) );
  buffer buf_n4157( .i (n4156), .o (n4157) );
  buffer buf_n4158( .i (n4157), .o (n4158) );
  buffer buf_n4159( .i (n4158), .o (n4159) );
  buffer buf_n4160( .i (n4159), .o (n4160) );
  buffer buf_n4161( .i (n4160), .o (n4161) );
  buffer buf_n4162( .i (n4161), .o (n4162) );
  buffer buf_n4163( .i (n4162), .o (n4163) );
  buffer buf_n4164( .i (n4163), .o (n4164) );
  buffer buf_n4165( .i (n4164), .o (n4165) );
  buffer buf_n4166( .i (n4165), .o (n4166) );
  buffer buf_n4167( .i (n4166), .o (n4167) );
  buffer buf_n4168( .i (n4167), .o (n4168) );
  buffer buf_n4169( .i (n4168), .o (n4169) );
  buffer buf_n4170( .i (n4169), .o (n4170) );
  buffer buf_n4171( .i (n4170), .o (n4171) );
  buffer buf_n4172( .i (n4171), .o (n4172) );
  buffer buf_n4173( .i (n4172), .o (n4173) );
  buffer buf_n4174( .i (n4173), .o (n4174) );
  buffer buf_n4175( .i (n4174), .o (n4175) );
  buffer buf_n4176( .i (n4175), .o (n4176) );
  buffer buf_n4177( .i (n4176), .o (n4177) );
  buffer buf_n4178( .i (n4177), .o (n4178) );
  buffer buf_n4179( .i (n4178), .o (n4179) );
  buffer buf_n4180( .i (n4179), .o (n4180) );
  buffer buf_n4181( .i (n4180), .o (n4181) );
  assign n4182 = ~n2426 & n4181 ;
  assign n4183 = n2426 & ~n4181 ;
  assign n4184 = ~n4182 & ~n4183 ;
  buffer buf_n2348( .i (n2347), .o (n2348) );
  buffer buf_n2349( .i (n2348), .o (n2349) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n1811( .i (n1810), .o (n1811) );
  assign n4185 = n1775 | n1811 ;
  buffer buf_n4186( .i (n4185), .o (n4186) );
  assign n4187 = n2349 & ~n4186 ;
  buffer buf_n4188( .i (n4187), .o (n4188) );
  assign n4189 = ~n2349 & n4186 ;
  buffer buf_n4190( .i (n4189), .o (n4190) );
  assign n4191 = ~n4188 & ~n4190 ;
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  assign n4192 = n407 & n2645 ;
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  assign n4193 = n412 | n2645 ;
  assign n4194 = ~n4192 & n4193 ;
  buffer buf_n4195( .i (n4194), .o (n4195) );
  assign n4196 = n290 & n4195 ;
  assign n4197 = n290 | n4195 ;
  assign n4198 = ~n4196 & n4197 ;
  buffer buf_n4199( .i (n4198), .o (n4199) );
  assign n4200 = n414 & n2645 ;
  buffer buf_n4201( .i (n4200), .o (n4201) );
  assign n4202 = n2647 & ~n4201 ;
  buffer buf_n4203( .i (n4202), .o (n4203) );
  buffer buf_n1918( .i (n1917), .o (n1918) );
  buffer buf_n1919( .i (n1918), .o (n1919) );
  buffer buf_n1920( .i (n1919), .o (n1920) );
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  assign n4204 = ~n1928 & n2347 ;
  buffer buf_n1969( .i (n1968), .o (n1969) );
  buffer buf_n1970( .i (n1969), .o (n1970) );
  buffer buf_n1971( .i (n1970), .o (n1971) );
  assign n4205 = ~n1971 & n2393 ;
  assign n4206 = n1971 & ~n2393 ;
  assign n4207 = n4205 | n4206 ;
  buffer buf_n4208( .i (n4207), .o (n4208) );
  buffer buf_n4209( .i (n4208), .o (n4209) );
  buffer buf_n4210( .i (n4209), .o (n4210) );
  buffer buf_n4211( .i (n4210), .o (n4211) );
  buffer buf_n4212( .i (n4211), .o (n4212) );
  buffer buf_n4213( .i (n4212), .o (n4213) );
  buffer buf_n4214( .i (n4213), .o (n4214) );
  assign n4215 = ~n4204 & n4214 ;
  assign n4216 = ~n2351 & ~n4215 ;
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n2379( .i (n2378), .o (n2379) );
  buffer buf_n2380( .i (n2379), .o (n2380) );
  buffer buf_n2381( .i (n2380), .o (n2381) );
  buffer buf_n2382( .i (n2381), .o (n2382) );
  buffer buf_n2383( .i (n2382), .o (n2383) );
  buffer buf_n2384( .i (n2383), .o (n2384) );
  buffer buf_n2385( .i (n2384), .o (n2385) );
  buffer buf_n2386( .i (n2385), .o (n2386) );
  buffer buf_n2387( .i (n2386), .o (n2387) );
  buffer buf_n2388( .i (n2387), .o (n2388) );
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  assign n4217 = n1820 | n1893 ;
  buffer buf_n4218( .i (n4217), .o (n4218) );
  buffer buf_n4219( .i (n4218), .o (n4219) );
  buffer buf_n4220( .i (n4219), .o (n4220) );
  buffer buf_n4221( .i (n4220), .o (n4221) );
  buffer buf_n4222( .i (n4221), .o (n4222) );
  buffer buf_n4223( .i (n4222), .o (n4223) );
  buffer buf_n4224( .i (n4223), .o (n4224) );
  buffer buf_n4225( .i (n4224), .o (n4225) );
  buffer buf_n4226( .i (n4225), .o (n4226) );
  buffer buf_n4227( .i (n4226), .o (n4227) );
  buffer buf_n4228( .i (n4227), .o (n4228) );
  buffer buf_n4229( .i (n4228), .o (n4229) );
  assign n4230 = n2347 & ~n4229 ;
  assign n4231 = n2390 | n4230 ;
  buffer buf_n4232( .i (n4231), .o (n4232) );
  assign n4233 = n1868 | n4232 ;
  assign n4234 = n1868 & n4232 ;
  assign n4235 = ~n4233 | n4234 ;
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1907( .i (n1906), .o (n1907) );
  buffer buf_n1908( .i (n1907), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n2355( .i (n2354), .o (n2355) );
  buffer buf_n2356( .i (n2355), .o (n2356) );
  buffer buf_n2357( .i (n2356), .o (n2357) );
  buffer buf_n2358( .i (n2357), .o (n2358) );
  buffer buf_n2359( .i (n2358), .o (n2359) );
  buffer buf_n2360( .i (n2359), .o (n2360) );
  buffer buf_n2361( .i (n2360), .o (n2361) );
  buffer buf_n2362( .i (n2361), .o (n2362) );
  buffer buf_n2363( .i (n2362), .o (n2363) );
  buffer buf_n2364( .i (n2363), .o (n2364) );
  buffer buf_n2365( .i (n2364), .o (n2365) );
  buffer buf_n2366( .i (n2365), .o (n2366) );
  buffer buf_n2367( .i (n2366), .o (n2367) );
  buffer buf_n2368( .i (n2367), .o (n2368) );
  buffer buf_n2369( .i (n2368), .o (n2369) );
  buffer buf_n2370( .i (n2369), .o (n2370) );
  buffer buf_n2371( .i (n2370), .o (n2371) );
  buffer buf_n2372( .i (n2371), .o (n2372) );
  buffer buf_n2373( .i (n2372), .o (n2373) );
  buffer buf_n2374( .i (n2373), .o (n2374) );
  assign n4236 = n1786 | n1813 ;
  buffer buf_n4237( .i (n4236), .o (n4237) );
  buffer buf_n4238( .i (n4237), .o (n4238) );
  buffer buf_n4239( .i (n4238), .o (n4239) );
  buffer buf_n4240( .i (n4239), .o (n4240) );
  buffer buf_n4241( .i (n4240), .o (n4241) );
  buffer buf_n4242( .i (n4241), .o (n4242) );
  buffer buf_n4243( .i (n4242), .o (n4243) );
  buffer buf_n4244( .i (n4243), .o (n4244) );
  buffer buf_n4245( .i (n4244), .o (n4245) );
  buffer buf_n4246( .i (n4245), .o (n4246) );
  buffer buf_n4247( .i (n4246), .o (n4247) );
  buffer buf_n4248( .i (n4247), .o (n4248) );
  buffer buf_n4249( .i (n4248), .o (n4249) );
  buffer buf_n4250( .i (n4249), .o (n4250) );
  buffer buf_n4251( .i (n4250), .o (n4251) );
  buffer buf_n4252( .i (n4251), .o (n4252) );
  buffer buf_n4253( .i (n4252), .o (n4253) );
  buffer buf_n4254( .i (n4253), .o (n4254) );
  buffer buf_n4255( .i (n4254), .o (n4255) );
  buffer buf_n4256( .i (n4255), .o (n4256) );
  buffer buf_n4257( .i (n4256), .o (n4257) );
  buffer buf_n4258( .i (n4257), .o (n4258) );
  assign n4261 = n4188 & ~n4258 ;
  assign n4262 = n2374 | n4261 ;
  buffer buf_n4263( .i (n4262), .o (n4263) );
  assign n4264 = n1913 & n4263 ;
  assign n4265 = n1913 | n4263 ;
  assign n4266 = n4264 | ~n4265 ;
  buffer buf_n4259( .i (n4258), .o (n4259) );
  buffer buf_n4260( .i (n4259), .o (n4260) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  assign n4267 = n1779 | n4188 ;
  buffer buf_n4268( .i (n4267), .o (n4268) );
  assign n4269 = n4260 | n4268 ;
  assign n4270 = n4260 & n4268 ;
  assign n4271 = ~n4269 | n4270 ;
  assign n4272 = n1476 | n1505 ;
  buffer buf_n4273( .i (n4272), .o (n4273) );
  buffer buf_n4274( .i (n4273), .o (n4274) );
  buffer buf_n4275( .i (n4274), .o (n4275) );
  buffer buf_n4276( .i (n4275), .o (n4276) );
  buffer buf_n4277( .i (n4276), .o (n4277) );
  buffer buf_n4278( .i (n4277), .o (n4278) );
  buffer buf_n4279( .i (n4278), .o (n4279) );
  buffer buf_n4280( .i (n4279), .o (n4280) );
  buffer buf_n4281( .i (n4280), .o (n4281) );
  buffer buf_n4282( .i (n4281), .o (n4282) );
  buffer buf_n4283( .i (n4282), .o (n4283) );
  buffer buf_n4284( .i (n4283), .o (n4284) );
  buffer buf_n4285( .i (n4284), .o (n4285) );
  buffer buf_n4286( .i (n4285), .o (n4286) );
  buffer buf_n4287( .i (n4286), .o (n4287) );
  buffer buf_n4288( .i (n4287), .o (n4288) );
  buffer buf_n4289( .i (n4288), .o (n4289) );
  buffer buf_n4290( .i (n4289), .o (n4290) );
  buffer buf_n4291( .i (n4290), .o (n4291) );
  buffer buf_n4292( .i (n4291), .o (n4292) );
  buffer buf_n4293( .i (n4292), .o (n4293) );
  buffer buf_n4294( .i (n4293), .o (n4294) );
  buffer buf_n4295( .i (n4294), .o (n4295) );
  buffer buf_n4296( .i (n4295), .o (n4296) );
  buffer buf_n4297( .i (n4296), .o (n4297) );
  assign n4298 = ~n2411 & n4297 ;
  assign n4299 = n2411 & ~n4297 ;
  assign n4300 = ~n4298 & ~n4299 ;
  assign n4301 = n1538 | n1546 ;
  buffer buf_n4302( .i (n4301), .o (n4302) );
  buffer buf_n4303( .i (n4302), .o (n4303) );
  buffer buf_n4304( .i (n4303), .o (n4304) );
  buffer buf_n4305( .i (n4304), .o (n4305) );
  buffer buf_n4306( .i (n4305), .o (n4306) );
  buffer buf_n4307( .i (n4306), .o (n4307) );
  buffer buf_n4308( .i (n4307), .o (n4308) );
  buffer buf_n4309( .i (n4308), .o (n4309) );
  buffer buf_n4310( .i (n4309), .o (n4310) );
  buffer buf_n4311( .i (n4310), .o (n4311) );
  buffer buf_n4312( .i (n4311), .o (n4312) );
  buffer buf_n4313( .i (n4312), .o (n4313) );
  buffer buf_n4314( .i (n4313), .o (n4314) );
  buffer buf_n4315( .i (n4314), .o (n4315) );
  buffer buf_n4316( .i (n4315), .o (n4316) );
  buffer buf_n4317( .i (n4316), .o (n4317) );
  buffer buf_n4318( .i (n4317), .o (n4318) );
  buffer buf_n4319( .i (n4318), .o (n4319) );
  buffer buf_n4320( .i (n4319), .o (n4320) );
  buffer buf_n4321( .i (n4320), .o (n4321) );
  buffer buf_n4322( .i (n4321), .o (n4322) );
  buffer buf_n4323( .i (n4322), .o (n4323) );
  buffer buf_n4324( .i (n4323), .o (n4324) );
  buffer buf_n4325( .i (n4324), .o (n4325) );
  buffer buf_n4326( .i (n4325), .o (n4326) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  assign n4327 = ~n1731 & n2405 ;
  assign n4328 = n1617 | n4327 ;
  buffer buf_n4329( .i (n4328), .o (n4329) );
  assign n4330 = n4326 | n4329 ;
  assign n4331 = n4326 & n4329 ;
  assign n4332 = ~n4330 | n4331 ;
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  buffer buf_n1658( .i (n1657), .o (n1658) );
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  assign n4333 = n1593 | n2405 ;
  assign n4334 = ~n1688 & n4333 ;
  buffer buf_n4335( .i (n4334), .o (n4335) );
  assign n4336 = n1662 & ~n4335 ;
  assign n4337 = ~n1662 & n4335 ;
  assign n4338 = ~n4336 & ~n4337 ;
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n2406( .i (n2405), .o (n2406) );
  buffer buf_n2407( .i (n2406), .o (n2407) );
  buffer buf_n2408( .i (n2407), .o (n2408) );
  assign n4339 = ~n1712 & n2408 ;
  assign n4340 = n1712 & ~n2408 ;
  assign n4341 = ~n4339 & ~n4340 ;
  assign n4342 = N242 & ~N5 ;
  inverter inv_n4343( .i (n4342), .o (n4343) );
  assign n4344 = N134 & ~N5 ;
  assign n4345 = N133 & n4344 ;
  inverter inv_n4346( .i (n4345), .o (n4346) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  assign n4347 = n1284 & n1317 ;
  buffer buf_n4348( .i (n4347), .o (n4348) );
  assign n4349 = n1354 & ~n4348 ;
  buffer buf_n4350( .i (n4349), .o (n4350) );
  buffer buf_n4351( .i (n4350), .o (n4351) );
  buffer buf_n4352( .i (n4351), .o (n4352) );
  buffer buf_n4353( .i (n4352), .o (n4353) );
  buffer buf_n4354( .i (n4353), .o (n4354) );
  buffer buf_n4355( .i (n4354), .o (n4355) );
  assign n4356 = n1241 & n4355 ;
  assign n4357 = n1241 | n4355 ;
  assign n4358 = ~n4356 & n4357 ;
  buffer buf_n4359( .i (n4358), .o (n4359) );
  assign n4360 = n1452 & ~n4359 ;
  buffer buf_n4361( .i (n4360), .o (n4361) );
  assign n4362 = ~n1215 & n3948 ;
  buffer buf_n4363( .i (n4362), .o (n4363) );
  assign n4364 = ~n1135 & n1282 ;
  assign n4365 = n1181 | n1282 ;
  assign n4366 = ~n4364 & n4365 ;
  buffer buf_n4367( .i (n4366), .o (n4367) );
  buffer buf_n4368( .i (n4367), .o (n4368) );
  buffer buf_n4369( .i (n4368), .o (n4369) );
  assign n4370 = n3915 & ~n4369 ;
  assign n4371 = ~n3915 & n4369 ;
  assign n4372 = n4370 | n4371 ;
  buffer buf_n4373( .i (n4372), .o (n4373) );
  buffer buf_n4374( .i (n4373), .o (n4374) );
  buffer buf_n4375( .i (n4374), .o (n4375) );
  assign n4376 = n4363 & ~n4375 ;
  assign n4377 = ~n4363 & n4375 ;
  assign n4378 = n4376 | n4377 ;
  buffer buf_n4379( .i (n4378), .o (n4379) );
  buffer buf_n4380( .i (n4379), .o (n4380) );
  buffer buf_n4381( .i (n4380), .o (n4381) );
  buffer buf_n4382( .i (n4381), .o (n4382) );
  assign n4383 = n4361 | n4382 ;
  assign n4384 = n4361 & n4382 ;
  assign n4385 = n4383 & ~n4384 ;
  buffer buf_n4386( .i (n4385), .o (n4386) );
  buffer buf_n4387( .i (n4386), .o (n4387) );
  buffer buf_n4388( .i (n4387), .o (n4388) );
  buffer buf_n4389( .i (n4388), .o (n4389) );
  buffer buf_n4390( .i (n4389), .o (n4390) );
  buffer buf_n4391( .i (n4390), .o (n4391) );
  buffer buf_n4392( .i (n4391), .o (n4392) );
  buffer buf_n4393( .i (n4392), .o (n4393) );
  buffer buf_n4394( .i (n4393), .o (n4394) );
  buffer buf_n4395( .i (n4394), .o (n4395) );
  buffer buf_n4396( .i (n4395), .o (n4396) );
  buffer buf_n4397( .i (n4396), .o (n4397) );
  buffer buf_n4398( .i (n4397), .o (n4398) );
  buffer buf_n4399( .i (n4398), .o (n4399) );
  buffer buf_n4400( .i (n4399), .o (n4400) );
  assign n4401 = n2418 & ~n4400 ;
  assign n4402 = n1135 | n1144 ;
  buffer buf_n4403( .i (n4402), .o (n4403) );
  assign n4404 = ~n1183 & n4403 ;
  buffer buf_n4405( .i (n4404), .o (n4405) );
  buffer buf_n4406( .i (n4405), .o (n4406) );
  assign n4407 = n3915 & n4406 ;
  buffer buf_n4408( .i (n3914), .o (n4408) );
  assign n4409 = n4406 | n4408 ;
  assign n4410 = ~n4407 & n4409 ;
  buffer buf_n4411( .i (n4410), .o (n4411) );
  assign n4412 = n1215 | n4411 ;
  buffer buf_n4413( .i (n1214), .o (n4413) );
  assign n4414 = n4411 & n4413 ;
  assign n4415 = n4412 & ~n4414 ;
  buffer buf_n4416( .i (n4415), .o (n4416) );
  buffer buf_n4417( .i (n4416), .o (n4417) );
  buffer buf_n4418( .i (n4417), .o (n4418) );
  buffer buf_n4419( .i (n4418), .o (n4419) );
  assign n4420 = n4359 & n4419 ;
  assign n4421 = n4359 | n4419 ;
  assign n4422 = ~n4420 & n4421 ;
  buffer buf_n4423( .i (n4422), .o (n4423) );
  buffer buf_n4424( .i (n4423), .o (n4424) );
  buffer buf_n4425( .i (n4424), .o (n4425) );
  buffer buf_n4426( .i (n4425), .o (n4426) );
  buffer buf_n4427( .i (n4426), .o (n4427) );
  buffer buf_n4428( .i (n4427), .o (n4428) );
  buffer buf_n4429( .i (n4428), .o (n4429) );
  buffer buf_n4430( .i (n4429), .o (n4430) );
  buffer buf_n4431( .i (n4430), .o (n4431) );
  buffer buf_n4432( .i (n4431), .o (n4432) );
  buffer buf_n4433( .i (n4432), .o (n4433) );
  buffer buf_n4434( .i (n4433), .o (n4434) );
  buffer buf_n4435( .i (n4434), .o (n4435) );
  buffer buf_n4436( .i (n4435), .o (n4436) );
  buffer buf_n4437( .i (n4436), .o (n4437) );
  buffer buf_n4438( .i (n4437), .o (n4438) );
  buffer buf_n4439( .i (n4438), .o (n4439) );
  assign n4440 = ~n2418 & n4439 ;
  assign n4441 = n4401 | n4440 ;
  buffer buf_n4442( .i (n4441), .o (n4442) );
  assign n4443 = n1381 & n1414 ;
  buffer buf_n4444( .i (n4443), .o (n4444) );
  assign n4445 = n1444 & ~n4444 ;
  buffer buf_n4446( .i (n4445), .o (n4446) );
  buffer buf_n4447( .i (n4446), .o (n4447) );
  buffer buf_n4448( .i (n4447), .o (n4448) );
  buffer buf_n4449( .i (n4448), .o (n4449) );
  buffer buf_n4450( .i (n4449), .o (n4450) );
  buffer buf_n4451( .i (n4450), .o (n4451) );
  buffer buf_n4452( .i (n4451), .o (n4452) );
  buffer buf_n4453( .i (n4452), .o (n4453) );
  buffer buf_n4454( .i (n4453), .o (n4454) );
  buffer buf_n4455( .i (n4454), .o (n4455) );
  buffer buf_n4456( .i (n4455), .o (n4456) );
  buffer buf_n4457( .i (n4456), .o (n4457) );
  buffer buf_n4458( .i (n4457), .o (n4458) );
  buffer buf_n4459( .i (n4458), .o (n4459) );
  buffer buf_n4460( .i (n4459), .o (n4460) );
  buffer buf_n4461( .i (n4460), .o (n4461) );
  buffer buf_n4462( .i (n4461), .o (n4462) );
  buffer buf_n4463( .i (n4462), .o (n4463) );
  buffer buf_n4464( .i (n4463), .o (n4464) );
  buffer buf_n4465( .i (n4464), .o (n4465) );
  buffer buf_n4466( .i (n4465), .o (n4466) );
  buffer buf_n4467( .i (n4466), .o (n4467) );
  buffer buf_n4468( .i (n4467), .o (n4468) );
  buffer buf_n4469( .i (n4468), .o (n4469) );
  buffer buf_n4470( .i (n4469), .o (n4470) );
  buffer buf_n4471( .i (n4470), .o (n4471) );
  buffer buf_n4472( .i (n4471), .o (n4472) );
  buffer buf_n4473( .i (n4472), .o (n4473) );
  buffer buf_n4474( .i (n4473), .o (n4474) );
  assign n4475 = n4442 & ~n4474 ;
  assign n4476 = ~n4442 & n4474 ;
  assign n4477 = n4475 | n4476 ;
  buffer buf_n4478( .i (n4477), .o (n4478) );
  buffer buf_n4479( .i (n4478), .o (n4479) );
  assign n4480 = n821 | n887 ;
  buffer buf_n4481( .i (n4480), .o (n4481) );
  assign n4482 = ~n916 & n4481 ;
  buffer buf_n4483( .i (n4482), .o (n4483) );
  buffer buf_n4484( .i (n4483), .o (n4484) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  assign n4485 = n843 & ~n974 ;
  assign n4486 = n944 & ~n4111 ;
  buffer buf_n4487( .i (n4486), .o (n4487) );
  assign n4488 = n4485 | n4487 ;
  buffer buf_n4489( .i (n4488), .o (n4489) );
  assign n4490 = ~n1003 & n4070 ;
  assign n4491 = n1003 & ~n4070 ;
  assign n4492 = n4490 | n4491 ;
  buffer buf_n4493( .i (n4492), .o (n4493) );
  assign n4494 = n4489 | n4493 ;
  assign n4495 = n4489 & n4493 ;
  assign n4496 = n4494 & ~n4495 ;
  buffer buf_n4497( .i (n4496), .o (n4497) );
  assign n4498 = ~n4484 & n4497 ;
  assign n4499 = n4484 & ~n4497 ;
  assign n4500 = n4498 | n4499 ;
  buffer buf_n4501( .i (n4500), .o (n4501) );
  buffer buf_n4502( .i (n4501), .o (n4502) );
  buffer buf_n4503( .i (n4502), .o (n4503) );
  buffer buf_n4504( .i (n4503), .o (n4504) );
  buffer buf_n4505( .i (n4504), .o (n4505) );
  buffer buf_n4506( .i (n4505), .o (n4506) );
  buffer buf_n4507( .i (n4506), .o (n4507) );
  buffer buf_n4508( .i (n4507), .o (n4508) );
  buffer buf_n4509( .i (n4508), .o (n4509) );
  buffer buf_n4510( .i (n4509), .o (n4510) );
  buffer buf_n4511( .i (n4510), .o (n4511) );
  buffer buf_n4512( .i (n4511), .o (n4512) );
  buffer buf_n4513( .i (n4512), .o (n4513) );
  buffer buf_n4514( .i (n4513), .o (n4514) );
  buffer buf_n4515( .i (n4514), .o (n4515) );
  buffer buf_n4516( .i (n4515), .o (n4516) );
  buffer buf_n4517( .i (n4516), .o (n4517) );
  buffer buf_n4518( .i (n4517), .o (n4518) );
  buffer buf_n4519( .i (n4518), .o (n4519) );
  buffer buf_n4520( .i (n4519), .o (n4520) );
  buffer buf_n4521( .i (n4520), .o (n4521) );
  buffer buf_n4522( .i (n4521), .o (n4522) );
  buffer buf_n4523( .i (n4522), .o (n4523) );
  buffer buf_n4524( .i (n4523), .o (n4524) );
  assign n4525 = n2426 & ~n4524 ;
  assign n4526 = n842 & n944 ;
  assign n4527 = n974 & ~n4526 ;
  buffer buf_n4528( .i (n4527), .o (n4528) );
  assign n4529 = ~n1005 & n4528 ;
  assign n4530 = n1005 & ~n4528 ;
  assign n4531 = n4529 | n4530 ;
  buffer buf_n4532( .i (n4531), .o (n4532) );
  buffer buf_n4533( .i (n4532), .o (n4533) );
  buffer buf_n4534( .i (n4533), .o (n4534) );
  buffer buf_n4535( .i (n4534), .o (n4535) );
  buffer buf_n4536( .i (n4535), .o (n4536) );
  buffer buf_n4537( .i (n4536), .o (n4537) );
  assign n4538 = n4113 | n4150 ;
  assign n4539 = ~n976 & n4538 ;
  buffer buf_n4540( .i (n4539), .o (n4540) );
  assign n4541 = n4074 & n4540 ;
  assign n4542 = n4074 | n4540 ;
  assign n4543 = ~n4541 & n4542 ;
  buffer buf_n4544( .i (n4543), .o (n4544) );
  assign n4545 = n1038 | n4544 ;
  assign n4546 = n1038 & n4544 ;
  assign n4547 = n4545 & ~n4546 ;
  buffer buf_n4548( .i (n4547), .o (n4548) );
  assign n4549 = n4537 & n4548 ;
  assign n4550 = n4537 | n4548 ;
  assign n4551 = ~n4549 & n4550 ;
  buffer buf_n4552( .i (n4551), .o (n4552) );
  buffer buf_n4553( .i (n4552), .o (n4553) );
  buffer buf_n4554( .i (n4553), .o (n4554) );
  buffer buf_n4555( .i (n4554), .o (n4555) );
  buffer buf_n4556( .i (n4555), .o (n4556) );
  buffer buf_n4557( .i (n4556), .o (n4557) );
  buffer buf_n4558( .i (n4557), .o (n4558) );
  buffer buf_n4559( .i (n4558), .o (n4559) );
  buffer buf_n4560( .i (n4559), .o (n4560) );
  buffer buf_n4561( .i (n4560), .o (n4561) );
  buffer buf_n4562( .i (n4561), .o (n4562) );
  buffer buf_n4563( .i (n4562), .o (n4563) );
  buffer buf_n4564( .i (n4563), .o (n4564) );
  buffer buf_n4565( .i (n4564), .o (n4565) );
  buffer buf_n4566( .i (n4565), .o (n4566) );
  buffer buf_n4567( .i (n4566), .o (n4567) );
  buffer buf_n4568( .i (n4567), .o (n4568) );
  buffer buf_n4569( .i (n4568), .o (n4569) );
  buffer buf_n4570( .i (n4569), .o (n4570) );
  buffer buf_n4571( .i (n4570), .o (n4571) );
  assign n4572 = ~n2426 & n4571 ;
  assign n4573 = n4525 | n4572 ;
  buffer buf_n4574( .i (n4573), .o (n4574) );
  assign n4575 = n4479 & ~n4574 ;
  assign n4576 = ~n4479 & n4574 ;
  assign n4577 = ~n4575 & ~n4576 ;
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n4578( .i (n2644), .o (n4578) );
  assign n4579 = n412 & n4578 ;
  assign n4580 = n408 | n4579 ;
  buffer buf_n4581( .i (n4580), .o (n4581) );
  assign n4582 = ~n688 & n2477 ;
  assign n4583 = n688 & ~n2477 ;
  assign n4584 = n4582 | n4583 ;
  buffer buf_n4585( .i (n4584), .o (n4585) );
  assign n4586 = ~n281 & n4585 ;
  assign n4587 = n281 & ~n4585 ;
  assign n4588 = n4586 | n4587 ;
  buffer buf_n4589( .i (n4588), .o (n4589) );
  assign n4590 = n2481 | n2523 ;
  buffer buf_n4591( .i (n4590), .o (n4591) );
  assign n4592 = ~n2569 & n4591 ;
  buffer buf_n4593( .i (n4592), .o (n4593) );
  buffer buf_n4594( .i (n4593), .o (n4594) );
  buffer buf_n4595( .i (n4594), .o (n4595) );
  buffer buf_n4596( .i (n4595), .o (n4596) );
  buffer buf_n4597( .i (n4596), .o (n4597) );
  buffer buf_n4598( .i (n4597), .o (n4598) );
  assign n4599 = n3996 & ~n4598 ;
  assign n4600 = ~n3996 & n4598 ;
  assign n4601 = n4599 | n4600 ;
  buffer buf_n4602( .i (n4601), .o (n4602) );
  assign n4603 = n655 & n2603 ;
  buffer buf_n4604( .i (n4603), .o (n4604) );
  buffer buf_n4605( .i (n4604), .o (n4605) );
  buffer buf_n4606( .i (n4605), .o (n4606) );
  buffer buf_n4607( .i (n4606), .o (n4607) );
  buffer buf_n4608( .i (n4607), .o (n4608) );
  buffer buf_n4609( .i (n4608), .o (n4609) );
  buffer buf_n4610( .i (n4609), .o (n4610) );
  assign n4611 = n4602 & ~n4610 ;
  buffer buf_n4612( .i (n4611), .o (n4612) );
  assign n4613 = n609 & ~n2605 ;
  buffer buf_n4614( .i (n4613), .o (n4614) );
  assign n4615 = n514 | n2479 ;
  assign n4616 = n568 & n2479 ;
  assign n4617 = n4615 & ~n4616 ;
  buffer buf_n4618( .i (n4617), .o (n4618) );
  assign n4619 = n692 & n4618 ;
  assign n4620 = n692 | n4618 ;
  assign n4621 = ~n4619 & n4620 ;
  buffer buf_n4622( .i (n4621), .o (n4622) );
  buffer buf_n4623( .i (n4622), .o (n4623) );
  buffer buf_n4624( .i (n4623), .o (n4624) );
  buffer buf_n4625( .i (n4624), .o (n4625) );
  buffer buf_n4626( .i (n4625), .o (n4626) );
  assign n4627 = ~n4614 & n4626 ;
  assign n4628 = n4614 & ~n4626 ;
  assign n4629 = n4627 | n4628 ;
  buffer buf_n4630( .i (n4629), .o (n4630) );
  buffer buf_n4631( .i (n4630), .o (n4631) );
  buffer buf_n4632( .i (n4631), .o (n4632) );
  buffer buf_n4633( .i (n4632), .o (n4633) );
  assign n4634 = n4612 & ~n4633 ;
  assign n4635 = ~n4612 & n4633 ;
  assign n4636 = n4634 | n4635 ;
  buffer buf_n4637( .i (n4636), .o (n4637) );
  buffer buf_n4638( .i (n4637), .o (n4638) );
  buffer buf_n4639( .i (n4638), .o (n4639) );
  buffer buf_n4640( .i (n4639), .o (n4640) );
  buffer buf_n4641( .i (n4640), .o (n4641) );
  buffer buf_n4642( .i (n4641), .o (n4642) );
  buffer buf_n4643( .i (n4642), .o (n4643) );
  buffer buf_n4644( .i (n4643), .o (n4644) );
  buffer buf_n4645( .i (n4644), .o (n4645) );
  buffer buf_n4646( .i (n4645), .o (n4646) );
  buffer buf_n4647( .i (n4646), .o (n4647) );
  buffer buf_n4648( .i (n4647), .o (n4648) );
  buffer buf_n4649( .i (n4648), .o (n4649) );
  buffer buf_n4650( .i (n4649), .o (n4650) );
  buffer buf_n4651( .i (n4650), .o (n4651) );
  buffer buf_n4652( .i (n4651), .o (n4652) );
  buffer buf_n4653( .i (n4652), .o (n4653) );
  buffer buf_n4654( .i (n4653), .o (n4654) );
  buffer buf_n4655( .i (n4654), .o (n4655) );
  buffer buf_n4656( .i (n4655), .o (n4656) );
  buffer buf_n4657( .i (n4656), .o (n4657) );
  buffer buf_n4658( .i (n4657), .o (n4658) );
  buffer buf_n4659( .i (n4658), .o (n4659) );
  buffer buf_n4660( .i (n4659), .o (n4660) );
  assign n4661 = n2438 | n4660 ;
  assign n4662 = n514 | n522 ;
  buffer buf_n4663( .i (n4662), .o (n4663) );
  assign n4664 = ~n570 & n4663 ;
  buffer buf_n4665( .i (n4664), .o (n4665) );
  assign n4666 = ~n693 & n4665 ;
  assign n4667 = n693 & ~n4665 ;
  assign n4668 = n4666 | n4667 ;
  buffer buf_n4669( .i (n4668), .o (n4669) );
  buffer buf_n4670( .i (n4669), .o (n4670) );
  assign n4671 = n609 | n4670 ;
  buffer buf_n4672( .i (n608), .o (n4672) );
  assign n4673 = n4670 & n4672 ;
  assign n4674 = n4671 & ~n4673 ;
  buffer buf_n4675( .i (n4674), .o (n4675) );
  buffer buf_n4676( .i (n4675), .o (n4676) );
  buffer buf_n4677( .i (n4676), .o (n4677) );
  buffer buf_n4678( .i (n4677), .o (n4678) );
  assign n4679 = n4602 & n4678 ;
  assign n4680 = n4602 | n4678 ;
  assign n4681 = ~n4679 & n4680 ;
  buffer buf_n4682( .i (n4681), .o (n4682) );
  buffer buf_n4683( .i (n4682), .o (n4683) );
  buffer buf_n4684( .i (n4683), .o (n4684) );
  buffer buf_n4685( .i (n4684), .o (n4685) );
  buffer buf_n4686( .i (n4685), .o (n4686) );
  buffer buf_n4687( .i (n4686), .o (n4687) );
  buffer buf_n4688( .i (n4687), .o (n4688) );
  buffer buf_n4689( .i (n4688), .o (n4689) );
  buffer buf_n4690( .i (n4689), .o (n4690) );
  buffer buf_n4691( .i (n4690), .o (n4691) );
  buffer buf_n4692( .i (n4691), .o (n4692) );
  buffer buf_n4693( .i (n4692), .o (n4693) );
  buffer buf_n4694( .i (n4693), .o (n4694) );
  buffer buf_n4695( .i (n4694), .o (n4695) );
  buffer buf_n4696( .i (n4695), .o (n4696) );
  buffer buf_n4697( .i (n4696), .o (n4697) );
  buffer buf_n4698( .i (n4697), .o (n4698) );
  buffer buf_n4699( .i (n4698), .o (n4699) );
  buffer buf_n4700( .i (n4699), .o (n4700) );
  buffer buf_n4701( .i (n4700), .o (n4701) );
  buffer buf_n4702( .i (n4701), .o (n4702) );
  buffer buf_n4703( .i (n4702), .o (n4703) );
  buffer buf_n4704( .i (n4703), .o (n4704) );
  buffer buf_n4705( .i (n4704), .o (n4705) );
  buffer buf_n4706( .i (n4705), .o (n4706) );
  buffer buf_n4707( .i (n4706), .o (n4707) );
  assign n4708 = n2438 & n4707 ;
  assign n4709 = n4661 & ~n4708 ;
  buffer buf_n4710( .i (n4709), .o (n4710) );
  assign n4711 = ~n4589 & n4710 ;
  assign n4712 = n4589 & ~n4710 ;
  assign n4713 = n4711 | n4712 ;
  buffer buf_n4714( .i (n4713), .o (n4714) );
  buffer buf_n4715( .i (n4714), .o (n4715) );
  buffer buf_n4716( .i (n4715), .o (n4716) );
  buffer buf_n4717( .i (n4716), .o (n4717) );
  assign n4718 = n4581 | n4717 ;
  assign n4719 = n4581 & n4717 ;
  assign n4720 = n4718 & ~n4719 ;
  assign n4721 = n1562 & n1570 ;
  buffer buf_n4722( .i (n4721), .o (n4722) );
  assign n4723 = n1595 & ~n4722 ;
  buffer buf_n4724( .i (n4723), .o (n4724) );
  assign n4725 = ~n1639 & n1667 ;
  assign n4726 = n4724 | n4725 ;
  buffer buf_n4727( .i (n4726), .o (n4727) );
  assign n4728 = ~n4274 & n4303 ;
  assign n4729 = n4274 & ~n4303 ;
  assign n4730 = n4728 | n4729 ;
  buffer buf_n4731( .i (n4730), .o (n4731) );
  assign n4732 = n4727 & ~n4731 ;
  assign n4733 = ~n4727 & n4731 ;
  assign n4734 = n4732 | n4733 ;
  buffer buf_n4735( .i (n4734), .o (n4735) );
  assign n4736 = n1734 & n4735 ;
  assign n4737 = n1734 | n4735 ;
  assign n4738 = ~n4736 & n4737 ;
  buffer buf_n4739( .i (n4738), .o (n4739) );
  buffer buf_n4740( .i (n4739), .o (n4740) );
  buffer buf_n4741( .i (n4740), .o (n4741) );
  buffer buf_n4742( .i (n4741), .o (n4742) );
  buffer buf_n4743( .i (n4742), .o (n4743) );
  buffer buf_n4744( .i (n4743), .o (n4744) );
  buffer buf_n4745( .i (n4744), .o (n4745) );
  buffer buf_n4746( .i (n4745), .o (n4746) );
  buffer buf_n4747( .i (n4746), .o (n4747) );
  buffer buf_n4748( .i (n4747), .o (n4748) );
  buffer buf_n4749( .i (n4748), .o (n4749) );
  buffer buf_n4750( .i (n4749), .o (n4750) );
  buffer buf_n4751( .i (n4750), .o (n4751) );
  buffer buf_n4752( .i (n4751), .o (n4752) );
  buffer buf_n4753( .i (n4752), .o (n4753) );
  assign n4754 = n2408 & ~n4753 ;
  buffer buf_n1551( .i (n1550), .o (n1551) );
  assign n4755 = n1542 | n1597 ;
  assign n4756 = ~n1551 & n4755 ;
  buffer buf_n4757( .i (n4756), .o (n4757) );
  assign n4758 = n1643 & ~n4757 ;
  assign n4759 = ~n1643 & n4757 ;
  assign n4760 = n4758 | n4759 ;
  buffer buf_n4761( .i (n4760), .o (n4761) );
  assign n4762 = n1597 & ~n1668 ;
  buffer buf_n1563( .i (n1562), .o (n1563) );
  assign n4763 = ~n1563 & n1665 ;
  buffer buf_n4764( .i (n4763), .o (n4764) );
  buffer buf_n4765( .i (n4764), .o (n4765) );
  buffer buf_n4766( .i (n4765), .o (n4766) );
  assign n4767 = n4762 | n4766 ;
  buffer buf_n4768( .i (n4767), .o (n4768) );
  assign n4769 = n4278 & ~n4768 ;
  assign n4770 = ~n4278 & n4768 ;
  assign n4771 = n4769 | n4770 ;
  buffer buf_n4772( .i (n4771), .o (n4772) );
  assign n4773 = n4761 | n4772 ;
  assign n4774 = n4761 & n4772 ;
  assign n4775 = n4773 & ~n4774 ;
  buffer buf_n4776( .i (n4775), .o (n4776) );
  buffer buf_n4777( .i (n4776), .o (n4777) );
  buffer buf_n4778( .i (n4777), .o (n4778) );
  buffer buf_n4779( .i (n4778), .o (n4779) );
  buffer buf_n4780( .i (n4779), .o (n4780) );
  buffer buf_n4781( .i (n4780), .o (n4781) );
  buffer buf_n4782( .i (n4781), .o (n4782) );
  buffer buf_n4783( .i (n4782), .o (n4783) );
  buffer buf_n4784( .i (n4783), .o (n4784) );
  buffer buf_n4785( .i (n4784), .o (n4785) );
  buffer buf_n4786( .i (n4785), .o (n4786) );
  buffer buf_n4787( .i (n4786), .o (n4787) );
  buffer buf_n4788( .i (n4787), .o (n4788) );
  buffer buf_n4789( .i (n4788), .o (n4789) );
  assign n4790 = n2408 | n4789 ;
  assign n4791 = ~n4754 & n4790 ;
  buffer buf_n4792( .i (n4791), .o (n4792) );
  assign n4793 = n1885 | n2354 ;
  buffer buf_n4794( .i (n4793), .o (n4794) );
  assign n4795 = ~n2376 & n4794 ;
  buffer buf_n4796( .i (n4795), .o (n4796) );
  assign n4797 = n1797 | n4240 ;
  assign n4798 = n1797 & n4240 ;
  assign n4799 = n4797 & ~n4798 ;
  buffer buf_n4800( .i (n4799), .o (n4800) );
  assign n4801 = n4796 & n4800 ;
  assign n4802 = n4796 | n4800 ;
  assign n4803 = ~n4801 & n4802 ;
  buffer buf_n4804( .i (n4803), .o (n4804) );
  buffer buf_n4805( .i (n4804), .o (n4805) );
  buffer buf_n4806( .i (n4805), .o (n4806) );
  buffer buf_n4807( .i (n4806), .o (n4807) );
  assign n4808 = n4208 | n4807 ;
  assign n4809 = n4208 & n4807 ;
  assign n4810 = n4808 & ~n4809 ;
  buffer buf_n4811( .i (n4810), .o (n4811) );
  buffer buf_n4812( .i (n4811), .o (n4812) );
  buffer buf_n4813( .i (n4812), .o (n4813) );
  buffer buf_n4814( .i (n4813), .o (n4814) );
  buffer buf_n4815( .i (n4814), .o (n4815) );
  assign n4816 = n2349 | n4815 ;
  assign n4817 = n1923 & n4208 ;
  assign n4818 = n1978 & ~n4817 ;
  buffer buf_n4819( .i (n4818), .o (n4819) );
  assign n4820 = ~n2378 & n4218 ;
  buffer buf_n4821( .i (n4820), .o (n4821) );
  assign n4822 = n1757 & ~n1814 ;
  buffer buf_n4823( .i (n4822), .o (n4823) );
  buffer buf_n4824( .i (n4823), .o (n4824) );
  buffer buf_n4825( .i (n4824), .o (n4825) );
  assign n4826 = ~n1790 & n1818 ;
  assign n4827 = n4825 | n4826 ;
  buffer buf_n4828( .i (n4827), .o (n4828) );
  buffer buf_n4829( .i (n4828), .o (n4829) );
  buffer buf_n4830( .i (n4829), .o (n4830) );
  buffer buf_n4831( .i (n4830), .o (n4831) );
  assign n4832 = n4821 | n4831 ;
  assign n4833 = n4821 & n4831 ;
  assign n4834 = n4832 & ~n4833 ;
  buffer buf_n4835( .i (n4834), .o (n4835) );
  buffer buf_n4836( .i (n4835), .o (n4836) );
  buffer buf_n4837( .i (n4836), .o (n4837) );
  buffer buf_n4838( .i (n4837), .o (n4838) );
  buffer buf_n4839( .i (n4838), .o (n4839) );
  assign n4840 = n4819 & ~n4839 ;
  assign n4841 = ~n4819 & n4839 ;
  assign n4842 = n4840 | n4841 ;
  buffer buf_n4843( .i (n4842), .o (n4843) );
  buffer buf_n4844( .i (n4843), .o (n4844) );
  assign n4845 = n2349 & n4844 ;
  assign n4846 = n4816 & ~n4845 ;
  buffer buf_n4847( .i (n4846), .o (n4847) );
  assign n4848 = n1851 & n1892 ;
  assign n4849 = n1915 & ~n4848 ;
  buffer buf_n4850( .i (n4849), .o (n4850) );
  buffer buf_n4851( .i (n4850), .o (n4851) );
  buffer buf_n4852( .i (n4851), .o (n4852) );
  buffer buf_n4853( .i (n4852), .o (n4853) );
  buffer buf_n4854( .i (n4853), .o (n4854) );
  buffer buf_n4855( .i (n4854), .o (n4855) );
  buffer buf_n4856( .i (n4855), .o (n4856) );
  buffer buf_n4857( .i (n4856), .o (n4857) );
  buffer buf_n4858( .i (n4857), .o (n4858) );
  buffer buf_n4859( .i (n4858), .o (n4859) );
  buffer buf_n4860( .i (n4859), .o (n4860) );
  buffer buf_n4861( .i (n4860), .o (n4861) );
  buffer buf_n4862( .i (n4861), .o (n4862) );
  buffer buf_n4863( .i (n4862), .o (n4863) );
  buffer buf_n4864( .i (n4863), .o (n4864) );
  buffer buf_n4865( .i (n4864), .o (n4865) );
  buffer buf_n4866( .i (n4865), .o (n4866) );
  assign n4867 = n4847 & ~n4866 ;
  assign n4868 = ~n4847 & n4866 ;
  assign n4869 = n4867 | n4868 ;
  buffer buf_n4870( .i (n4869), .o (n4870) );
  buffer buf_n4871( .i (n4870), .o (n4871) );
  buffer buf_n4872( .i (n4871), .o (n4872) );
  assign n4873 = ~n4792 & n4872 ;
  assign n4874 = n4792 & ~n4872 ;
  assign n4875 = n4873 | n4874 ;
  assign n4876 = n2059 | n2260 ;
  assign n4877 = n2030 & n2257 ;
  buffer buf_n4878( .i (n4877), .o (n4878) );
  buffer buf_n4879( .i (n4878), .o (n4879) );
  buffer buf_n4880( .i (n4879), .o (n4880) );
  assign n4881 = n4876 & ~n4880 ;
  buffer buf_n4882( .i (n4881), .o (n4882) );
  buffer buf_n4883( .i (n4882), .o (n4883) );
  buffer buf_n4884( .i (n4883), .o (n4884) );
  assign n4885 = n2080 | n4884 ;
  assign n4886 = n2080 & n4884 ;
  assign n4887 = n4885 & ~n4886 ;
  buffer buf_n4888( .i (n4887), .o (n4888) );
  assign n4889 = n2295 & n2316 ;
  assign n4890 = n2333 & ~n4889 ;
  buffer buf_n4891( .i (n4890), .o (n4891) );
  assign n4896 = n2242 & ~n4891 ;
  assign n4897 = ~n2242 & n4891 ;
  assign n4898 = n4896 | n4897 ;
  buffer buf_n4899( .i (n4898), .o (n4899) );
  buffer buf_n4900( .i (n4899), .o (n4900) );
  assign n4901 = n4888 & n4900 ;
  assign n4902 = n4888 | n4900 ;
  assign n4903 = ~n4901 & n4902 ;
  buffer buf_n4904( .i (n4903), .o (n4904) );
  assign n4905 = n2232 & ~n4904 ;
  buffer buf_n4906( .i (n4905), .o (n4906) );
  buffer buf_n4892( .i (n4891), .o (n4892) );
  buffer buf_n4893( .i (n4892), .o (n4893) );
  buffer buf_n4894( .i (n4893), .o (n4894) );
  buffer buf_n4895( .i (n4894), .o (n4895) );
  assign n4907 = n2028 & ~n2039 ;
  buffer buf_n2031( .i (n2030), .o (n2031) );
  assign n4908 = n2031 & n2039 ;
  assign n4909 = n4907 | n4908 ;
  buffer buf_n4910( .i (n4909), .o (n4910) );
  buffer buf_n4911( .i (n4910), .o (n4911) );
  assign n4912 = n2291 & ~n4911 ;
  buffer buf_n4913( .i (n4912), .o (n4913) );
  buffer buf_n4914( .i (n4913), .o (n4914) );
  assign n4915 = n2080 & n4914 ;
  assign n4916 = n3345 & ~n4913 ;
  buffer buf_n4917( .i (n2079), .o (n4917) );
  assign n4918 = n4916 & ~n4917 ;
  assign n4919 = n4915 | n4918 ;
  buffer buf_n4920( .i (n4919), .o (n4920) );
  assign n4921 = ~n4895 & n4920 ;
  assign n4922 = n4895 & ~n4920 ;
  assign n4923 = n4921 | n4922 ;
  buffer buf_n4924( .i (n4923), .o (n4924) );
  assign n4925 = n2232 | n4924 ;
  assign n4926 = N367 & n4925 ;
  assign n4927 = ~n4906 & n4926 ;
  assign n4928 = ~n2201 & n4904 ;
  assign n4929 = ~N367 & n2199 ;
  buffer buf_n4930( .i (n4929), .o (n4930) );
  assign n4931 = n4924 & n4930 ;
  assign n4932 = n4928 | n4931 ;
  buffer buf_n4933( .i (n4932), .o (n4933) );
  assign n4934 = n4927 | n4933 ;
  buffer buf_n4935( .i (n4934), .o (n4935) );
  buffer buf_n4936( .i (n4935), .o (n4936) );
  buffer buf_n4937( .i (n4936), .o (n4937) );
  buffer buf_n4938( .i (n4937), .o (n4938) );
  assign n4939 = ~n2144 & n2188 ;
  buffer buf_n4940( .i (n4939), .o (n4940) );
  assign n4941 = n2193 & ~n4940 ;
  buffer buf_n4942( .i (n4941), .o (n4942) );
  buffer buf_n4943( .i (n4942), .o (n4943) );
  buffer buf_n4944( .i (n4943), .o (n4944) );
  buffer buf_n4945( .i (n4944), .o (n4945) );
  assign n4946 = ~n2177 & n3332 ;
  buffer buf_n4947( .i (n4946), .o (n4947) );
  buffer buf_n4948( .i (n4947), .o (n4948) );
  buffer buf_n4949( .i (n4948), .o (n4949) );
  buffer buf_n4950( .i (n4949), .o (n4950) );
  buffer buf_n4951( .i (n4950), .o (n4951) );
  buffer buf_n4952( .i (n4951), .o (n4952) );
  assign n4953 = n227 & n2208 ;
  buffer buf_n4954( .i (n4953), .o (n4954) );
  assign n4955 = n2212 & ~n4954 ;
  buffer buf_n4956( .i (n4955), .o (n4956) );
  assign n4957 = n3312 & n4956 ;
  assign n4958 = n3312 | n4956 ;
  assign n4959 = ~n4957 & n4958 ;
  buffer buf_n4960( .i (n4959), .o (n4960) );
  assign n4963 = ~n4952 & n4960 ;
  assign n4964 = n4952 & ~n4960 ;
  assign n4965 = n4963 | n4964 ;
  buffer buf_n4966( .i (n4965), .o (n4966) );
  assign n4967 = n4945 & ~n4966 ;
  buffer buf_n4968( .i (n4967), .o (n4968) );
  assign n4969 = ~n4945 & n4966 ;
  assign n4970 = N367 | n4969 ;
  assign n4971 = n4968 | n4970 ;
  buffer buf_n4972( .i (n4971), .o (n4972) );
  buffer buf_n4973( .i (n4972), .o (n4973) );
  assign n4974 = ~n2189 & n2214 ;
  buffer buf_n4975( .i (n4974), .o (n4975) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  assign n4976 = n220 | n2172 ;
  buffer buf_n4977( .i (n4976), .o (n4977) );
  buffer buf_n4978( .i (n4977), .o (n4978) );
  buffer buf_n4979( .i (n4978), .o (n4979) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n2182( .i (n2181), .o (n2182) );
  buffer buf_n2183( .i (n2182), .o (n2183) );
  assign n4980 = n2177 | n2183 ;
  assign n4981 = n223 & ~n4980 ;
  assign n4982 = n4979 & ~n4981 ;
  buffer buf_n4983( .i (n4982), .o (n4983) );
  buffer buf_n4984( .i (n4983), .o (n4984) );
  buffer buf_n4985( .i (n4984), .o (n4985) );
  assign n4986 = ~n4975 & n4985 ;
  assign n4987 = n4975 & ~n4985 ;
  assign n4988 = n4986 | n4987 ;
  buffer buf_n4989( .i (n4988), .o (n4989) );
  buffer buf_n4990( .i (n4989), .o (n4990) );
  buffer buf_n4991( .i (n4990), .o (n4991) );
  buffer buf_n4992( .i (n4991), .o (n4992) );
  buffer buf_n4961( .i (n4960), .o (n4961) );
  buffer buf_n4962( .i (n4961), .o (n4962) );
  assign n4993 = n2229 & ~n4962 ;
  assign n4994 = ~n2229 & n4962 ;
  assign n4995 = n4993 | n4994 ;
  buffer buf_n4996( .i (n4995), .o (n4996) );
  assign n4997 = n4992 & n4996 ;
  buffer buf_n4998( .i (n4997), .o (n4998) );
  assign n4999 = n4992 | n4996 ;
  assign n5000 = N367 & n4999 ;
  assign n5001 = ~n4998 & n5000 ;
  assign n5002 = n4973 & ~n5001 ;
  buffer buf_n5003( .i (n5002), .o (n5003) );
  assign n5004 = n2204 & n2217 ;
  assign n5005 = n2204 | n2217 ;
  assign n5006 = ~n5004 & n5005 ;
  buffer buf_n5007( .i (n5006), .o (n5007) );
  buffer buf_n5008( .i (n5007), .o (n5008) );
  buffer buf_n5009( .i (n5008), .o (n5009) );
  buffer buf_n5010( .i (n5009), .o (n5010) );
  buffer buf_n5011( .i (n5010), .o (n5011) );
  buffer buf_n5012( .i (n5011), .o (n5012) );
  buffer buf_n5013( .i (n5012), .o (n5013) );
  buffer buf_n5014( .i (n5013), .o (n5014) );
  buffer buf_n5015( .i (n5014), .o (n5015) );
  buffer buf_n5016( .i (n5015), .o (n5016) );
  buffer buf_n5017( .i (n5016), .o (n5017) );
  buffer buf_n5018( .i (n5017), .o (n5018) );
  buffer buf_n5019( .i (n5018), .o (n5019) );
  buffer buf_n5020( .i (n5019), .o (n5020) );
  assign n5021 = n5003 | n5020 ;
  assign n5022 = n5003 & n5020 ;
  assign n5023 = n5021 & ~n5022 ;
  buffer buf_n5024( .i (n5023), .o (n5024) );
  assign n5025 = n4938 | n5024 ;
  assign n5026 = n4938 & n5024 ;
  assign n5027 = n5025 & ~n5026 ;
  assign n5028 = N1 & N163 ;
  assign n5029 = N5 | N57 ;
  inverter inv_n5033( .i (n4050), .o (n5033) );
  inverter inv_n5034( .i (n4054), .o (n5034) );
  inverter inv_n5035( .i (n4059), .o (n5035) );
  inverter inv_n5036( .i (n4063), .o (n5036) );
  assign N10025 = n232 ;
  assign N10101 = n2650 ;
  assign N10102 = n3306 ;
  assign N10103 = n3306 ;
  assign N10104 = n2650 ;
  assign N10109 = n3325 ;
  assign N10110 = n3330 ;
  assign N10111 = n3338 ;
  assign N10112 = n3343 ;
  assign N10350 = n3360 ;
  assign N10351 = n3368 ;
  assign N10352 = n3373 ;
  assign N10353 = n3376 ;
  assign N10574 = n5030 ;
  assign N10575 = n5031 ;
  assign N10576 = n5032 ;
  assign N10628 = n3306 ;
  assign N10632 = n3907 ;
  assign N10641 = n3912 ;
  assign N10704 = n2972 ;
  assign N10706 = n2650 ;
  assign N10711 = n3977 ;
  assign N10712 = n3982 ;
  assign N10713 = n3988 ;
  assign N10714 = n3993 ;
  assign N10715 = n4030 ;
  assign N10716 = n4035 ;
  assign N10717 = n4041 ;
  assign N10718 = n4046 ;
  assign N10729 = n4068 ;
  assign N10759 = n2650 ;
  assign N10760 = n4103 ;
  assign N10761 = n4109 ;
  assign N10762 = n4148 ;
  assign N10763 = n4184 ;
  assign N10827 = n4191 ;
  assign N10837 = n4199 ;
  assign N10838 = n4199 ;
  assign N10839 = n4203 ;
  assign N10840 = n4203 ;
  assign N10868 = n4216 ;
  assign N10869 = n4235 ;
  assign N10870 = n4266 ;
  assign N10871 = n4271 ;
  assign N10905 = n4300 ;
  assign N10906 = n4332 ;
  assign N10907 = n4338 ;
  assign N10908 = n4341 ;
  assign N1110 = n4343 ;
  assign N1111 = ~N15 ;
  assign N1112 = n4343 ;
  assign N1113 = n4346 ;
  assign N1114 = ~N15 ;
  assign N11333 = n4577 ;
  assign N11334 = n4720 ;
  assign N11340 = n4875 ;
  assign N11342 = n5027 ;
  assign N1489 = n4346 ;
  assign N1490 = N1 ;
  assign N1781 = n5028 ;
  assign N241_O = N241_I ;
  assign N387 = N1 ;
  assign N388 = N1 ;
  assign N478 = N248 ;
  assign N482 = N254 ;
  assign N484 = N257 ;
  assign N486 = N260 ;
  assign N489 = N263 ;
  assign N492 = N267 ;
  assign N501 = N274 ;
  assign N505 = N280 ;
  assign N507 = N283 ;
  assign N509 = N286 ;
  assign N511 = N289 ;
  assign N513 = N293 ;
  assign N515 = N296 ;
  assign N517 = N299 ;
  assign N519 = N303 ;
  assign N535 = N307 ;
  assign N537 = N310 ;
  assign N539 = N313 ;
  assign N541 = N316 ;
  assign N543 = N319 ;
  assign N545 = N322 ;
  assign N547 = N325 ;
  assign N549 = N328 ;
  assign N551 = N331 ;
  assign N553 = N334 ;
  assign N556 = N337 ;
  assign N559 = N343 ;
  assign N561 = N346 ;
  assign N563 = N349 ;
  assign N565 = N352 ;
  assign N567 = N355 ;
  assign N569 = N358 ;
  assign N571 = N361 ;
  assign N573 = N364 ;
  assign N582 = ~N15 ;
  assign N643 = N251 ;
  assign N707 = N277 ;
  assign N813 = N340 ;
  assign N881 = n5029 ;
  assign N882 = n5033 ;
  assign N883 = n5034 ;
  assign N884 = n5035 ;
  assign N885 = n5036 ;
  assign N889 = N1 ;
  assign N945 = N106 ;
endmodule
