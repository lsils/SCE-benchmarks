module ALU32(io_in2_1_,io_in1_7_,io_in2_4_,io_in2_16_,io_in1_11_,io_in2_26_,io_fn_0_,io_in2_12_,io_in2_21_,io_in2_14_,io_in1_3_,io_in1_17_,io_in1_20_,io_in1_6_,io_in1_5_,io_in1_18_,io_in2_27_,io_in2_28_,io_in2_25_,io_in1_14_,io_in2_17_,io_in1_25_,io_in1_2_,io_in1_15_,io_in2_22_,io_in1_8_,io_in1_21_,io_in2_23_,io_in1_19_,io_in2_6_,io_in2_9_,io_in2_3_,io_in1_13_,io_in1_23_,io_in2_13_,io_in1_12_,io_in1_0_,io_in2_15_,io_fn_2_,io_in1_28_,io_in2_8_,io_in1_31_,io_in2_0_,io_in2_20_,io_in2_5_,io_in2_29_,io_in2_31_,io_in2_18_,io_in1_16_,io_in1_1_,io_in1_29_,io_in2_24_,io_in2_30_,io_in1_9_,io_in1_30_,io_in2_19_,io_in2_7_,io_in2_2_,io_in1_27_,io_in2_11_,io_in1_24_,io_fn_3_,io_in2_10_,io_fn_1_,io_in1_4_,io_in1_26_,io_in1_10_,io_in1_22_,io_out_22_,io_adder_out_22_,io_out_7_,io_test_adder_Cout,io_adder_out_17_,io_adder_out_26_,io_adder_out_1_,io_adder_out_23_,io_out_1_,io_adder_out_8_,io_adder_out_0_,io_adder_out_7_,io_out_15_,io_out_31_,io_adder_out_10_,io_out_25_,io_out_10_,io_out_14_,io_out_24_,io_adder_out_5_,io_out_12_,io_adder_out_9_,io_adder_out_30_,io_adder_out_12_,io_adder_out_13_,io_out_13_,io_out_21_,io_adder_out_16_,io_out_30_,io_adder_out_2_,io_out_2_,io_adder_out_31_,io_adder_out_14_,io_out_26_,io_out_17_,io_adder_out_6_,io_out_18_,io_out_0_,io_out_4_,io_out_19_,io_adder_out_19_,io_out_23_,io_out_8_,io_adder_out_20_,io_out_20_,io_adder_out_25_,io_adder_out_29_,io_adder_out_15_,io_out_3_,io_out_28_,io_out_27_,io_adder_out_11_,io_out_5_,io_adder_out_4_,io_out_9_,io_adder_out_28_,io_adder_out_21_,io_adder_out_24_,io_out_29_,io_adder_out_27_,io_out_16_,io_out_11_,io_out_6_,io_adder_out_3_,io_adder_out_18_);
    wire jinkela_wire_0;
    wire jinkela_wire_1;
    wire jinkela_wire_2;
    wire jinkela_wire_3;
    wire jinkela_wire_4;
    wire jinkela_wire_5;
    wire jinkela_wire_6;
    wire jinkela_wire_7;
    wire jinkela_wire_8;
    wire jinkela_wire_9;
    wire jinkela_wire_10;
    wire jinkela_wire_11;
    wire jinkela_wire_12;
    wire jinkela_wire_13;
    wire jinkela_wire_14;
    wire jinkela_wire_15;
    wire jinkela_wire_16;
    wire jinkela_wire_17;
    wire jinkela_wire_18;
    wire jinkela_wire_19;
    wire jinkela_wire_20;
    wire jinkela_wire_21;
    wire jinkela_wire_22;
    wire jinkela_wire_23;
    wire jinkela_wire_24;
    wire jinkela_wire_25;
    wire jinkela_wire_26;
    wire jinkela_wire_27;
    wire jinkela_wire_28;
    wire jinkela_wire_29;
    wire jinkela_wire_30;
    wire jinkela_wire_31;
    wire jinkela_wire_32;
    wire jinkela_wire_33;
    wire jinkela_wire_34;
    wire jinkela_wire_35;
    wire jinkela_wire_36;
    wire jinkela_wire_37;
    wire jinkela_wire_38;
    wire jinkela_wire_39;
    wire jinkela_wire_40;
    wire jinkela_wire_41;
    wire jinkela_wire_42;
    wire jinkela_wire_43;
    wire jinkela_wire_44;
    wire jinkela_wire_45;
    wire jinkela_wire_46;
    wire jinkela_wire_47;
    wire jinkela_wire_48;
    wire jinkela_wire_49;
    wire jinkela_wire_50;
    wire jinkela_wire_51;
    wire jinkela_wire_52;
    wire jinkela_wire_53;
    wire jinkela_wire_54;
    wire jinkela_wire_55;
    wire jinkela_wire_56;
    wire jinkela_wire_57;
    wire jinkela_wire_58;
    wire jinkela_wire_59;
    wire jinkela_wire_60;
    wire jinkela_wire_61;
    wire jinkela_wire_62;
    wire jinkela_wire_63;
    wire jinkela_wire_64;
    wire jinkela_wire_65;
    wire jinkela_wire_66;
    wire jinkela_wire_67;
    wire jinkela_wire_68;
    wire jinkela_wire_69;
    wire jinkela_wire_70;
    wire jinkela_wire_71;
    wire jinkela_wire_72;
    wire jinkela_wire_73;
    wire jinkela_wire_74;
    wire jinkela_wire_75;
    wire jinkela_wire_76;
    wire jinkela_wire_77;
    wire jinkela_wire_78;
    wire jinkela_wire_79;
    wire jinkela_wire_80;
    wire jinkela_wire_81;
    wire jinkela_wire_82;
    wire jinkela_wire_83;
    wire jinkela_wire_84;
    wire jinkela_wire_85;
    wire jinkela_wire_86;
    wire jinkela_wire_87;
    wire jinkela_wire_88;
    wire jinkela_wire_89;
    wire jinkela_wire_90;
    wire jinkela_wire_91;
    wire jinkela_wire_92;
    wire jinkela_wire_93;
    wire jinkela_wire_94;
    wire jinkela_wire_95;
    wire jinkela_wire_96;
    wire jinkela_wire_97;
    wire jinkela_wire_98;
    wire jinkela_wire_99;
    wire jinkela_wire_100;
    wire jinkela_wire_101;
    wire jinkela_wire_102;
    wire jinkela_wire_103;
    wire jinkela_wire_104;
    wire jinkela_wire_105;
    wire jinkela_wire_106;
    wire jinkela_wire_107;
    wire jinkela_wire_108;
    wire jinkela_wire_109;
    wire jinkela_wire_110;
    wire jinkela_wire_111;
    wire jinkela_wire_112;
    wire jinkela_wire_113;
    wire jinkela_wire_114;
    wire jinkela_wire_115;
    wire jinkela_wire_116;
    wire jinkela_wire_117;
    wire jinkela_wire_118;
    wire jinkela_wire_119;
    wire jinkela_wire_120;
    wire jinkela_wire_121;
    wire jinkela_wire_122;
    wire jinkela_wire_123;
    wire jinkela_wire_124;
    wire jinkela_wire_125;
    wire jinkela_wire_126;
    wire jinkela_wire_127;
    wire jinkela_wire_128;
    wire jinkela_wire_129;
    wire jinkela_wire_130;
    wire jinkela_wire_131;
    wire jinkela_wire_132;
    wire jinkela_wire_133;
    wire jinkela_wire_134;
    wire jinkela_wire_135;
    wire jinkela_wire_136;
    wire jinkela_wire_137;
    wire jinkela_wire_138;
    wire jinkela_wire_139;
    wire jinkela_wire_140;
    wire jinkela_wire_141;
    wire jinkela_wire_142;
    wire jinkela_wire_143;
    wire jinkela_wire_144;
    wire jinkela_wire_145;
    wire jinkela_wire_146;
    wire jinkela_wire_147;
    wire jinkela_wire_148;
    wire jinkela_wire_149;
    wire jinkela_wire_150;
    wire jinkela_wire_151;
    wire jinkela_wire_152;
    wire jinkela_wire_153;
    wire jinkela_wire_154;
    wire jinkela_wire_155;
    wire jinkela_wire_156;
    wire jinkela_wire_157;
    wire jinkela_wire_158;
    wire jinkela_wire_159;
    wire jinkela_wire_160;
    wire jinkela_wire_161;
    wire jinkela_wire_162;
    wire jinkela_wire_163;
    wire jinkela_wire_164;
    wire jinkela_wire_165;
    wire jinkela_wire_166;
    wire jinkela_wire_167;
    wire jinkela_wire_168;
    wire jinkela_wire_169;
    wire jinkela_wire_170;
    wire jinkela_wire_171;
    wire jinkela_wire_172;
    wire jinkela_wire_173;
    wire jinkela_wire_174;
    wire jinkela_wire_175;
    wire jinkela_wire_176;
    wire jinkela_wire_177;
    wire jinkela_wire_178;
    wire jinkela_wire_179;
    wire jinkela_wire_180;
    wire jinkela_wire_181;
    wire jinkela_wire_182;
    wire jinkela_wire_183;
    wire jinkela_wire_184;
    wire jinkela_wire_185;
    wire jinkela_wire_186;
    wire jinkela_wire_187;
    wire jinkela_wire_188;
    wire jinkela_wire_189;
    wire jinkela_wire_190;
    wire jinkela_wire_191;
    wire jinkela_wire_192;
    wire jinkela_wire_193;
    wire jinkela_wire_194;
    wire jinkela_wire_195;
    wire jinkela_wire_196;
    wire jinkela_wire_197;
    wire jinkela_wire_198;
    wire jinkela_wire_199;
    wire jinkela_wire_200;
    wire jinkela_wire_201;
    wire jinkela_wire_202;
    wire jinkela_wire_203;
    wire jinkela_wire_204;
    wire jinkela_wire_205;
    wire jinkela_wire_206;
    wire jinkela_wire_207;
    wire jinkela_wire_208;
    wire jinkela_wire_209;
    wire jinkela_wire_210;
    wire jinkela_wire_211;
    wire jinkela_wire_212;
    wire jinkela_wire_213;
    wire jinkela_wire_214;
    wire jinkela_wire_215;
    wire jinkela_wire_216;
    wire jinkela_wire_217;
    wire jinkela_wire_218;
    wire jinkela_wire_219;
    wire jinkela_wire_220;
    wire jinkela_wire_221;
    wire jinkela_wire_222;
    wire jinkela_wire_223;
    wire jinkela_wire_224;
    wire jinkela_wire_225;
    wire jinkela_wire_226;
    wire jinkela_wire_227;
    wire jinkela_wire_228;
    wire jinkela_wire_229;
    wire jinkela_wire_230;
    wire jinkela_wire_231;
    wire jinkela_wire_232;
    wire jinkela_wire_233;
    wire jinkela_wire_234;
    wire jinkela_wire_235;
    wire jinkela_wire_236;
    wire jinkela_wire_237;
    wire jinkela_wire_238;
    wire jinkela_wire_239;
    wire jinkela_wire_240;
    wire jinkela_wire_241;
    wire jinkela_wire_242;
    wire jinkela_wire_243;
    wire jinkela_wire_244;
    wire jinkela_wire_245;
    wire jinkela_wire_246;
    wire jinkela_wire_247;
    wire jinkela_wire_248;
    wire jinkela_wire_249;
    wire jinkela_wire_250;
    wire jinkela_wire_251;
    wire jinkela_wire_252;
    wire jinkela_wire_253;
    wire jinkela_wire_254;
    wire jinkela_wire_255;
    wire jinkela_wire_256;
    wire jinkela_wire_257;
    wire jinkela_wire_258;
    wire jinkela_wire_259;
    wire jinkela_wire_260;
    wire jinkela_wire_261;
    wire jinkela_wire_262;
    wire jinkela_wire_263;
    wire jinkela_wire_264;
    wire jinkela_wire_265;
    wire jinkela_wire_266;
    wire jinkela_wire_267;
    wire jinkela_wire_268;
    wire jinkela_wire_269;
    wire jinkela_wire_270;
    wire jinkela_wire_271;
    wire jinkela_wire_272;
    wire jinkela_wire_273;
    wire jinkela_wire_274;
    wire jinkela_wire_275;
    wire jinkela_wire_276;
    wire jinkela_wire_277;
    wire jinkela_wire_278;
    wire jinkela_wire_279;
    wire jinkela_wire_280;
    wire jinkela_wire_281;
    wire jinkela_wire_282;
    wire jinkela_wire_283;
    wire jinkela_wire_284;
    wire jinkela_wire_285;
    wire jinkela_wire_286;
    wire jinkela_wire_287;
    wire jinkela_wire_288;
    wire jinkela_wire_289;
    wire jinkela_wire_290;
    wire jinkela_wire_291;
    wire jinkela_wire_292;
    wire jinkela_wire_293;
    wire jinkela_wire_294;
    wire jinkela_wire_295;
    wire jinkela_wire_296;
    wire jinkela_wire_297;
    wire jinkela_wire_298;
    wire jinkela_wire_299;
    wire jinkela_wire_300;
    wire jinkela_wire_301;
    wire jinkela_wire_302;
    wire jinkela_wire_303;
    wire jinkela_wire_304;
    wire jinkela_wire_305;
    wire jinkela_wire_306;
    wire jinkela_wire_307;
    wire jinkela_wire_308;
    wire jinkela_wire_309;
    wire jinkela_wire_310;
    wire jinkela_wire_311;
    wire jinkela_wire_312;
    wire jinkela_wire_313;
    wire jinkela_wire_314;
    wire jinkela_wire_315;
    wire jinkela_wire_316;
    wire jinkela_wire_317;
    wire jinkela_wire_318;
    wire jinkela_wire_319;
    wire jinkela_wire_320;
    wire jinkela_wire_321;
    wire jinkela_wire_322;
    wire jinkela_wire_323;
    wire jinkela_wire_324;
    wire jinkela_wire_325;
    wire jinkela_wire_326;
    wire jinkela_wire_327;
    wire jinkela_wire_328;
    wire jinkela_wire_329;
    wire jinkela_wire_330;
    wire jinkela_wire_331;
    wire jinkela_wire_332;
    wire jinkela_wire_333;
    wire jinkela_wire_334;
    wire jinkela_wire_335;
    wire jinkela_wire_336;
    wire jinkela_wire_337;
    wire jinkela_wire_338;
    wire jinkela_wire_339;
    wire jinkela_wire_340;
    wire jinkela_wire_341;
    wire jinkela_wire_342;
    wire jinkela_wire_343;
    wire jinkela_wire_344;
    wire jinkela_wire_345;
    wire jinkela_wire_346;
    wire jinkela_wire_347;
    wire jinkela_wire_348;
    wire jinkela_wire_349;
    wire jinkela_wire_350;
    wire jinkela_wire_351;
    wire jinkela_wire_352;
    wire jinkela_wire_353;
    wire jinkela_wire_354;
    wire jinkela_wire_355;
    wire jinkela_wire_356;
    wire jinkela_wire_357;
    wire jinkela_wire_358;
    wire jinkela_wire_359;
    wire jinkela_wire_360;
    wire jinkela_wire_361;
    wire jinkela_wire_362;
    wire jinkela_wire_363;
    wire jinkela_wire_364;
    wire jinkela_wire_365;
    wire jinkela_wire_366;
    wire jinkela_wire_367;
    wire jinkela_wire_368;
    wire jinkela_wire_369;
    wire jinkela_wire_370;
    wire jinkela_wire_371;
    wire jinkela_wire_372;
    wire jinkela_wire_373;
    wire jinkela_wire_374;
    wire jinkela_wire_375;
    wire jinkela_wire_376;
    wire jinkela_wire_377;
    wire jinkela_wire_378;
    wire jinkela_wire_379;
    wire jinkela_wire_380;
    wire jinkela_wire_381;
    wire jinkela_wire_382;
    wire jinkela_wire_383;
    wire jinkela_wire_384;
    wire jinkela_wire_385;
    wire jinkela_wire_386;
    wire jinkela_wire_387;
    wire jinkela_wire_388;
    wire jinkela_wire_389;
    wire jinkela_wire_390;
    wire jinkela_wire_391;
    wire jinkela_wire_392;
    wire jinkela_wire_393;
    wire jinkela_wire_394;
    wire jinkela_wire_395;
    wire jinkela_wire_396;
    wire jinkela_wire_397;
    wire jinkela_wire_398;
    wire jinkela_wire_399;
    wire jinkela_wire_400;
    wire jinkela_wire_401;
    wire jinkela_wire_402;
    wire jinkela_wire_403;
    wire jinkela_wire_404;
    wire jinkela_wire_405;
    wire jinkela_wire_406;
    wire jinkela_wire_407;
    wire jinkela_wire_408;
    wire jinkela_wire_409;
    wire jinkela_wire_410;
    wire jinkela_wire_411;
    wire jinkela_wire_412;
    wire jinkela_wire_413;
    wire jinkela_wire_414;
    wire jinkela_wire_415;
    wire jinkela_wire_416;
    wire jinkela_wire_417;
    wire jinkela_wire_418;
    wire jinkela_wire_419;
    wire jinkela_wire_420;
    wire jinkela_wire_421;
    wire jinkela_wire_422;
    wire jinkela_wire_423;
    wire jinkela_wire_424;
    wire jinkela_wire_425;
    wire jinkela_wire_426;
    wire jinkela_wire_427;
    wire jinkela_wire_428;
    wire jinkela_wire_429;
    wire jinkela_wire_430;
    wire jinkela_wire_431;
    wire jinkela_wire_432;
    wire jinkela_wire_433;
    wire jinkela_wire_434;
    wire jinkela_wire_435;
    wire jinkela_wire_436;
    wire jinkela_wire_437;
    wire jinkela_wire_438;
    wire jinkela_wire_439;
    wire jinkela_wire_440;
    wire jinkela_wire_441;
    wire jinkela_wire_442;
    wire jinkela_wire_443;
    wire jinkela_wire_444;
    wire jinkela_wire_445;
    wire jinkela_wire_446;
    wire jinkela_wire_447;
    wire jinkela_wire_448;
    wire jinkela_wire_449;
    wire jinkela_wire_450;
    wire jinkela_wire_451;
    wire jinkela_wire_452;
    wire jinkela_wire_453;
    wire jinkela_wire_454;
    wire jinkela_wire_455;
    wire jinkela_wire_456;
    wire jinkela_wire_457;
    wire jinkela_wire_458;
    wire jinkela_wire_459;
    wire jinkela_wire_460;
    wire jinkela_wire_461;
    wire jinkela_wire_462;
    wire jinkela_wire_463;
    wire jinkela_wire_464;
    wire jinkela_wire_465;
    wire jinkela_wire_466;
    wire jinkela_wire_467;
    wire jinkela_wire_468;
    wire jinkela_wire_469;
    wire jinkela_wire_470;
    wire jinkela_wire_471;
    wire jinkela_wire_472;
    wire jinkela_wire_473;
    wire jinkela_wire_474;
    wire jinkela_wire_475;
    wire jinkela_wire_476;
    wire jinkela_wire_477;
    wire jinkela_wire_478;
    wire jinkela_wire_479;
    wire jinkela_wire_480;
    wire jinkela_wire_481;
    wire jinkela_wire_482;
    wire jinkela_wire_483;
    wire jinkela_wire_484;
    wire jinkela_wire_485;
    wire jinkela_wire_486;
    wire jinkela_wire_487;
    wire jinkela_wire_488;
    wire jinkela_wire_489;
    wire jinkela_wire_490;
    wire jinkela_wire_491;
    wire jinkela_wire_492;
    wire jinkela_wire_493;
    wire jinkela_wire_494;
    wire jinkela_wire_495;
    wire jinkela_wire_496;
    wire jinkela_wire_497;
    wire jinkela_wire_498;
    wire jinkela_wire_499;
    wire jinkela_wire_500;
    wire jinkela_wire_501;
    wire jinkela_wire_502;
    wire jinkela_wire_503;
    wire jinkela_wire_504;
    wire jinkela_wire_505;
    wire jinkela_wire_506;
    wire jinkela_wire_507;
    wire jinkela_wire_508;
    wire jinkela_wire_509;
    wire jinkela_wire_510;
    wire jinkela_wire_511;
    wire jinkela_wire_512;
    wire jinkela_wire_513;
    wire jinkela_wire_514;
    wire jinkela_wire_515;
    wire jinkela_wire_516;
    wire jinkela_wire_517;
    wire jinkela_wire_518;
    wire jinkela_wire_519;
    wire jinkela_wire_520;
    wire jinkela_wire_521;
    wire jinkela_wire_522;
    wire jinkela_wire_523;
    wire jinkela_wire_524;
    wire jinkela_wire_525;
    wire jinkela_wire_526;
    wire jinkela_wire_527;
    wire jinkela_wire_528;
    wire jinkela_wire_529;
    wire jinkela_wire_530;
    wire jinkela_wire_531;
    wire jinkela_wire_532;
    wire jinkela_wire_533;
    wire jinkela_wire_534;
    wire jinkela_wire_535;
    wire jinkela_wire_536;
    wire jinkela_wire_537;
    wire jinkela_wire_538;
    wire jinkela_wire_539;
    wire jinkela_wire_540;
    wire jinkela_wire_541;
    wire jinkela_wire_542;
    wire jinkela_wire_543;
    wire jinkela_wire_544;
    wire jinkela_wire_545;
    wire jinkela_wire_546;
    wire jinkela_wire_547;
    wire jinkela_wire_548;
    wire jinkela_wire_549;
    wire jinkela_wire_550;
    wire jinkela_wire_551;
    wire jinkela_wire_552;
    wire jinkela_wire_553;
    wire jinkela_wire_554;
    wire jinkela_wire_555;
    wire jinkela_wire_556;
    wire jinkela_wire_557;
    wire jinkela_wire_558;
    wire jinkela_wire_559;
    wire jinkela_wire_560;
    wire jinkela_wire_561;
    wire jinkela_wire_562;
    wire jinkela_wire_563;
    wire jinkela_wire_564;
    wire jinkela_wire_565;
    wire jinkela_wire_566;
    wire jinkela_wire_567;
    wire jinkela_wire_568;
    wire jinkela_wire_569;
    wire jinkela_wire_570;
    wire jinkela_wire_571;
    wire jinkela_wire_572;
    wire jinkela_wire_573;
    wire jinkela_wire_574;
    wire jinkela_wire_575;
    wire jinkela_wire_576;
    wire jinkela_wire_577;
    wire jinkela_wire_578;
    wire jinkela_wire_579;
    wire jinkela_wire_580;
    wire jinkela_wire_581;
    wire jinkela_wire_582;
    wire jinkela_wire_583;
    wire jinkela_wire_584;
    wire jinkela_wire_585;
    wire jinkela_wire_586;
    wire jinkela_wire_587;
    wire jinkela_wire_588;
    wire jinkela_wire_589;
    wire jinkela_wire_590;
    wire jinkela_wire_591;
    wire jinkela_wire_592;
    wire jinkela_wire_593;
    wire jinkela_wire_594;
    wire jinkela_wire_595;
    wire jinkela_wire_596;
    wire jinkela_wire_597;
    wire jinkela_wire_598;
    wire jinkela_wire_599;
    wire jinkela_wire_600;
    wire jinkela_wire_601;
    wire jinkela_wire_602;
    wire jinkela_wire_603;
    wire jinkela_wire_604;
    wire jinkela_wire_605;
    wire jinkela_wire_606;
    wire jinkela_wire_607;
    wire jinkela_wire_608;
    wire jinkela_wire_609;
    wire jinkela_wire_610;
    wire jinkela_wire_611;
    wire jinkela_wire_612;
    wire jinkela_wire_613;
    wire jinkela_wire_614;
    wire jinkela_wire_615;
    wire jinkela_wire_616;
    wire jinkela_wire_617;
    wire jinkela_wire_618;
    wire jinkela_wire_619;
    wire jinkela_wire_620;
    wire jinkela_wire_621;
    wire jinkela_wire_622;
    wire jinkela_wire_623;
    wire jinkela_wire_624;
    wire jinkela_wire_625;
    wire jinkela_wire_626;
    wire jinkela_wire_627;
    wire jinkela_wire_628;
    wire jinkela_wire_629;
    wire jinkela_wire_630;
    wire jinkela_wire_631;
    wire jinkela_wire_632;
    wire jinkela_wire_633;
    wire jinkela_wire_634;
    wire jinkela_wire_635;
    wire jinkela_wire_636;
    wire jinkela_wire_637;
    wire jinkela_wire_638;
    wire jinkela_wire_639;
    wire jinkela_wire_640;
    wire jinkela_wire_641;
    wire jinkela_wire_642;
    wire jinkela_wire_643;
    wire jinkela_wire_644;
    wire jinkela_wire_645;
    wire jinkela_wire_646;
    wire jinkela_wire_647;
    wire jinkela_wire_648;
    wire jinkela_wire_649;
    wire jinkela_wire_650;
    wire jinkela_wire_651;
    wire jinkela_wire_652;
    wire jinkela_wire_653;
    wire jinkela_wire_654;
    wire jinkela_wire_655;
    wire jinkela_wire_656;
    wire jinkela_wire_657;
    wire jinkela_wire_658;
    wire jinkela_wire_659;
    wire jinkela_wire_660;
    wire jinkela_wire_661;
    wire jinkela_wire_662;
    wire jinkela_wire_663;
    wire jinkela_wire_664;
    wire jinkela_wire_665;
    wire jinkela_wire_666;
    wire jinkela_wire_667;
    wire jinkela_wire_668;
    wire jinkela_wire_669;
    wire jinkela_wire_670;
    wire jinkela_wire_671;
    wire jinkela_wire_672;
    wire jinkela_wire_673;
    wire jinkela_wire_674;
    wire jinkela_wire_675;
    wire jinkela_wire_676;
    wire jinkela_wire_677;
    wire jinkela_wire_678;
    wire jinkela_wire_679;
    wire jinkela_wire_680;
    wire jinkela_wire_681;
    wire jinkela_wire_682;
    wire jinkela_wire_683;
    wire jinkela_wire_684;
    wire jinkela_wire_685;
    wire jinkela_wire_686;
    wire jinkela_wire_687;
    wire jinkela_wire_688;
    wire jinkela_wire_689;
    wire jinkela_wire_690;
    wire jinkela_wire_691;
    wire jinkela_wire_692;
    wire jinkela_wire_693;
    wire jinkela_wire_694;
    wire jinkela_wire_695;
    wire jinkela_wire_696;
    wire jinkela_wire_697;
    wire jinkela_wire_698;
    wire jinkela_wire_699;
    wire jinkela_wire_700;
    wire jinkela_wire_701;
    wire jinkela_wire_702;
    wire jinkela_wire_703;
    wire jinkela_wire_704;
    wire jinkela_wire_705;
    wire jinkela_wire_706;
    wire jinkela_wire_707;
    wire jinkela_wire_708;
    wire jinkela_wire_709;
    wire jinkela_wire_710;
    wire jinkela_wire_711;
    wire jinkela_wire_712;
    wire jinkela_wire_713;
    wire jinkela_wire_714;
    wire jinkela_wire_715;
    wire jinkela_wire_716;
    wire jinkela_wire_717;
    wire jinkela_wire_718;
    wire jinkela_wire_719;
    wire jinkela_wire_720;
    wire jinkela_wire_721;
    wire jinkela_wire_722;
    wire jinkela_wire_723;
    wire jinkela_wire_724;
    wire jinkela_wire_725;
    wire jinkela_wire_726;
    wire jinkela_wire_727;
    wire jinkela_wire_728;
    wire jinkela_wire_729;
    wire jinkela_wire_730;
    wire jinkela_wire_731;
    wire jinkela_wire_732;
    wire jinkela_wire_733;
    wire jinkela_wire_734;
    wire jinkela_wire_735;
    wire jinkela_wire_736;
    wire jinkela_wire_737;
    wire jinkela_wire_738;
    wire jinkela_wire_739;
    wire jinkela_wire_740;
    wire jinkela_wire_741;
    wire jinkela_wire_742;
    wire jinkela_wire_743;
    wire jinkela_wire_744;
    wire jinkela_wire_745;
    wire jinkela_wire_746;
    wire jinkela_wire_747;
    wire jinkela_wire_748;
    wire jinkela_wire_749;
    wire jinkela_wire_750;
    wire jinkela_wire_751;
    wire jinkela_wire_752;
    wire jinkela_wire_753;
    wire jinkela_wire_754;
    wire jinkela_wire_755;
    wire jinkela_wire_756;
    wire jinkela_wire_757;
    wire jinkela_wire_758;
    wire jinkela_wire_759;
    wire jinkela_wire_760;
    wire jinkela_wire_761;
    wire jinkela_wire_762;
    wire jinkela_wire_763;
    wire jinkela_wire_764;
    wire jinkela_wire_765;
    wire jinkela_wire_766;
    wire jinkela_wire_767;
    wire jinkela_wire_768;
    wire jinkela_wire_769;
    wire jinkela_wire_770;
    wire jinkela_wire_771;
    wire jinkela_wire_772;
    wire jinkela_wire_773;
    wire jinkela_wire_774;
    wire jinkela_wire_775;
    wire jinkela_wire_776;
    wire jinkela_wire_777;
    wire jinkela_wire_778;
    wire jinkela_wire_779;
    wire jinkela_wire_780;
    wire jinkela_wire_781;
    wire jinkela_wire_782;
    wire jinkela_wire_783;
    wire jinkela_wire_784;
    wire jinkela_wire_785;
    wire jinkela_wire_786;
    wire jinkela_wire_787;
    wire jinkela_wire_788;
    wire jinkela_wire_789;
    wire jinkela_wire_790;
    wire jinkela_wire_791;
    wire jinkela_wire_792;
    wire jinkela_wire_793;
    wire jinkela_wire_794;
    wire jinkela_wire_795;
    wire jinkela_wire_796;
    wire jinkela_wire_797;
    wire jinkela_wire_798;
    wire jinkela_wire_799;
    wire jinkela_wire_800;
    wire jinkela_wire_801;
    wire jinkela_wire_802;
    wire jinkela_wire_803;
    wire jinkela_wire_804;
    wire jinkela_wire_805;
    wire jinkela_wire_806;
    wire jinkela_wire_807;
    wire jinkela_wire_808;
    wire jinkela_wire_809;
    wire jinkela_wire_810;
    wire jinkela_wire_811;
    wire jinkela_wire_812;
    wire jinkela_wire_813;
    wire jinkela_wire_814;
    wire jinkela_wire_815;
    wire jinkela_wire_816;
    wire jinkela_wire_817;
    wire jinkela_wire_818;
    wire jinkela_wire_819;
    wire jinkela_wire_820;
    wire jinkela_wire_821;
    wire jinkela_wire_822;
    wire jinkela_wire_823;
    wire jinkela_wire_824;
    wire jinkela_wire_825;
    wire jinkela_wire_826;
    wire jinkela_wire_827;
    wire jinkela_wire_828;
    wire jinkela_wire_829;
    wire jinkela_wire_830;
    wire jinkela_wire_831;
    wire jinkela_wire_832;
    wire jinkela_wire_833;
    wire jinkela_wire_834;
    wire jinkela_wire_835;
    wire jinkela_wire_836;
    wire jinkela_wire_837;
    wire jinkela_wire_838;
    wire jinkela_wire_839;
    wire jinkela_wire_840;
    wire jinkela_wire_841;
    wire jinkela_wire_842;
    wire jinkela_wire_843;
    wire jinkela_wire_844;
    wire jinkela_wire_845;
    wire jinkela_wire_846;
    wire jinkela_wire_847;
    wire jinkela_wire_848;
    wire jinkela_wire_849;
    wire jinkela_wire_850;
    wire jinkela_wire_851;
    wire jinkela_wire_852;
    wire jinkela_wire_853;
    wire jinkela_wire_854;
    wire jinkela_wire_855;
    wire jinkela_wire_856;
    wire jinkela_wire_857;
    wire jinkela_wire_858;
    wire jinkela_wire_859;
    wire jinkela_wire_860;
    wire jinkela_wire_861;
    wire jinkela_wire_862;
    wire jinkela_wire_863;
    wire jinkela_wire_864;
    wire jinkela_wire_865;
    wire jinkela_wire_866;
    wire jinkela_wire_867;
    wire jinkela_wire_868;
    wire jinkela_wire_869;
    wire jinkela_wire_870;
    wire jinkela_wire_871;
    wire jinkela_wire_872;
    wire jinkela_wire_873;
    wire jinkela_wire_874;
    wire jinkela_wire_875;
    wire jinkela_wire_876;
    wire jinkela_wire_877;
    wire jinkela_wire_878;
    wire jinkela_wire_879;
    wire jinkela_wire_880;
    wire jinkela_wire_881;
    wire jinkela_wire_882;
    wire jinkela_wire_883;
    wire jinkela_wire_884;
    wire jinkela_wire_885;
    wire jinkela_wire_886;
    wire jinkela_wire_887;
    wire jinkela_wire_888;
    wire jinkela_wire_889;
    wire jinkela_wire_890;
    wire jinkela_wire_891;
    wire jinkela_wire_892;
    wire jinkela_wire_893;
    wire jinkela_wire_894;
    wire jinkela_wire_895;
    wire jinkela_wire_896;
    wire jinkela_wire_897;
    wire jinkela_wire_898;
    wire jinkela_wire_899;
    wire jinkela_wire_900;
    wire jinkela_wire_901;
    wire jinkela_wire_902;
    wire jinkela_wire_903;
    wire jinkela_wire_904;
    wire jinkela_wire_905;
    wire jinkela_wire_906;
    wire jinkela_wire_907;
    wire jinkela_wire_908;
    wire jinkela_wire_909;
    wire jinkela_wire_910;
    wire jinkela_wire_911;
    wire jinkela_wire_912;
    wire jinkela_wire_913;
    wire jinkela_wire_914;
    wire jinkela_wire_915;
    wire jinkela_wire_916;
    wire jinkela_wire_917;
    wire jinkela_wire_918;
    wire jinkela_wire_919;
    wire jinkela_wire_920;
    wire jinkela_wire_921;
    wire jinkela_wire_922;
    wire jinkela_wire_923;
    wire jinkela_wire_924;
    wire jinkela_wire_925;
    wire jinkela_wire_926;
    wire jinkela_wire_927;
    wire jinkela_wire_928;
    wire jinkela_wire_929;
    wire jinkela_wire_930;
    wire jinkela_wire_931;
    wire jinkela_wire_932;
    wire jinkela_wire_933;
    wire jinkela_wire_934;
    wire jinkela_wire_935;
    wire jinkela_wire_936;
    wire jinkela_wire_937;
    wire jinkela_wire_938;
    wire jinkela_wire_939;
    wire jinkela_wire_940;
    wire jinkela_wire_941;
    wire jinkela_wire_942;
    wire jinkela_wire_943;
    wire jinkela_wire_944;
    wire jinkela_wire_945;
    wire jinkela_wire_946;
    wire jinkela_wire_947;
    wire jinkela_wire_948;
    wire jinkela_wire_949;
    wire jinkela_wire_950;
    wire jinkela_wire_951;
    wire jinkela_wire_952;
    wire jinkela_wire_953;
    wire jinkela_wire_954;
    wire jinkela_wire_955;
    wire jinkela_wire_956;
    wire jinkela_wire_957;
    wire jinkela_wire_958;
    wire jinkela_wire_959;
    wire jinkela_wire_960;
    wire jinkela_wire_961;
    wire jinkela_wire_962;
    wire jinkela_wire_963;
    wire jinkela_wire_964;
    wire jinkela_wire_965;
    wire jinkela_wire_966;
    wire jinkela_wire_967;
    wire jinkela_wire_968;
    wire jinkela_wire_969;
    wire jinkela_wire_970;
    wire jinkela_wire_971;
    wire jinkela_wire_972;
    wire jinkela_wire_973;
    wire jinkela_wire_974;
    wire jinkela_wire_975;
    wire jinkela_wire_976;
    wire jinkela_wire_977;
    wire jinkela_wire_978;
    wire jinkela_wire_979;
    wire jinkela_wire_980;
    wire jinkela_wire_981;
    wire jinkela_wire_982;
    wire jinkela_wire_983;
    wire jinkela_wire_984;
    wire jinkela_wire_985;
    wire jinkela_wire_986;
    wire jinkela_wire_987;
    wire jinkela_wire_988;
    wire jinkela_wire_989;
    wire jinkela_wire_990;
    wire jinkela_wire_991;
    wire jinkela_wire_992;
    wire jinkela_wire_993;
    wire jinkela_wire_994;
    wire jinkela_wire_995;
    wire jinkela_wire_996;
    wire jinkela_wire_997;
    wire jinkela_wire_998;
    wire jinkela_wire_999;
    wire jinkela_wire_1000;
    wire jinkela_wire_1001;
    wire jinkela_wire_1002;
    wire jinkela_wire_1003;
    wire jinkela_wire_1004;
    wire jinkela_wire_1005;
    wire jinkela_wire_1006;
    wire jinkela_wire_1007;
    wire jinkela_wire_1008;
    wire jinkela_wire_1009;
    wire jinkela_wire_1010;
    wire jinkela_wire_1011;
    wire jinkela_wire_1012;
    wire jinkela_wire_1013;
    wire jinkela_wire_1014;
    wire jinkela_wire_1015;
    wire jinkela_wire_1016;
    wire jinkela_wire_1017;
    wire jinkela_wire_1018;
    wire jinkela_wire_1019;
    wire jinkela_wire_1020;
    wire jinkela_wire_1021;
    wire jinkela_wire_1022;
    wire jinkela_wire_1023;
    wire jinkela_wire_1024;
    wire jinkela_wire_1025;
    wire jinkela_wire_1026;
    wire jinkela_wire_1027;
    wire jinkela_wire_1028;
    wire jinkela_wire_1029;
    wire jinkela_wire_1030;
    wire jinkela_wire_1031;
    wire jinkela_wire_1032;
    wire jinkela_wire_1033;
    wire jinkela_wire_1034;
    wire jinkela_wire_1035;
    wire jinkela_wire_1036;
    wire jinkela_wire_1037;
    wire jinkela_wire_1038;
    wire jinkela_wire_1039;
    wire jinkela_wire_1040;
    wire jinkela_wire_1041;
    wire jinkela_wire_1042;
    wire jinkela_wire_1043;
    wire jinkela_wire_1044;
    wire jinkela_wire_1045;
    wire jinkela_wire_1046;
    wire jinkela_wire_1047;
    wire jinkela_wire_1048;
    wire jinkela_wire_1049;
    wire jinkela_wire_1050;
    wire jinkela_wire_1051;
    wire jinkela_wire_1052;
    wire jinkela_wire_1053;
    wire jinkela_wire_1054;
    wire jinkela_wire_1055;
    wire jinkela_wire_1056;
    wire jinkela_wire_1057;
    wire jinkela_wire_1058;
    wire jinkela_wire_1059;
    wire jinkela_wire_1060;
    wire jinkela_wire_1061;
    wire jinkela_wire_1062;
    wire jinkela_wire_1063;
    wire jinkela_wire_1064;
    wire jinkela_wire_1065;
    wire jinkela_wire_1066;
    wire jinkela_wire_1067;
    wire jinkela_wire_1068;
    wire jinkela_wire_1069;
    wire jinkela_wire_1070;
    wire jinkela_wire_1071;
    wire jinkela_wire_1072;
    wire jinkela_wire_1073;
    wire jinkela_wire_1074;
    wire jinkela_wire_1075;
    wire jinkela_wire_1076;
    wire jinkela_wire_1077;
    wire jinkela_wire_1078;
    wire jinkela_wire_1079;
    wire jinkela_wire_1080;
    wire jinkela_wire_1081;
    wire jinkela_wire_1082;
    wire jinkela_wire_1083;
    wire jinkela_wire_1084;
    wire jinkela_wire_1085;
    wire jinkela_wire_1086;
    wire jinkela_wire_1087;
    wire jinkela_wire_1088;
    wire jinkela_wire_1089;
    wire jinkela_wire_1090;
    wire jinkela_wire_1091;
    wire jinkela_wire_1092;
    wire jinkela_wire_1093;
    wire jinkela_wire_1094;
    wire jinkela_wire_1095;
    wire jinkela_wire_1096;
    wire jinkela_wire_1097;
    wire jinkela_wire_1098;
    wire jinkela_wire_1099;
    wire jinkela_wire_1100;
    wire jinkela_wire_1101;
    wire jinkela_wire_1102;
    wire jinkela_wire_1103;
    wire jinkela_wire_1104;
    wire jinkela_wire_1105;
    wire jinkela_wire_1106;
    wire jinkela_wire_1107;
    wire jinkela_wire_1108;
    wire jinkela_wire_1109;
    wire jinkela_wire_1110;
    wire jinkela_wire_1111;
    wire jinkela_wire_1112;
    wire jinkela_wire_1113;
    wire jinkela_wire_1114;
    wire jinkela_wire_1115;
    wire jinkela_wire_1116;
    wire jinkela_wire_1117;
    wire jinkela_wire_1118;
    wire jinkela_wire_1119;
    wire jinkela_wire_1120;
    wire jinkela_wire_1121;
    wire jinkela_wire_1122;
    wire jinkela_wire_1123;
    wire jinkela_wire_1124;
    wire jinkela_wire_1125;
    wire jinkela_wire_1126;
    wire jinkela_wire_1127;
    wire jinkela_wire_1128;
    wire jinkela_wire_1129;
    wire jinkela_wire_1130;
    wire jinkela_wire_1131;
    wire jinkela_wire_1132;
    wire jinkela_wire_1133;
    wire jinkela_wire_1134;
    wire jinkela_wire_1135;
    wire jinkela_wire_1136;
    wire jinkela_wire_1137;
    wire jinkela_wire_1138;
    wire jinkela_wire_1139;
    wire jinkela_wire_1140;
    wire jinkela_wire_1141;
    wire jinkela_wire_1142;
    wire jinkela_wire_1143;
    wire jinkela_wire_1144;
    wire jinkela_wire_1145;
    wire jinkela_wire_1146;
    wire jinkela_wire_1147;
    wire jinkela_wire_1148;
    wire jinkela_wire_1149;
    wire jinkela_wire_1150;
    wire jinkela_wire_1151;
    wire jinkela_wire_1152;
    wire jinkela_wire_1153;
    wire jinkela_wire_1154;
    wire jinkela_wire_1155;
    wire jinkela_wire_1156;
    wire jinkela_wire_1157;
    wire jinkela_wire_1158;
    wire jinkela_wire_1159;
    wire jinkela_wire_1160;
    wire jinkela_wire_1161;
    wire jinkela_wire_1162;
    wire jinkela_wire_1163;
    wire jinkela_wire_1164;
    wire jinkela_wire_1165;
    wire jinkela_wire_1166;
    wire jinkela_wire_1167;
    wire jinkela_wire_1168;
    wire jinkela_wire_1169;
    wire jinkela_wire_1170;
    wire jinkela_wire_1171;
    wire jinkela_wire_1172;
    wire jinkela_wire_1173;
    wire jinkela_wire_1174;
    wire jinkela_wire_1175;
    wire jinkela_wire_1176;
    wire jinkela_wire_1177;
    wire jinkela_wire_1178;
    wire jinkela_wire_1179;
    wire jinkela_wire_1180;
    wire jinkela_wire_1181;
    wire jinkela_wire_1182;
    wire jinkela_wire_1183;
    wire jinkela_wire_1184;
    wire jinkela_wire_1185;
    wire jinkela_wire_1186;
    wire jinkela_wire_1187;
    wire jinkela_wire_1188;
    wire jinkela_wire_1189;
    wire jinkela_wire_1190;
    wire jinkela_wire_1191;
    wire jinkela_wire_1192;
    wire jinkela_wire_1193;
    wire jinkela_wire_1194;
    wire jinkela_wire_1195;
    wire jinkela_wire_1196;
    wire jinkela_wire_1197;
    wire jinkela_wire_1198;
    wire jinkela_wire_1199;
    wire jinkela_wire_1200;
    wire jinkela_wire_1201;
    wire jinkela_wire_1202;
    wire jinkela_wire_1203;
    wire jinkela_wire_1204;
    wire jinkela_wire_1205;
    wire jinkela_wire_1206;
    wire jinkela_wire_1207;
    wire jinkela_wire_1208;
    wire jinkela_wire_1209;
    wire jinkela_wire_1210;
    wire jinkela_wire_1211;
    wire jinkela_wire_1212;
    wire jinkela_wire_1213;
    wire jinkela_wire_1214;
    wire jinkela_wire_1215;
    wire jinkela_wire_1216;
    wire jinkela_wire_1217;
    wire jinkela_wire_1218;
    wire jinkela_wire_1219;
    wire jinkela_wire_1220;
    wire jinkela_wire_1221;
    wire jinkela_wire_1222;
    wire jinkela_wire_1223;
    wire jinkela_wire_1224;
    wire jinkela_wire_1225;
    wire jinkela_wire_1226;
    wire jinkela_wire_1227;
    wire jinkela_wire_1228;
    wire jinkela_wire_1229;
    wire jinkela_wire_1230;
    wire jinkela_wire_1231;
    wire jinkela_wire_1232;
    wire jinkela_wire_1233;
    wire jinkela_wire_1234;
    wire jinkela_wire_1235;
    wire jinkela_wire_1236;
    wire jinkela_wire_1237;
    wire jinkela_wire_1238;
    wire jinkela_wire_1239;
    wire jinkela_wire_1240;
    wire jinkela_wire_1241;
    wire jinkela_wire_1242;
    wire jinkela_wire_1243;
    wire jinkela_wire_1244;
    wire jinkela_wire_1245;
    wire jinkela_wire_1246;
    wire jinkela_wire_1247;
    wire jinkela_wire_1248;
    wire jinkela_wire_1249;
    wire jinkela_wire_1250;
    wire jinkela_wire_1251;
    wire jinkela_wire_1252;
    wire jinkela_wire_1253;
    wire jinkela_wire_1254;
    wire jinkela_wire_1255;
    wire jinkela_wire_1256;
    wire jinkela_wire_1257;
    wire jinkela_wire_1258;
    wire jinkela_wire_1259;
    wire jinkela_wire_1260;
    wire jinkela_wire_1261;
    wire jinkela_wire_1262;
    wire jinkela_wire_1263;
    wire jinkela_wire_1264;
    wire jinkela_wire_1265;
    wire jinkela_wire_1266;
    wire jinkela_wire_1267;
    wire jinkela_wire_1268;
    wire jinkela_wire_1269;
    wire jinkela_wire_1270;
    wire jinkela_wire_1271;
    wire jinkela_wire_1272;
    wire jinkela_wire_1273;
    wire jinkela_wire_1274;
    wire jinkela_wire_1275;
    wire jinkela_wire_1276;
    wire jinkela_wire_1277;
    wire jinkela_wire_1278;
    wire jinkela_wire_1279;
    wire jinkela_wire_1280;
    wire jinkela_wire_1281;
    wire jinkela_wire_1282;
    wire jinkela_wire_1283;
    wire jinkela_wire_1284;
    wire jinkela_wire_1285;
    wire jinkela_wire_1286;
    wire jinkela_wire_1287;
    wire jinkela_wire_1288;
    wire jinkela_wire_1289;
    wire jinkela_wire_1290;
    wire jinkela_wire_1291;
    wire jinkela_wire_1292;
    wire jinkela_wire_1293;
    wire jinkela_wire_1294;
    wire jinkela_wire_1295;
    wire jinkela_wire_1296;
    wire jinkela_wire_1297;
    wire jinkela_wire_1298;
    wire jinkela_wire_1299;
    wire jinkela_wire_1300;
    wire jinkela_wire_1301;
    wire jinkela_wire_1302;
    wire jinkela_wire_1303;
    wire jinkela_wire_1304;
    wire jinkela_wire_1305;
    wire jinkela_wire_1306;
    wire jinkela_wire_1307;
    wire jinkela_wire_1308;
    wire jinkela_wire_1309;
    wire jinkela_wire_1310;
    wire jinkela_wire_1311;
    wire jinkela_wire_1312;
    wire jinkela_wire_1313;
    wire jinkela_wire_1314;
    wire jinkela_wire_1315;
    wire jinkela_wire_1316;
    wire jinkela_wire_1317;
    wire jinkela_wire_1318;
    wire jinkela_wire_1319;
    wire jinkela_wire_1320;
    wire jinkela_wire_1321;
    wire jinkela_wire_1322;
    wire jinkela_wire_1323;
    wire jinkela_wire_1324;
    wire jinkela_wire_1325;
    wire jinkela_wire_1326;
    wire jinkela_wire_1327;
    wire jinkela_wire_1328;
    wire jinkela_wire_1329;
    wire jinkela_wire_1330;
    wire jinkela_wire_1331;
    wire jinkela_wire_1332;
    wire jinkela_wire_1333;
    wire jinkela_wire_1334;
    wire jinkela_wire_1335;
    wire jinkela_wire_1336;
    wire jinkela_wire_1337;
    wire jinkela_wire_1338;
    wire jinkela_wire_1339;
    wire jinkela_wire_1340;
    wire jinkela_wire_1341;
    wire jinkela_wire_1342;
    wire jinkela_wire_1343;
    wire jinkela_wire_1344;
    wire jinkela_wire_1345;
    wire jinkela_wire_1346;
    wire jinkela_wire_1347;
    wire jinkela_wire_1348;
    wire jinkela_wire_1349;
    wire jinkela_wire_1350;
    wire jinkela_wire_1351;
    wire jinkela_wire_1352;
    wire jinkela_wire_1353;
    wire jinkela_wire_1354;
    wire jinkela_wire_1355;
    wire jinkela_wire_1356;
    wire jinkela_wire_1357;
    wire jinkela_wire_1358;
    wire jinkela_wire_1359;
    wire jinkela_wire_1360;
    wire jinkela_wire_1361;
    wire jinkela_wire_1362;
    wire jinkela_wire_1363;
    wire jinkela_wire_1364;
    wire jinkela_wire_1365;
    wire jinkela_wire_1366;
    wire jinkela_wire_1367;
    wire jinkela_wire_1368;
    wire jinkela_wire_1369;
    wire jinkela_wire_1370;
    wire jinkela_wire_1371;
    wire jinkela_wire_1372;
    wire jinkela_wire_1373;
    wire jinkela_wire_1374;
    wire jinkela_wire_1375;
    wire jinkela_wire_1376;
    wire jinkela_wire_1377;
    wire jinkela_wire_1378;
    wire jinkela_wire_1379;
    wire jinkela_wire_1380;
    wire jinkela_wire_1381;
    wire jinkela_wire_1382;
    wire jinkela_wire_1383;
    wire jinkela_wire_1384;
    wire jinkela_wire_1385;
    wire jinkela_wire_1386;
    wire jinkela_wire_1387;
    wire jinkela_wire_1388;
    wire jinkela_wire_1389;
    wire jinkela_wire_1390;
    wire jinkela_wire_1391;
    wire jinkela_wire_1392;
    wire jinkela_wire_1393;
    wire jinkela_wire_1394;
    wire jinkela_wire_1395;
    wire jinkela_wire_1396;
    wire jinkela_wire_1397;
    wire jinkela_wire_1398;
    wire jinkela_wire_1399;
    wire jinkela_wire_1400;
    wire jinkela_wire_1401;
    wire jinkela_wire_1402;
    wire jinkela_wire_1403;
    wire jinkela_wire_1404;
    wire jinkela_wire_1405;
    wire jinkela_wire_1406;
    wire jinkela_wire_1407;
    wire jinkela_wire_1408;
    wire jinkela_wire_1409;
    wire jinkela_wire_1410;
    wire jinkela_wire_1411;
    wire jinkela_wire_1412;
    wire jinkela_wire_1413;
    wire jinkela_wire_1414;
    wire jinkela_wire_1415;
    wire jinkela_wire_1416;
    wire jinkela_wire_1417;
    wire jinkela_wire_1418;
    wire jinkela_wire_1419;
    wire jinkela_wire_1420;
    wire jinkela_wire_1421;
    wire jinkela_wire_1422;
    wire jinkela_wire_1423;
    wire jinkela_wire_1424;
    wire jinkela_wire_1425;
    wire jinkela_wire_1426;
    wire jinkela_wire_1427;
    wire jinkela_wire_1428;
    wire jinkela_wire_1429;
    wire jinkela_wire_1430;
    wire jinkela_wire_1431;
    wire jinkela_wire_1432;
    wire jinkela_wire_1433;
    wire jinkela_wire_1434;
    wire jinkela_wire_1435;
    wire jinkela_wire_1436;
    wire jinkela_wire_1437;
    wire jinkela_wire_1438;
    wire jinkela_wire_1439;
    wire jinkela_wire_1440;
    wire jinkela_wire_1441;
    wire jinkela_wire_1442;
    wire jinkela_wire_1443;
    wire jinkela_wire_1444;
    wire jinkela_wire_1445;
    wire jinkela_wire_1446;
    wire jinkela_wire_1447;
    wire jinkela_wire_1448;
    wire jinkela_wire_1449;
    wire jinkela_wire_1450;
    wire jinkela_wire_1451;
    wire jinkela_wire_1452;
    wire jinkela_wire_1453;
    wire jinkela_wire_1454;
    wire jinkela_wire_1455;
    wire jinkela_wire_1456;
    wire jinkela_wire_1457;
    wire jinkela_wire_1458;
    wire jinkela_wire_1459;
    wire jinkela_wire_1460;
    wire jinkela_wire_1461;
    wire jinkela_wire_1462;
    wire jinkela_wire_1463;
    wire jinkela_wire_1464;
    wire jinkela_wire_1465;
    wire jinkela_wire_1466;
    wire jinkela_wire_1467;
    wire jinkela_wire_1468;
    wire jinkela_wire_1469;
    wire jinkela_wire_1470;
    wire jinkela_wire_1471;
    wire jinkela_wire_1472;
    wire jinkela_wire_1473;
    wire jinkela_wire_1474;
    wire jinkela_wire_1475;
    wire jinkela_wire_1476;
    wire jinkela_wire_1477;
    wire jinkela_wire_1478;
    wire jinkela_wire_1479;
    wire jinkela_wire_1480;
    wire jinkela_wire_1481;
    wire jinkela_wire_1482;
    wire jinkela_wire_1483;
    wire jinkela_wire_1484;
    wire jinkela_wire_1485;
    wire jinkela_wire_1486;
    wire jinkela_wire_1487;
    wire jinkela_wire_1488;
    wire jinkela_wire_1489;
    wire jinkela_wire_1490;
    wire jinkela_wire_1491;
    wire jinkela_wire_1492;
    wire jinkela_wire_1493;
    wire jinkela_wire_1494;
    wire jinkela_wire_1495;
    wire jinkela_wire_1496;
    wire jinkela_wire_1497;
    wire jinkela_wire_1498;
    wire jinkela_wire_1499;
    wire jinkela_wire_1500;
    wire jinkela_wire_1501;
    wire jinkela_wire_1502;
    wire jinkela_wire_1503;
    wire jinkela_wire_1504;
    wire jinkela_wire_1505;
    wire jinkela_wire_1506;
    wire jinkela_wire_1507;
    wire jinkela_wire_1508;
    wire jinkela_wire_1509;
    wire jinkela_wire_1510;
    wire jinkela_wire_1511;
    wire jinkela_wire_1512;
    wire jinkela_wire_1513;
    wire jinkela_wire_1514;
    wire jinkela_wire_1515;
    wire jinkela_wire_1516;
    wire jinkela_wire_1517;
    input io_in2_1_;
    input io_in1_7_;
    input io_in2_4_;
    input io_in2_16_;
    input io_in1_11_;
    input io_in2_26_;
    input io_fn_0_;
    input io_in2_12_;
    input io_in2_21_;
    input io_in2_14_;
    input io_in1_3_;
    input io_in1_17_;
    input io_in1_20_;
    input io_in1_6_;
    input io_in1_5_;
    input io_in1_18_;
    input io_in2_27_;
    input io_in2_28_;
    input io_in2_25_;
    input io_in1_14_;
    input io_in2_17_;
    input io_in1_25_;
    input io_in1_2_;
    input io_in1_15_;
    input io_in2_22_;
    input io_in1_8_;
    input io_in1_21_;
    input io_in2_23_;
    input io_in1_19_;
    input io_in2_6_;
    input io_in2_9_;
    input io_in2_3_;
    input io_in1_13_;
    input io_in1_23_;
    input io_in2_13_;
    input io_in1_12_;
    input io_in1_0_;
    input io_in2_15_;
    input io_fn_2_;
    input io_in1_28_;
    input io_in2_8_;
    input io_in1_31_;
    input io_in2_0_;
    input io_in2_20_;
    input io_in2_5_;
    input io_in2_29_;
    input io_in2_31_;
    input io_in2_18_;
    input io_in1_16_;
    input io_in1_1_;
    input io_in1_29_;
    input io_in2_24_;
    input io_in2_30_;
    input io_in1_9_;
    input io_in1_30_;
    input io_in2_19_;
    input io_in2_7_;
    input io_in2_2_;
    input io_in1_27_;
    input io_in2_11_;
    input io_in1_24_;
    input io_fn_3_;
    input io_in2_10_;
    input io_fn_1_;
    input io_in1_4_;
    input io_in1_26_;
    input io_in1_10_;
    input io_in1_22_;
    output io_out_22_;
    output io_adder_out_22_;
    output io_out_7_;
    output io_test_adder_Cout;
    output io_adder_out_17_;
    output io_adder_out_26_;
    output io_adder_out_1_;
    output io_adder_out_23_;
    output io_out_1_;
    output io_adder_out_8_;
    output io_adder_out_0_;
    output io_adder_out_7_;
    output io_out_15_;
    output io_out_31_;
    output io_adder_out_10_;
    output io_out_25_;
    output io_out_10_;
    output io_out_14_;
    output io_out_24_;
    output io_adder_out_5_;
    output io_out_12_;
    output io_adder_out_9_;
    output io_adder_out_30_;
    output io_adder_out_12_;
    output io_adder_out_13_;
    output io_out_13_;
    output io_out_21_;
    output io_adder_out_16_;
    output io_out_30_;
    output io_adder_out_2_;
    output io_out_2_;
    output io_adder_out_31_;
    output io_adder_out_14_;
    output io_out_26_;
    output io_out_17_;
    output io_adder_out_6_;
    output io_out_18_;
    output io_out_0_;
    output io_out_4_;
    output io_out_19_;
    output io_adder_out_19_;
    output io_out_23_;
    output io_out_8_;
    output io_adder_out_20_;
    output io_out_20_;
    output io_adder_out_25_;
    output io_adder_out_29_;
    output io_adder_out_15_;
    output io_out_3_;
    output io_out_28_;
    output io_out_27_;
    output io_adder_out_11_;
    output io_out_5_;
    output io_adder_out_4_;
    output io_out_9_;
    output io_adder_out_28_;
    output io_adder_out_21_;
    output io_adder_out_24_;
    output io_out_29_;
    output io_adder_out_27_;
    output io_out_16_;
    output io_out_11_;
    output io_out_6_;
    output io_adder_out_3_;
    output io_adder_out_18_;

    or_bb _2706_ (
        .b(jinkela_wire_718),
        .a(jinkela_wire_936),
        .c(io_out_10_)
    );

    and_bi _2707_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_11_),
        .c(jinkela_wire_1346)
    );

    and_bi _2708_ (
        .b(io_in2_4_),
        .a(jinkela_wire_731),
        .c(jinkela_wire_1097)
    );

    and_bi _2709_ (
        .b(jinkela_wire_1097),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_815)
    );

    and_bi _2710_ (
        .b(jinkela_wire_815),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_1104)
    );

    and_bi _2711_ (
        .b(jinkela_wire_347),
        .a(io_in1_11_),
        .c(jinkela_wire_365)
    );

    and_bi _2712_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_719),
        .c(jinkela_wire_1147)
    );

    and_bi _2713_ (
        .b(jinkela_wire_1147),
        .a(io_in2_11_),
        .c(jinkela_wire_332)
    );

    or_bb _2714_ (
        .b(jinkela_wire_365),
        .a(jinkela_wire_332),
        .c(jinkela_wire_1019)
    );

    and_bi _2715_ (
        .b(jinkela_wire_126),
        .a(jinkela_wire_349),
        .c(jinkela_wire_639)
    );

    and_bb _2716_ (
        .b(jinkela_wire_365),
        .a(jinkela_wire_639),
        .c(jinkela_wire_1202)
    );

    or_bb _2717_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_1202),
        .c(jinkela_wire_824)
    );

    and_bi _2718_ (
        .b(jinkela_wire_824),
        .a(jinkela_wire_1019),
        .c(jinkela_wire_736)
    );

    or_bb _2719_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_736),
        .c(jinkela_wire_1283)
    );

    or_bb _2720_ (
        .b(jinkela_wire_1104),
        .a(jinkela_wire_1283),
        .c(jinkela_wire_691)
    );

    and_bi _2721_ (
        .b(jinkela_wire_1406),
        .a(jinkela_wire_804),
        .c(jinkela_wire_460)
    );

    and_bi _2722_ (
        .b(jinkela_wire_1115),
        .a(io_in2_3_),
        .c(jinkela_wire_886)
    );

    or_bb _2723_ (
        .b(io_in2_4_),
        .a(jinkela_wire_886),
        .c(jinkela_wire_330)
    );

    or_bb _2724_ (
        .b(jinkela_wire_460),
        .a(jinkela_wire_330),
        .c(jinkela_wire_416)
    );

    and_bi _2725_ (
        .b(jinkela_wire_1248),
        .a(jinkela_wire_107),
        .c(jinkela_wire_1362)
    );

    or_bi _2726_ (
        .b(jinkela_wire_416),
        .a(jinkela_wire_1362),
        .c(jinkela_wire_64)
    );

    and_bb _2727_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_64),
        .c(jinkela_wire_997)
    );

    or_bb _2728_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_997),
        .c(jinkela_wire_302)
    );

    and_bi _2729_ (
        .b(jinkela_wire_302),
        .a(jinkela_wire_691),
        .c(jinkela_wire_900)
    );

    or_bb _2730_ (
        .b(jinkela_wire_1346),
        .a(jinkela_wire_900),
        .c(io_out_11_)
    );

    and_bi _2731_ (
        .b(jinkela_wire_1162),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_595)
    );

    and_bi _2732_ (
        .b(jinkela_wire_595),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_340)
    );

    and_bi _2733_ (
        .b(jinkela_wire_340),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_229)
    );

    and_bi _2734_ (
        .b(jinkela_wire_347),
        .a(io_in1_12_),
        .c(jinkela_wire_1120)
    );

    and_bi _2735_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_374),
        .c(jinkela_wire_534)
    );

    and_bi _2736_ (
        .b(jinkela_wire_534),
        .a(io_in2_12_),
        .c(jinkela_wire_671)
    );

    or_bb _2737_ (
        .b(jinkela_wire_1120),
        .a(jinkela_wire_671),
        .c(jinkela_wire_689)
    );

    and_bb _2738_ (
        .b(io_in2_12_),
        .a(jinkela_wire_349),
        .c(jinkela_wire_662)
    );

    and_bb _2739_ (
        .b(jinkela_wire_1120),
        .a(jinkela_wire_662),
        .c(jinkela_wire_116)
    );

    or_bb _2740_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_116),
        .c(jinkela_wire_1223)
    );

    and_bi _2741_ (
        .b(jinkela_wire_1223),
        .a(jinkela_wire_689),
        .c(jinkela_wire_1306)
    );

    or_bb _2742_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1306),
        .c(jinkela_wire_1383)
    );

    or_bb _2743_ (
        .b(jinkela_wire_229),
        .a(jinkela_wire_1383),
        .c(jinkela_wire_57)
    );

    and_bi _2744_ (
        .b(jinkela_wire_757),
        .a(jinkela_wire_804),
        .c(jinkela_wire_721)
    );

    and_bi _2745_ (
        .b(jinkela_wire_376),
        .a(io_in2_3_),
        .c(jinkela_wire_636)
    );

    or_bb _2746_ (
        .b(jinkela_wire_721),
        .a(jinkela_wire_636),
        .c(jinkela_wire_506)
    );

    and_bi _2747_ (
        .b(jinkela_wire_506),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_19)
    );

    and_bi _1989_ (
        .b(io_in1_31_),
        .a(io_in2_31_),
        .c(jinkela_wire_1270)
    );

    and_bi _2535_ (
        .b(jinkela_wire_624),
        .a(jinkela_wire_102),
        .c(jinkela_wire_577)
    );

    or_bb _1990_ (
        .b(jinkela_wire_159),
        .a(jinkela_wire_1270),
        .c(jinkela_wire_344)
    );

    and_bi _2536_ (
        .b(jinkela_wire_577),
        .a(jinkela_wire_804),
        .c(jinkela_wire_1043)
    );

    and_bi _2604_ (
        .b(jinkela_wire_1490),
        .a(jinkela_wire_349),
        .c(jinkela_wire_147)
    );

    or_bi _1991_ (
        .b(io_adder_out_31_),
        .a(jinkela_wire_344),
        .c(jinkela_wire_951)
    );

    and_bi _2537_ (
        .b(jinkela_wire_937),
        .a(jinkela_wire_158),
        .c(jinkela_wire_578)
    );

    or_ii _1992_ (
        .b(io_fn_1_),
        .a(jinkela_wire_1187),
        .c(jinkela_wire_968)
    );

    and_bi _2538_ (
        .b(jinkela_wire_647),
        .a(io_in2_2_),
        .c(jinkela_wire_351)
    );

    or_bb _1993_ (
        .b(jinkela_wire_1270),
        .a(jinkela_wire_968),
        .c(jinkela_wire_1388)
    );

    or_bb _2539_ (
        .b(jinkela_wire_578),
        .a(jinkela_wire_351),
        .c(jinkela_wire_77)
    );

    and_bi _1994_ (
        .b(jinkela_wire_159),
        .a(jinkela_wire_968),
        .c(jinkela_wire_941)
    );

    and_bi _2540_ (
        .b(jinkela_wire_77),
        .a(io_in2_3_),
        .c(jinkela_wire_1090)
    );

    and_bi _1995_ (
        .b(jinkela_wire_941),
        .a(jinkela_wire_1388),
        .c(jinkela_wire_1445)
    );

    or_bb _2541_ (
        .b(jinkela_wire_1043),
        .a(jinkela_wire_1090),
        .c(jinkela_wire_1160)
    );

    and_bi _1996_ (
        .b(jinkela_wire_1445),
        .a(jinkela_wire_951),
        .c(jinkela_wire_488)
    );

    and_bi _2542_ (
        .b(jinkela_wire_1160),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_980)
    );

    and_bi _2605_ (
        .b(jinkela_wire_489),
        .a(jinkela_wire_147),
        .c(jinkela_wire_1242)
    );

    or_bi _1997_ (
        .b(jinkela_wire_1187),
        .a(jinkela_wire_488),
        .c(jinkela_wire_649)
    );

    and_bi _2543_ (
        .b(jinkela_wire_804),
        .a(jinkela_wire_830),
        .c(jinkela_wire_969)
    );

    or_bb _1670_ (
        .b(jinkela_wire_503),
        .a(jinkela_wire_1284),
        .c(jinkela_wire_101)
    );

    and_bi _1998_ (
        .b(io_fn_1_),
        .a(io_fn_0_),
        .c(jinkela_wire_728)
    );

    and_bi _2544_ (
        .b(jinkela_wire_745),
        .a(jinkela_wire_158),
        .c(jinkela_wire_540)
    );

    and_bi _1999_ (
        .b(io_fn_3_),
        .a(io_fn_2_),
        .c(jinkela_wire_527)
    );

    and_bi _2545_ (
        .b(jinkela_wire_1066),
        .a(io_in2_2_),
        .c(jinkela_wire_960)
    );

    or_ii _1671_ (
        .b(jinkela_wire_719),
        .a(jinkela_wire_101),
        .c(jinkela_wire_1326)
    );

    and_bb _2000_ (
        .b(jinkela_wire_728),
        .a(jinkela_wire_527),
        .c(jinkela_wire_1292)
    );

    or_bb _2546_ (
        .b(jinkela_wire_540),
        .a(jinkela_wire_960),
        .c(jinkela_wire_1369)
    );

    and_bi _1669_ (
        .b(jinkela_wire_232),
        .a(jinkela_wire_889),
        .c(jinkela_wire_1284)
    );

    and_bi _2001_ (
        .b(io_fn_2_),
        .a(io_fn_3_),
        .c(jinkela_wire_554)
    );

    and_bi _2547_ (
        .b(jinkela_wire_1369),
        .a(jinkela_wire_804),
        .c(jinkela_wire_1413)
    );

    or_ii _2002_ (
        .b(io_fn_0_),
        .a(io_fn_1_),
        .c(jinkela_wire_305)
    );

    or_bb _2548_ (
        .b(jinkela_wire_969),
        .a(jinkela_wire_1413),
        .c(jinkela_wire_1503)
    );

    and_bi _2003_ (
        .b(jinkela_wire_305),
        .a(jinkela_wire_554),
        .c(jinkela_wire_916)
    );

    and_bi _2549_ (
        .b(jinkela_wire_1503),
        .a(io_in2_4_),
        .c(jinkela_wire_1368)
    );

    or_bb _2004_ (
        .b(jinkela_wire_1292),
        .a(jinkela_wire_916),
        .c(jinkela_wire_188)
    );

    or_bb _2550_ (
        .b(jinkela_wire_980),
        .a(jinkela_wire_1368),
        .c(jinkela_wire_1449)
    );

    inv _2005_ (
        .din(io_in2_4_),
        .dout(jinkela_wire_1248)
    );

    and_bi _2551_ (
        .b(jinkela_wire_1449),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1042)
    );

    or_bb _2606_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_1242),
        .c(jinkela_wire_1444)
    );

    or_bb _2006_ (
        .b(jinkela_wire_268),
        .a(jinkela_wire_188),
        .c(jinkela_wire_589)
    );

    or_bb _2552_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1042),
        .c(jinkela_wire_157)
    );

    and_bi _2007_ (
        .b(jinkela_wire_391),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1141)
    );

    and_bi _2553_ (
        .b(jinkela_wire_157),
        .a(jinkela_wire_981),
        .c(jinkela_wire_1394)
    );

    and_bi _2008_ (
        .b(jinkela_wire_1141),
        .a(jinkela_wire_589),
        .c(jinkela_wire_737)
    );

    or_bb _2554_ (
        .b(jinkela_wire_32),
        .a(jinkela_wire_1394),
        .c(io_out_5_)
    );

    or_bb _2009_ (
        .b(io_in2_0_),
        .a(jinkela_wire_737),
        .c(jinkela_wire_203)
    );

    and_bi _2555_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_6_),
        .c(jinkela_wire_975)
    );

    or_bb _2010_ (
        .b(jinkela_wire_278),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1464)
    );

    and_bi _2556_ (
        .b(jinkela_wire_740),
        .a(jinkela_wire_804),
        .c(jinkela_wire_155)
    );

    and_bi _2011_ (
        .b(jinkela_wire_293),
        .a(jinkela_wire_188),
        .c(jinkela_wire_952)
    );

    and_bi _2557_ (
        .b(jinkela_wire_155),
        .a(jinkela_wire_1269),
        .c(jinkela_wire_883)
    );

    and_bi _2012_ (
        .b(jinkela_wire_952),
        .a(jinkela_wire_1464),
        .c(jinkela_wire_895)
    );

    and_bi _2558_ (
        .b(jinkela_wire_883),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_1150)
    );

    and_bi _2013_ (
        .b(jinkela_wire_895),
        .a(io_in2_0_),
        .c(jinkela_wire_1262)
    );

    and_bi _2559_ (
        .b(jinkela_wire_1150),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_799)
    );

    and_bi _2014_ (
        .b(jinkela_wire_1262),
        .a(jinkela_wire_203),
        .c(jinkela_wire_267)
    );

    and_bi _2560_ (
        .b(jinkela_wire_799),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_1301)
    );

    or_bb _2015_ (
        .b(io_in2_1_),
        .a(jinkela_wire_267),
        .c(jinkela_wire_568)
    );

    and_bb _2561_ (
        .b(io_in2_6_),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_459)
    );

    or_bb _2016_ (
        .b(jinkela_wire_1253),
        .a(jinkela_wire_188),
        .c(jinkela_wire_809)
    );

    or_bb _2562_ (
        .b(io_in1_6_),
        .a(jinkela_wire_459),
        .c(jinkela_wire_1414)
    );

    and_bi _2017_ (
        .b(jinkela_wire_217),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1391)
    );

    and_bb _2563_ (
        .b(io_in1_6_),
        .a(io_in2_6_),
        .c(jinkela_wire_1165)
    );

    and_bi _2018_ (
        .b(jinkela_wire_1391),
        .a(jinkela_wire_809),
        .c(jinkela_wire_202)
    );

    and_bb _2564_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_1165),
        .c(jinkela_wire_1166)
    );

    or_bb _2019_ (
        .b(io_in2_0_),
        .a(jinkela_wire_202),
        .c(jinkela_wire_1067)
    );

    and_bi _2565_ (
        .b(jinkela_wire_1166),
        .a(jinkela_wire_1414),
        .c(jinkela_wire_450)
    );

    or_bb _2020_ (
        .b(jinkela_wire_1329),
        .a(jinkela_wire_188),
        .c(jinkela_wire_913)
    );

    or_bb _2566_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_450),
        .c(jinkela_wire_1048)
    );

    and_bi _2021_ (
        .b(jinkela_wire_719),
        .a(jinkela_wire_188),
        .c(jinkela_wire_16)
    );

    and_bi _2567_ (
        .b(jinkela_wire_1165),
        .a(jinkela_wire_347),
        .c(jinkela_wire_693)
    );

    and_bi _2022_ (
        .b(jinkela_wire_16),
        .a(jinkela_wire_913),
        .c(jinkela_wire_1205)
    );

    or_bb _2568_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_693),
        .c(jinkela_wire_849)
    );

    and_bi _2023_ (
        .b(jinkela_wire_1205),
        .a(io_in2_0_),
        .c(jinkela_wire_52)
    );

    and_bi _2569_ (
        .b(jinkela_wire_849),
        .a(jinkela_wire_1048),
        .c(jinkela_wire_1055)
    );

    and_bi _2024_ (
        .b(jinkela_wire_52),
        .a(jinkela_wire_1067),
        .c(jinkela_wire_1386)
    );

    or_bb _2570_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1055),
        .c(jinkela_wire_328)
    );

    and_bi _2025_ (
        .b(jinkela_wire_1386),
        .a(io_in2_1_),
        .c(jinkela_wire_422)
    );

    or_bb _2571_ (
        .b(jinkela_wire_1301),
        .a(jinkela_wire_328),
        .c(jinkela_wire_290)
    );

    and_bi _2026_ (
        .b(jinkela_wire_422),
        .a(jinkela_wire_568),
        .c(jinkela_wire_976)
    );

    or_bb _2572_ (
        .b(io_in2_2_),
        .a(jinkela_wire_138),
        .c(jinkela_wire_558)
    );

    and_bi _2027_ (
        .b(jinkela_wire_976),
        .a(jinkela_wire_158),
        .c(jinkela_wire_840)
    );

    and_bi _2573_ (
        .b(jinkela_wire_1507),
        .a(io_in2_2_),
        .c(jinkela_wire_424)
    );

    or_bb _2028_ (
        .b(jinkela_wire_842),
        .a(jinkela_wire_188),
        .c(jinkela_wire_25)
    );

    and_bi _2574_ (
        .b(jinkela_wire_424),
        .a(jinkela_wire_558),
        .c(jinkela_wire_989)
    );

    and_bi _2029_ (
        .b(jinkela_wire_374),
        .a(jinkela_wire_188),
        .c(jinkela_wire_132)
    );

    and_bi _2575_ (
        .b(jinkela_wire_989),
        .a(jinkela_wire_804),
        .c(jinkela_wire_377)
    );

    and_bi _2030_ (
        .b(jinkela_wire_132),
        .a(jinkela_wire_25),
        .c(jinkela_wire_911)
    );

    and_bi _2576_ (
        .b(jinkela_wire_457),
        .a(jinkela_wire_158),
        .c(jinkela_wire_531)
    );

    or_bb _1821_ (
        .b(jinkela_wire_1234),
        .a(jinkela_wire_591),
        .c(jinkela_wire_1471)
    );

    or_bb _1822_ (
        .b(jinkela_wire_1424),
        .a(jinkela_wire_1224),
        .c(jinkela_wire_1012)
    );

    or_bb _1823_ (
        .b(io_in2_27_),
        .a(jinkela_wire_1012),
        .c(jinkela_wire_555)
    );

    or_ii _1824_ (
        .b(io_in2_27_),
        .a(jinkela_wire_1012),
        .c(jinkela_wire_313)
    );

    or_ii _1825_ (
        .b(jinkela_wire_555),
        .a(jinkela_wire_313),
        .c(jinkela_wire_255)
    );

    and_bi _1826_ (
        .b(jinkela_wire_255),
        .a(jinkela_wire_1471),
        .c(jinkela_wire_1062)
    );

    and_bi _1827_ (
        .b(jinkela_wire_1062),
        .a(jinkela_wire_61),
        .c(jinkela_wire_1515)
    );

    or_ii _1828_ (
        .b(io_in1_28_),
        .a(jinkela_wire_1515),
        .c(jinkela_wire_227)
    );

    or_bb _1829_ (
        .b(io_in1_28_),
        .a(jinkela_wire_1515),
        .c(jinkela_wire_1196)
    );

    and_bi _1830_ (
        .b(jinkela_wire_1195),
        .a(io_in2_28_),
        .c(jinkela_wire_120)
    );

    or_bb _1831_ (
        .b(jinkela_wire_308),
        .a(jinkela_wire_120),
        .c(jinkela_wire_1491)
    );

    and_bi _1832_ (
        .b(jinkela_wire_1491),
        .a(jinkela_wire_1196),
        .c(jinkela_wire_186)
    );

    and_bi _1833_ (
        .b(jinkela_wire_186),
        .a(jinkela_wire_227),
        .c(jinkela_wire_103)
    );

    and_bi _1834_ (
        .b(io_in1_29_),
        .a(jinkela_wire_103),
        .c(jinkela_wire_281)
    );

    inv _1835_ (
        .din(io_in1_29_),
        .dout(jinkela_wire_1493)
    );

    or_bb _1836_ (
        .b(jinkela_wire_1493),
        .a(jinkela_wire_103),
        .c(jinkela_wire_1364)
    );

    and_bi _1837_ (
        .b(jinkela_wire_262),
        .a(jinkela_wire_1014),
        .c(jinkela_wire_686)
    );

    or_bb _1838_ (
        .b(jinkela_wire_1411),
        .a(jinkela_wire_686),
        .c(jinkela_wire_627)
    );

    inv _1839_ (
        .din(jinkela_wire_627),
        .dout(jinkela_wire_580)
    );

    and_bi _1840_ (
        .b(jinkela_wire_580),
        .a(jinkela_wire_1364),
        .c(jinkela_wire_1129)
    );

    or_bb _1841_ (
        .b(jinkela_wire_281),
        .a(jinkela_wire_1129),
        .c(jinkela_wire_615)
    );

    or_bb _1842_ (
        .b(jinkela_wire_964),
        .a(jinkela_wire_615),
        .c(jinkela_wire_1191)
    );

    and_bi _1843_ (
        .b(io_in1_30_),
        .a(jinkela_wire_615),
        .c(jinkela_wire_546)
    );

    and_bi _1844_ (
        .b(jinkela_wire_559),
        .a(io_in2_30_),
        .c(jinkela_wire_1119)
    );

    and_bi _1845_ (
        .b(io_in2_30_),
        .a(jinkela_wire_559),
        .c(jinkela_wire_1420)
    );

    or_bb _1846_ (
        .b(jinkela_wire_1119),
        .a(jinkela_wire_1420),
        .c(jinkela_wire_1072)
    );

    inv _1847_ (
        .din(jinkela_wire_1072),
        .dout(jinkela_wire_584)
    );

    and_bi _1848_ (
        .b(jinkela_wire_546),
        .a(jinkela_wire_584),
        .c(jinkela_wire_350)
    );

    or_bi _1849_ (
        .b(jinkela_wire_1191),
        .a(jinkela_wire_350),
        .c(jinkela_wire_1339)
    );

    and_bi _1850_ (
        .b(jinkela_wire_80),
        .a(jinkela_wire_1339),
        .c(jinkela_wire_542)
    );

    and_bi _1851_ (
        .b(jinkela_wire_1339),
        .a(jinkela_wire_80),
        .c(jinkela_wire_1243)
    );

    or_bb _1852_ (
        .b(jinkela_wire_542),
        .a(jinkela_wire_1243),
        .c(io_adder_out_31_)
    );

    and_bi _1853_ (
        .b(jinkela_wire_546),
        .a(jinkela_wire_1191),
        .c(jinkela_wire_729)
    );

    or_bb _1854_ (
        .b(jinkela_wire_584),
        .a(jinkela_wire_729),
        .c(jinkela_wire_1221)
    );

    and_bb _1855_ (
        .b(jinkela_wire_1191),
        .a(jinkela_wire_350),
        .c(jinkela_wire_1071)
    );

    and_bi _1856_ (
        .b(jinkela_wire_1071),
        .a(jinkela_wire_1221),
        .c(io_adder_out_30_)
    );

    and_bi _1857_ (
        .b(jinkela_wire_281),
        .a(jinkela_wire_1364),
        .c(jinkela_wire_556)
    );

    and_bi _1858_ (
        .b(jinkela_wire_556),
        .a(jinkela_wire_580),
        .c(jinkela_wire_204)
    );

    and_bi _1859_ (
        .b(jinkela_wire_580),
        .a(jinkela_wire_556),
        .c(jinkela_wire_918)
    );

    or_bb _1860_ (
        .b(jinkela_wire_204),
        .a(jinkela_wire_918),
        .c(io_adder_out_29_)
    );

    and_bb _1861_ (
        .b(jinkela_wire_227),
        .a(jinkela_wire_1196),
        .c(jinkela_wire_312)
    );

    and_bi _1862_ (
        .b(jinkela_wire_312),
        .a(jinkela_wire_1491),
        .c(jinkela_wire_1332)
    );

    or_bb _3084_ (
        .b(jinkela_wire_794),
        .a(jinkela_wire_1289),
        .c(io_out_30_)
    );

    or_bb _1650_ (
        .b(jinkela_wire_609),
        .a(jinkela_wire_199),
        .c(jinkela_wire_837)
    );

    or_bb _2367_ (
        .b(io_in2_2_),
        .a(jinkela_wire_1045),
        .c(jinkela_wire_963)
    );

    and_bi _3085_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_31_),
        .c(jinkela_wire_412)
    );

    and_bi _1651_ (
        .b(io_in1_9_),
        .a(jinkela_wire_837),
        .c(jinkela_wire_264)
    );

    and_bi _2368_ (
        .b(jinkela_wire_963),
        .a(jinkela_wire_335),
        .c(jinkela_wire_1004)
    );

    and_bi _3086_ (
        .b(jinkela_wire_44),
        .a(jinkela_wire_1214),
        .c(jinkela_wire_1181)
    );

    inv _1652_ (
        .din(io_in1_9_),
        .dout(jinkela_wire_293)
    );

    and_bi _2369_ (
        .b(jinkela_wire_18),
        .a(jinkela_wire_15),
        .c(jinkela_wire_1384)
    );

    and_bb _3087_ (
        .b(io_in1_31_),
        .a(io_in2_31_),
        .c(jinkela_wire_1082)
    );

    or_bb _1653_ (
        .b(jinkela_wire_293),
        .a(jinkela_wire_837),
        .c(jinkela_wire_994)
    );

    and_bi _2370_ (
        .b(jinkela_wire_267),
        .a(io_in2_1_),
        .c(jinkela_wire_451)
    );

    and_bi _3088_ (
        .b(jinkela_wire_1082),
        .a(jinkela_wire_347),
        .c(jinkela_wire_1351)
    );

    inv _1654_ (
        .din(io_in2_9_),
        .dout(jinkela_wire_567)
    );

    or_bb _2371_ (
        .b(jinkela_wire_1384),
        .a(jinkela_wire_451),
        .c(jinkela_wire_138)
    );

    and_bi _3089_ (
        .b(jinkela_wire_1351),
        .a(jinkela_wire_44),
        .c(jinkela_wire_1041)
    );

    and_bi _1655_ (
        .b(jinkela_wire_870),
        .a(io_fn_3_),
        .c(jinkela_wire_1111)
    );

    and_bi _2372_ (
        .b(jinkela_wire_138),
        .a(io_in2_2_),
        .c(jinkela_wire_304)
    );

    or_bb _3090_ (
        .b(jinkela_wire_560),
        .a(jinkela_wire_349),
        .c(jinkela_wire_256)
    );

    or_bb _2373_ (
        .b(jinkela_wire_1004),
        .a(jinkela_wire_304),
        .c(jinkela_wire_552)
    );

    and_bi _1656_ (
        .b(jinkela_wire_567),
        .a(jinkela_wire_1111),
        .c(jinkela_wire_418)
    );

    and_bb _3091_ (
        .b(jinkela_wire_1270),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_524)
    );

    and_bi _2374_ (
        .b(jinkela_wire_552),
        .a(jinkela_wire_804),
        .c(jinkela_wire_419)
    );

    and_bi _1657_ (
        .b(jinkela_wire_1111),
        .a(jinkela_wire_567),
        .c(jinkela_wire_942)
    );

    or_bb _3092_ (
        .b(jinkela_wire_159),
        .a(jinkela_wire_524),
        .c(jinkela_wire_714)
    );

    and_bi _2375_ (
        .b(jinkela_wire_1386),
        .a(jinkela_wire_15),
        .c(jinkela_wire_1456)
    );

    or_bb _1658_ (
        .b(jinkela_wire_418),
        .a(jinkela_wire_942),
        .c(jinkela_wire_484)
    );

    and_bi _3093_ (
        .b(jinkela_wire_714),
        .a(jinkela_wire_256),
        .c(jinkela_wire_343)
    );

    and_bi _2376_ (
        .b(jinkela_wire_844),
        .a(io_in2_1_),
        .c(jinkela_wire_600)
    );

    inv _1659_ (
        .din(jinkela_wire_484),
        .dout(jinkela_wire_630)
    );

    and_bi _3094_ (
        .b(jinkela_wire_343),
        .a(jinkela_wire_1041),
        .c(jinkela_wire_608)
    );

    or_bb _2377_ (
        .b(jinkela_wire_1456),
        .a(jinkela_wire_600),
        .c(jinkela_wire_1507)
    );

    and_bi _1660_ (
        .b(jinkela_wire_630),
        .a(jinkela_wire_994),
        .c(jinkela_wire_292)
    );

    or_bb _3095_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_608),
        .c(jinkela_wire_173)
    );

    or_ii _2378_ (
        .b(jinkela_wire_158),
        .a(jinkela_wire_1507),
        .c(jinkela_wire_1081)
    );

    or_bb _1661_ (
        .b(jinkela_wire_264),
        .a(jinkela_wire_292),
        .c(jinkela_wire_587)
    );

    or_bb _3096_ (
        .b(jinkela_wire_1181),
        .a(jinkela_wire_173),
        .c(jinkela_wire_528)
    );

    or_bb _2379_ (
        .b(io_in2_1_),
        .a(jinkela_wire_1152),
        .c(jinkela_wire_863)
    );

    and_bi _1662_ (
        .b(io_in1_10_),
        .a(jinkela_wire_587),
        .c(jinkela_wire_503)
    );

    and_bb _3097_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1341),
        .c(jinkela_wire_1037)
    );

    and_bi _2380_ (
        .b(jinkela_wire_45),
        .a(io_in2_1_),
        .c(jinkela_wire_645)
    );

    inv _1663_ (
        .din(io_in1_10_),
        .dout(jinkela_wire_217)
    );

    or_bb _3098_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1037),
        .c(jinkela_wire_1358)
    );

    and_bi _2381_ (
        .b(jinkela_wire_645),
        .a(jinkela_wire_863),
        .c(jinkela_wire_457)
    );

    or_bb _1664_ (
        .b(jinkela_wire_217),
        .a(jinkela_wire_587),
        .c(jinkela_wire_889)
    );

    and_bi _3099_ (
        .b(jinkela_wire_1358),
        .a(jinkela_wire_528),
        .c(jinkela_wire_827)
    );

    and_bi _2382_ (
        .b(jinkela_wire_457),
        .a(io_in2_2_),
        .c(jinkela_wire_908)
    );

    and_bi _1665_ (
        .b(jinkela_wire_667),
        .a(io_fn_3_),
        .c(jinkela_wire_1015)
    );

    or_bb _3100_ (
        .b(jinkela_wire_412),
        .a(jinkela_wire_827),
        .c(io_out_31_)
    );

    and_bi _2383_ (
        .b(jinkela_wire_908),
        .a(jinkela_wire_1081),
        .c(jinkela_wire_962)
    );

    and_bi _1666_ (
        .b(io_in2_10_),
        .a(jinkela_wire_1015),
        .c(jinkela_wire_110)
    );

    and_bi _2384_ (
        .b(jinkela_wire_962),
        .a(io_in2_3_),
        .c(jinkela_wire_196)
    );

    and_bi _1667_ (
        .b(jinkela_wire_1015),
        .a(io_in2_10_),
        .c(jinkela_wire_283)
    );

    or_bb _2385_ (
        .b(io_in2_4_),
        .a(jinkela_wire_196),
        .c(jinkela_wire_547)
    );

    or_bb _1668_ (
        .b(jinkela_wire_110),
        .a(jinkela_wire_283),
        .c(jinkela_wire_232)
    );

    or_bb _2386_ (
        .b(jinkela_wire_419),
        .a(jinkela_wire_547),
        .c(jinkela_wire_910)
    );

    or_bb _1672_ (
        .b(jinkela_wire_719),
        .a(jinkela_wire_101),
        .c(jinkela_wire_153)
    );

    or_bb _2387_ (
        .b(io_in2_1_),
        .a(jinkela_wire_1077),
        .c(jinkela_wire_797)
    );

    and_bi _1673_ (
        .b(jinkela_wire_652),
        .a(io_fn_3_),
        .c(jinkela_wire_835)
    );

    and_bi _2388_ (
        .b(jinkela_wire_735),
        .a(io_in2_1_),
        .c(jinkela_wire_384)
    );

    or_ii _1674_ (
        .b(io_in2_11_),
        .a(jinkela_wire_835),
        .c(jinkela_wire_51)
    );

    and_bi _2389_ (
        .b(jinkela_wire_384),
        .a(jinkela_wire_797),
        .c(jinkela_wire_1099)
    );

    inv _1675_ (
        .din(io_in2_11_),
        .dout(jinkela_wire_126)
    );

    or_bb _2390_ (
        .b(io_in2_2_),
        .a(jinkela_wire_1099),
        .c(jinkela_wire_20)
    );

    and_bi _1676_ (
        .b(jinkela_wire_835),
        .a(jinkela_wire_126),
        .c(jinkela_wire_1201)
    );

    or_bb _2391_ (
        .b(io_in2_1_),
        .a(jinkela_wire_10),
        .c(jinkela_wire_663)
    );

    and_bi _1677_ (
        .b(jinkela_wire_1201),
        .a(jinkela_wire_51),
        .c(jinkela_wire_1177)
    );

    and_bi _2392_ (
        .b(jinkela_wire_1052),
        .a(io_in2_1_),
        .c(jinkela_wire_1059)
    );

    and_bi _1678_ (
        .b(jinkela_wire_1177),
        .a(jinkela_wire_153),
        .c(jinkela_wire_993)
    );

    and_bi _2393_ (
        .b(jinkela_wire_1059),
        .a(jinkela_wire_663),
        .c(jinkela_wire_144)
    );

    or_bi _1679_ (
        .b(jinkela_wire_1326),
        .a(jinkela_wire_993),
        .c(jinkela_wire_383)
    );

    and_bi _2394_ (
        .b(jinkela_wire_144),
        .a(io_in2_2_),
        .c(jinkela_wire_465)
    );

    and_bi _1680_ (
        .b(io_in1_12_),
        .a(jinkela_wire_383),
        .c(jinkela_wire_1506)
    );

    and_bi _2395_ (
        .b(jinkela_wire_465),
        .a(jinkela_wire_20),
        .c(jinkela_wire_998)
    );

    inv _1681_ (
        .din(io_in1_12_),
        .dout(jinkela_wire_374)
    );

    and_bi _2396_ (
        .b(jinkela_wire_998),
        .a(jinkela_wire_804),
        .c(jinkela_wire_249)
    );

    or_bb _1682_ (
        .b(jinkela_wire_374),
        .a(jinkela_wire_383),
        .c(jinkela_wire_669)
    );

    and_bi _2397_ (
        .b(jinkela_wire_158),
        .a(jinkela_wire_588),
        .c(jinkela_wire_1308)
    );

    and_bi _1683_ (
        .b(jinkela_wire_598),
        .a(io_fn_3_),
        .c(jinkela_wire_1033)
    );

    and_bi _2398_ (
        .b(jinkela_wire_572),
        .a(jinkela_wire_15),
        .c(jinkela_wire_1484)
    );

    and_bi _1684_ (
        .b(io_in2_12_),
        .a(jinkela_wire_1033),
        .c(jinkela_wire_1344)
    );

    and_bi _2399_ (
        .b(jinkela_wire_922),
        .a(io_in2_1_),
        .c(jinkela_wire_1451)
    );

    and_bi _1685_ (
        .b(jinkela_wire_1033),
        .a(io_in2_12_),
        .c(jinkela_wire_1235)
    );

    or_bb _2400_ (
        .b(jinkela_wire_1484),
        .a(jinkela_wire_1451),
        .c(jinkela_wire_944)
    );

    or_bb _1686_ (
        .b(jinkela_wire_1344),
        .a(jinkela_wire_1235),
        .c(jinkela_wire_634)
    );

    and_bi _2401_ (
        .b(jinkela_wire_944),
        .a(jinkela_wire_158),
        .c(jinkela_wire_463)
    );

    and_bi _1687_ (
        .b(jinkela_wire_634),
        .a(jinkela_wire_669),
        .c(jinkela_wire_323)
    );

    or_bb _2402_ (
        .b(jinkela_wire_1308),
        .a(jinkela_wire_463),
        .c(jinkela_wire_650)
    );

    or_bb _1688_ (
        .b(jinkela_wire_1506),
        .a(jinkela_wire_323),
        .c(jinkela_wire_586)
    );

    and_bi _2403_ (
        .b(jinkela_wire_650),
        .a(io_in2_3_),
        .c(jinkela_wire_1302)
    );

    or_ii _1689_ (
        .b(jinkela_wire_78),
        .a(jinkela_wire_586),
        .c(jinkela_wire_1251)
    );

    or_bb _2404_ (
        .b(jinkela_wire_249),
        .a(jinkela_wire_1302),
        .c(jinkela_wire_930)
    );

    or_bb _1690_ (
        .b(jinkela_wire_78),
        .a(jinkela_wire_586),
        .c(jinkela_wire_1029)
    );

    and_bi _2405_ (
        .b(jinkela_wire_930),
        .a(io_in2_4_),
        .c(jinkela_wire_987)
    );

    and_bi _1691_ (
        .b(jinkela_wire_333),
        .a(io_fn_3_),
        .c(jinkela_wire_337)
    );

    or_bi _2406_ (
        .b(jinkela_wire_910),
        .a(jinkela_wire_987),
        .c(jinkela_wire_68)
    );

    or_ii _1692_ (
        .b(io_in2_13_),
        .a(jinkela_wire_337),
        .c(jinkela_wire_877)
    );

    and_bb _2407_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_68),
        .c(jinkela_wire_368)
    );

    inv _1693_ (
        .din(io_in2_13_),
        .dout(jinkela_wire_1517)
    );

    and_bi _1694_ (
        .b(jinkela_wire_337),
        .a(jinkela_wire_1517),
        .c(jinkela_wire_1005)
    );

    or_bb _2408_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_368),
        .c(jinkela_wire_626)
    );

    and_bi _2916_ (
        .b(jinkela_wire_628),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_817)
    );

    or_bi _2199_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1214),
        .c(jinkela_wire_1423)
    );

    and_bi _2917_ (
        .b(jinkela_wire_244),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_277)
    );

    and_bi _2200_ (
        .b(jinkela_wire_1226),
        .a(jinkela_wire_728),
        .c(jinkela_wire_1131)
    );

    or_bb _2918_ (
        .b(io_in1_21_),
        .a(jinkela_wire_277),
        .c(jinkela_wire_1455)
    );

    inv _2201_ (
        .din(jinkela_wire_1131),
        .dout(jinkela_wire_44)
    );

    and_bb _2919_ (
        .b(io_in1_21_),
        .a(io_in2_21_),
        .c(jinkela_wire_1393)
    );

    and_bi _2202_ (
        .b(jinkela_wire_1405),
        .a(jinkela_wire_1424),
        .c(jinkela_wire_1140)
    );

    and_bb _2920_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_1393),
        .c(jinkela_wire_501)
    );

    or_bi _2203_ (
        .b(jinkela_wire_618),
        .a(jinkela_wire_1140),
        .c(jinkela_wire_1341)
    );

    and_bi _2921_ (
        .b(jinkela_wire_501),
        .a(jinkela_wire_1455),
        .c(jinkela_wire_1396)
    );

    or_bb _2204_ (
        .b(jinkela_wire_44),
        .a(jinkela_wire_1341),
        .c(jinkela_wire_1286)
    );

    or_bb _2922_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_1396),
        .c(jinkela_wire_1313)
    );

    and_bi _2205_ (
        .b(jinkela_wire_1064),
        .a(jinkela_wire_527),
        .c(jinkela_wire_349)
    );

    and_bi _2923_ (
        .b(jinkela_wire_1393),
        .a(jinkela_wire_347),
        .c(jinkela_wire_954)
    );

    and_bb _2206_ (
        .b(jinkela_wire_394),
        .a(jinkela_wire_349),
        .c(jinkela_wire_282)
    );

    or_bb _2924_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_954),
        .c(jinkela_wire_183)
    );

    and_bi _2207_ (
        .b(io_fn_0_),
        .a(jinkela_wire_527),
        .c(jinkela_wire_1345)
    );

    and_bi _2925_ (
        .b(jinkela_wire_183),
        .a(jinkela_wire_1313),
        .c(jinkela_wire_934)
    );

    and_bi _2208_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_1300),
        .c(jinkela_wire_1229)
    );

    or_bb _2926_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_934),
        .c(jinkela_wire_1025)
    );

    and_bi _2209_ (
        .b(jinkela_wire_305),
        .a(jinkela_wire_527),
        .c(jinkela_wire_347)
    );

    or_bb _2927_ (
        .b(jinkela_wire_817),
        .a(jinkela_wire_1025),
        .c(jinkela_wire_407)
    );

    or_bb _2210_ (
        .b(jinkela_wire_276),
        .a(jinkela_wire_347),
        .c(jinkela_wire_1108)
    );

    and_bb _2928_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_770),
        .c(jinkela_wire_1440)
    );

    or_bb _2211_ (
        .b(jinkela_wire_1229),
        .a(jinkela_wire_1108),
        .c(jinkela_wire_874)
    );

    or_bb _2929_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1440),
        .c(jinkela_wire_1401)
    );

    or_bb _2212_ (
        .b(jinkela_wire_282),
        .a(jinkela_wire_874),
        .c(jinkela_wire_130)
    );

    and_bi _2930_ (
        .b(jinkela_wire_1401),
        .a(jinkela_wire_407),
        .c(jinkela_wire_1161)
    );

    and_bi _2213_ (
        .b(jinkela_wire_1192),
        .a(jinkela_wire_347),
        .c(jinkela_wire_1304)
    );

    or_bb _2931_ (
        .b(jinkela_wire_518),
        .a(jinkela_wire_1161),
        .c(io_out_21_)
    );

    and_bi _2214_ (
        .b(jinkela_wire_1304),
        .a(jinkela_wire_130),
        .c(jinkela_wire_726)
    );

    and_bi _2932_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_22_),
        .c(jinkela_wire_91)
    );

    and_bi _2215_ (
        .b(jinkela_wire_726),
        .a(jinkela_wire_44),
        .c(jinkela_wire_129)
    );

    and_bi _2933_ (
        .b(jinkela_wire_21),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_89)
    );

    or_bb _2216_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_129),
        .c(jinkela_wire_738)
    );

    or_bb _2934_ (
        .b(jinkela_wire_278),
        .a(jinkela_wire_347),
        .c(jinkela_wire_177)
    );

    and_bi _2217_ (
        .b(jinkela_wire_738),
        .a(jinkela_wire_1286),
        .c(jinkela_wire_1182)
    );

    inv _2935_ (
        .din(io_in2_22_),
        .dout(jinkela_wire_453)
    );

    or_bb _2218_ (
        .b(jinkela_wire_1187),
        .a(jinkela_wire_1182),
        .c(jinkela_wire_1450)
    );

    and_bi _2936_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_278),
        .c(jinkela_wire_1447)
    );

    and_bi _2219_ (
        .b(jinkela_wire_1450),
        .a(jinkela_wire_1423),
        .c(jinkela_wire_0)
    );

    or_bb _2937_ (
        .b(jinkela_wire_453),
        .a(jinkela_wire_1447),
        .c(jinkela_wire_777)
    );

    or_bi _2220_ (
        .b(jinkela_wire_1389),
        .a(jinkela_wire_0),
        .c(jinkela_wire_242)
    );

    or_ii _2938_ (
        .b(jinkela_wire_177),
        .a(jinkela_wire_777),
        .c(jinkela_wire_1477)
    );

    and_bi _2221_ (
        .b(jinkela_wire_242),
        .a(jinkela_wire_649),
        .c(jinkela_wire_1084)
    );

    and_bi _2939_ (
        .b(jinkela_wire_453),
        .a(jinkela_wire_349),
        .c(jinkela_wire_446)
    );

    and_bi _2222_ (
        .b(jinkela_wire_1084),
        .a(jinkela_wire_1175),
        .c(io_out_0_)
    );

    and_bi _2940_ (
        .b(jinkela_wire_177),
        .a(jinkela_wire_446),
        .c(jinkela_wire_651)
    );

    and_bi _2223_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_1_),
        .c(jinkela_wire_432)
    );

    or_bb _2941_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_651),
        .c(jinkela_wire_415)
    );

    or_ii _2224_ (
        .b(io_fn_3_),
        .a(jinkela_wire_618),
        .c(jinkela_wire_931)
    );

    and_bi _2942_ (
        .b(jinkela_wire_415),
        .a(jinkela_wire_1477),
        .c(jinkela_wire_143)
    );

    and_bi _2225_ (
        .b(jinkela_wire_931),
        .a(io_in2_4_),
        .c(jinkela_wire_369)
    );

    or_bb _2943_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_143),
        .c(jinkela_wire_316)
    );

    inv _2226_ (
        .din(jinkela_wire_369),
        .dout(jinkela_wire_1268)
    );

    or_bb _2944_ (
        .b(jinkela_wire_89),
        .a(jinkela_wire_316),
        .c(jinkela_wire_594)
    );

    or_bb _2227_ (
        .b(jinkela_wire_804),
        .a(jinkela_wire_931),
        .c(jinkela_wire_1269)
    );

    and_bb _2945_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_885),
        .c(jinkela_wire_1068)
    );

    and_bi _2228_ (
        .b(jinkela_wire_931),
        .a(io_in2_2_),
        .c(jinkela_wire_1080)
    );

    or_bb _2946_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1068),
        .c(jinkela_wire_248)
    );

    inv _2229_ (
        .din(jinkela_wire_1080),
        .dout(jinkela_wire_970)
    );

    and_bi _2947_ (
        .b(jinkela_wire_248),
        .a(jinkela_wire_594),
        .c(jinkela_wire_907)
    );

    and_bi _2230_ (
        .b(jinkela_wire_15),
        .a(jinkela_wire_931),
        .c(jinkela_wire_1407)
    );

    or_bb _2948_ (
        .b(jinkela_wire_91),
        .a(jinkela_wire_907),
        .c(io_out_22_)
    );

    and_bi _2231_ (
        .b(jinkela_wire_4),
        .a(jinkela_wire_15),
        .c(jinkela_wire_1212)
    );

    and_bi _2949_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_23_),
        .c(jinkela_wire_852)
    );

    or_bb _2232_ (
        .b(jinkela_wire_1407),
        .a(jinkela_wire_1212),
        .c(jinkela_wire_588)
    );

    and_bi _2950_ (
        .b(jinkela_wire_44),
        .a(jinkela_wire_1366),
        .c(jinkela_wire_700)
    );

    and_bi _2233_ (
        .b(jinkela_wire_588),
        .a(jinkela_wire_158),
        .c(jinkela_wire_1415)
    );

    and_bi _2951_ (
        .b(jinkela_wire_535),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_1492)
    );

    and_bi _2234_ (
        .b(jinkela_wire_1415),
        .a(jinkela_wire_970),
        .c(jinkela_wire_1331)
    );

    or_bb _2952_ (
        .b(io_in1_23_),
        .a(jinkela_wire_1492),
        .c(jinkela_wire_1259)
    );

    and_bi _2235_ (
        .b(jinkela_wire_1331),
        .a(jinkela_wire_804),
        .c(jinkela_wire_140)
    );

    and_bb _2953_ (
        .b(io_in1_23_),
        .a(io_in2_23_),
        .c(jinkela_wire_776)
    );

    and_bi _2236_ (
        .b(jinkela_wire_140),
        .a(jinkela_wire_1269),
        .c(jinkela_wire_98)
    );

    and_bb _2954_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_776),
        .c(jinkela_wire_739)
    );

    and_bi _2237_ (
        .b(jinkela_wire_98),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_440)
    );

    and_bi _2955_ (
        .b(jinkela_wire_739),
        .a(jinkela_wire_1259),
        .c(jinkela_wire_680)
    );

    and_bi _2238_ (
        .b(jinkela_wire_440),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_1499)
    );

    or_bb _2956_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_680),
        .c(jinkela_wire_375)
    );

    and_bi _2239_ (
        .b(jinkela_wire_1499),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_37)
    );

    and_bi _2957_ (
        .b(jinkela_wire_776),
        .a(jinkela_wire_347),
        .c(jinkela_wire_1427)
    );

    and_bi _2240_ (
        .b(jinkela_wire_15),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_213)
    );

    and_bi _2748_ (
        .b(jinkela_wire_752),
        .a(io_in2_4_),
        .c(jinkela_wire_810)
    );

    or_bb _2031_ (
        .b(io_in2_0_),
        .a(jinkela_wire_911),
        .c(jinkela_wire_438)
    );

    or_bb _2749_ (
        .b(jinkela_wire_19),
        .a(jinkela_wire_810),
        .c(jinkela_wire_1296)
    );

    inv _2032_ (
        .din(io_in1_18_),
        .dout(jinkela_wire_865)
    );

    and_bi _2750_ (
        .b(jinkela_wire_1296),
        .a(jinkela_wire_188),
        .c(jinkela_wire_214)
    );

    or_bb _2033_ (
        .b(jinkela_wire_865),
        .a(jinkela_wire_188),
        .c(jinkela_wire_156)
    );

    or_bb _2751_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_214),
        .c(jinkela_wire_1397)
    );

    and_bi _2034_ (
        .b(jinkela_wire_78),
        .a(jinkela_wire_188),
        .c(jinkela_wire_903)
    );

    and_bi _2752_ (
        .b(jinkela_wire_1397),
        .a(jinkela_wire_57),
        .c(jinkela_wire_1102)
    );

    and_bi _2035_ (
        .b(jinkela_wire_903),
        .a(jinkela_wire_156),
        .c(jinkela_wire_772)
    );

    and_bi _2753_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_12_),
        .c(jinkela_wire_1281)
    );

    and_bi _2036_ (
        .b(jinkela_wire_772),
        .a(io_in2_0_),
        .c(jinkela_wire_373)
    );

    or_bb _2754_ (
        .b(jinkela_wire_1102),
        .a(jinkela_wire_1281),
        .c(io_out_12_)
    );

    and_bi _2037_ (
        .b(jinkela_wire_373),
        .a(jinkela_wire_438),
        .c(jinkela_wire_844)
    );

    and_bi _2755_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_13_),
        .c(jinkela_wire_697)
    );

    or_bb _2038_ (
        .b(io_in2_1_),
        .a(jinkela_wire_844),
        .c(jinkela_wire_657)
    );

    and_bi _2756_ (
        .b(io_in2_4_),
        .a(jinkela_wire_930),
        .c(jinkela_wire_677)
    );

    or_bb _2039_ (
        .b(jinkela_wire_899),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1417)
    );

    and_bi _2757_ (
        .b(jinkela_wire_677),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_543)
    );

    and_bi _2040_ (
        .b(jinkela_wire_1073),
        .a(jinkela_wire_188),
        .c(jinkela_wire_362)
    );

    and_bi _2758_ (
        .b(jinkela_wire_543),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_822)
    );

    and_bi _2041_ (
        .b(jinkela_wire_362),
        .a(jinkela_wire_1417),
        .c(jinkela_wire_200)
    );

    or_bb _2759_ (
        .b(jinkela_wire_78),
        .a(jinkela_wire_347),
        .c(jinkela_wire_246)
    );

    or_bb _2042_ (
        .b(io_in2_0_),
        .a(jinkela_wire_200),
        .c(jinkela_wire_798)
    );

    and_bi _2760_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_78),
        .c(jinkela_wire_823)
    );

    inv _2043_ (
        .din(io_in2_0_),
        .dout(jinkela_wire_915)
    );

    or_bb _2761_ (
        .b(jinkela_wire_1517),
        .a(jinkela_wire_823),
        .c(jinkela_wire_352)
    );

    and_bi _2044_ (
        .b(jinkela_wire_188),
        .a(io_in1_16_),
        .c(jinkela_wire_190)
    );

    or_ii _2762_ (
        .b(jinkela_wire_246),
        .a(jinkela_wire_352),
        .c(jinkela_wire_1278)
    );

    and_bi _2045_ (
        .b(jinkela_wire_224),
        .a(jinkela_wire_188),
        .c(jinkela_wire_461)
    );

    and_bi _2763_ (
        .b(jinkela_wire_1517),
        .a(jinkela_wire_349),
        .c(jinkela_wire_683)
    );

    or_bb _2046_ (
        .b(jinkela_wire_190),
        .a(jinkela_wire_461),
        .c(jinkela_wire_288)
    );

    and_bi _2764_ (
        .b(jinkela_wire_246),
        .a(jinkela_wire_683),
        .c(jinkela_wire_1360)
    );

    and_bi _2047_ (
        .b(jinkela_wire_915),
        .a(jinkela_wire_288),
        .c(jinkela_wire_784)
    );

    or_bb _2765_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_1360),
        .c(jinkela_wire_300)
    );

    and_bi _2048_ (
        .b(jinkela_wire_784),
        .a(jinkela_wire_798),
        .c(jinkela_wire_1152)
    );

    and_bi _2766_ (
        .b(jinkela_wire_300),
        .a(jinkela_wire_1278),
        .c(jinkela_wire_602)
    );

    and_bi _2049_ (
        .b(jinkela_wire_1152),
        .a(io_in2_1_),
        .c(jinkela_wire_192)
    );

    or_bb _2767_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_602),
        .c(jinkela_wire_136)
    );

    and_bi _2050_ (
        .b(jinkela_wire_192),
        .a(jinkela_wire_657),
        .c(jinkela_wire_1275)
    );

    or_bb _2768_ (
        .b(jinkela_wire_822),
        .a(jinkela_wire_136),
        .c(jinkela_wire_617)
    );

    and_bi _2051_ (
        .b(jinkela_wire_1275),
        .a(io_in2_2_),
        .c(jinkela_wire_1343)
    );

    and_bi _2769_ (
        .b(jinkela_wire_77),
        .a(jinkela_wire_804),
        .c(jinkela_wire_1267)
    );

    or_bb _2052_ (
        .b(jinkela_wire_840),
        .a(jinkela_wire_1343),
        .c(jinkela_wire_1107)
    );

    and_bi _2770_ (
        .b(jinkela_wire_1369),
        .a(io_in2_3_),
        .c(jinkela_wire_321)
    );

    or_ii _2053_ (
        .b(io_in2_3_),
        .a(jinkela_wire_1107),
        .c(jinkela_wire_467)
    );

    or_bb _2771_ (
        .b(jinkela_wire_1267),
        .a(jinkela_wire_321),
        .c(jinkela_wire_825)
    );

    inv _2054_ (
        .din(io_in2_1_),
        .dout(jinkela_wire_15)
    );

    and_bi _2772_ (
        .b(jinkela_wire_825),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_187)
    );

    or_bb _2055_ (
        .b(jinkela_wire_1234),
        .a(jinkela_wire_188),
        .c(jinkela_wire_401)
    );

    and_bi _2773_ (
        .b(jinkela_wire_1392),
        .a(io_in2_4_),
        .c(jinkela_wire_285)
    );

    and_bi _2056_ (
        .b(jinkela_wire_1174),
        .a(jinkela_wire_188),
        .c(jinkela_wire_881)
    );

    or_bb _2774_ (
        .b(jinkela_wire_187),
        .a(jinkela_wire_285),
        .c(jinkela_wire_1228)
    );

    and_bi _2057_ (
        .b(jinkela_wire_881),
        .a(jinkela_wire_401),
        .c(jinkela_wire_436)
    );

    and_bi _2775_ (
        .b(jinkela_wire_1228),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1317)
    );

    or_bb _2058_ (
        .b(io_in2_0_),
        .a(jinkela_wire_436),
        .c(jinkela_wire_1154)
    );

    or_bb _2776_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1317),
        .c(jinkela_wire_13)
    );

    or_bb _2059_ (
        .b(jinkela_wire_562),
        .a(jinkela_wire_188),
        .c(jinkela_wire_434)
    );

    and_bi _2777_ (
        .b(jinkela_wire_13),
        .a(jinkela_wire_617),
        .c(jinkela_wire_448)
    );

    and_bi _2060_ (
        .b(jinkela_wire_1137),
        .a(jinkela_wire_188),
        .c(jinkela_wire_166)
    );

    or_bb _2778_ (
        .b(jinkela_wire_697),
        .a(jinkela_wire_448),
        .c(io_out_13_)
    );

    and_bi _2061_ (
        .b(jinkela_wire_166),
        .a(jinkela_wire_434),
        .c(jinkela_wire_317)
    );

    and_bi _2779_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_14_),
        .c(jinkela_wire_93)
    );

    and_bi _2062_ (
        .b(jinkela_wire_317),
        .a(io_in2_0_),
        .c(jinkela_wire_341)
    );

    and_bi _2780_ (
        .b(jinkela_wire_456),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_747)
    );

    and_bi _2063_ (
        .b(jinkela_wire_341),
        .a(jinkela_wire_1154),
        .c(jinkela_wire_775)
    );

    and_bi _2781_ (
        .b(jinkela_wire_747),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_991)
    );

    and_bi _2064_ (
        .b(jinkela_wire_775),
        .a(jinkela_wire_15),
        .c(jinkela_wire_1074)
    );

    and_bi _2782_ (
        .b(jinkela_wire_991),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_311)
    );

    or_bb _2065_ (
        .b(jinkela_wire_1241),
        .a(jinkela_wire_188),
        .c(jinkela_wire_470)
    );

    and_bb _2783_ (
        .b(io_in2_14_),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_1425)
    );

    and_bi _2066_ (
        .b(jinkela_wire_561),
        .a(jinkela_wire_188),
        .c(jinkela_wire_135)
    );

    or_bb _2784_ (
        .b(io_in1_14_),
        .a(jinkela_wire_1425),
        .c(jinkela_wire_1060)
    );

    and_bi _2067_ (
        .b(jinkela_wire_135),
        .a(jinkela_wire_470),
        .c(jinkela_wire_236)
    );

    and_bb _2785_ (
        .b(io_in1_14_),
        .a(io_in2_14_),
        .c(jinkela_wire_1121)
    );

    or_bb _2068_ (
        .b(io_in2_0_),
        .a(jinkela_wire_236),
        .c(jinkela_wire_538)
    );

    and_bb _2786_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_1121),
        .c(jinkela_wire_530)
    );

    or_bb _2069_ (
        .b(jinkela_wire_251),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1117)
    );

    and_bi _2787_ (
        .b(jinkela_wire_530),
        .a(jinkela_wire_1060),
        .c(jinkela_wire_597)
    );

    and_bi _2070_ (
        .b(jinkela_wire_95),
        .a(jinkela_wire_188),
        .c(jinkela_wire_487)
    );

    or_bb _2788_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_597),
        .c(jinkela_wire_1330)
    );

    and_bi _2071_ (
        .b(jinkela_wire_487),
        .a(jinkela_wire_1117),
        .c(jinkela_wire_955)
    );

    and_bi _2789_ (
        .b(jinkela_wire_1121),
        .a(jinkela_wire_347),
        .c(jinkela_wire_3)
    );

    and_bi _2072_ (
        .b(jinkela_wire_955),
        .a(io_in2_0_),
        .c(jinkela_wire_643)
    );

    and_bi _2577_ (
        .b(jinkela_wire_1099),
        .a(io_in2_2_),
        .c(jinkela_wire_170)
    );

    or_bb _2578_ (
        .b(jinkela_wire_531),
        .a(jinkela_wire_170),
        .c(jinkela_wire_761)
    );

    and_bi _2579_ (
        .b(jinkela_wire_761),
        .a(io_in2_3_),
        .c(jinkela_wire_1335)
    );

    or_bb _2580_ (
        .b(jinkela_wire_377),
        .a(jinkela_wire_1335),
        .c(jinkela_wire_79)
    );

    and_bi _2581_ (
        .b(jinkela_wire_79),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_1508)
    );

    and_bi _2582_ (
        .b(jinkela_wire_804),
        .a(jinkela_wire_1331),
        .c(jinkela_wire_28)
    );

    and_bi _2583_ (
        .b(jinkela_wire_144),
        .a(jinkela_wire_158),
        .c(jinkela_wire_1225)
    );

    and_bi _2584_ (
        .b(jinkela_wire_158),
        .a(jinkela_wire_944),
        .c(jinkela_wire_1208)
    );

    or_bb _2585_ (
        .b(jinkela_wire_1225),
        .a(jinkela_wire_1208),
        .c(jinkela_wire_1347)
    );

    and_bi _2586_ (
        .b(jinkela_wire_1347),
        .a(jinkela_wire_804),
        .c(jinkela_wire_1238)
    );

    or_bb _2587_ (
        .b(jinkela_wire_28),
        .a(jinkela_wire_1238),
        .c(jinkela_wire_787)
    );

    and_bi _2588_ (
        .b(jinkela_wire_787),
        .a(io_in2_4_),
        .c(jinkela_wire_1076)
    );

    or_bb _2589_ (
        .b(jinkela_wire_1508),
        .a(jinkela_wire_1076),
        .c(jinkela_wire_1340)
    );

    and_bi _2590_ (
        .b(jinkela_wire_1340),
        .a(jinkela_wire_188),
        .c(jinkela_wire_928)
    );

    or_bb _2591_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_928),
        .c(jinkela_wire_508)
    );

    and_bi _2592_ (
        .b(jinkela_wire_508),
        .a(jinkela_wire_290),
        .c(jinkela_wire_53)
    );

    or_bb _2593_ (
        .b(jinkela_wire_975),
        .a(jinkela_wire_53),
        .c(io_out_6_)
    );

    and_bi _2594_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_7_),
        .c(jinkela_wire_1197)
    );

    and_bi _2595_ (
        .b(jinkela_wire_1158),
        .a(jinkela_wire_804),
        .c(jinkela_wire_1496)
    );

    and_bi _2596_ (
        .b(jinkela_wire_1496),
        .a(jinkela_wire_1269),
        .c(jinkela_wire_566)
    );

    and_bi _2597_ (
        .b(jinkela_wire_566),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_84)
    );

    and_bi _2598_ (
        .b(jinkela_wire_84),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_646)
    );

    and_bi _2599_ (
        .b(jinkela_wire_646),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_387)
    );

    or_bb _2600_ (
        .b(jinkela_wire_95),
        .a(jinkela_wire_347),
        .c(jinkela_wire_489)
    );

    and_bi _2601_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_95),
        .c(jinkela_wire_1403)
    );

    or_bb _2602_ (
        .b(jinkela_wire_1490),
        .a(jinkela_wire_1403),
        .c(jinkela_wire_118)
    );

    or_ii _2603_ (
        .b(jinkela_wire_489),
        .a(jinkela_wire_118),
        .c(jinkela_wire_1432)
    );

    and_bi _2607_ (
        .b(jinkela_wire_1444),
        .a(jinkela_wire_1432),
        .c(jinkela_wire_1476)
    );

    or_bb _2608_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1476),
        .c(jinkela_wire_1280)
    );

    or_bb _2609_ (
        .b(jinkela_wire_387),
        .a(jinkela_wire_1280),
        .c(jinkela_wire_252)
    );

    or_bb _2610_ (
        .b(io_in2_2_),
        .a(jinkela_wire_363),
        .c(jinkela_wire_263)
    );

    and_bi _2611_ (
        .b(jinkela_wire_724),
        .a(io_in2_2_),
        .c(jinkela_wire_1310)
    );

    and_bi _2612_ (
        .b(jinkela_wire_1310),
        .a(jinkela_wire_263),
        .c(jinkela_wire_935)
    );

    and_bi _2613_ (
        .b(jinkela_wire_935),
        .a(jinkela_wire_804),
        .c(jinkela_wire_1167)
    );

    and_bi _2614_ (
        .b(jinkela_wire_1482),
        .a(jinkela_wire_158),
        .c(jinkela_wire_455)
    );

    and_bi _2615_ (
        .b(jinkela_wire_479),
        .a(io_in2_2_),
        .c(jinkela_wire_660)
    );

    or_bb _2616_ (
        .b(jinkela_wire_455),
        .a(jinkela_wire_660),
        .c(jinkela_wire_1246)
    );

    and_bi _2617_ (
        .b(jinkela_wire_804),
        .a(jinkela_wire_1246),
        .c(jinkela_wire_709)
    );

    or_bb _2618_ (
        .b(jinkela_wire_1167),
        .a(jinkela_wire_709),
        .c(jinkela_wire_1442)
    );

    and_bi _2619_ (
        .b(jinkela_wire_1442),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_1312)
    );

    or_bb _2620_ (
        .b(io_in2_2_),
        .a(jinkela_wire_1010),
        .c(jinkela_wire_748)
    );

    and_bi _2621_ (
        .b(jinkela_wire_158),
        .a(jinkela_wire_12),
        .c(jinkela_wire_56)
    );

    or_ii _1863_ (
        .b(jinkela_wire_227),
        .a(jinkela_wire_186),
        .c(jinkela_wire_1416)
    );

    and_bi _1864_ (
        .b(jinkela_wire_1332),
        .a(jinkela_wire_1416),
        .c(io_adder_out_28_)
    );

    and_bb _1865_ (
        .b(jinkela_wire_61),
        .a(jinkela_wire_1471),
        .c(jinkela_wire_805)
    );

    and_bi _1866_ (
        .b(jinkela_wire_805),
        .a(jinkela_wire_255),
        .c(jinkela_wire_36)
    );

    and_bb _1867_ (
        .b(jinkela_wire_61),
        .a(jinkela_wire_1062),
        .c(jinkela_wire_69)
    );

    or_bb _1868_ (
        .b(jinkela_wire_36),
        .a(jinkela_wire_69),
        .c(io_adder_out_27_)
    );

    and_bb _1869_ (
        .b(jinkela_wire_814),
        .a(jinkela_wire_516),
        .c(jinkela_wire_167)
    );

    or_ii _1870_ (
        .b(jinkela_wire_8),
        .a(jinkela_wire_167),
        .c(jinkela_wire_666)
    );

    or_bb _1871_ (
        .b(jinkela_wire_8),
        .a(jinkela_wire_167),
        .c(jinkela_wire_58)
    );

    or_ii _1872_ (
        .b(jinkela_wire_666),
        .a(jinkela_wire_58),
        .c(io_adder_out_26_)
    );

    and_bi _1873_ (
        .b(jinkela_wire_1468),
        .a(jinkela_wire_342),
        .c(jinkela_wire_393)
    );

    or_bb _1874_ (
        .b(jinkela_wire_228),
        .a(jinkela_wire_393),
        .c(jinkela_wire_1215)
    );

    and_bb _1875_ (
        .b(jinkela_wire_228),
        .a(jinkela_wire_393),
        .c(jinkela_wire_1348)
    );

    and_bi _1876_ (
        .b(jinkela_wire_1348),
        .a(jinkela_wire_1215),
        .c(io_adder_out_25_)
    );

    and_bi _1877_ (
        .b(jinkela_wire_856),
        .a(jinkela_wire_299),
        .c(jinkela_wire_1116)
    );

    or_bb _1878_ (
        .b(jinkela_wire_1319),
        .a(jinkela_wire_1116),
        .c(jinkela_wire_1008)
    );

    and_bb _1879_ (
        .b(jinkela_wire_1319),
        .a(jinkela_wire_1116),
        .c(jinkela_wire_326)
    );

    and_bi _1880_ (
        .b(jinkela_wire_326),
        .a(jinkela_wire_1008),
        .c(io_adder_out_24_)
    );

    and_bi _1881_ (
        .b(jinkela_wire_1245),
        .a(jinkela_wire_165),
        .c(jinkela_wire_1148)
    );

    and_bi _1882_ (
        .b(jinkela_wire_180),
        .a(jinkela_wire_1148),
        .c(jinkela_wire_1435)
    );

    and_bi _1883_ (
        .b(jinkela_wire_1148),
        .a(jinkela_wire_180),
        .c(jinkela_wire_88)
    );

    or_bb _1884_ (
        .b(jinkela_wire_1435),
        .a(jinkela_wire_88),
        .c(io_adder_out_23_)
    );

    and_bi _1885_ (
        .b(jinkela_wire_1096),
        .a(jinkela_wire_834),
        .c(jinkela_wire_1130)
    );

    or_bb _1886_ (
        .b(jinkela_wire_420),
        .a(jinkela_wire_1130),
        .c(jinkela_wire_428)
    );

    and_bb _1887_ (
        .b(jinkela_wire_420),
        .a(jinkela_wire_1130),
        .c(jinkela_wire_245)
    );

    and_bi _1888_ (
        .b(jinkela_wire_245),
        .a(jinkela_wire_428),
        .c(io_adder_out_22_)
    );

    and_bi _1889_ (
        .b(jinkela_wire_1230),
        .a(jinkela_wire_684),
        .c(jinkela_wire_946)
    );

    and_bi _1890_ (
        .b(jinkela_wire_946),
        .a(jinkela_wire_1244),
        .c(jinkela_wire_1454)
    );

    and_bi _1891_ (
        .b(jinkela_wire_1244),
        .a(jinkela_wire_946),
        .c(jinkela_wire_1249)
    );

    or_bb _1892_ (
        .b(jinkela_wire_1454),
        .a(jinkela_wire_1249),
        .c(io_adder_out_21_)
    );

    and_bi _1893_ (
        .b(jinkela_wire_270),
        .a(jinkela_wire_656),
        .c(jinkela_wire_966)
    );

    or_bb _1894_ (
        .b(jinkela_wire_847),
        .a(jinkela_wire_966),
        .c(jinkela_wire_672)
    );

    and_bb _1895_ (
        .b(jinkela_wire_847),
        .a(jinkela_wire_966),
        .c(jinkela_wire_1163)
    );

    and_bi _1896_ (
        .b(jinkela_wire_1163),
        .a(jinkela_wire_672),
        .c(io_adder_out_20_)
    );

    and_bi _1897_ (
        .b(jinkela_wire_1114),
        .a(jinkela_wire_1264),
        .c(jinkela_wire_723)
    );

    and_bi _1898_ (
        .b(jinkela_wire_237),
        .a(jinkela_wire_723),
        .c(jinkela_wire_146)
    );

    and_bi _1899_ (
        .b(jinkela_wire_723),
        .a(jinkela_wire_237),
        .c(jinkela_wire_851)
    );

    or_bb _1900_ (
        .b(jinkela_wire_146),
        .a(jinkela_wire_851),
        .c(io_adder_out_19_)
    );

    and_bb _1901_ (
        .b(jinkela_wire_271),
        .a(jinkela_wire_983),
        .c(jinkela_wire_841)
    );

    and_bi _1902_ (
        .b(jinkela_wire_1086),
        .a(jinkela_wire_841),
        .c(jinkela_wire_813)
    );

    and_bi _1903_ (
        .b(jinkela_wire_841),
        .a(jinkela_wire_1086),
        .c(jinkela_wire_66)
    );

    or_bb _1904_ (
        .b(jinkela_wire_813),
        .a(jinkela_wire_66),
        .c(io_adder_out_18_)
    );

    and_bi _2409_ (
        .b(jinkela_wire_626),
        .a(jinkela_wire_544),
        .c(jinkela_wire_629)
    );

    or_bb _2410_ (
        .b(jinkela_wire_574),
        .a(jinkela_wire_629),
        .c(io_out_2_)
    );

    and_bi _2411_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_3_),
        .c(jinkela_wire_640)
    );

    and_bi _2412_ (
        .b(jinkela_wire_1418),
        .a(jinkela_wire_158),
        .c(jinkela_wire_1357)
    );

    or_bb _2413_ (
        .b(jinkela_wire_1080),
        .a(jinkela_wire_1357),
        .c(jinkela_wire_1036)
    );

    and_bi _2414_ (
        .b(io_in2_3_),
        .a(jinkela_wire_1036),
        .c(jinkela_wire_631)
    );

    and_bi _2415_ (
        .b(jinkela_wire_631),
        .a(jinkela_wire_1269),
        .c(jinkela_wire_752)
    );

    and_bi _2416_ (
        .b(jinkela_wire_752),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_85)
    );

    and_bi _2417_ (
        .b(jinkela_wire_85),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_1381)
    );

    and_bi _2418_ (
        .b(jinkela_wire_1381),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_1183)
    );

    or_ii _2419_ (
        .b(io_in1_3_),
        .a(io_in2_3_),
        .c(jinkela_wire_81)
    );

    or_bi _2420_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_81),
        .c(jinkela_wire_1093)
    );

    and_bi _2421_ (
        .b(jinkela_wire_804),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_536)
    );

    or_bb _2422_ (
        .b(io_in1_3_),
        .a(jinkela_wire_536),
        .c(jinkela_wire_279)
    );

    and_bi _2423_ (
        .b(jinkela_wire_81),
        .a(jinkela_wire_349),
        .c(jinkela_wire_348)
    );

    or_bb _2424_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_348),
        .c(jinkela_wire_444)
    );

    and_bi _2425_ (
        .b(jinkela_wire_444),
        .a(jinkela_wire_279),
        .c(jinkela_wire_1164)
    );

    and_bi _2426_ (
        .b(jinkela_wire_1164),
        .a(jinkela_wire_1093),
        .c(jinkela_wire_447)
    );

    and_bi _2427_ (
        .b(jinkela_wire_447),
        .a(jinkela_wire_44),
        .c(jinkela_wire_1486)
    );

    or_bb _2428_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1486),
        .c(jinkela_wire_398)
    );

    or_bb _2429_ (
        .b(jinkela_wire_1183),
        .a(jinkela_wire_398),
        .c(jinkela_wire_273)
    );

    or_bb _2430_ (
        .b(jinkela_wire_15),
        .a(jinkela_wire_1473),
        .c(jinkela_wire_751)
    );

    and_bi _2431_ (
        .b(jinkela_wire_1040),
        .a(jinkela_wire_15),
        .c(jinkela_wire_1065)
    );

    and_bi _2432_ (
        .b(jinkela_wire_1065),
        .a(jinkela_wire_751),
        .c(jinkela_wire_676)
    );

    or_bb _2433_ (
        .b(io_in2_2_),
        .a(jinkela_wire_676),
        .c(jinkela_wire_1047)
    );

    or_bb _2434_ (
        .b(io_in2_1_),
        .a(jinkela_wire_258),
        .c(jinkela_wire_257)
    );

    and_bi _2435_ (
        .b(jinkela_wire_1433),
        .a(io_in2_1_),
        .c(jinkela_wire_151)
    );

    and_bi _2436_ (
        .b(jinkela_wire_151),
        .a(jinkela_wire_257),
        .c(jinkela_wire_363)
    );

    and_bi _2437_ (
        .b(jinkela_wire_363),
        .a(io_in2_2_),
        .c(jinkela_wire_1122)
    );

    and_bi _2438_ (
        .b(jinkela_wire_1122),
        .a(jinkela_wire_1047),
        .c(jinkela_wire_806)
    );

    or_bb _2439_ (
        .b(io_in2_3_),
        .a(jinkela_wire_806),
        .c(jinkela_wire_296)
    );

    or_bb _2440_ (
        .b(io_in2_1_),
        .a(jinkela_wire_1419),
        .c(jinkela_wire_286)
    );

    and_bi _2441_ (
        .b(jinkela_wire_750),
        .a(io_in2_1_),
        .c(jinkela_wire_694)
    );

    and_bi _2442_ (
        .b(jinkela_wire_694),
        .a(jinkela_wire_286),
        .c(jinkela_wire_724)
    );

    or_bb _2443_ (
        .b(io_in2_2_),
        .a(jinkela_wire_724),
        .c(jinkela_wire_795)
    );

    or_bb _2444_ (
        .b(io_in2_1_),
        .a(jinkela_wire_621),
        .c(jinkela_wire_833)
    );

    and_bi _2445_ (
        .b(jinkela_wire_811),
        .a(io_in2_1_),
        .c(jinkela_wire_1404)
    );

    and_bi _2446_ (
        .b(jinkela_wire_1404),
        .a(jinkela_wire_833),
        .c(jinkela_wire_1482)
    );

    and_bi _2447_ (
        .b(jinkela_wire_1482),
        .a(io_in2_2_),
        .c(jinkela_wire_1054)
    );

    and_bi _2448_ (
        .b(jinkela_wire_1054),
        .a(jinkela_wire_795),
        .c(jinkela_wire_1406)
    );

    and_bi _2449_ (
        .b(jinkela_wire_1406),
        .a(io_in2_3_),
        .c(jinkela_wire_1261)
    );

    and_bi _2450_ (
        .b(jinkela_wire_1261),
        .a(jinkela_wire_296),
        .c(jinkela_wire_610)
    );

    and_bi _1695_ (
        .b(jinkela_wire_1005),
        .a(jinkela_wire_877),
        .c(jinkela_wire_395)
    );

    and_bi _1696_ (
        .b(jinkela_wire_395),
        .a(jinkela_wire_1029),
        .c(jinkela_wire_789)
    );

    or_bi _1697_ (
        .b(jinkela_wire_1251),
        .a(jinkela_wire_789),
        .c(jinkela_wire_206)
    );

    and_bi _1698_ (
        .b(io_in1_14_),
        .a(jinkela_wire_206),
        .c(jinkela_wire_1446)
    );

    inv _1699_ (
        .din(io_in1_14_),
        .dout(jinkela_wire_1073)
    );

    or_bb _1700_ (
        .b(jinkela_wire_1073),
        .a(jinkela_wire_206),
        .c(jinkela_wire_893)
    );

    and_bi _1701_ (
        .b(jinkela_wire_1475),
        .a(io_fn_3_),
        .c(jinkela_wire_1069)
    );

    and_bi _1702_ (
        .b(io_in2_14_),
        .a(jinkela_wire_1069),
        .c(jinkela_wire_1210)
    );

    and_bi _1703_ (
        .b(jinkela_wire_1069),
        .a(io_in2_14_),
        .c(jinkela_wire_661)
    );

    or_bb _1704_ (
        .b(jinkela_wire_1210),
        .a(jinkela_wire_661),
        .c(jinkela_wire_790)
    );

    and_bi _1705_ (
        .b(jinkela_wire_790),
        .a(jinkela_wire_893),
        .c(jinkela_wire_760)
    );

    or_bb _1706_ (
        .b(jinkela_wire_1446),
        .a(jinkela_wire_760),
        .c(jinkela_wire_1159)
    );

    and_bi _1707_ (
        .b(io_in1_15_),
        .a(jinkela_wire_1159),
        .c(jinkela_wire_222)
    );

    inv _1708_ (
        .din(io_in1_15_),
        .dout(jinkela_wire_224)
    );

    or_bb _1709_ (
        .b(jinkela_wire_224),
        .a(jinkela_wire_1159),
        .c(jinkela_wire_30)
    );

    inv _1710_ (
        .din(io_in2_15_),
        .dout(jinkela_wire_301)
    );

    and_bi _1711_ (
        .b(jinkela_wire_971),
        .a(io_fn_3_),
        .c(jinkela_wire_575)
    );

    and_bi _1712_ (
        .b(jinkela_wire_301),
        .a(jinkela_wire_575),
        .c(jinkela_wire_1265)
    );

    and_bi _1713_ (
        .b(jinkela_wire_575),
        .a(jinkela_wire_301),
        .c(jinkela_wire_441)
    );

    or_bb _1714_ (
        .b(jinkela_wire_1265),
        .a(jinkela_wire_441),
        .c(jinkela_wire_1470)
    );

    inv _1715_ (
        .din(jinkela_wire_1470),
        .dout(jinkela_wire_563)
    );

    and_bi _1716_ (
        .b(jinkela_wire_563),
        .a(jinkela_wire_30),
        .c(jinkela_wire_853)
    );

    or_bb _1717_ (
        .b(jinkela_wire_222),
        .a(jinkela_wire_853),
        .c(jinkela_wire_678)
    );

    and_bi _1718_ (
        .b(jinkela_wire_678),
        .a(io_in1_16_),
        .c(jinkela_wire_409)
    );

    inv _1719_ (
        .din(io_in1_16_),
        .dout(jinkela_wire_7)
    );

    or_ii _1720_ (
        .b(jinkela_wire_7),
        .a(jinkela_wire_678),
        .c(jinkela_wire_545)
    );

    and_bi _1721_ (
        .b(jinkela_wire_421),
        .a(io_fn_3_),
        .c(jinkela_wire_41)
    );

    and_bi _1722_ (
        .b(io_in2_16_),
        .a(jinkela_wire_41),
        .c(jinkela_wire_557)
    );

    and_bi _1723_ (
        .b(jinkela_wire_41),
        .a(io_in2_16_),
        .c(jinkela_wire_902)
    );

    or_bb _1724_ (
        .b(jinkela_wire_557),
        .a(jinkela_wire_902),
        .c(jinkela_wire_1481)
    );

    and_bb _1725_ (
        .b(jinkela_wire_545),
        .a(jinkela_wire_1481),
        .c(jinkela_wire_541)
    );

    or_bb _1726_ (
        .b(jinkela_wire_409),
        .a(jinkela_wire_541),
        .c(jinkela_wire_539)
    );

    and_bi _1727_ (
        .b(jinkela_wire_899),
        .a(jinkela_wire_539),
        .c(jinkela_wire_1441)
    );

    or_bb _1728_ (
        .b(io_in1_17_),
        .a(jinkela_wire_539),
        .c(jinkela_wire_606)
    );

    inv _1729_ (
        .din(io_in2_17_),
        .dout(jinkela_wire_34)
    );

    and_bi _1730_ (
        .b(jinkela_wire_887),
        .a(io_fn_3_),
        .c(jinkela_wire_1039)
    );

    and_bi _1731_ (
        .b(jinkela_wire_34),
        .a(jinkela_wire_1039),
        .c(jinkela_wire_443)
    );

    and_bi _1732_ (
        .b(jinkela_wire_1039),
        .a(jinkela_wire_34),
        .c(jinkela_wire_1157)
    );

    inv _1521_ (
        .din(io_in2_29_),
        .dout(jinkela_wire_262)
    );

    inv _1519_ (
        .din(io_in2_31_),
        .dout(jinkela_wire_231)
    );

    or_bb _1733_ (
        .b(jinkela_wire_443),
        .a(jinkela_wire_1157),
        .c(jinkela_wire_243)
    );

    inv _1520_ (
        .din(io_fn_3_),
        .dout(jinkela_wire_1424)
    );

    and_bi _1734_ (
        .b(jinkela_wire_243),
        .a(jinkela_wire_606),
        .c(jinkela_wire_607)
    );

    or_bb _1735_ (
        .b(jinkela_wire_1441),
        .a(jinkela_wire_607),
        .c(jinkela_wire_984)
    );

    inv _1518_ (
        .din(io_in1_31_),
        .dout(jinkela_wire_560)
    );

    inv _1522_ (
        .din(io_in2_2_),
        .dout(jinkela_wire_158)
    );

    or_ii _1736_ (
        .b(io_in1_18_),
        .a(jinkela_wire_984),
        .c(jinkela_wire_271)
    );

    or_bb _1523_ (
        .b(io_in2_0_),
        .a(io_in2_1_),
        .c(jinkela_wire_1038)
    );

    or_bb _2958_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_1427),
        .c(jinkela_wire_614)
    );

    and_bi _1524_ (
        .b(jinkela_wire_1038),
        .a(jinkela_wire_158),
        .c(jinkela_wire_1338)
    );

    or_bb _2241_ (
        .b(io_in1_1_),
        .a(jinkela_wire_213),
        .c(jinkela_wire_1390)
    );

    and_bi _2959_ (
        .b(jinkela_wire_614),
        .a(jinkela_wire_375),
        .c(jinkela_wire_517)
    );

    and_bi _1525_ (
        .b(io_in2_3_),
        .a(jinkela_wire_1338),
        .c(jinkela_wire_29)
    );

    and_bb _2242_ (
        .b(io_in1_1_),
        .a(io_in2_1_),
        .c(jinkela_wire_725)
    );

    or_bb _2960_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_517),
        .c(jinkela_wire_1502)
    );

    and_bi _1526_ (
        .b(io_in2_4_),
        .a(jinkela_wire_29),
        .c(jinkela_wire_1405)
    );

    and_bb _2243_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_725),
        .c(jinkela_wire_1276)
    );

    or_bb _2961_ (
        .b(jinkela_wire_700),
        .a(jinkela_wire_1502),
        .c(jinkela_wire_1199)
    );

    and_bi _1527_ (
        .b(io_in2_5_),
        .a(jinkela_wire_1405),
        .c(jinkela_wire_1168)
    );

    and_bi _2244_ (
        .b(jinkela_wire_1276),
        .a(jinkela_wire_1390),
        .c(jinkela_wire_808)
    );

    and_bb _2962_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1309),
        .c(jinkela_wire_717)
    );

    and_bi _1528_ (
        .b(io_in2_6_),
        .a(jinkela_wire_1168),
        .c(jinkela_wire_1079)
    );

    or_bb _2245_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_808),
        .c(jinkela_wire_707)
    );

    or_bb _2963_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_717),
        .c(jinkela_wire_1431)
    );

    and_bi _1529_ (
        .b(io_in2_7_),
        .a(jinkela_wire_1079),
        .c(jinkela_wire_100)
    );

    and_bi _2246_ (
        .b(jinkela_wire_725),
        .a(jinkela_wire_347),
        .c(jinkela_wire_1179)
    );

    and_bi _2964_ (
        .b(jinkela_wire_1431),
        .a(jinkela_wire_1199),
        .c(jinkela_wire_511)
    );

    and_bi _1530_ (
        .b(io_in2_8_),
        .a(jinkela_wire_100),
        .c(jinkela_wire_870)
    );

    or_bb _2247_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_1179),
        .c(jinkela_wire_495)
    );

    or_bb _2965_ (
        .b(jinkela_wire_852),
        .a(jinkela_wire_511),
        .c(io_out_23_)
    );

    and_bi _1531_ (
        .b(io_in2_9_),
        .a(jinkela_wire_870),
        .c(jinkela_wire_667)
    );

    and_bi _2248_ (
        .b(jinkela_wire_495),
        .a(jinkela_wire_707),
        .c(jinkela_wire_1489)
    );

    and_bi _2966_ (
        .b(jinkela_wire_866),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_653)
    );

    and_bi _1532_ (
        .b(io_in2_10_),
        .a(jinkela_wire_667),
        .c(jinkela_wire_652)
    );

    or_bb _2249_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1489),
        .c(jinkela_wire_17)
    );

    and_bb _2967_ (
        .b(io_in2_24_),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_1220)
    );

    and_bi _1533_ (
        .b(io_in2_11_),
        .a(jinkela_wire_652),
        .c(jinkela_wire_598)
    );

    or_bb _2250_ (
        .b(jinkela_wire_37),
        .a(jinkela_wire_17),
        .c(jinkela_wire_986)
    );

    or_bb _2968_ (
        .b(io_in1_24_),
        .a(jinkela_wire_1220),
        .c(jinkela_wire_774)
    );

    and_bi _1534_ (
        .b(io_in2_12_),
        .a(jinkela_wire_598),
        .c(jinkela_wire_333)
    );

    or_bb _2251_ (
        .b(io_in2_0_),
        .a(jinkela_wire_895),
        .c(jinkela_wire_861)
    );

    and_bb _2969_ (
        .b(io_in1_24_),
        .a(io_in2_24_),
        .c(jinkela_wire_31)
    );

    and_bi _1535_ (
        .b(io_in2_13_),
        .a(jinkela_wire_333),
        .c(jinkela_wire_1475)
    );

    and_bi _2252_ (
        .b(jinkela_wire_202),
        .a(io_in2_0_),
        .c(jinkela_wire_124)
    );

    and_bb _2970_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_31),
        .c(jinkela_wire_150)
    );

    and_bi _1536_ (
        .b(io_in2_14_),
        .a(jinkela_wire_1475),
        .c(jinkela_wire_971)
    );

    and_bi _2253_ (
        .b(jinkela_wire_124),
        .a(jinkela_wire_861),
        .c(jinkela_wire_1433)
    );

    and_bi _2971_ (
        .b(jinkela_wire_150),
        .a(jinkela_wire_774),
        .c(jinkela_wire_641)
    );

    and_bi _1537_ (
        .b(io_in2_15_),
        .a(jinkela_wire_971),
        .c(jinkela_wire_421)
    );

    and_bi _2254_ (
        .b(jinkela_wire_1433),
        .a(jinkela_wire_15),
        .c(jinkela_wire_42)
    );

    or_bb _2972_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_641),
        .c(jinkela_wire_1089)
    );

    and_bi _1538_ (
        .b(io_in2_16_),
        .a(jinkela_wire_421),
        .c(jinkela_wire_887)
    );

    or_bb _2255_ (
        .b(io_in2_0_),
        .a(jinkela_wire_1205),
        .c(jinkela_wire_1257)
    );

    and_bi _2973_ (
        .b(jinkela_wire_31),
        .a(jinkela_wire_347),
        .c(jinkela_wire_168)
    );

    and_bi _1539_ (
        .b(io_in2_17_),
        .a(jinkela_wire_887),
        .c(jinkela_wire_145)
    );

    and_bi _2256_ (
        .b(jinkela_wire_911),
        .a(io_in2_0_),
        .c(jinkela_wire_995)
    );

    or_bb _2974_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_168),
        .c(jinkela_wire_884)
    );

    and_bi _1540_ (
        .b(io_in2_18_),
        .a(jinkela_wire_145),
        .c(jinkela_wire_957)
    );

    and_bi _2257_ (
        .b(jinkela_wire_995),
        .a(jinkela_wire_1257),
        .c(jinkela_wire_1419)
    );

    and_bi _2975_ (
        .b(jinkela_wire_884),
        .a(jinkela_wire_1089),
        .c(jinkela_wire_792)
    );

    and_bi _1541_ (
        .b(io_in2_19_),
        .a(jinkela_wire_957),
        .c(jinkela_wire_1186)
    );

    and_bi _2258_ (
        .b(jinkela_wire_1419),
        .a(io_in2_1_),
        .c(jinkela_wire_431)
    );

    or_bb _2976_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_792),
        .c(jinkela_wire_74)
    );

    and_bi _1542_ (
        .b(io_in2_20_),
        .a(jinkela_wire_1186),
        .c(jinkela_wire_154)
    );

    or_bb _2259_ (
        .b(jinkela_wire_42),
        .a(jinkela_wire_431),
        .c(jinkela_wire_137)
    );

    or_bb _2977_ (
        .b(jinkela_wire_653),
        .a(jinkela_wire_74),
        .c(jinkela_wire_838)
    );

    and_bi _1543_ (
        .b(io_in2_21_),
        .a(jinkela_wire_154),
        .c(jinkela_wire_1359)
    );

    or_ii _2260_ (
        .b(jinkela_wire_158),
        .a(jinkela_wire_137),
        .c(jinkela_wire_1250)
    );

    and_bb _2978_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_646),
        .c(jinkela_wire_766)
    );

    and_bi _1544_ (
        .b(io_in2_22_),
        .a(jinkela_wire_1359),
        .c(jinkela_wire_839)
    );

    or_bb _2261_ (
        .b(io_in2_0_),
        .a(jinkela_wire_772),
        .c(jinkela_wire_331)
    );

    or_bb _2979_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_766),
        .c(jinkela_wire_999)
    );

    and_bi _1545_ (
        .b(io_in2_23_),
        .a(jinkela_wire_839),
        .c(jinkela_wire_1128)
    );

    and_bi _2262_ (
        .b(jinkela_wire_200),
        .a(io_in2_0_),
        .c(jinkela_wire_226)
    );

    and_bi _2980_ (
        .b(jinkela_wire_999),
        .a(jinkela_wire_838),
        .c(jinkela_wire_439)
    );

    and_bi _1546_ (
        .b(io_in2_24_),
        .a(jinkela_wire_1128),
        .c(jinkela_wire_923)
    );

    and_bi _2263_ (
        .b(jinkela_wire_226),
        .a(jinkela_wire_331),
        .c(jinkela_wire_750)
    );

    and_bi _2981_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_24_),
        .c(jinkela_wire_1290)
    );

    and_bi _1547_ (
        .b(io_in2_25_),
        .a(jinkela_wire_923),
        .c(jinkela_wire_1058)
    );

    or_bb _2264_ (
        .b(io_in2_1_),
        .a(jinkela_wire_750),
        .c(jinkela_wire_933)
    );

    or_bb _2982_ (
        .b(jinkela_wire_439),
        .a(jinkela_wire_1290),
        .c(io_out_24_)
    );

    and_bi _1548_ (
        .b(io_in2_26_),
        .a(jinkela_wire_1058),
        .c(jinkela_wire_1224)
    );

    and_bi _2265_ (
        .b(jinkela_wire_1087),
        .a(io_in2_0_),
        .c(jinkela_wire_1355)
    );

    and_bi _2983_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_25_),
        .c(jinkela_wire_1185)
    );

    and_bi _1549_ (
        .b(io_in2_27_),
        .a(jinkela_wire_1224),
        .c(jinkela_wire_117)
    );

    and_bi _2266_ (
        .b(jinkela_wire_288),
        .a(jinkela_wire_915),
        .c(jinkela_wire_486)
    );

    and_bi _2984_ (
        .b(jinkela_wire_44),
        .a(jinkela_wire_1340),
        .c(jinkela_wire_496)
    );

    or_bb _1550_ (
        .b(jinkela_wire_1424),
        .a(jinkela_wire_117),
        .c(jinkela_wire_1195)
    );

    or_bb _2267_ (
        .b(jinkela_wire_1355),
        .a(jinkela_wire_486),
        .c(jinkela_wire_621)
    );

    and_bb _2985_ (
        .b(io_in2_25_),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_1105)
    );

    and_bi _1551_ (
        .b(io_in2_28_),
        .a(jinkela_wire_1195),
        .c(jinkela_wire_308)
    );

    and_bi _2268_ (
        .b(jinkela_wire_621),
        .a(io_in2_1_),
        .c(jinkela_wire_802)
    );

    or_bb _2986_ (
        .b(io_in1_25_),
        .a(jinkela_wire_1105),
        .c(jinkela_wire_1421)
    );

    and_bi _1552_ (
        .b(jinkela_wire_308),
        .a(io_fn_3_),
        .c(jinkela_wire_1014)
    );

    and_bi _2269_ (
        .b(jinkela_wire_802),
        .a(jinkela_wire_933),
        .c(jinkela_wire_937)
    );

    and_bb _2987_ (
        .b(io_in1_25_),
        .a(io_in2_25_),
        .c(jinkela_wire_967)
    );

    and_bi _1553_ (
        .b(jinkela_wire_1014),
        .a(jinkela_wire_262),
        .c(jinkela_wire_1411)
    );

    and_bi _2270_ (
        .b(jinkela_wire_937),
        .a(io_in2_2_),
        .c(jinkela_wire_1500)
    );

    and_bb _2988_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_967),
        .c(jinkela_wire_612)
    );

    or_bb _1554_ (
        .b(jinkela_wire_1424),
        .a(jinkela_wire_1411),
        .c(jinkela_wire_559)
    );

    and_bi _2271_ (
        .b(jinkela_wire_1500),
        .a(jinkela_wire_1250),
        .c(jinkela_wire_635)
    );

    and_bi _2989_ (
        .b(jinkela_wire_612),
        .a(jinkela_wire_1421),
        .c(jinkela_wire_50)
    );

    and_bb _1555_ (
        .b(io_fn_3_),
        .a(io_in2_30_),
        .c(jinkela_wire_239)
    );

    or_bb _2272_ (
        .b(jinkela_wire_804),
        .a(jinkela_wire_635),
        .c(jinkela_wire_507)
    );

    or_bb _2990_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_50),
        .c(jinkela_wire_139)
    );

    and_bi _1556_ (
        .b(jinkela_wire_239),
        .a(jinkela_wire_559),
        .c(jinkela_wire_515)
    );

    or_bb _2273_ (
        .b(io_in2_0_),
        .a(jinkela_wire_871),
        .c(jinkela_wire_685)
    );

    and_bi _2991_ (
        .b(jinkela_wire_967),
        .a(jinkela_wire_347),
        .c(jinkela_wire_39)
    );

    and_bi _1557_ (
        .b(jinkela_wire_515),
        .a(jinkela_wire_231),
        .c(jinkela_wire_820)
    );

    and_bi _2274_ (
        .b(jinkela_wire_436),
        .a(io_in2_0_),
        .c(jinkela_wire_974)
    );

    or_bb _2992_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_39),
        .c(jinkela_wire_675)
    );

    and_bi _1558_ (
        .b(jinkela_wire_231),
        .a(jinkela_wire_515),
        .c(jinkela_wire_1260)
    );

    and_bi _2275_ (
        .b(jinkela_wire_974),
        .a(jinkela_wire_685),
        .c(jinkela_wire_1040)
    );

    and_bi _2993_ (
        .b(jinkela_wire_675),
        .a(jinkela_wire_139),
        .c(jinkela_wire_265)
    );

    or_bb _1559_ (
        .b(jinkela_wire_820),
        .a(jinkela_wire_1260),
        .c(jinkela_wire_925)
    );

    or_bb _2276_ (
        .b(jinkela_wire_15),
        .a(jinkela_wire_1040),
        .c(jinkela_wire_1334)
    );

    or_bb _2994_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_265),
        .c(jinkela_wire_1395)
    );

    and_bi _1560_ (
        .b(jinkela_wire_560),
        .a(jinkela_wire_925),
        .c(jinkela_wire_338)
    );

    and_bb _2277_ (
        .b(jinkela_wire_1288),
        .a(jinkela_wire_201),
        .c(jinkela_wire_1430)
    );

    or_bb _2995_ (
        .b(jinkela_wire_496),
        .a(jinkela_wire_1395),
        .c(jinkela_wire_1145)
    );

    inv _1561_ (
        .din(jinkela_wire_338),
        .dout(jinkela_wire_882)
    );

    or_bb _2278_ (
        .b(jinkela_wire_1038),
        .a(jinkela_wire_905),
        .c(jinkela_wire_247)
    );

    and_bb _2996_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_799),
        .c(jinkela_wire_864)
    );

    and_bi _1562_ (
        .b(jinkela_wire_925),
        .a(jinkela_wire_560),
        .c(jinkela_wire_785)
    );

    or_ii _2279_ (
        .b(jinkela_wire_158),
        .a(jinkela_wire_247),
        .c(jinkela_wire_22)
    );

    or_bb _2997_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_864),
        .c(jinkela_wire_550)
    );

    and_bi _1563_ (
        .b(jinkela_wire_785),
        .a(jinkela_wire_882),
        .c(jinkela_wire_80)
    );

    or_bb _2280_ (
        .b(jinkela_wire_1430),
        .a(jinkela_wire_22),
        .c(jinkela_wire_452)
    );

    and_bi _2998_ (
        .b(jinkela_wire_550),
        .a(jinkela_wire_1145),
        .c(jinkela_wire_1314)
    );

    inv _1564_ (
        .din(io_in1_30_),
        .dout(jinkela_wire_964)
    );

    and_bi _2281_ (
        .b(jinkela_wire_452),
        .a(jinkela_wire_1334),
        .c(jinkela_wire_1514)
    );

    or_bb _2999_ (
        .b(jinkela_wire_1185),
        .a(jinkela_wire_1314),
        .c(io_out_25_)
    );

    inv _1565_ (
        .din(io_in1_27_),
        .dout(jinkela_wire_1234)
    );

    or_bb _2282_ (
        .b(io_in2_0_),
        .a(jinkela_wire_317),
        .c(jinkela_wire_590)
    );

    or_bb _2790_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_3),
        .c(jinkela_wire_193)
    );

    and_bi _2073_ (
        .b(jinkela_wire_643),
        .a(jinkela_wire_538),
        .c(jinkela_wire_18)
    );

    and_bi _2791_ (
        .b(jinkela_wire_193),
        .a(jinkela_wire_1330),
        .c(jinkela_wire_82)
    );

    and_bi _2074_ (
        .b(jinkela_wire_18),
        .a(io_in2_1_),
        .c(jinkela_wire_620)
    );

    or_bb _2792_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_82),
        .c(jinkela_wire_1236)
    );

    or_bb _2075_ (
        .b(jinkela_wire_1074),
        .a(jinkela_wire_620),
        .c(jinkela_wire_648)
    );

    or_bb _2793_ (
        .b(jinkela_wire_311),
        .a(jinkela_wire_1236),
        .c(jinkela_wire_655)
    );

    and_bi _2076_ (
        .b(jinkela_wire_648),
        .a(io_in2_2_),
        .c(jinkela_wire_1374)
    );

    and_bi _2794_ (
        .b(jinkela_wire_761),
        .a(jinkela_wire_804),
        .c(jinkela_wire_205)
    );

    and_bi _2077_ (
        .b(jinkela_wire_188),
        .a(io_in1_29_),
        .c(jinkela_wire_2)
    );

    and_bi _2795_ (
        .b(jinkela_wire_1347),
        .a(io_in2_3_),
        .c(jinkela_wire_408)
    );

    and_bi _2078_ (
        .b(jinkela_wire_958),
        .a(jinkela_wire_188),
        .c(jinkela_wire_570)
    );

    or_bb _2796_ (
        .b(jinkela_wire_205),
        .a(jinkela_wire_408),
        .c(jinkela_wire_1110)
    );

    or_bb _2079_ (
        .b(jinkela_wire_2),
        .a(jinkela_wire_570),
        .c(jinkela_wire_1288)
    );

    and_bi _2797_ (
        .b(jinkela_wire_1110),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_1026)
    );

    or_ii _2080_ (
        .b(jinkela_wire_915),
        .a(jinkela_wire_1288),
        .c(jinkela_wire_346)
    );

    and_bi _2798_ (
        .b(jinkela_wire_98),
        .a(io_in2_4_),
        .c(jinkela_wire_800)
    );

    inv _2081_ (
        .din(io_in1_28_),
        .dout(jinkela_wire_1091)
    );

    or_bb _2799_ (
        .b(jinkela_wire_1026),
        .a(jinkela_wire_800),
        .c(jinkela_wire_992)
    );

    or_bb _2082_ (
        .b(jinkela_wire_1091),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1353)
    );

    and_bi _2800_ (
        .b(jinkela_wire_992),
        .a(jinkela_wire_188),
        .c(jinkela_wire_33)
    );

    and_bi _2083_ (
        .b(jinkela_wire_111),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1382)
    );

    or_bb _2801_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_33),
        .c(jinkela_wire_1437)
    );

    and_bi _2084_ (
        .b(jinkela_wire_1382),
        .a(jinkela_wire_1353),
        .c(jinkela_wire_871)
    );

    and_bi _2802_ (
        .b(jinkela_wire_1437),
        .a(jinkela_wire_655),
        .c(jinkela_wire_427)
    );

    and_bi _2085_ (
        .b(jinkela_wire_871),
        .a(io_in2_0_),
        .c(jinkela_wire_216)
    );

    or_bb _2803_ (
        .b(jinkela_wire_93),
        .a(jinkela_wire_427),
        .c(io_out_14_)
    );

    and_bi _2086_ (
        .b(jinkela_wire_216),
        .a(jinkela_wire_346),
        .c(jinkela_wire_551)
    );

    and_bi _2804_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_15_),
        .c(jinkela_wire_169)
    );

    or_bb _2087_ (
        .b(jinkela_wire_15),
        .a(jinkela_wire_551),
        .c(jinkela_wire_510)
    );

    and_bi _2805_ (
        .b(jinkela_wire_846),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_414)
    );

    and_bi _2088_ (
        .b(io_in2_1_),
        .a(io_in2_0_),
        .c(jinkela_wire_201)
    );

    and_bi _2806_ (
        .b(jinkela_wire_414),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_435)
    );

    or_bb _2089_ (
        .b(jinkela_wire_964),
        .a(jinkela_wire_188),
        .c(jinkela_wire_182)
    );

    and_bi _2807_ (
        .b(jinkela_wire_435),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_901)
    );

    and_bi _2090_ (
        .b(jinkela_wire_746),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1020)
    );

    and_bi _2808_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_224),
        .c(jinkela_wire_1453)
    );

    and_bi _2091_ (
        .b(jinkela_wire_1020),
        .a(jinkela_wire_182),
        .c(jinkela_wire_905)
    );

    and_bi _2809_ (
        .b(jinkela_wire_347),
        .a(io_in1_15_),
        .c(jinkela_wire_1510)
    );

    and_bi _2092_ (
        .b(jinkela_wire_905),
        .a(jinkela_wire_201),
        .c(jinkela_wire_269)
    );

    or_bb _2810_ (
        .b(jinkela_wire_301),
        .a(jinkela_wire_1510),
        .c(jinkela_wire_404)
    );

    and_bi _2093_ (
        .b(jinkela_wire_269),
        .a(jinkela_wire_510),
        .c(jinkela_wire_1016)
    );

    or_bb _2811_ (
        .b(jinkela_wire_1453),
        .a(jinkela_wire_404),
        .c(jinkela_wire_392)
    );

    or_ii _2094_ (
        .b(jinkela_wire_1300),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1372)
    );

    and_bi _2812_ (
        .b(jinkela_wire_301),
        .a(jinkela_wire_349),
        .c(jinkela_wire_325)
    );

    and_bi _2095_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_560),
        .c(jinkela_wire_985)
    );

    and_bi _2813_ (
        .b(jinkela_wire_325),
        .a(jinkela_wire_1510),
        .c(jinkela_wire_1438)
    );

    or_bb _2096_ (
        .b(jinkela_wire_1038),
        .a(jinkela_wire_985),
        .c(jinkela_wire_142)
    );

    and_bi _2814_ (
        .b(jinkela_wire_1438),
        .a(jinkela_wire_392),
        .c(jinkela_wire_1352)
    );

    and_bi _2097_ (
        .b(jinkela_wire_142),
        .a(jinkela_wire_1372),
        .c(jinkela_wire_1216)
    );

    and_bi _2815_ (
        .b(jinkela_wire_1352),
        .a(jinkela_wire_44),
        .c(jinkela_wire_522)
    );

    or_bb _2098_ (
        .b(io_in2_2_),
        .a(jinkela_wire_1216),
        .c(jinkela_wire_131)
    );

    or_bb _2816_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_522),
        .c(jinkela_wire_466)
    );

    and_bi _2099_ (
        .b(jinkela_wire_131),
        .a(jinkela_wire_1016),
        .c(jinkela_wire_1254)
    );

    or_bb _2817_ (
        .b(jinkela_wire_901),
        .a(jinkela_wire_466),
        .c(jinkela_wire_1452)
    );

    or_bb _2100_ (
        .b(jinkela_wire_1374),
        .a(jinkela_wire_1254),
        .c(jinkela_wire_592)
    );

    and_bi _2818_ (
        .b(jinkela_wire_29),
        .a(jinkela_wire_1424),
        .c(jinkela_wire_1113)
    );

    and_bi _2101_ (
        .b(jinkela_wire_592),
        .a(jinkela_wire_804),
        .c(jinkela_wire_1448)
    );

    and_bi _2819_ (
        .b(jinkela_wire_1113),
        .a(io_in2_4_),
        .c(jinkela_wire_537)
    );

    and_bi _2102_ (
        .b(jinkela_wire_1448),
        .a(jinkela_wire_467),
        .c(jinkela_wire_961)
    );

    or_ii _2820_ (
        .b(jinkela_wire_618),
        .a(jinkela_wire_537),
        .c(jinkela_wire_644)
    );

    and_bi _2103_ (
        .b(jinkela_wire_961),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_318)
    );

    or_ii _2821_ (
        .b(io_in2_3_),
        .a(jinkela_wire_596),
        .c(jinkela_wire_576)
    );

    and_bi _2104_ (
        .b(jinkela_wire_188),
        .a(io_in1_15_),
        .c(jinkela_wire_765)
    );

    and_bi _2822_ (
        .b(jinkela_wire_1246),
        .a(jinkela_wire_804),
        .c(jinkela_wire_360)
    );

    and_bi _2105_ (
        .b(jinkela_wire_7),
        .a(jinkela_wire_188),
        .c(jinkela_wire_324)
    );

    or_bb _2823_ (
        .b(io_in2_4_),
        .a(jinkela_wire_360),
        .c(jinkela_wire_1011)
    );

    or_bb _2106_ (
        .b(jinkela_wire_765),
        .a(jinkela_wire_324),
        .c(jinkela_wire_1087)
    );

    and_bi _2824_ (
        .b(jinkela_wire_1011),
        .a(jinkela_wire_576),
        .c(jinkela_wire_38)
    );

    or_ii _2107_ (
        .b(jinkela_wire_915),
        .a(jinkela_wire_1087),
        .c(jinkela_wire_1184)
    );

    and_bi _2825_ (
        .b(jinkela_wire_38),
        .a(jinkela_wire_644),
        .c(jinkela_wire_1028)
    );

    or_bb _2108_ (
        .b(jinkela_wire_1073),
        .a(jinkela_wire_188),
        .c(jinkela_wire_890)
    );

    and_bb _2826_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1028),
        .c(jinkela_wire_533)
    );

    and_bi _2109_ (
        .b(jinkela_wire_899),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1101)
    );

    or_bb _2827_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_533),
        .c(jinkela_wire_208)
    );

    and_bi _2110_ (
        .b(jinkela_wire_1101),
        .a(jinkela_wire_890),
        .c(jinkela_wire_378)
    );

    and_bi _2828_ (
        .b(jinkela_wire_208),
        .a(jinkela_wire_1452),
        .c(jinkela_wire_704)
    );

    and_bi _2111_ (
        .b(jinkela_wire_378),
        .a(io_in2_0_),
        .c(jinkela_wire_1032)
    );

    or_bb _2829_ (
        .b(jinkela_wire_169),
        .a(jinkela_wire_704),
        .c(io_out_15_)
    );

    and_bi _2112_ (
        .b(jinkela_wire_1032),
        .a(jinkela_wire_1184),
        .c(jinkela_wire_45)
    );

    and_bi _2830_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_16_),
        .c(jinkela_wire_1027)
    );

    or_bb _2113_ (
        .b(io_in2_1_),
        .a(jinkela_wire_45),
        .c(jinkela_wire_386)
    );

    and_bi _2831_ (
        .b(jinkela_wire_1028),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_1063)
    );

    or_bb _2114_ (
        .b(jinkela_wire_78),
        .a(jinkela_wire_188),
        .c(jinkela_wire_481)
    );

    and_bi _2622_ (
        .b(jinkela_wire_56),
        .a(jinkela_wire_748),
        .c(jinkela_wire_596)
    );

    and_bi _1905_ (
        .b(jinkela_wire_1441),
        .a(jinkela_wire_606),
        .c(jinkela_wire_1126)
    );

    and_bi _2623_ (
        .b(jinkela_wire_596),
        .a(jinkela_wire_804),
        .c(jinkela_wire_673)
    );

    or_ii _1906_ (
        .b(jinkela_wire_243),
        .a(jinkela_wire_1126),
        .c(jinkela_wire_1075)
    );

    and_bi _2624_ (
        .b(jinkela_wire_1338),
        .a(jinkela_wire_1424),
        .c(jinkela_wire_1457)
    );

    or_bb _1907_ (
        .b(jinkela_wire_243),
        .a(jinkela_wire_1126),
        .c(jinkela_wire_730)
    );

    or_bb _2625_ (
        .b(jinkela_wire_804),
        .a(jinkela_wire_1457),
        .c(jinkela_wire_682)
    );

    or_ii _1908_ (
        .b(jinkela_wire_1075),
        .a(jinkela_wire_730),
        .c(io_adder_out_17_)
    );

    and_bi _2626_ (
        .b(jinkela_wire_682),
        .a(jinkela_wire_618),
        .c(jinkela_wire_1297)
    );

    and_bi _1909_ (
        .b(jinkela_wire_409),
        .a(jinkela_wire_545),
        .c(jinkela_wire_389)
    );

    or_bb _2627_ (
        .b(jinkela_wire_673),
        .a(jinkela_wire_1297),
        .c(jinkela_wire_894)
    );

    or_bb _1910_ (
        .b(jinkela_wire_1481),
        .a(jinkela_wire_389),
        .c(jinkela_wire_261)
    );

    and_bi _2628_ (
        .b(jinkela_wire_894),
        .a(io_in2_4_),
        .c(jinkela_wire_413)
    );

    and_bb _1911_ (
        .b(jinkela_wire_1481),
        .a(jinkela_wire_389),
        .c(jinkela_wire_1106)
    );

    or_bb _2629_ (
        .b(jinkela_wire_1312),
        .a(jinkela_wire_413),
        .c(jinkela_wire_866)
    );

    and_bi _1912_ (
        .b(jinkela_wire_1106),
        .a(jinkela_wire_261),
        .c(io_adder_out_16_)
    );

    and_bb _2630_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_866),
        .c(jinkela_wire_1188)
    );

    and_bi _1913_ (
        .b(jinkela_wire_222),
        .a(jinkela_wire_30),
        .c(jinkela_wire_357)
    );

    or_bb _2631_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1188),
        .c(jinkela_wire_1263)
    );

    and_bi _1914_ (
        .b(jinkela_wire_357),
        .a(jinkela_wire_563),
        .c(jinkela_wire_1050)
    );

    and_bi _2632_ (
        .b(jinkela_wire_1263),
        .a(jinkela_wire_252),
        .c(jinkela_wire_1034)
    );

    and_bi _1915_ (
        .b(jinkela_wire_563),
        .a(jinkela_wire_357),
        .c(jinkela_wire_1169)
    );

    or_bb _2633_ (
        .b(jinkela_wire_1197),
        .a(jinkela_wire_1034),
        .c(io_out_7_)
    );

    or_bb _1916_ (
        .b(jinkela_wire_1050),
        .a(jinkela_wire_1169),
        .c(io_adder_out_15_)
    );

    and_bi _2634_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_8_),
        .c(jinkela_wire_55)
    );

    and_bi _1917_ (
        .b(jinkela_wire_1446),
        .a(jinkela_wire_893),
        .c(jinkela_wire_696)
    );

    and_bi _2635_ (
        .b(io_in2_4_),
        .a(jinkela_wire_894),
        .c(jinkela_wire_668)
    );

    or_ii _1918_ (
        .b(jinkela_wire_790),
        .a(jinkela_wire_696),
        .c(jinkela_wire_742)
    );

    and_bi _2636_ (
        .b(jinkela_wire_668),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_1309)
    );

    or_bb _1919_ (
        .b(jinkela_wire_790),
        .a(jinkela_wire_696),
        .c(jinkela_wire_1092)
    );

    and_bi _2637_ (
        .b(jinkela_wire_1309),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_60)
    );

    and_bb _1920_ (
        .b(jinkela_wire_742),
        .a(jinkela_wire_1092),
        .c(io_adder_out_14_)
    );

    and_bi _2638_ (
        .b(jinkela_wire_347),
        .a(io_in1_8_),
        .c(jinkela_wire_99)
    );

    and_bb _1921_ (
        .b(jinkela_wire_1251),
        .a(jinkela_wire_789),
        .c(jinkela_wire_1293)
    );

    and_bi _2639_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_391),
        .c(jinkela_wire_1370)
    );

    and_bb _1922_ (
        .b(jinkela_wire_1251),
        .a(jinkela_wire_1029),
        .c(jinkela_wire_6)
    );

    and_bi _2640_ (
        .b(jinkela_wire_1370),
        .a(io_in2_8_),
        .c(jinkela_wire_843)
    );

    and_bi _1923_ (
        .b(jinkela_wire_6),
        .a(jinkela_wire_395),
        .c(jinkela_wire_715)
    );

    or_bb _2641_ (
        .b(jinkela_wire_99),
        .a(jinkela_wire_843),
        .c(jinkela_wire_86)
    );

    or_bb _1924_ (
        .b(jinkela_wire_1293),
        .a(jinkela_wire_715),
        .c(io_adder_out_13_)
    );

    and_bb _2642_ (
        .b(io_in2_8_),
        .a(jinkela_wire_349),
        .c(jinkela_wire_164)
    );

    and_bi _1925_ (
        .b(jinkela_wire_1506),
        .a(jinkela_wire_669),
        .c(jinkela_wire_11)
    );

    and_bb _2643_ (
        .b(jinkela_wire_99),
        .a(jinkela_wire_164),
        .c(jinkela_wire_76)
    );

    or_ii _1926_ (
        .b(jinkela_wire_634),
        .a(jinkela_wire_11),
        .c(jinkela_wire_819)
    );

    or_bb _2644_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_76),
        .c(jinkela_wire_906)
    );

    or_bb _1927_ (
        .b(jinkela_wire_634),
        .a(jinkela_wire_11),
        .c(jinkela_wire_1376)
    );

    and_bi _2645_ (
        .b(jinkela_wire_906),
        .a(jinkela_wire_86),
        .c(jinkela_wire_1155)
    );

    and_bb _1928_ (
        .b(jinkela_wire_819),
        .a(jinkela_wire_1376),
        .c(io_adder_out_12_)
    );

    or_bb _2646_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1155),
        .c(jinkela_wire_1255)
    );

    and_bb _1929_ (
        .b(jinkela_wire_1326),
        .a(jinkela_wire_993),
        .c(jinkela_wire_956)
    );

    or_bb _2647_ (
        .b(jinkela_wire_60),
        .a(jinkela_wire_1255),
        .c(jinkela_wire_471)
    );

    and_bb _1930_ (
        .b(jinkela_wire_1326),
        .a(jinkela_wire_153),
        .c(jinkela_wire_845)
    );

    and_bi _2648_ (
        .b(jinkela_wire_1107),
        .a(jinkela_wire_804),
        .c(jinkela_wire_513)
    );

    and_bi _1931_ (
        .b(jinkela_wire_845),
        .a(jinkela_wire_1177),
        .c(jinkela_wire_1321)
    );

    and_bi _2649_ (
        .b(jinkela_wire_1399),
        .a(io_in2_3_),
        .c(jinkela_wire_1194)
    );

    or_bb _1932_ (
        .b(jinkela_wire_956),
        .a(jinkela_wire_1321),
        .c(io_adder_out_11_)
    );

    or_bb _2650_ (
        .b(jinkela_wire_513),
        .a(jinkela_wire_1194),
        .c(jinkela_wire_83)
    );

    and_bi _1933_ (
        .b(jinkela_wire_503),
        .a(jinkela_wire_889),
        .c(jinkela_wire_695)
    );

    and_bi _2651_ (
        .b(jinkela_wire_83),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_720)
    );

    or_bb _1934_ (
        .b(jinkela_wire_232),
        .a(jinkela_wire_695),
        .c(jinkela_wire_741)
    );

    and_bi _2652_ (
        .b(jinkela_wire_566),
        .a(io_in2_4_),
        .c(jinkela_wire_654)
    );

    and_bb _1935_ (
        .b(jinkela_wire_232),
        .a(jinkela_wire_695),
        .c(jinkela_wire_289)
    );

    or_bb _2653_ (
        .b(jinkela_wire_720),
        .a(jinkela_wire_654),
        .c(jinkela_wire_1366)
    );

    and_bi _1936_ (
        .b(jinkela_wire_289),
        .a(jinkela_wire_741),
        .c(io_adder_out_10_)
    );

    and_bi _2654_ (
        .b(jinkela_wire_1366),
        .a(jinkela_wire_188),
        .c(jinkela_wire_571)
    );

    and_bi _1937_ (
        .b(jinkela_wire_264),
        .a(jinkela_wire_994),
        .c(jinkela_wire_426)
    );

    or_bb _2655_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_571),
        .c(jinkela_wire_585)
    );

    and_bi _1938_ (
        .b(jinkela_wire_426),
        .a(jinkela_wire_630),
        .c(jinkela_wire_891)
    );

    and_bi _2656_ (
        .b(jinkela_wire_585),
        .a(jinkela_wire_471),
        .c(jinkela_wire_1218)
    );

    and_bi _1939_ (
        .b(jinkela_wire_630),
        .a(jinkela_wire_426),
        .c(jinkela_wire_796)
    );

    or_bb _2657_ (
        .b(jinkela_wire_55),
        .a(jinkela_wire_1218),
        .c(io_out_8_)
    );

    or_bb _1940_ (
        .b(jinkela_wire_891),
        .a(jinkela_wire_796),
        .c(io_adder_out_9_)
    );

    and_bi _2658_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_9_),
        .c(jinkela_wire_850)
    );

    and_bi _1941_ (
        .b(jinkela_wire_609),
        .a(jinkela_wire_807),
        .c(jinkela_wire_681)
    );

    and_bi _2659_ (
        .b(jinkela_wire_787),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_1439)
    );

    or_bb _1942_ (
        .b(jinkela_wire_1463),
        .a(jinkela_wire_681),
        .c(jinkela_wire_1013)
    );

    and_bi _2660_ (
        .b(jinkela_wire_1439),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_885)
    );

    and_bb _1943_ (
        .b(jinkela_wire_1463),
        .a(jinkela_wire_681),
        .c(jinkela_wire_73)
    );

    and_bi _2661_ (
        .b(jinkela_wire_885),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_23)
    );

    and_bi _1944_ (
        .b(jinkela_wire_73),
        .a(jinkela_wire_1013),
        .c(io_adder_out_8_)
    );

    and_bi _2662_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_293),
        .c(jinkela_wire_191)
    );

    and_bi _1945_ (
        .b(jinkela_wire_1462),
        .a(jinkela_wire_148),
        .c(jinkela_wire_1410)
    );

    and_bi _2663_ (
        .b(jinkela_wire_347),
        .a(io_in1_9_),
        .c(jinkela_wire_141)
    );

    and_bi _1946_ (
        .b(jinkela_wire_1479),
        .a(jinkela_wire_1410),
        .c(jinkela_wire_593)
    );

    and_bi _2451_ (
        .b(jinkela_wire_610),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_390)
    );

    or_bb _2452_ (
        .b(io_in2_1_),
        .a(jinkela_wire_1088),
        .c(jinkela_wire_403)
    );

    and_bi _2453_ (
        .b(jinkela_wire_1287),
        .a(io_in2_1_),
        .c(jinkela_wire_1200)
    );

    and_bi _2454_ (
        .b(jinkela_wire_1200),
        .a(jinkela_wire_403),
        .c(jinkela_wire_479)
    );

    or_bb _2455_ (
        .b(io_in2_2_),
        .a(jinkela_wire_479),
        .c(jinkela_wire_803)
    );

    or_bb _2456_ (
        .b(io_in2_1_),
        .a(jinkela_wire_160),
        .c(jinkela_wire_1035)
    );

    and_bi _2457_ (
        .b(jinkela_wire_361),
        .a(io_in2_1_),
        .c(jinkela_wire_788)
    );

    and_bi _2458_ (
        .b(jinkela_wire_788),
        .a(jinkela_wire_1035),
        .c(jinkela_wire_1010)
    );

    and_bi _2459_ (
        .b(jinkela_wire_1010),
        .a(io_in2_2_),
        .c(jinkela_wire_924)
    );

    and_bi _2460_ (
        .b(jinkela_wire_924),
        .a(jinkela_wire_803),
        .c(jinkela_wire_1115)
    );

    or_bb _2461_ (
        .b(io_in2_3_),
        .a(jinkela_wire_1115),
        .c(jinkela_wire_1400)
    );

    and_bi _2462_ (
        .b(io_fn_3_),
        .a(jinkela_wire_1038),
        .c(jinkela_wire_1204)
    );

    and_bi _2463_ (
        .b(jinkela_wire_1204),
        .a(jinkela_wire_618),
        .c(jinkela_wire_909)
    );

    and_bi _2464_ (
        .b(jinkela_wire_909),
        .a(io_in2_2_),
        .c(jinkela_wire_174)
    );

    and_bi _2465_ (
        .b(jinkela_wire_1387),
        .a(jinkela_wire_15),
        .c(jinkela_wire_209)
    );

    and_bi _2466_ (
        .b(jinkela_wire_15),
        .a(jinkela_wire_929),
        .c(jinkela_wire_927)
    );

    or_bb _2467_ (
        .b(jinkela_wire_209),
        .a(jinkela_wire_927),
        .c(jinkela_wire_12)
    );

    and_bi _2468_ (
        .b(jinkela_wire_12),
        .a(jinkela_wire_158),
        .c(jinkela_wire_1127)
    );

    or_bb _2469_ (
        .b(jinkela_wire_174),
        .a(jinkela_wire_1127),
        .c(jinkela_wire_92)
    );

    and_bi _2470_ (
        .b(jinkela_wire_92),
        .a(io_in2_3_),
        .c(jinkela_wire_734)
    );

    and_bi _2471_ (
        .b(jinkela_wire_734),
        .a(jinkela_wire_1400),
        .c(jinkela_wire_1162)
    );

    and_bi _2472_ (
        .b(jinkela_wire_1162),
        .a(io_in2_4_),
        .c(jinkela_wire_253)
    );

    or_bb _2473_ (
        .b(jinkela_wire_390),
        .a(jinkela_wire_253),
        .c(jinkela_wire_291)
    );

    and_bi _2474_ (
        .b(jinkela_wire_291),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1378)
    );

    or_bb _2475_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1378),
        .c(jinkela_wire_499)
    );

    and_bi _2476_ (
        .b(jinkela_wire_499),
        .a(jinkela_wire_273),
        .c(jinkela_wire_104)
    );

    or_bb _2477_ (
        .b(jinkela_wire_640),
        .a(jinkela_wire_104),
        .c(io_out_3_)
    );

    and_bi _2478_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_4_),
        .c(jinkela_wire_1349)
    );

    and_bi _2479_ (
        .b(jinkela_wire_92),
        .a(jinkela_wire_804),
        .c(jinkela_wire_1315)
    );

    and_bi _2480_ (
        .b(jinkela_wire_1315),
        .a(jinkela_wire_1269),
        .c(jinkela_wire_107)
    );

    and_bi _2481_ (
        .b(jinkela_wire_107),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_134)
    );

    and_bi _2482_ (
        .b(jinkela_wire_134),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_476)
    );

    and_bi _2483_ (
        .b(jinkela_wire_476),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_382)
    );

    and_bi _2484_ (
        .b(jinkela_wire_1248),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_449)
    );

    or_bb _2485_ (
        .b(io_in1_4_),
        .a(jinkela_wire_449),
        .c(jinkela_wire_514)
    );

    and_bb _2486_ (
        .b(io_in1_4_),
        .a(io_in2_4_),
        .c(jinkela_wire_548)
    );

    and_bb _2487_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_548),
        .c(jinkela_wire_105)
    );

    and_bi _2488_ (
        .b(jinkela_wire_105),
        .a(jinkela_wire_514),
        .c(jinkela_wire_896)
    );

    or_bb _2489_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_896),
        .c(jinkela_wire_275)
    );

    and_bi _2490_ (
        .b(jinkela_wire_548),
        .a(jinkela_wire_347),
        .c(jinkela_wire_477)
    );

    or_bb _2491_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_477),
        .c(jinkela_wire_425)
    );

    and_bi _2492_ (
        .b(jinkela_wire_425),
        .a(jinkela_wire_275),
        .c(jinkela_wire_1504)
    );

    inv _1566_ (
        .din(io_in1_26_),
        .dout(jinkela_wire_562)
    );

    or_bb _1737_ (
        .b(io_in1_18_),
        .a(jinkela_wire_984),
        .c(jinkela_wire_983)
    );

    and_bi _2283_ (
        .b(jinkela_wire_236),
        .a(io_in2_0_),
        .c(jinkela_wire_462)
    );

    inv _1567_ (
        .din(io_in1_25_),
        .dout(jinkela_wire_1241)
    );

    and_bi _1738_ (
        .b(jinkela_wire_145),
        .a(io_fn_3_),
        .c(jinkela_wire_260)
    );

    and_bi _2284_ (
        .b(jinkela_wire_462),
        .a(jinkela_wire_590),
        .c(jinkela_wire_1473)
    );

    inv _1568_ (
        .din(io_in1_23_),
        .dout(jinkela_wire_268)
    );

    and_bi _1739_ (
        .b(io_in2_18_),
        .a(jinkela_wire_260),
        .c(jinkela_wire_106)
    );

    and_bi _2285_ (
        .b(jinkela_wire_1473),
        .a(jinkela_wire_15),
        .c(jinkela_wire_498)
    );

    inv _1569_ (
        .din(io_in1_17_),
        .dout(jinkela_wire_899)
    );

    and_bi _1740_ (
        .b(jinkela_wire_260),
        .a(io_in2_18_),
        .c(jinkela_wire_320)
    );

    or_bb _2286_ (
        .b(io_in2_0_),
        .a(jinkela_wire_955),
        .c(jinkela_wire_1402)
    );

    inv _1570_ (
        .din(io_in1_13_),
        .dout(jinkela_wire_78)
    );

    or_bb _1741_ (
        .b(jinkela_wire_106),
        .a(jinkela_wire_320),
        .c(jinkela_wire_1086)
    );

    and_bi _2287_ (
        .b(jinkela_wire_737),
        .a(io_in2_0_),
        .c(jinkela_wire_194)
    );

    inv _1571_ (
        .din(io_in1_11_),
        .dout(jinkela_wire_719)
    );

    and_bb _1742_ (
        .b(jinkela_wire_983),
        .a(jinkela_wire_1086),
        .c(jinkela_wire_623)
    );

    and_bi _2288_ (
        .b(jinkela_wire_194),
        .a(jinkela_wire_1402),
        .c(jinkela_wire_258)
    );

    inv _1572_ (
        .din(io_in1_7_),
        .dout(jinkela_wire_95)
    );

    and_bi _1743_ (
        .b(jinkela_wire_623),
        .a(jinkela_wire_271),
        .c(jinkela_wire_1083)
    );

    and_bi _2289_ (
        .b(jinkela_wire_258),
        .a(io_in2_1_),
        .c(jinkela_wire_943)
    );

    inv _1573_ (
        .din(io_in1_1_),
        .dout(jinkela_wire_746)
    );

    and_bi _1744_ (
        .b(io_in1_19_),
        .a(jinkela_wire_1083),
        .c(jinkela_wire_1114)
    );

    or_bb _2290_ (
        .b(jinkela_wire_498),
        .a(jinkela_wire_943),
        .c(jinkela_wire_1294)
    );

    and_bb _1574_ (
        .b(io_in1_0_),
        .a(io_in2_0_),
        .c(jinkela_wire_394)
    );

    inv _1745_ (
        .din(io_in1_19_),
        .dout(jinkela_wire_842)
    );

    and_bi _2291_ (
        .b(jinkela_wire_1294),
        .a(io_in2_2_),
        .c(jinkela_wire_197)
    );

    and_bi _1575_ (
        .b(jinkela_wire_394),
        .a(jinkela_wire_746),
        .c(jinkela_wire_115)
    );

    or_bb _1746_ (
        .b(jinkela_wire_842),
        .a(jinkela_wire_1083),
        .c(jinkela_wire_1264)
    );

    or_bb _2292_ (
        .b(jinkela_wire_1514),
        .a(jinkela_wire_197),
        .c(jinkela_wire_1023)
    );

    or_ii _1576_ (
        .b(io_in1_1_),
        .a(jinkela_wire_394),
        .c(jinkela_wire_119)
    );

    inv _1747_ (
        .din(io_in2_19_),
        .dout(jinkela_wire_616)
    );

    and_bi _2293_ (
        .b(jinkela_wire_1023),
        .a(jinkela_wire_804),
        .c(jinkela_wire_1373)
    );

    and_bi _1577_ (
        .b(io_fn_3_),
        .a(io_in2_1_),
        .c(jinkela_wire_1143)
    );

    and_bi _1748_ (
        .b(jinkela_wire_957),
        .a(io_fn_3_),
        .c(jinkela_wire_1322)
    );

    and_bi _2294_ (
        .b(jinkela_wire_1373),
        .a(jinkela_wire_507),
        .c(jinkela_wire_122)
    );

    or_ii _1578_ (
        .b(io_in2_0_),
        .a(io_in2_1_),
        .c(jinkela_wire_642)
    );

    and_bi _1749_ (
        .b(jinkela_wire_616),
        .a(jinkela_wire_1322),
        .c(jinkela_wire_670)
    );

    and_bi _2295_ (
        .b(jinkela_wire_122),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_762)
    );

    or_ii _1579_ (
        .b(io_fn_3_),
        .a(jinkela_wire_1038),
        .c(jinkela_wire_14)
    );

    and_bi _1750_ (
        .b(jinkela_wire_1322),
        .a(jinkela_wire_616),
        .c(jinkela_wire_1501)
    );

    or_bb _2296_ (
        .b(io_in2_0_),
        .a(jinkela_wire_378),
        .c(jinkela_wire_430)
    );

    and_bi _1580_ (
        .b(jinkela_wire_14),
        .a(jinkela_wire_642),
        .c(jinkela_wire_475)
    );

    or_bb _1751_ (
        .b(jinkela_wire_670),
        .a(jinkela_wire_1501),
        .c(jinkela_wire_1211)
    );

    and_bi _2297_ (
        .b(jinkela_wire_1256),
        .a(io_in2_0_),
        .c(jinkela_wire_914)
    );

    or_bb _1581_ (
        .b(jinkela_wire_1143),
        .a(jinkela_wire_475),
        .c(jinkela_wire_1509)
    );

    inv _1752_ (
        .din(jinkela_wire_1211),
        .dout(jinkela_wire_237)
    );

    and_bi _2298_ (
        .b(jinkela_wire_914),
        .a(jinkela_wire_430),
        .c(jinkela_wire_811)
    );

    and_bi _1582_ (
        .b(jinkela_wire_1509),
        .a(jinkela_wire_119),
        .c(jinkela_wire_364)
    );

    and_bi _1753_ (
        .b(jinkela_wire_237),
        .a(jinkela_wire_1264),
        .c(jinkela_wire_1488)
    );

    or_bb _2299_ (
        .b(io_in2_1_),
        .a(jinkela_wire_811),
        .c(jinkela_wire_230)
    );

    or_bb _1583_ (
        .b(jinkela_wire_115),
        .a(jinkela_wire_364),
        .c(jinkela_wire_234)
    );

    or_bb _1754_ (
        .b(jinkela_wire_1114),
        .a(jinkela_wire_1488),
        .c(jinkela_wire_1354)
    );

    or_bb _2300_ (
        .b(io_in2_0_),
        .a(jinkela_wire_353),
        .c(jinkela_wire_108)
    );

    and_bi _1584_ (
        .b(io_in1_2_),
        .a(jinkela_wire_234),
        .c(jinkela_wire_127)
    );

    and_bi _1755_ (
        .b(io_in1_20_),
        .a(jinkela_wire_1354),
        .c(jinkela_wire_270)
    );

    and_bi _2301_ (
        .b(jinkela_wire_1494),
        .a(io_in2_0_),
        .c(jinkela_wire_225)
    );

    inv _1585_ (
        .din(io_in1_2_),
        .dout(jinkela_wire_958)
    );

    inv _1756_ (
        .din(io_in1_20_),
        .dout(jinkela_wire_1329)
    );

    and_bi _2302_ (
        .b(jinkela_wire_225),
        .a(jinkela_wire_108),
        .c(jinkela_wire_1088)
    );

    or_bb _1586_ (
        .b(jinkela_wire_958),
        .a(jinkela_wire_234),
        .c(jinkela_wire_779)
    );

    or_bb _1757_ (
        .b(jinkela_wire_1329),
        .a(jinkela_wire_1354),
        .c(jinkela_wire_656)
    );

    and_bi _2303_ (
        .b(jinkela_wire_1088),
        .a(io_in2_1_),
        .c(jinkela_wire_1467)
    );

    and_bi _1587_ (
        .b(jinkela_wire_14),
        .a(jinkela_wire_158),
        .c(jinkela_wire_519)
    );

    and_bi _1758_ (
        .b(jinkela_wire_1186),
        .a(io_fn_3_),
        .c(jinkela_wire_1017)
    );

    and_bi _2304_ (
        .b(jinkela_wire_1467),
        .a(jinkela_wire_230),
        .c(jinkela_wire_647)
    );

    and_bi _1588_ (
        .b(jinkela_wire_158),
        .a(jinkela_wire_14),
        .c(jinkela_wire_329)
    );

    and_bi _1759_ (
        .b(io_in2_20_),
        .a(jinkela_wire_1017),
        .c(jinkela_wire_1030)
    );

    or_bb _2305_ (
        .b(io_in2_2_),
        .a(jinkela_wire_647),
        .c(jinkela_wire_128)
    );

    or_bb _1589_ (
        .b(jinkela_wire_519),
        .a(jinkela_wire_329),
        .c(jinkela_wire_755)
    );

    and_bi _1760_ (
        .b(jinkela_wire_1017),
        .a(io_in2_20_),
        .c(jinkela_wire_1318)
    );

    or_bb _2306_ (
        .b(io_in2_0_),
        .a(jinkela_wire_179),
        .c(jinkela_wire_613)
    );

    and_bi _1590_ (
        .b(jinkela_wire_755),
        .a(jinkela_wire_779),
        .c(jinkela_wire_171)
    );

    or_bb _1761_ (
        .b(jinkela_wire_1030),
        .a(jinkela_wire_1318),
        .c(jinkela_wire_847)
    );

    and_bi _2307_ (
        .b(jinkela_wire_1171),
        .a(io_in2_0_),
        .c(jinkela_wire_692)
    );

    or_bb _1591_ (
        .b(jinkela_wire_127),
        .a(jinkela_wire_171),
        .c(jinkela_wire_1190)
    );

    and_bi _1762_ (
        .b(jinkela_wire_847),
        .a(jinkela_wire_656),
        .c(jinkela_wire_1298)
    );

    and_bi _2308_ (
        .b(jinkela_wire_692),
        .a(jinkela_wire_613),
        .c(jinkela_wire_1287)
    );

    and_bi _1592_ (
        .b(io_in1_3_),
        .a(jinkela_wire_1190),
        .c(jinkela_wire_1061)
    );

    or_bb _1763_ (
        .b(jinkela_wire_270),
        .a(jinkela_wire_1298),
        .c(jinkela_wire_711)
    );

    or_bb _2309_ (
        .b(io_in2_1_),
        .a(jinkela_wire_1287),
        .c(jinkela_wire_710)
    );

    inv _1593_ (
        .din(io_in1_3_),
        .dout(jinkela_wire_111)
    );

    and_bi _1764_ (
        .b(io_in1_21_),
        .a(jinkela_wire_711),
        .c(jinkela_wire_1230)
    );

    or_bb _2310_ (
        .b(io_in2_0_),
        .a(jinkela_wire_356),
        .c(jinkela_wire_469)
    );

    or_bb _1594_ (
        .b(jinkela_wire_111),
        .a(jinkela_wire_1190),
        .c(jinkela_wire_310)
    );

    inv _1765_ (
        .din(io_in1_21_),
        .dout(jinkela_wire_1253)
    );

    and_bi _2311_ (
        .b(jinkela_wire_1134),
        .a(io_in2_0_),
        .c(jinkela_wire_1203)
    );

    inv _1595_ (
        .din(io_in2_3_),
        .dout(jinkela_wire_804)
    );

    or_bb _1766_ (
        .b(jinkela_wire_1253),
        .a(jinkela_wire_711),
        .c(jinkela_wire_684)
    );

    and_bi _2312_ (
        .b(jinkela_wire_1203),
        .a(jinkela_wire_469),
        .c(jinkela_wire_160)
    );

    and_bi _1596_ (
        .b(jinkela_wire_1338),
        .a(io_fn_3_),
        .c(jinkela_wire_778)
    );

    inv _1767_ (
        .din(io_in2_21_),
        .dout(jinkela_wire_244)
    );

    and_bi _2313_ (
        .b(jinkela_wire_160),
        .a(io_in2_1_),
        .c(jinkela_wire_1282)
    );

    and_bi _1597_ (
        .b(jinkela_wire_804),
        .a(jinkela_wire_778),
        .c(jinkela_wire_309)
    );

    and_bi _1768_ (
        .b(jinkela_wire_154),
        .a(io_fn_3_),
        .c(jinkela_wire_221)
    );

    and_bi _2314_ (
        .b(jinkela_wire_1282),
        .a(jinkela_wire_710),
        .c(jinkela_wire_745)
    );

    and_bi _1598_ (
        .b(jinkela_wire_778),
        .a(jinkela_wire_804),
        .c(jinkela_wire_62)
    );

    and_bi _1769_ (
        .b(jinkela_wire_244),
        .a(jinkela_wire_221),
        .c(jinkela_wire_702)
    );

    and_bi _2315_ (
        .b(jinkela_wire_745),
        .a(io_in2_2_),
        .c(jinkela_wire_297)
    );

    or_bb _1599_ (
        .b(jinkela_wire_309),
        .a(jinkela_wire_62),
        .c(jinkela_wire_888)
    );

    and_bi _1770_ (
        .b(jinkela_wire_221),
        .a(jinkela_wire_244),
        .c(jinkela_wire_743)
    );

    and_bi _2316_ (
        .b(jinkela_wire_297),
        .a(jinkela_wire_128),
        .c(jinkela_wire_1461)
    );

    inv _1600_ (
        .din(jinkela_wire_888),
        .dout(jinkela_wire_24)
    );

    or_bb _1771_ (
        .b(jinkela_wire_702),
        .a(jinkela_wire_743),
        .c(jinkela_wire_665)
    );

    or_bb _2317_ (
        .b(io_in2_3_),
        .a(jinkela_wire_1461),
        .c(jinkela_wire_123)
    );

    and_bi _1601_ (
        .b(jinkela_wire_24),
        .a(jinkela_wire_310),
        .c(jinkela_wire_1109)
    );

    inv _1772_ (
        .din(jinkela_wire_665),
        .dout(jinkela_wire_1244)
    );

    or_bb _2318_ (
        .b(io_in2_0_),
        .a(jinkela_wire_274),
        .c(jinkela_wire_771)
    );

    or_bb _1602_ (
        .b(jinkela_wire_1061),
        .a(jinkela_wire_1109),
        .c(jinkela_wire_454)
    );

    and_bi _1773_ (
        .b(jinkela_wire_1244),
        .a(jinkela_wire_684),
        .c(jinkela_wire_854)
    );

    and_bi _2319_ (
        .b(jinkela_wire_1336),
        .a(io_in2_0_),
        .c(jinkela_wire_1426)
    );

    and_bi _2320_ (
        .b(jinkela_wire_1426),
        .a(jinkela_wire_771),
        .c(jinkela_wire_361)
    );

    and_bi _1603_ (
        .b(io_in1_4_),
        .a(jinkela_wire_454),
        .c(jinkela_wire_1103)
    );

    or_bb _1774_ (
        .b(jinkela_wire_1230),
        .a(jinkela_wire_854),
        .c(jinkela_wire_27)
    );

    or_bb _2321_ (
        .b(io_in2_1_),
        .a(jinkela_wire_361),
        .c(jinkela_wire_1443)
    );

    inv _1604_ (
        .din(io_in1_4_),
        .dout(jinkela_wire_1174)
    );

    and_bi _1775_ (
        .b(jinkela_wire_27),
        .a(io_in1_22_),
        .c(jinkela_wire_1096)
    );

    or_bb _2322_ (
        .b(io_in2_0_),
        .a(jinkela_wire_1325),
        .c(jinkela_wire_339)
    );

    or_bb _1605_ (
        .b(jinkela_wire_1174),
        .a(jinkela_wire_454),
        .c(jinkela_wire_26)
    );

    inv _1776_ (
        .din(io_in1_22_),
        .dout(jinkela_wire_278)
    );

    and_bi _2323_ (
        .b(jinkela_wire_1144),
        .a(io_in2_0_),
        .c(jinkela_wire_1125)
    );

    or_ii _1777_ (
        .b(jinkela_wire_278),
        .a(jinkela_wire_27),
        .c(jinkela_wire_834)
    );

    and_bi _1606_ (
        .b(jinkela_wire_29),
        .a(io_fn_3_),
        .c(jinkela_wire_565)
    );

    and_bi _1778_ (
        .b(jinkela_wire_1359),
        .a(io_fn_3_),
        .c(jinkela_wire_926)
    );

    and_bi _1607_ (
        .b(io_in2_4_),
        .a(jinkela_wire_565),
        .c(jinkela_wire_525)
    );

    and_bi _2324_ (
        .b(jinkela_wire_1125),
        .a(jinkela_wire_339),
        .c(jinkela_wire_1387)
    );

    and_bi _3000_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_26_),
        .c(jinkela_wire_1356)
    );

    and_bi _3001_ (
        .b(jinkela_wire_44),
        .a(jinkela_wire_1449),
        .c(jinkela_wire_423)
    );

    or_bb _3002_ (
        .b(jinkela_wire_562),
        .a(jinkela_wire_347),
        .c(jinkela_wire_1002)
    );

    inv _3003_ (
        .din(io_in2_26_),
        .dout(jinkela_wire_1478)
    );

    and_bi _3004_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_562),
        .c(jinkela_wire_988)
    );

    or_bb _3005_ (
        .b(jinkela_wire_1478),
        .a(jinkela_wire_988),
        .c(jinkela_wire_1206)
    );

    or_ii _3006_ (
        .b(jinkela_wire_1002),
        .a(jinkela_wire_1206),
        .c(jinkela_wire_633)
    );

    and_bi _3007_ (
        .b(jinkela_wire_1478),
        .a(jinkela_wire_349),
        .c(jinkela_wire_1070)
    );

    and_bi _3008_ (
        .b(jinkela_wire_1002),
        .a(jinkela_wire_1070),
        .c(jinkela_wire_1240)
    );

    or_bb _3009_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_1240),
        .c(jinkela_wire_912)
    );

    and_bi _3010_ (
        .b(jinkela_wire_912),
        .a(jinkela_wire_633),
        .c(jinkela_wire_298)
    );

    or_bb _3011_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_298),
        .c(jinkela_wire_371)
    );

    or_bb _3012_ (
        .b(jinkela_wire_423),
        .a(jinkela_wire_371),
        .c(jinkela_wire_990)
    );

    and_bb _3013_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_295),
        .c(jinkela_wire_599)
    );

    or_bb _3014_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_599),
        .c(jinkela_wire_1371)
    );

    and_bi _3015_ (
        .b(jinkela_wire_1371),
        .a(jinkela_wire_990),
        .c(jinkela_wire_482)
    );

    or_bb _3016_ (
        .b(jinkela_wire_1356),
        .a(jinkela_wire_482),
        .c(io_out_26_)
    );

    and_bi _3017_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_27_),
        .c(jinkela_wire_699)
    );

    and_bi _3018_ (
        .b(jinkela_wire_1232),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_72)
    );

    and_bb _3019_ (
        .b(io_in2_27_),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_1512)
    );

    or_bb _3020_ (
        .b(io_in1_27_),
        .a(jinkela_wire_1512),
        .c(jinkela_wire_1436)
    );

    and_bb _3021_ (
        .b(io_in1_27_),
        .a(io_in2_27_),
        .c(jinkela_wire_1173)
    );

    and_bb _3022_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_1173),
        .c(jinkela_wire_241)
    );

    and_bi _3023_ (
        .b(jinkela_wire_241),
        .a(jinkela_wire_1436),
        .c(jinkela_wire_1006)
    );

    or_bb _3024_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_1006),
        .c(jinkela_wire_358)
    );

    and_bi _3025_ (
        .b(jinkela_wire_1173),
        .a(jinkela_wire_347),
        .c(jinkela_wire_411)
    );

    or_bb _3026_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_411),
        .c(jinkela_wire_1009)
    );

    and_bi _3027_ (
        .b(jinkela_wire_1009),
        .a(jinkela_wire_358),
        .c(jinkela_wire_1132)
    );

    or_bb _3028_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1132),
        .c(jinkela_wire_996)
    );

    or_bb _3029_ (
        .b(jinkela_wire_72),
        .a(jinkela_wire_996),
        .c(jinkela_wire_1367)
    );

    and_bb _3030_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_476),
        .c(jinkela_wire_184)
    );

    or_bb _3031_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_184),
        .c(jinkela_wire_493)
    );

    and_bi _3032_ (
        .b(jinkela_wire_493),
        .a(jinkela_wire_1367),
        .c(jinkela_wire_473)
    );

    or_bb _3033_ (
        .b(jinkela_wire_699),
        .a(jinkela_wire_473),
        .c(io_out_27_)
    );

    and_bi _3034_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_28_),
        .c(jinkela_wire_1118)
    );

    and_bi _3035_ (
        .b(jinkela_wire_44),
        .a(jinkela_wire_291),
        .c(jinkela_wire_605)
    );

    and_bb _3036_ (
        .b(io_in2_28_),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_48)
    );

    or_bb _3037_ (
        .b(io_in1_28_),
        .a(jinkela_wire_48),
        .c(jinkela_wire_1516)
    );

    and_bb _3038_ (
        .b(io_in1_28_),
        .a(io_in2_28_),
        .c(jinkela_wire_523)
    );

    and_bb _3039_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_523),
        .c(jinkela_wire_873)
    );

    and_bi _3040_ (
        .b(jinkela_wire_873),
        .a(jinkela_wire_1516),
        .c(jinkela_wire_1151)
    );

    or_bb _3041_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_1151),
        .c(jinkela_wire_485)
    );

    and_bb _2832_ (
        .b(io_in2_16_),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_1258)
    );

    or_bb _2833_ (
        .b(io_in1_16_),
        .a(jinkela_wire_1258),
        .c(jinkela_wire_979)
    );

    and_bb _2834_ (
        .b(io_in1_16_),
        .a(io_in2_16_),
        .c(jinkela_wire_1375)
    );

    and_bb _2835_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_1375),
        .c(jinkela_wire_480)
    );

    and_bi _2836_ (
        .b(jinkela_wire_480),
        .a(jinkela_wire_979),
        .c(jinkela_wire_1513)
    );

    or_bb _2837_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_1513),
        .c(jinkela_wire_857)
    );

    and_bi _2838_ (
        .b(jinkela_wire_1375),
        .a(jinkela_wire_347),
        .c(jinkela_wire_1483)
    );

    or_bb _2839_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_1483),
        .c(jinkela_wire_1153)
    );

    and_bi _2840_ (
        .b(jinkela_wire_1153),
        .a(jinkela_wire_857),
        .c(jinkela_wire_1044)
    );

    or_bb _2841_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1044),
        .c(jinkela_wire_464)
    );

    or_bb _2842_ (
        .b(jinkela_wire_1063),
        .a(jinkela_wire_464),
        .c(jinkela_wire_579)
    );

    and_bb _2843_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_435),
        .c(jinkela_wire_826)
    );

    or_bb _2844_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_826),
        .c(jinkela_wire_836)
    );

    and_bi _2845_ (
        .b(jinkela_wire_836),
        .a(jinkela_wire_579),
        .c(jinkela_wire_125)
    );

    or_bb _2846_ (
        .b(jinkela_wire_1027),
        .a(jinkela_wire_125),
        .c(io_out_16_)
    );

    and_bi _2847_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_17_),
        .c(jinkela_wire_732)
    );

    and_bi _2848_ (
        .b(jinkela_wire_44),
        .a(jinkela_wire_992),
        .c(jinkela_wire_569)
    );

    and_bi _2849_ (
        .b(jinkela_wire_34),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_1031)
    );

    or_bb _2850_ (
        .b(io_in1_17_),
        .a(jinkela_wire_1031),
        .c(jinkela_wire_220)
    );

    and_bb _2851_ (
        .b(io_in1_17_),
        .a(io_in2_17_),
        .c(jinkela_wire_1274)
    );

    and_bb _2852_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_1274),
        .c(jinkela_wire_526)
    );

    and_bi _2853_ (
        .b(jinkela_wire_526),
        .a(jinkela_wire_220),
        .c(jinkela_wire_500)
    );

    or_bb _2854_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_500),
        .c(jinkela_wire_948)
    );

    and_bi _2855_ (
        .b(jinkela_wire_1274),
        .a(jinkela_wire_347),
        .c(jinkela_wire_659)
    );

    or_bb _2856_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_659),
        .c(jinkela_wire_294)
    );

    and_bi _2857_ (
        .b(jinkela_wire_294),
        .a(jinkela_wire_948),
        .c(jinkela_wire_953)
    );

    or_bb _2858_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_953),
        .c(jinkela_wire_512)
    );

    or_bb _2859_ (
        .b(jinkela_wire_569),
        .a(jinkela_wire_512),
        .c(jinkela_wire_687)
    );

    and_bb _2860_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_991),
        .c(jinkela_wire_133)
    );

    or_bb _2861_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_133),
        .c(jinkela_wire_862)
    );

    and_bi _2862_ (
        .b(jinkela_wire_862),
        .a(jinkela_wire_687),
        .c(jinkela_wire_879)
    );

    or_bb _2863_ (
        .b(jinkela_wire_732),
        .a(jinkela_wire_879),
        .c(io_out_17_)
    );

    and_bi _2864_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_18_),
        .c(jinkela_wire_674)
    );

    and_bi _2865_ (
        .b(jinkela_wire_44),
        .a(jinkela_wire_1228),
        .c(jinkela_wire_722)
    );

    and_bb _2866_ (
        .b(io_in2_18_),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_163)
    );

    or_bb _2867_ (
        .b(io_in1_18_),
        .a(jinkela_wire_163),
        .c(jinkela_wire_1498)
    );

    and_bb _2868_ (
        .b(io_in1_18_),
        .a(io_in2_18_),
        .c(jinkela_wire_212)
    );

    and_bb _2869_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_212),
        .c(jinkela_wire_860)
    );

    and_bi _2870_ (
        .b(jinkela_wire_860),
        .a(jinkela_wire_1498),
        .c(jinkela_wire_816)
    );

    or_bb _2871_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_816),
        .c(jinkela_wire_1213)
    );

    and_bi _2872_ (
        .b(jinkela_wire_212),
        .a(jinkela_wire_347),
        .c(jinkela_wire_786)
    );

    or_bb _2873_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_786),
        .c(jinkela_wire_783)
    );

    and_bi _2115_ (
        .b(jinkela_wire_865),
        .a(jinkela_wire_188),
        .c(jinkela_wire_497)
    );

    and_bi _2116_ (
        .b(jinkela_wire_497),
        .a(jinkela_wire_481),
        .c(jinkela_wire_1256)
    );

    or_bb _2117_ (
        .b(io_in2_0_),
        .a(jinkela_wire_1256),
        .c(jinkela_wire_327)
    );

    or_bb _2118_ (
        .b(jinkela_wire_374),
        .a(jinkela_wire_188),
        .c(jinkela_wire_781)
    );

    and_bi _2119_ (
        .b(jinkela_wire_842),
        .a(jinkela_wire_188),
        .c(jinkela_wire_71)
    );

    and_bi _2120_ (
        .b(jinkela_wire_71),
        .a(jinkela_wire_781),
        .c(jinkela_wire_353)
    );

    and_bi _2121_ (
        .b(jinkela_wire_353),
        .a(io_in2_0_),
        .c(jinkela_wire_973)
    );

    and_bi _2122_ (
        .b(jinkela_wire_973),
        .a(jinkela_wire_327),
        .c(jinkela_wire_1077)
    );

    and_bi _2123_ (
        .b(jinkela_wire_1077),
        .a(io_in2_1_),
        .c(jinkela_wire_54)
    );

    and_bi _2124_ (
        .b(jinkela_wire_54),
        .a(jinkela_wire_386),
        .c(jinkela_wire_1219)
    );

    and_bi _2125_ (
        .b(jinkela_wire_1219),
        .a(jinkela_wire_158),
        .c(jinkela_wire_1324)
    );

    or_bb _2126_ (
        .b(jinkela_wire_719),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1057)
    );

    and_bi _2127_ (
        .b(jinkela_wire_1329),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1207)
    );

    and_bi _2128_ (
        .b(jinkela_wire_1207),
        .a(jinkela_wire_1057),
        .c(jinkela_wire_1494)
    );

    or_bb _2129_ (
        .b(io_in2_0_),
        .a(jinkela_wire_1494),
        .c(jinkela_wire_1511)
    );

    or_bb _2130_ (
        .b(jinkela_wire_217),
        .a(jinkela_wire_188),
        .c(jinkela_wire_855)
    );

    and_bi _2131_ (
        .b(jinkela_wire_1253),
        .a(jinkela_wire_188),
        .c(jinkela_wire_632)
    );

    and_bi _2132_ (
        .b(jinkela_wire_632),
        .a(jinkela_wire_855),
        .c(jinkela_wire_179)
    );

    and_bi _2133_ (
        .b(jinkela_wire_179),
        .a(io_in2_0_),
        .c(jinkela_wire_397)
    );

    and_bi _2134_ (
        .b(jinkela_wire_397),
        .a(jinkela_wire_1511),
        .c(jinkela_wire_735)
    );

    or_bb _2135_ (
        .b(io_in2_1_),
        .a(jinkela_wire_735),
        .c(jinkela_wire_831)
    );

    or_bb _2136_ (
        .b(jinkela_wire_293),
        .a(jinkela_wire_188),
        .c(jinkela_wire_97)
    );

    and_bi _2137_ (
        .b(jinkela_wire_278),
        .a(jinkela_wire_188),
        .c(jinkela_wire_379)
    );

    and_bi _2138_ (
        .b(jinkela_wire_379),
        .a(jinkela_wire_97),
        .c(jinkela_wire_1171)
    );

    or_bb _2139_ (
        .b(io_in2_0_),
        .a(jinkela_wire_1171),
        .c(jinkela_wire_366)
    );

    or_bb _2140_ (
        .b(jinkela_wire_391),
        .a(jinkela_wire_188),
        .c(jinkela_wire_897)
    );

    and_bi _2141_ (
        .b(jinkela_wire_268),
        .a(jinkela_wire_188),
        .c(jinkela_wire_549)
    );

    and_bi _2142_ (
        .b(jinkela_wire_549),
        .a(jinkela_wire_897),
        .c(jinkela_wire_356)
    );

    and_bi _2143_ (
        .b(jinkela_wire_356),
        .a(io_in2_0_),
        .c(jinkela_wire_1291)
    );

    and_bi _2144_ (
        .b(jinkela_wire_1291),
        .a(jinkela_wire_366),
        .c(jinkela_wire_10)
    );

    and_bi _2145_ (
        .b(jinkela_wire_10),
        .a(io_in2_1_),
        .c(jinkela_wire_869)
    );

    and_bi _2146_ (
        .b(jinkela_wire_869),
        .a(jinkela_wire_831),
        .c(jinkela_wire_272)
    );

    and_bi _2147_ (
        .b(jinkela_wire_272),
        .a(io_in2_2_),
        .c(jinkela_wire_801)
    );

    or_bb _2148_ (
        .b(jinkela_wire_1324),
        .a(jinkela_wire_801),
        .c(jinkela_wire_1399)
    );

    or_ii _2149_ (
        .b(jinkela_wire_804),
        .a(jinkela_wire_1399),
        .c(jinkela_wire_1189)
    );

    or_bb _2150_ (
        .b(jinkela_wire_95),
        .a(jinkela_wire_188),
        .c(jinkela_wire_189)
    );

    and_bi _2151_ (
        .b(jinkela_wire_251),
        .a(jinkela_wire_188),
        .c(jinkela_wire_491)
    );

    and_bi _2152_ (
        .b(jinkela_wire_491),
        .a(jinkela_wire_189),
        .c(jinkela_wire_1134)
    );

    or_bb _2153_ (
        .b(io_in2_0_),
        .a(jinkela_wire_1134),
        .c(jinkela_wire_176)
    );

    or_bb _2154_ (
        .b(jinkela_wire_561),
        .a(jinkela_wire_188),
        .c(jinkela_wire_698)
    );

    and_bi _2155_ (
        .b(jinkela_wire_1241),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1305)
    );

    and_bi _2156_ (
        .b(jinkela_wire_1305),
        .a(jinkela_wire_698),
        .c(jinkela_wire_274)
    );

    or_bb _2664_ (
        .b(jinkela_wire_567),
        .a(jinkela_wire_141),
        .c(jinkela_wire_266)
    );

    and_bi _1947_ (
        .b(jinkela_wire_1410),
        .a(jinkela_wire_1479),
        .c(jinkela_wire_1085)
    );

    or_bb _2665_ (
        .b(jinkela_wire_191),
        .a(jinkela_wire_266),
        .c(jinkela_wire_1193)
    );

    or_bb _1948_ (
        .b(jinkela_wire_593),
        .a(jinkela_wire_1085),
        .c(io_adder_out_7_)
    );

    and_bi _2666_ (
        .b(jinkela_wire_567),
        .a(jinkela_wire_349),
        .c(jinkela_wire_198)
    );

    and_bi _1949_ (
        .b(jinkela_wire_1123),
        .a(jinkela_wire_442),
        .c(jinkela_wire_478)
    );

    and_bi _2667_ (
        .b(jinkela_wire_198),
        .a(jinkela_wire_141),
        .c(jinkela_wire_658)
    );

    or_bb _1950_ (
        .b(jinkela_wire_195),
        .a(jinkela_wire_478),
        .c(jinkela_wire_152)
    );

    and_bi _2668_ (
        .b(jinkela_wire_658),
        .a(jinkela_wire_1193),
        .c(jinkela_wire_287)
    );

    and_bb _1951_ (
        .b(jinkela_wire_195),
        .a(jinkela_wire_478),
        .c(jinkela_wire_1049)
    );

    and_bi _2669_ (
        .b(jinkela_wire_287),
        .a(jinkela_wire_44),
        .c(jinkela_wire_334)
    );

    and_bi _1952_ (
        .b(jinkela_wire_1049),
        .a(jinkela_wire_152),
        .c(io_adder_out_6_)
    );

    or_bb _2670_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_334),
        .c(jinkela_wire_1377)
    );

    and_bi _1953_ (
        .b(jinkela_wire_1408),
        .a(jinkela_wire_1327),
        .c(jinkela_wire_706)
    );

    or_bb _2671_ (
        .b(jinkela_wire_23),
        .a(jinkela_wire_1377),
        .c(jinkela_wire_1139)
    );

    and_bi _1954_ (
        .b(jinkela_wire_706),
        .a(jinkela_wire_793),
        .c(jinkela_wire_113)
    );

    and_bi _2672_ (
        .b(jinkela_wire_635),
        .a(jinkela_wire_804),
        .c(jinkela_wire_59)
    );

    and_bi _1955_ (
        .b(jinkela_wire_793),
        .a(jinkela_wire_706),
        .c(jinkela_wire_1000)
    );

    and_bi _2673_ (
        .b(jinkela_wire_1461),
        .a(io_in2_3_),
        .c(jinkela_wire_982)
    );

    or_bb _1956_ (
        .b(jinkela_wire_113),
        .a(jinkela_wire_1000),
        .c(io_adder_out_5_)
    );

    or_bb _2674_ (
        .b(io_in2_4_),
        .a(jinkela_wire_982),
        .c(jinkela_wire_381)
    );

    and_bi _1957_ (
        .b(jinkela_wire_1103),
        .a(jinkela_wire_26),
        .c(jinkela_wire_875)
    );

    or_bb _2675_ (
        .b(jinkela_wire_59),
        .a(jinkela_wire_381),
        .c(jinkela_wire_1385)
    );

    or_bb _1958_ (
        .b(jinkela_wire_70),
        .a(jinkela_wire_875),
        .c(jinkela_wire_9)
    );

    and_bi _2676_ (
        .b(jinkela_wire_1248),
        .a(jinkela_wire_883),
        .c(jinkela_wire_701)
    );

    and_bb _1959_ (
        .b(jinkela_wire_70),
        .a(jinkela_wire_875),
        .c(jinkela_wire_1172)
    );

    or_bi _2677_ (
        .b(jinkela_wire_1385),
        .a(jinkela_wire_701),
        .c(jinkela_wire_21)
    );

    and_bi _1960_ (
        .b(jinkela_wire_1172),
        .a(jinkela_wire_9),
        .c(io_adder_out_4_)
    );

    and_bb _2678_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_21),
        .c(jinkela_wire_1237)
    );

    and_bi _1961_ (
        .b(jinkela_wire_1061),
        .a(jinkela_wire_310),
        .c(jinkela_wire_1227)
    );

    or_bb _2679_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1237),
        .c(jinkela_wire_859)
    );

    and_bi _1962_ (
        .b(jinkela_wire_1227),
        .a(jinkela_wire_24),
        .c(jinkela_wire_303)
    );

    and_bi _2680_ (
        .b(jinkela_wire_859),
        .a(jinkela_wire_1139),
        .c(jinkela_wire_716)
    );

    and_bi _1963_ (
        .b(jinkela_wire_24),
        .a(jinkela_wire_1227),
        .c(jinkela_wire_284)
    );

    or_bb _2681_ (
        .b(jinkela_wire_850),
        .a(jinkela_wire_716),
        .c(io_out_9_)
    );

    or_bb _1964_ (
        .b(jinkela_wire_303),
        .a(jinkela_wire_284),
        .c(io_adder_out_3_)
    );

    and_bi _2682_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_10_),
        .c(jinkela_wire_718)
    );

    and_bi _1965_ (
        .b(jinkela_wire_127),
        .a(jinkela_wire_779),
        .c(jinkela_wire_832)
    );

    and_bi _2683_ (
        .b(jinkela_wire_1503),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_529)
    );

    and_bi _1966_ (
        .b(jinkela_wire_832),
        .a(jinkela_wire_755),
        .c(jinkela_wire_1112)
    );

    and_bi _2684_ (
        .b(jinkela_wire_529),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_770)
    );

    and_bi _1967_ (
        .b(jinkela_wire_755),
        .a(jinkela_wire_832),
        .c(jinkela_wire_336)
    );

    and_bi _2685_ (
        .b(jinkela_wire_770),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_35)
    );

    or_bb _1968_ (
        .b(jinkela_wire_1112),
        .a(jinkela_wire_336),
        .c(io_adder_out_2_)
    );

    and_bi _2686_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_217),
        .c(jinkela_wire_1046)
    );

    and_bi _1969_ (
        .b(jinkela_wire_115),
        .a(jinkela_wire_119),
        .c(jinkela_wire_149)
    );

    inv _2687_ (
        .din(io_in2_10_),
        .dout(jinkela_wire_950)
    );

    or_bb _1970_ (
        .b(jinkela_wire_1509),
        .a(jinkela_wire_149),
        .c(jinkela_wire_898)
    );

    and_bi _2688_ (
        .b(jinkela_wire_347),
        .a(io_in1_10_),
        .c(jinkela_wire_1176)
    );

    and_bb _1971_ (
        .b(jinkela_wire_1509),
        .a(jinkela_wire_149),
        .c(jinkela_wire_417)
    );

    or_bb _2689_ (
        .b(jinkela_wire_950),
        .a(jinkela_wire_1176),
        .c(jinkela_wire_1024)
    );

    and_bi _1972_ (
        .b(jinkela_wire_417),
        .a(jinkela_wire_898),
        .c(io_adder_out_1_)
    );

    or_bb _2690_ (
        .b(jinkela_wire_1046),
        .a(jinkela_wire_1024),
        .c(jinkela_wire_1434)
    );

    inv _1973_ (
        .din(jinkela_wire_394),
        .dout(jinkela_wire_1192)
    );

    and_bi _2691_ (
        .b(jinkela_wire_950),
        .a(jinkela_wire_349),
        .c(jinkela_wire_821)
    );

    inv _1974_ (
        .din(io_in1_0_),
        .dout(jinkela_wire_1300)
    );

    and_bi _2692_ (
        .b(jinkela_wire_821),
        .a(jinkela_wire_1176),
        .c(jinkela_wire_733)
    );

    and_bi _1975_ (
        .b(io_in2_0_),
        .a(jinkela_wire_1300),
        .c(jinkela_wire_276)
    );

    and_bi _2693_ (
        .b(jinkela_wire_733),
        .a(jinkela_wire_1434),
        .c(jinkela_wire_240)
    );

    and_bi _1976_ (
        .b(jinkela_wire_276),
        .a(jinkela_wire_1192),
        .c(io_adder_out_0_)
    );

    and_bi _2694_ (
        .b(jinkela_wire_240),
        .a(jinkela_wire_44),
        .c(jinkela_wire_1323)
    );

    or_bb _1977_ (
        .b(jinkela_wire_338),
        .a(jinkela_wire_1339),
        .c(jinkela_wire_828)
    );

    or_bb _2695_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1323),
        .c(jinkela_wire_940)
    );

    and_bi _1978_ (
        .b(jinkela_wire_785),
        .a(jinkela_wire_828),
        .c(io_test_adder_Cout)
    );

    or_bb _2696_ (
        .b(jinkela_wire_35),
        .a(jinkela_wire_940),
        .c(jinkela_wire_49)
    );

    or_bi _1979_ (
        .b(io_fn_3_),
        .a(io_fn_0_),
        .c(jinkela_wire_218)
    );

    and_bi _2697_ (
        .b(jinkela_wire_962),
        .a(jinkela_wire_804),
        .c(jinkela_wire_818)
    );

    or_bi _1980_ (
        .b(io_fn_1_),
        .a(io_fn_2_),
        .c(jinkela_wire_109)
    );

    and_bi _2698_ (
        .b(jinkela_wire_998),
        .a(io_in2_3_),
        .c(jinkela_wire_892)
    );

    or_bb _1981_ (
        .b(jinkela_wire_218),
        .a(jinkela_wire_109),
        .c(jinkela_wire_947)
    );

    or_bb _2699_ (
        .b(io_in2_4_),
        .a(jinkela_wire_892),
        .c(jinkela_wire_410)
    );

    or_bb _1982_ (
        .b(io_fn_3_),
        .a(io_fn_2_),
        .c(jinkela_wire_1226)
    );

    or_bb _2700_ (
        .b(jinkela_wire_818),
        .a(jinkela_wire_410),
        .c(jinkela_wire_521)
    );

    or_bb _1983_ (
        .b(io_fn_0_),
        .a(io_fn_1_),
        .c(jinkela_wire_1064)
    );

    and_bi _2701_ (
        .b(jinkela_wire_1248),
        .a(jinkela_wire_259),
        .c(jinkela_wire_472)
    );

    or_bb _1984_ (
        .b(jinkela_wire_1226),
        .a(jinkela_wire_1064),
        .c(jinkela_wire_483)
    );

    or_bi _2702_ (
        .b(jinkela_wire_521),
        .a(jinkela_wire_472),
        .c(jinkela_wire_628)
    );

    and_bb _1985_ (
        .b(jinkela_wire_947),
        .a(jinkela_wire_483),
        .c(jinkela_wire_1389)
    );

    and_bb _2703_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_628),
        .c(jinkela_wire_532)
    );

    or_bb _1986_ (
        .b(io_adder_out_0_),
        .a(jinkela_wire_1389),
        .c(jinkela_wire_1175)
    );

    or_bb _2704_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_532),
        .c(jinkela_wire_1135)
    );

    and_bi _1987_ (
        .b(jinkela_wire_218),
        .a(io_fn_2_),
        .c(jinkela_wire_1187)
    );

    and_bi _2705_ (
        .b(jinkela_wire_1135),
        .a(jinkela_wire_49),
        .c(jinkela_wire_936)
    );

    and_bi _1988_ (
        .b(io_in2_31_),
        .a(io_in1_31_),
        .c(jinkela_wire_159)
    );

    and_bi _1779_ (
        .b(io_in2_22_),
        .a(jinkela_wire_926),
        .c(jinkela_wire_1480)
    );

    or_bb _2493_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1504),
        .c(jinkela_wire_1239)
    );

    and_bi _1780_ (
        .b(jinkela_wire_926),
        .a(io_in2_22_),
        .c(jinkela_wire_372)
    );

    or_bb _2494_ (
        .b(jinkela_wire_382),
        .a(jinkela_wire_1239),
        .c(jinkela_wire_1222)
    );

    or_bb _1781_ (
        .b(jinkela_wire_1480),
        .a(jinkela_wire_372),
        .c(jinkela_wire_420)
    );

    or_bb _2495_ (
        .b(jinkela_wire_804),
        .a(jinkela_wire_1036),
        .c(jinkela_wire_938)
    );

    and_bb _1782_ (
        .b(jinkela_wire_834),
        .a(jinkela_wire_420),
        .c(jinkela_wire_385)
    );

    and_bi _2496_ (
        .b(jinkela_wire_272),
        .a(jinkela_wire_158),
        .c(jinkela_wire_876)
    );

    or_bb _1783_ (
        .b(jinkela_wire_1096),
        .a(jinkela_wire_385),
        .c(jinkela_wire_1124)
    );

    and_bi _2497_ (
        .b(jinkela_wire_1136),
        .a(io_in2_2_),
        .c(jinkela_wire_175)
    );

    and_bi _1784_ (
        .b(jinkela_wire_1124),
        .a(jinkela_wire_268),
        .c(jinkela_wire_1245)
    );

    or_bb _2498_ (
        .b(jinkela_wire_876),
        .a(jinkela_wire_175),
        .c(jinkela_wire_376)
    );

    or_ii _1785_ (
        .b(io_in1_23_),
        .a(jinkela_wire_1124),
        .c(jinkela_wire_165)
    );

    and_bi _2499_ (
        .b(jinkela_wire_376),
        .a(jinkela_wire_804),
        .c(jinkela_wire_504)
    );

    inv _1786_ (
        .din(io_in2_23_),
        .dout(jinkela_wire_535)
    );

    and_bi _2500_ (
        .b(jinkela_wire_504),
        .a(jinkela_wire_938),
        .c(jinkela_wire_731)
    );

    and_bi _1787_ (
        .b(jinkela_wire_839),
        .a(io_fn_3_),
        .c(jinkela_wire_767)
    );

    and_bi _2501_ (
        .b(jinkela_wire_731),
        .a(io_in2_4_),
        .c(jinkela_wire_114)
    );

    and_bi _1788_ (
        .b(jinkela_wire_535),
        .a(jinkela_wire_767),
        .c(jinkela_wire_945)
    );

    or_ii _2502_ (
        .b(jinkela_wire_158),
        .a(jinkela_wire_648),
        .c(jinkela_wire_768)
    );

    and_bi _1789_ (
        .b(jinkela_wire_767),
        .a(jinkela_wire_535),
        .c(jinkela_wire_1078)
    );

    and_bi _2503_ (
        .b(jinkela_wire_976),
        .a(io_in2_2_),
        .c(jinkela_wire_402)
    );

    or_bb _1790_ (
        .b(jinkela_wire_945),
        .a(jinkela_wire_1078),
        .c(jinkela_wire_1380)
    );

    and_bi _2504_ (
        .b(jinkela_wire_402),
        .a(jinkela_wire_768),
        .c(jinkela_wire_396)
    );

    inv _1791_ (
        .din(jinkela_wire_1380),
        .dout(jinkela_wire_180)
    );

    and_bi _2505_ (
        .b(jinkela_wire_396),
        .a(jinkela_wire_804),
        .c(jinkela_wire_172)
    );

    and_bi _1792_ (
        .b(jinkela_wire_180),
        .a(jinkela_wire_165),
        .c(jinkela_wire_315)
    );

    and_bi _2506_ (
        .b(jinkela_wire_1275),
        .a(jinkela_wire_158),
        .c(jinkela_wire_917)
    );

    or_bb _1793_ (
        .b(jinkela_wire_1245),
        .a(jinkela_wire_315),
        .c(jinkela_wire_1361)
    );

    and_bi _2507_ (
        .b(jinkela_wire_1219),
        .a(io_in2_2_),
        .c(jinkela_wire_210)
    );

    and_bi _1794_ (
        .b(jinkela_wire_1361),
        .a(io_in1_24_),
        .c(jinkela_wire_856)
    );

    or_bb _2508_ (
        .b(jinkela_wire_917),
        .a(jinkela_wire_210),
        .c(jinkela_wire_757)
    );

    inv _1795_ (
        .din(io_in1_24_),
        .dout(jinkela_wire_251)
    );

    and_bi _2509_ (
        .b(jinkela_wire_804),
        .a(jinkela_wire_757),
        .c(jinkela_wire_1018)
    );

    or_ii _1796_ (
        .b(jinkela_wire_251),
        .a(jinkela_wire_1361),
        .c(jinkela_wire_299)
    );

    or_bb _2510_ (
        .b(jinkela_wire_172),
        .a(jinkela_wire_1018),
        .c(jinkela_wire_1412)
    );

    and_bi _1797_ (
        .b(jinkela_wire_1128),
        .a(io_fn_3_),
        .c(jinkela_wire_429)
    );

    and_bi _2511_ (
        .b(jinkela_wire_1412),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_306)
    );

    and_bi _1798_ (
        .b(io_in2_24_),
        .a(jinkela_wire_429),
        .c(jinkela_wire_1156)
    );

    or_bb _2512_ (
        .b(jinkela_wire_114),
        .a(jinkela_wire_306),
        .c(jinkela_wire_1232)
    );

    and_bi _1799_ (
        .b(jinkela_wire_429),
        .a(io_in2_24_),
        .c(jinkela_wire_1487)
    );

    and_bb _2513_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1232),
        .c(jinkela_wire_1149)
    );

    or_bb _1800_ (
        .b(jinkela_wire_1156),
        .a(jinkela_wire_1487),
        .c(jinkela_wire_1319)
    );

    or_bb _2514_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1149),
        .c(jinkela_wire_181)
    );

    and_bb _1801_ (
        .b(jinkela_wire_299),
        .a(jinkela_wire_1319),
        .c(jinkela_wire_1051)
    );

    and_bi _2515_ (
        .b(jinkela_wire_181),
        .a(jinkela_wire_1222),
        .c(jinkela_wire_161)
    );

    or_bb _1802_ (
        .b(jinkela_wire_856),
        .a(jinkela_wire_1051),
        .c(jinkela_wire_445)
    );

    or_bb _2516_ (
        .b(jinkela_wire_1349),
        .a(jinkela_wire_161),
        .c(io_out_4_)
    );

    and_bi _1803_ (
        .b(jinkela_wire_1241),
        .a(jinkela_wire_445),
        .c(jinkela_wire_1468)
    );

    and_bi _2517_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_5_),
        .c(jinkela_wire_32)
    );

    inv _1804_ (
        .din(jinkela_wire_1468),
        .dout(jinkela_wire_712)
    );

    and_bi _2518_ (
        .b(jinkela_wire_650),
        .a(jinkela_wire_804),
        .c(jinkela_wire_1233)
    );

    or_bb _1805_ (
        .b(io_in1_25_),
        .a(jinkela_wire_445),
        .c(jinkela_wire_342)
    );

    and_bi _2519_ (
        .b(jinkela_wire_1233),
        .a(jinkela_wire_1269),
        .c(jinkela_wire_259)
    );

    and_bi _1806_ (
        .b(jinkela_wire_923),
        .a(io_fn_3_),
        .c(jinkela_wire_235)
    );

    and_bi _2520_ (
        .b(jinkela_wire_259),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_1337)
    );

    and_bi _1807_ (
        .b(jinkela_wire_235),
        .a(io_in2_25_),
        .c(jinkela_wire_474)
    );

    and_bi _2521_ (
        .b(jinkela_wire_1337),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_295)
    );

    and_bi _1808_ (
        .b(io_in2_25_),
        .a(jinkela_wire_235),
        .c(jinkela_wire_1022)
    );

    and_bi _2522_ (
        .b(jinkela_wire_295),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_1460)
    );

    or_bb _1809_ (
        .b(jinkela_wire_474),
        .a(jinkela_wire_1022),
        .c(jinkela_wire_228)
    );

    and_bi _2523_ (
        .b(jinkela_wire_347),
        .a(io_in1_5_),
        .c(jinkela_wire_112)
    );

    and_bb _1810_ (
        .b(jinkela_wire_342),
        .a(jinkela_wire_228),
        .c(jinkela_wire_688)
    );

    and_bi _2524_ (
        .b(jinkela_wire_921),
        .a(jinkela_wire_349),
        .c(jinkela_wire_1271)
    );

    and_bi _1811_ (
        .b(jinkela_wire_688),
        .a(jinkela_wire_712),
        .c(jinkela_wire_713)
    );

    and_bi _2525_ (
        .b(jinkela_wire_1271),
        .a(jinkela_wire_112),
        .c(jinkela_wire_1100)
    );

    or_bb _1812_ (
        .b(jinkela_wire_562),
        .a(jinkela_wire_713),
        .c(jinkela_wire_814)
    );

    and_bi _2526_ (
        .b(jinkela_wire_112),
        .a(io_in2_5_),
        .c(jinkela_wire_611)
    );

    or_ii _1813_ (
        .b(jinkela_wire_562),
        .a(jinkela_wire_713),
        .c(jinkela_wire_516)
    );

    or_bb _2527_ (
        .b(jinkela_wire_1100),
        .a(jinkela_wire_611),
        .c(jinkela_wire_63)
    );

    or_bb _1814_ (
        .b(jinkela_wire_1424),
        .a(jinkela_wire_1058),
        .c(jinkela_wire_604)
    );

    and_bi _2528_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_1137),
        .c(jinkela_wire_1178)
    );

    and_bi _1815_ (
        .b(jinkela_wire_604),
        .a(io_in2_26_),
        .c(jinkela_wire_754)
    );

    or_bb _2529_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_1178),
        .c(jinkela_wire_319)
    );

    and_bi _1816_ (
        .b(io_in2_26_),
        .a(jinkela_wire_604),
        .c(jinkela_wire_758)
    );

    and_bi _2530_ (
        .b(jinkela_wire_319),
        .a(jinkela_wire_63),
        .c(jinkela_wire_509)
    );

    or_bb _1817_ (
        .b(jinkela_wire_754),
        .a(jinkela_wire_758),
        .c(jinkela_wire_8)
    );

    or_bb _2531_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_509),
        .c(jinkela_wire_433)
    );

    and_bi _1818_ (
        .b(jinkela_wire_8),
        .a(jinkela_wire_516),
        .c(jinkela_wire_1277)
    );

    or_bb _2532_ (
        .b(jinkela_wire_1460),
        .a(jinkela_wire_433),
        .c(jinkela_wire_981)
    );

    and_bi _1819_ (
        .b(jinkela_wire_1277),
        .a(jinkela_wire_814),
        .c(jinkela_wire_591)
    );

    or_bb _2533_ (
        .b(io_in2_2_),
        .a(jinkela_wire_1294),
        .c(jinkela_wire_102)
    );

    or_ii _1820_ (
        .b(jinkela_wire_1234),
        .a(jinkela_wire_591),
        .c(jinkela_wire_61)
    );

    and_bi _2534_ (
        .b(jinkela_wire_137),
        .a(io_in2_2_),
        .c(jinkela_wire_624)
    );

    and_bi _3042_ (
        .b(jinkela_wire_523),
        .a(jinkela_wire_347),
        .c(jinkela_wire_1295)
    );

    and_bi _1608_ (
        .b(jinkela_wire_565),
        .a(io_in2_4_),
        .c(jinkela_wire_1266)
    );

    and_bi _2325_ (
        .b(jinkela_wire_1387),
        .a(io_in2_1_),
        .c(jinkela_wire_703)
    );

    or_bb _3043_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_1295),
        .c(jinkela_wire_1217)
    );

    or_bb _1609_ (
        .b(jinkela_wire_525),
        .a(jinkela_wire_1266),
        .c(jinkela_wire_70)
    );

    and_bi _2326_ (
        .b(jinkela_wire_703),
        .a(jinkela_wire_1443),
        .c(jinkela_wire_1066)
    );

    and_bi _3044_ (
        .b(jinkela_wire_1217),
        .a(jinkela_wire_485),
        .c(jinkela_wire_219)
    );

    and_bi _1610_ (
        .b(jinkela_wire_70),
        .a(jinkela_wire_26),
        .c(jinkela_wire_1365)
    );

    or_bb _2327_ (
        .b(io_in2_2_),
        .a(jinkela_wire_1066),
        .c(jinkela_wire_1350)
    );

    or_bb _3045_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_219),
        .c(jinkela_wire_972)
    );

    or_bb _1611_ (
        .b(jinkela_wire_1103),
        .a(jinkela_wire_1365),
        .c(jinkela_wire_1007)
    );

    and_bi _2328_ (
        .b(io_in2_0_),
        .a(jinkela_wire_618),
        .c(jinkela_wire_581)
    );

    or_bb _3046_ (
        .b(jinkela_wire_605),
        .a(jinkela_wire_972),
        .c(jinkela_wire_769)
    );

    and_bi _1612_ (
        .b(io_in1_5_),
        .a(jinkela_wire_1007),
        .c(jinkela_wire_1408)
    );

    and_bi _2329_ (
        .b(jinkela_wire_581),
        .a(jinkela_wire_1407),
        .c(jinkela_wire_505)
    );

    and_bb _3047_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1381),
        .c(jinkela_wire_1272)
    );

    inv _1613_ (
        .din(io_in1_5_),
        .dout(jinkela_wire_1137)
    );

    and_bi _2330_ (
        .b(jinkela_wire_1466),
        .a(jinkela_wire_915),
        .c(jinkela_wire_47)
    );

    or_bb _3048_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1272),
        .c(jinkela_wire_1133)
    );

    or_bb _1614_ (
        .b(jinkela_wire_1137),
        .a(jinkela_wire_1007),
        .c(jinkela_wire_1327)
    );

    and_bi _2331_ (
        .b(jinkela_wire_1497),
        .a(io_in2_0_),
        .c(jinkela_wire_1021)
    );

    and_bi _3049_ (
        .b(jinkela_wire_1133),
        .a(jinkela_wire_769),
        .c(jinkela_wire_1465)
    );

    inv _1615_ (
        .din(io_in2_5_),
        .dout(jinkela_wire_921)
    );

    or_bb _2332_ (
        .b(jinkela_wire_47),
        .a(jinkela_wire_1021),
        .c(jinkela_wire_929)
    );

    or_bb _3050_ (
        .b(jinkela_wire_1118),
        .a(jinkela_wire_1465),
        .c(io_out_28_)
    );

    and_bi _1616_ (
        .b(jinkela_wire_1405),
        .a(io_fn_3_),
        .c(jinkela_wire_564)
    );

    and_bi _2333_ (
        .b(jinkela_wire_929),
        .a(jinkela_wire_15),
        .c(jinkela_wire_1458)
    );

    and_bi _3051_ (
        .b(jinkela_wire_68),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_637)
    );

    or_bb _2334_ (
        .b(jinkela_wire_505),
        .a(jinkela_wire_1458),
        .c(jinkela_wire_782)
    );

    and_bi _1617_ (
        .b(jinkela_wire_921),
        .a(jinkela_wire_564),
        .c(jinkela_wire_215)
    );

    and_bi _3052_ (
        .b(jinkela_wire_262),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_250)
    );

    and_bi _2335_ (
        .b(jinkela_wire_782),
        .a(io_in2_2_),
        .c(jinkela_wire_1307)
    );

    and_bi _1618_ (
        .b(jinkela_wire_564),
        .a(jinkela_wire_921),
        .c(jinkela_wire_238)
    );

    or_bb _3053_ (
        .b(io_in1_29_),
        .a(jinkela_wire_250),
        .c(jinkela_wire_1485)
    );

    and_bi _2336_ (
        .b(jinkela_wire_1307),
        .a(jinkela_wire_1350),
        .c(jinkela_wire_740)
    );

    or_bb _1619_ (
        .b(jinkela_wire_215),
        .a(jinkela_wire_238),
        .c(jinkela_wire_1342)
    );

    and_bb _3054_ (
        .b(io_in1_29_),
        .a(io_in2_29_),
        .c(jinkela_wire_664)
    );

    and_bi _2337_ (
        .b(jinkela_wire_740),
        .a(io_in2_3_),
        .c(jinkela_wire_1398)
    );

    inv _1620_ (
        .din(jinkela_wire_1342),
        .dout(jinkela_wire_793)
    );

    and_bb _3055_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_664),
        .c(jinkela_wire_1409)
    );

    and_bi _2338_ (
        .b(jinkela_wire_1398),
        .a(jinkela_wire_123),
        .c(jinkela_wire_456)
    );

    and_bi _1621_ (
        .b(jinkela_wire_793),
        .a(jinkela_wire_1327),
        .c(jinkela_wire_490)
    );

    and_bi _3056_ (
        .b(jinkela_wire_1409),
        .a(jinkela_wire_1485),
        .c(jinkela_wire_858)
    );

    and_bi _2339_ (
        .b(jinkela_wire_456),
        .a(io_in2_4_),
        .c(jinkela_wire_87)
    );

    or_bb _1622_ (
        .b(jinkela_wire_1408),
        .a(jinkela_wire_490),
        .c(jinkela_wire_1053)
    );

    or_bb _3057_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_858),
        .c(jinkela_wire_920)
    );

    or_bb _2340_ (
        .b(jinkela_wire_762),
        .a(jinkela_wire_87),
        .c(jinkela_wire_583)
    );

    and_bi _1623_ (
        .b(jinkela_wire_1053),
        .a(io_in1_6_),
        .c(jinkela_wire_1123)
    );

    and_bi _3058_ (
        .b(jinkela_wire_664),
        .a(jinkela_wire_347),
        .c(jinkela_wire_502)
    );

    and_bi _2341_ (
        .b(jinkela_wire_583),
        .a(jinkela_wire_188),
        .c(jinkela_wire_458)
    );

    inv _1624_ (
        .din(io_in1_6_),
        .dout(jinkela_wire_561)
    );

    or_bb _3059_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_502),
        .c(jinkela_wire_1311)
    );

    or_bi _2342_ (
        .b(jinkela_wire_1389),
        .a(jinkela_wire_1187),
        .c(jinkela_wire_625)
    );

    or_ii _1625_ (
        .b(jinkela_wire_561),
        .a(jinkela_wire_1053),
        .c(jinkela_wire_442)
    );

    and_bi _3060_ (
        .b(jinkela_wire_1311),
        .a(jinkela_wire_920),
        .c(jinkela_wire_1198)
    );

    or_bb _2343_ (
        .b(jinkela_wire_458),
        .a(jinkela_wire_625),
        .c(jinkela_wire_932)
    );

    and_bi _1626_ (
        .b(jinkela_wire_1168),
        .a(io_fn_3_),
        .c(jinkela_wire_75)
    );

    or_bb _3061_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1198),
        .c(jinkela_wire_65)
    );

    and_bi _2344_ (
        .b(jinkela_wire_932),
        .a(jinkela_wire_986),
        .c(jinkela_wire_1252)
    );

    and_bi _1627_ (
        .b(io_in2_6_),
        .a(jinkela_wire_75),
        .c(jinkela_wire_965)
    );

    or_bb _3062_ (
        .b(jinkela_wire_637),
        .a(jinkela_wire_65),
        .c(jinkela_wire_367)
    );

    or_bb _2345_ (
        .b(jinkela_wire_432),
        .a(jinkela_wire_1252),
        .c(io_out_1_)
    );

    and_bi _1628_ (
        .b(jinkela_wire_75),
        .a(io_in2_6_),
        .c(jinkela_wire_727)
    );

    and_bb _3063_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_868),
        .c(jinkela_wire_1170)
    );

    and_bi _2346_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_2_),
        .c(jinkela_wire_574)
    );

    or_bb _1629_ (
        .b(jinkela_wire_965),
        .a(jinkela_wire_727),
        .c(jinkela_wire_195)
    );

    or_bb _3064_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1170),
        .c(jinkela_wire_1285)
    );

    and_bi _2347_ (
        .b(jinkela_wire_782),
        .a(jinkela_wire_158),
        .c(jinkela_wire_1320)
    );

    and_bb _1630_ (
        .b(jinkela_wire_442),
        .a(jinkela_wire_195),
        .c(jinkela_wire_1429)
    );

    and_bi _3065_ (
        .b(jinkela_wire_1285),
        .a(jinkela_wire_367),
        .c(jinkela_wire_1098)
    );

    and_bi _2348_ (
        .b(jinkela_wire_1320),
        .a(jinkela_wire_970),
        .c(jinkela_wire_830)
    );

    or_bb _1631_ (
        .b(jinkela_wire_1123),
        .a(jinkela_wire_1429),
        .c(jinkela_wire_791)
    );

    and_bi _3066_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_29_),
        .c(jinkela_wire_622)
    );

    and_bi _2349_ (
        .b(jinkela_wire_830),
        .a(jinkela_wire_804),
        .c(jinkela_wire_380)
    );

    and_bi _1632_ (
        .b(jinkela_wire_791),
        .a(jinkela_wire_95),
        .c(jinkela_wire_1462)
    );

    or_bb _3067_ (
        .b(jinkela_wire_1098),
        .a(jinkela_wire_622),
        .c(io_out_29_)
    );

    and_bi _2350_ (
        .b(jinkela_wire_380),
        .a(jinkela_wire_1269),
        .c(jinkela_wire_1392)
    );

    or_ii _1633_ (
        .b(io_in1_7_),
        .a(jinkela_wire_791),
        .c(jinkela_wire_148)
    );

    and_bi _3068_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_30_),
        .c(jinkela_wire_794)
    );

    and_bi _2351_ (
        .b(jinkela_wire_1392),
        .a(jinkela_wire_1248),
        .c(jinkela_wire_812)
    );

    inv _1634_ (
        .din(io_in2_7_),
        .dout(jinkela_wire_1490)
    );

    and_bi _3069_ (
        .b(jinkela_wire_44),
        .a(jinkela_wire_583),
        .c(jinkela_wire_90)
    );

    and_bi _2352_ (
        .b(jinkela_wire_812),
        .a(jinkela_wire_1268),
        .c(jinkela_wire_868)
    );

    and_bi _1635_ (
        .b(jinkela_wire_1079),
        .a(io_fn_3_),
        .c(jinkela_wire_1428)
    );

    and_bi _3070_ (
        .b(jinkela_wire_1345),
        .a(jinkela_wire_964),
        .c(jinkela_wire_1273)
    );

    and_bi _2353_ (
        .b(jinkela_wire_868),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_94)
    );

    and_bi _1636_ (
        .b(jinkela_wire_1490),
        .a(jinkela_wire_1428),
        .c(jinkela_wire_468)
    );

    inv _3071_ (
        .din(io_in2_30_),
        .dout(jinkela_wire_919)
    );

    and_bi _2354_ (
        .b(jinkela_wire_158),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_1146)
    );

    and_bi _1637_ (
        .b(jinkela_wire_1428),
        .a(jinkela_wire_1490),
        .c(jinkela_wire_405)
    );

    and_bi _3072_ (
        .b(jinkela_wire_347),
        .a(io_in1_30_),
        .c(jinkela_wire_756)
    );

    or_bb _2355_ (
        .b(io_in1_2_),
        .a(jinkela_wire_1146),
        .c(jinkela_wire_1505)
    );

    or_bb _1638_ (
        .b(jinkela_wire_468),
        .a(jinkela_wire_405),
        .c(jinkela_wire_780)
    );

    or_bb _3073_ (
        .b(jinkela_wire_919),
        .a(jinkela_wire_756),
        .c(jinkela_wire_406)
    );

    and_bb _2356_ (
        .b(io_in1_2_),
        .a(io_in2_2_),
        .c(jinkela_wire_233)
    );

    inv _1639_ (
        .din(jinkela_wire_780),
        .dout(jinkela_wire_1479)
    );

    or_bb _3074_ (
        .b(jinkela_wire_1273),
        .a(jinkela_wire_406),
        .c(jinkela_wire_978)
    );

    and_bb _2357_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_233),
        .c(jinkela_wire_959)
    );

    and_bi _1640_ (
        .b(jinkela_wire_1479),
        .a(jinkela_wire_148),
        .c(jinkela_wire_520)
    );

    and_bi _3075_ (
        .b(jinkela_wire_919),
        .a(jinkela_wire_349),
        .c(jinkela_wire_400)
    );

    and_bi _2358_ (
        .b(jinkela_wire_959),
        .a(jinkela_wire_1505),
        .c(jinkela_wire_848)
    );

    or_bb _1641_ (
        .b(jinkela_wire_1462),
        .a(jinkela_wire_520),
        .c(jinkela_wire_708)
    );

    and_bi _3076_ (
        .b(jinkela_wire_400),
        .a(jinkela_wire_756),
        .c(jinkela_wire_829)
    );

    or_bb _2359_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_848),
        .c(jinkela_wire_679)
    );

    and_bi _1642_ (
        .b(io_in1_8_),
        .a(jinkela_wire_708),
        .c(jinkela_wire_609)
    );

    and_bi _3077_ (
        .b(jinkela_wire_829),
        .a(jinkela_wire_978),
        .c(jinkela_wire_977)
    );

    and_bi _2360_ (
        .b(jinkela_wire_233),
        .a(jinkela_wire_347),
        .c(jinkela_wire_1495)
    );

    inv _1643_ (
        .din(io_in1_8_),
        .dout(jinkela_wire_391)
    );

    and_bi _3078_ (
        .b(jinkela_wire_977),
        .a(jinkela_wire_44),
        .c(jinkela_wire_1474)
    );

    or_bb _2361_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_1495),
        .c(jinkela_wire_307)
    );

    or_bb _1644_ (
        .b(jinkela_wire_391),
        .a(jinkela_wire_708),
        .c(jinkela_wire_807)
    );

    or_bb _3079_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1474),
        .c(jinkela_wire_773)
    );

    and_bi _2362_ (
        .b(jinkela_wire_307),
        .a(jinkela_wire_679),
        .c(jinkela_wire_370)
    );

    and_bi _1645_ (
        .b(jinkela_wire_100),
        .a(io_fn_3_),
        .c(jinkela_wire_207)
    );

    or_bb _3080_ (
        .b(jinkela_wire_90),
        .a(jinkela_wire_773),
        .c(jinkela_wire_904)
    );

    or_bb _2363_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_370),
        .c(jinkela_wire_1459)
    );

    and_bi _1646_ (
        .b(io_in2_8_),
        .a(jinkela_wire_207),
        .c(jinkela_wire_1422)
    );

    and_bb _3081_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1499),
        .c(jinkela_wire_1247)
    );

    or_bb _2364_ (
        .b(jinkela_wire_94),
        .a(jinkela_wire_1459),
        .c(jinkela_wire_544)
    );

    and_bi _1647_ (
        .b(jinkela_wire_207),
        .a(io_in2_8_),
        .c(jinkela_wire_880)
    );

    or_bb _3082_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1247),
        .c(jinkela_wire_1363)
    );

    or_bb _2365_ (
        .b(io_in2_1_),
        .a(jinkela_wire_551),
        .c(jinkela_wire_335)
    );

    or_bb _1648_ (
        .b(jinkela_wire_1422),
        .a(jinkela_wire_880),
        .c(jinkela_wire_1463)
    );

    and_bi _3083_ (
        .b(jinkela_wire_1363),
        .a(jinkela_wire_904),
        .c(jinkela_wire_1289)
    );

    and_bi _1649_ (
        .b(jinkela_wire_1463),
        .a(jinkela_wire_807),
        .c(jinkela_wire_199)
    );

    and_bi _2366_ (
        .b(jinkela_wire_775),
        .a(io_in2_1_),
        .c(jinkela_wire_1045)
    );

    and_bi _2874_ (
        .b(jinkela_wire_783),
        .a(jinkela_wire_1213),
        .c(jinkela_wire_603)
    );

    and_bi _2157_ (
        .b(jinkela_wire_274),
        .a(io_in2_0_),
        .c(jinkela_wire_354)
    );

    or_bb _2875_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_603),
        .c(jinkela_wire_314)
    );

    and_bi _2158_ (
        .b(jinkela_wire_354),
        .a(jinkela_wire_176),
        .c(jinkela_wire_1052)
    );

    or_bb _2876_ (
        .b(jinkela_wire_722),
        .a(jinkela_wire_314),
        .c(jinkela_wire_254)
    );

    or_bb _2159_ (
        .b(io_in2_1_),
        .a(jinkela_wire_1052),
        .c(jinkela_wire_359)
    );

    and_bb _2877_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_543),
        .c(jinkela_wire_67)
    );

    or_bb _2160_ (
        .b(jinkela_wire_1137),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1333)
    );

    or_bb _2878_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_67),
        .c(jinkela_wire_939)
    );

    and_bi _2161_ (
        .b(jinkela_wire_562),
        .a(jinkela_wire_188),
        .c(jinkela_wire_619)
    );

    and_bi _2879_ (
        .b(jinkela_wire_939),
        .a(jinkela_wire_254),
        .c(jinkela_wire_355)
    );

    and_bi _2162_ (
        .b(jinkela_wire_619),
        .a(jinkela_wire_1333),
        .c(jinkela_wire_1336)
    );

    or_bb _2880_ (
        .b(jinkela_wire_674),
        .a(jinkela_wire_355),
        .c(io_out_18_)
    );

    or_bb _2163_ (
        .b(io_in2_0_),
        .a(jinkela_wire_1336),
        .c(jinkela_wire_40)
    );

    and_bi _2881_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_19_),
        .c(jinkela_wire_1180)
    );

    or_bb _2164_ (
        .b(jinkela_wire_1174),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1328)
    );

    and_bi _2882_ (
        .b(jinkela_wire_44),
        .a(jinkela_wire_1296),
        .c(jinkela_wire_399)
    );

    and_bi _2165_ (
        .b(jinkela_wire_1234),
        .a(jinkela_wire_188),
        .c(jinkela_wire_223)
    );

    and_bi _2883_ (
        .b(jinkela_wire_616),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_492)
    );

    and_bi _2166_ (
        .b(jinkela_wire_223),
        .a(jinkela_wire_1328),
        .c(jinkela_wire_1325)
    );

    or_bb _2884_ (
        .b(io_in1_19_),
        .a(jinkela_wire_492),
        .c(jinkela_wire_1142)
    );

    and_bi _2167_ (
        .b(jinkela_wire_1325),
        .a(io_in2_0_),
        .c(jinkela_wire_43)
    );

    and_bb _2885_ (
        .b(io_in1_19_),
        .a(io_in2_19_),
        .c(jinkela_wire_322)
    );

    and_bi _2168_ (
        .b(jinkela_wire_43),
        .a(jinkela_wire_40),
        .c(jinkela_wire_572)
    );

    and_bb _2886_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_322),
        .c(jinkela_wire_1)
    );

    and_bi _2169_ (
        .b(jinkela_wire_572),
        .a(io_in2_1_),
        .c(jinkela_wire_5)
    );

    and_bi _2887_ (
        .b(jinkela_wire_1),
        .a(jinkela_wire_1142),
        .c(jinkela_wire_744)
    );

    and_bi _2170_ (
        .b(jinkela_wire_5),
        .a(jinkela_wire_359),
        .c(jinkela_wire_1136)
    );

    or_bb _2888_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_744),
        .c(jinkela_wire_867)
    );

    or_bb _2171_ (
        .b(io_in2_2_),
        .a(jinkela_wire_1136),
        .c(jinkela_wire_1138)
    );

    and_bi _2889_ (
        .b(jinkela_wire_322),
        .a(jinkela_wire_347),
        .c(jinkela_wire_690)
    );

    or_bb _2172_ (
        .b(jinkela_wire_111),
        .a(jinkela_wire_188),
        .c(jinkela_wire_494)
    );

    or_bb _2890_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_690),
        .c(jinkela_wire_1056)
    );

    and_bi _2173_ (
        .b(jinkela_wire_1091),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1303)
    );

    and_bi _2891_ (
        .b(jinkela_wire_1056),
        .a(jinkela_wire_867),
        .c(jinkela_wire_1094)
    );

    and_bi _2174_ (
        .b(jinkela_wire_1303),
        .a(jinkela_wire_494),
        .c(jinkela_wire_1144)
    );

    or_bb _2892_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_1094),
        .c(jinkela_wire_1316)
    );

    or_bb _2175_ (
        .b(io_in2_0_),
        .a(jinkela_wire_1144),
        .c(jinkela_wire_638)
    );

    or_bb _2893_ (
        .b(jinkela_wire_399),
        .a(jinkela_wire_1316),
        .c(jinkela_wire_759)
    );

    or_bb _2176_ (
        .b(jinkela_wire_958),
        .a(jinkela_wire_188),
        .c(jinkela_wire_46)
    );

    and_bb _2894_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_340),
        .c(jinkela_wire_1469)
    );

    and_bi _2177_ (
        .b(jinkela_wire_1493),
        .a(jinkela_wire_188),
        .c(jinkela_wire_749)
    );

    or_bb _2895_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1469),
        .c(jinkela_wire_949)
    );

    and_bi _2178_ (
        .b(jinkela_wire_749),
        .a(jinkela_wire_46),
        .c(jinkela_wire_1466)
    );

    and_bi _2896_ (
        .b(jinkela_wire_949),
        .a(jinkela_wire_759),
        .c(jinkela_wire_872)
    );

    and_bi _2179_ (
        .b(jinkela_wire_1466),
        .a(io_in2_0_),
        .c(jinkela_wire_1209)
    );

    or_bb _2897_ (
        .b(jinkela_wire_1180),
        .a(jinkela_wire_872),
        .c(io_out_19_)
    );

    and_bi _2180_ (
        .b(jinkela_wire_1209),
        .a(jinkela_wire_638),
        .c(jinkela_wire_922)
    );

    and_bi _2898_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_20_),
        .c(jinkela_wire_162)
    );

    or_bb _2181_ (
        .b(io_in2_1_),
        .a(jinkela_wire_922),
        .c(jinkela_wire_1001)
    );

    and_bi _2899_ (
        .b(jinkela_wire_64),
        .a(jinkela_wire_1131),
        .c(jinkela_wire_185)
    );

    or_bb _2182_ (
        .b(jinkela_wire_746),
        .a(jinkela_wire_188),
        .c(jinkela_wire_1472)
    );

    and_bb _2900_ (
        .b(io_in2_20_),
        .a(jinkela_wire_1345),
        .c(jinkela_wire_1379)
    );

    and_bi _2183_ (
        .b(jinkela_wire_964),
        .a(jinkela_wire_188),
        .c(jinkela_wire_764)
    );

    or_bb _2901_ (
        .b(io_in1_20_),
        .a(jinkela_wire_1379),
        .c(jinkela_wire_582)
    );

    and_bi _2184_ (
        .b(jinkela_wire_764),
        .a(jinkela_wire_1472),
        .c(jinkela_wire_1497)
    );

    and_bb _2902_ (
        .b(io_in1_20_),
        .a(io_in2_20_),
        .c(jinkela_wire_878)
    );

    and_bi _2185_ (
        .b(jinkela_wire_1497),
        .a(jinkela_wire_915),
        .c(jinkela_wire_96)
    );

    and_bb _2903_ (
        .b(jinkela_wire_349),
        .a(jinkela_wire_878),
        .c(jinkela_wire_1279)
    );

    and_bi _2186_ (
        .b(jinkela_wire_188),
        .a(io_in1_0_),
        .c(jinkela_wire_705)
    );

    and_bi _2904_ (
        .b(jinkela_wire_1279),
        .a(jinkela_wire_582),
        .c(jinkela_wire_178)
    );

    and_bi _2187_ (
        .b(jinkela_wire_560),
        .a(jinkela_wire_188),
        .c(jinkela_wire_573)
    );

    or_bb _2905_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_178),
        .c(jinkela_wire_1003)
    );

    or_bb _2188_ (
        .b(jinkela_wire_705),
        .a(jinkela_wire_573),
        .c(jinkela_wire_618)
    );

    and_bi _2906_ (
        .b(jinkela_wire_878),
        .a(jinkela_wire_347),
        .c(jinkela_wire_763)
    );

    and_bi _2189_ (
        .b(jinkela_wire_915),
        .a(jinkela_wire_618),
        .c(jinkela_wire_553)
    );

    or_bb _2907_ (
        .b(jinkela_wire_1131),
        .a(jinkela_wire_763),
        .c(jinkela_wire_211)
    );

    or_bb _2190_ (
        .b(jinkela_wire_96),
        .a(jinkela_wire_553),
        .c(jinkela_wire_4)
    );

    and_bi _2908_ (
        .b(jinkela_wire_211),
        .a(jinkela_wire_1003),
        .c(jinkela_wire_388)
    );

    and_bi _2191_ (
        .b(jinkela_wire_15),
        .a(jinkela_wire_4),
        .c(jinkela_wire_1299)
    );

    or_bb _2909_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_388),
        .c(jinkela_wire_753)
    );

    and_bi _2192_ (
        .b(jinkela_wire_1299),
        .a(jinkela_wire_1001),
        .c(jinkela_wire_1418)
    );

    or_bb _2910_ (
        .b(jinkela_wire_185),
        .a(jinkela_wire_753),
        .c(jinkela_wire_601)
    );

    and_bi _2193_ (
        .b(jinkela_wire_1418),
        .a(io_in2_2_),
        .c(jinkela_wire_121)
    );

    and_bb _2911_ (
        .b(jinkela_wire_188),
        .a(jinkela_wire_815),
        .c(jinkela_wire_1231)
    );

    and_bi _2194_ (
        .b(jinkela_wire_121),
        .a(jinkela_wire_1138),
        .c(jinkela_wire_1158)
    );

    or_bb _2912_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_1231),
        .c(jinkela_wire_280)
    );

    and_bi _2195_ (
        .b(jinkela_wire_1158),
        .a(io_in2_3_),
        .c(jinkela_wire_1095)
    );

    and_bi _2913_ (
        .b(jinkela_wire_280),
        .a(jinkela_wire_601),
        .c(jinkela_wire_345)
    );

    and_bi _2196_ (
        .b(jinkela_wire_1095),
        .a(jinkela_wire_1189),
        .c(jinkela_wire_846)
    );

    or_bb _2914_ (
        .b(jinkela_wire_162),
        .a(jinkela_wire_345),
        .c(io_out_20_)
    );

    and_bi _2197_ (
        .b(jinkela_wire_846),
        .a(io_in2_4_),
        .c(jinkela_wire_437)
    );

    and_bi _2915_ (
        .b(jinkela_wire_1389),
        .a(io_adder_out_21_),
        .c(jinkela_wire_518)
    );

    or_bb _2198_ (
        .b(jinkela_wire_318),
        .a(jinkela_wire_437),
        .c(jinkela_wire_1214)
    );

endmodule
