module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 ;
  buffer buf_n69( .i (x4), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n82( .i (x5), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n97( .i (x6), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n38( .i (x2), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n53( .i (x3), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  assign n111 = n42 & n57 ;
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n23( .i (x1), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  assign n115 = n29 | n103 ;
  assign n116 = ( n104 & n113 ) | ( n104 & n115 ) | ( n113 & n115 ) ;
  buffer buf_n8( .i (x0), .o (n8) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  assign n117 = n12 & n86 ;
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  assign n121 = ( n90 & n116 ) | ( n90 & n120 ) | ( n116 & n120 ) ;
  assign n122 = n78 & n121 ;
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  assign n128 = ( n14 & n29 ) | ( n14 & n103 ) | ( n29 & n103 ) ;
  assign n129 = ~n113 & n128 ;
  assign n130 = ( n105 & n114 ) | ( n105 & n129 ) | ( n114 & n129 ) ;
  assign n131 = n91 & n130 ;
  assign n132 = n79 | n131 ;
  assign n133 = ~n123 & n132 ;
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  assign n137 = ( n29 & n103 ) | ( n29 & ~n112 ) | ( n103 & ~n112 ) ;
  buffer buf_n138( .i (n102), .o (n138) );
  assign n139 = ( n75 & n112 ) | ( n75 & n138 ) | ( n112 & n138 ) ;
  assign n140 = n137 & ~n139 ;
  assign n141 = ( n31 & n105 ) | ( n31 & ~n140 ) | ( n105 & ~n140 ) ;
  assign n142 = n17 | n141 ;
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  assign n145 = n108 & n143 ;
  assign n146 = ( n81 & n144 ) | ( n81 & n145 ) | ( n144 & n145 ) ;
  assign n147 = n95 & ~n146 ;
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  assign n148 = ( n30 & n45 ) | ( n30 & ~n76 ) | ( n45 & ~n76 ) ;
  assign n149 = n40 & n99 ;
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  assign n155 = ( n77 & n148 ) | ( n77 & n154 ) | ( n148 & n154 ) ;
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n156( .i (n28), .o (n156) );
  assign n157 = ( ~n59 & n75 ) | ( ~n59 & n156 ) | ( n75 & n156 ) ;
  assign n158 = n138 & n156 ;
  assign n159 = ( n60 & n157 ) | ( n60 & n158 ) | ( n157 & n158 ) ;
  assign n160 = n16 & n159 ;
  assign n161 = ( n17 & n155 ) | ( n17 & n160 ) | ( n155 & n160 ) ;
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  assign n164 = n108 | n162 ;
  assign n165 = ( n81 & n163 ) | ( n81 & n164 ) | ( n163 & n164 ) ;
  assign n166 = n95 | n165 ;
  assign n167 = ( ~n96 & n147 ) | ( ~n96 & n166 ) | ( n147 & n166 ) ;
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n18( .i (n17), .o (n18) );
  assign n168 = ( n12 & ~n42 ) | ( n12 & n57 ) | ( ~n42 & n57 ) ;
  assign n169 = ( n12 & n42 ) | ( n12 & n86 ) | ( n42 & n86 ) ;
  assign n170 = ~n168 & n169 ;
  assign n171 = ( n14 & n59 ) | ( n14 & n170 ) | ( n59 & n170 ) ;
  assign n172 = n30 & n171 ;
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  assign n175 = n91 | n173 ;
  assign n176 = ( n18 & n174 ) | ( n18 & n175 ) | ( n174 & n175 ) ;
  assign n177 = ~n80 & n176 ;
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n46( .i (n45), .o (n46) );
  assign n178 = ( n46 & ~n61 ) | ( n46 & n90 ) | ( ~n61 & n90 ) ;
  assign n179 = n16 | n46 ;
  assign n180 = ( n62 & n178 ) | ( n62 & n179 ) | ( n178 & n179 ) ;
  buffer buf_n181( .i (n11), .o (n181) );
  assign n182 = n57 | n181 ;
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n187 = n16 & n31 ;
  assign n188 = ( n91 & n186 ) | ( n91 & n187 ) | ( n186 & n187 ) ;
  assign n189 = n180 & n188 ;
  assign n190 = n80 & ~n189 ;
  assign n191 = n177 | n190 ;
  buffer buf_n19( .i (n18), .o (n19) );
  assign n192 = n61 & n90 ;
  assign n193 = n78 & n192 ;
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n47( .i (n46), .o (n47) );
  assign n194 = ~n32 & n47 ;
  assign n195 = ( n18 & n193 ) | ( n18 & n194 ) | ( n193 & n194 ) ;
  assign n196 = ~n19 & n195 ;
  buffer buf_n197( .i (n196), .o (n197) );
  assign n198 = ( ~n110 & n191 ) | ( ~n110 & n197 ) | ( n191 & n197 ) ;
  buffer buf_n199( .i (n15), .o (n199) );
  buffer buf_n200( .i (n89), .o (n200) );
  assign n201 = ( ~n31 & n199 ) | ( ~n31 & n200 ) | ( n199 & n200 ) ;
  buffer buf_n202( .i (n30), .o (n202) );
  assign n203 = ( n46 & n199 ) | ( n46 & n202 ) | ( n199 & n202 ) ;
  assign n204 = n201 & ~n203 ;
  assign n205 = ( n18 & n92 ) | ( n18 & ~n204 ) | ( n92 & ~n204 ) ;
  assign n206 = n80 & n205 ;
  assign n207 = ( n44 & n118 ) | ( n44 & n183 ) | ( n118 & n183 ) ;
  buffer buf_n208( .i (n156), .o (n208) );
  assign n209 = n207 | n208 ;
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n200), .o (n212) );
  assign n213 = n210 & n212 ;
  buffer buf_n214( .i (n17), .o (n214) );
  assign n215 = ( n211 & n213 ) | ( n211 & n214 ) | ( n213 & n214 ) ;
  buffer buf_n216( .i (n79), .o (n216) );
  assign n217 = n215 & ~n216 ;
  assign n218 = ( n81 & ~n206 ) | ( n81 & n217 ) | ( ~n206 & n217 ) ;
  assign n219 = ( n110 & n197 ) | ( n110 & ~n218 ) | ( n197 & ~n218 ) ;
  assign n220 = n198 | n219 ;
  assign n221 = ~n199 & n200 ;
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  assign n224 = ( ~n15 & n89 ) | ( ~n15 & n104 ) | ( n89 & n104 ) ;
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  assign n227 = ( n62 & n212 ) | ( n62 & n225 ) | ( n212 & n225 ) ;
  assign n228 = n226 | n227 ;
  assign n229 = ~n223 & n228 ;
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  assign n232 = ~n36 & n230 ;
  assign n233 = ~n34 & n108 ;
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  assign n234 = n61 & ~n199 ;
  assign n235 = ~n212 & n234 ;
  assign n236 = ( n92 & ~n222 ) | ( n92 & n235 ) | ( ~n222 & n235 ) ;
  assign n237 = n49 & n236 ;
  assign n238 = ( n35 & n233 ) | ( n35 & n237 ) | ( n233 & n237 ) ;
  assign n239 = ( ~n47 & n62 ) | ( ~n47 & n212 ) | ( n62 & n212 ) ;
  assign n240 = ( n48 & n214 ) | ( n48 & ~n239 ) | ( n214 & ~n239 ) ;
  assign n241 = ( ~n49 & n223 ) | ( ~n49 & n240 ) | ( n223 & n240 ) ;
  assign n242 = n15 | n89 ;
  assign n243 = ( n86 & n150 ) | ( n86 & n181 ) | ( n150 & n181 ) ;
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  assign n246 = ( n14 & n59 ) | ( n14 & n244 ) | ( n59 & n244 ) ;
  assign n247 = n245 & n246 ;
  assign n248 = n242 & ~n247 ;
  assign n249 = ~n32 & n248 ;
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n107), .o (n252) );
  assign n253 = ~n250 & n252 ;
  assign n254 = ( n241 & n251 ) | ( n241 & ~n253 ) | ( n251 & ~n253 ) ;
  assign n255 = n238 | n254 ;
  assign n256 = ( n231 & ~n232 ) | ( n231 & n255 ) | ( ~n232 & n255 ) ;
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n257( .i (n13), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n60), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  assign n263 = ( n47 & n260 ) | ( n47 & n262 ) | ( n260 & n262 ) ;
  buffer buf_n264( .i (n263), .o (n264) );
  assign n265 = n252 & ~n264 ;
  assign n266 = ~n252 & n264 ;
  assign n267 = n265 | n266 ;
  assign n268 = n36 & ~n267 ;
  buffer buf_n269( .i (n45), .o (n269) );
  assign n270 = n259 & n269 ;
  buffer buf_n271( .i (n269), .o (n271) );
  assign n272 = ( n262 & n270 ) | ( n262 & n271 ) | ( n270 & n271 ) ;
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  assign n275 = n252 | n273 ;
  buffer buf_n276( .i (n107), .o (n276) );
  assign n277 = n273 & ~n276 ;
  assign n278 = ( ~n274 & n275 ) | ( ~n274 & n277 ) | ( n275 & n277 ) ;
  assign n279 = n36 | n278 ;
  assign n280 = ( ~n37 & n268 ) | ( ~n37 & n279 ) | ( n268 & n279 ) ;
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  assign n281 = n34 & n64 ;
  buffer buf_n282( .i (n281), .o (n282) );
  assign n283 = ( ~n19 & n49 ) | ( ~n19 & n64 ) | ( n49 & n64 ) ;
  buffer buf_n284( .i (n283), .o (n284) );
  assign n285 = ( ~n66 & n282 ) | ( ~n66 & n284 ) | ( n282 & n284 ) ;
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  assign n286 = ( n51 & n282 ) | ( n51 & ~n284 ) | ( n282 & ~n284 ) ;
  assign n287 = ( n22 & n285 ) | ( n22 & ~n286 ) | ( n285 & ~n286 ) ;
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n288( .i (n48), .o (n288) );
  assign n289 = n64 | n288 ;
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n292( .i (n35), .o (n292) );
  assign n293 = ( n51 & n290 ) | ( n51 & ~n292 ) | ( n290 & ~n292 ) ;
  assign n294 = ( n51 & ~n290 ) | ( n51 & n292 ) | ( ~n290 & n292 ) ;
  assign n295 = ( ~n52 & n293 ) | ( ~n52 & n294 ) | ( n293 & n294 ) ;
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n296( .i (n50), .o (n296) );
  assign n297 = ~n66 & n296 ;
  assign n298 = ( ~n52 & n291 ) | ( ~n52 & n297 ) | ( n291 & n297 ) ;
  buffer buf_n67( .i (n66), .o (n67) );
  inverter inv_n68( .i (n67), .o (n68) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  assign y0 = n136 ;
  assign y1 = n167 ;
  assign y2 = n220 ;
  assign y3 = n256 ;
  assign y4 = n280 ;
  assign y5 = n287 ;
  assign y6 = n295 ;
  assign y7 = n298 ;
  assign y8 = n68 ;
  assign y9 = n127 ;
endmodule
