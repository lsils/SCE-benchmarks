module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( in_15_ , in_0_ , in_4_ , in_29_ , in_38_ , in_53_ , in_42_ , in_11_ , in_59_ , in_48_ , in_54_ , in_16_ , in_43_ , in_37_ , in_61_ , in_14_ , in_62_ , in_60_ , in_40_ , in_5_ , in_28_ , in_7_ , in_6_ , in_34_ , in_57_ , in_3_ , in_56_ , in_45_ , in_10_ , in_27_ , in_21_ , in_25_ , in_22_ , in_12_ , in_58_ , in_36_ , in_51_ , in_18_ , in_9_ , in_39_ , in_24_ , in_26_ , in_8_ , in_41_ , in_55_ , in_2_ , in_49_ , in_19_ , in_35_ , in_50_ , in_32_ , in_30_ , in_33_ , in_17_ , in_31_ , in_44_ , in_1_ , in_23_ , in_52_ , in_20_ , in_46_ , in_13_ , in_63_ , in_47_ , out_1_ , out_3_ , out_6_ , out_2_ , out_0_ , out_4_ , out_5_ );
  input in_15_ , in_0_ , in_4_ , in_29_ , in_38_ , in_53_ , in_42_ , in_11_ , in_59_ , in_48_ , in_54_ , in_16_ , in_43_ , in_37_ , in_61_ , in_14_ , in_62_ , in_60_ , in_40_ , in_5_ , in_28_ , in_7_ , in_6_ , in_34_ , in_57_ , in_3_ , in_56_ , in_45_ , in_10_ , in_27_ , in_21_ , in_25_ , in_22_ , in_12_ , in_58_ , in_36_ , in_51_ , in_18_ , in_9_ , in_39_ , in_24_ , in_26_ , in_8_ , in_41_ , in_55_ , in_2_ , in_49_ , in_19_ , in_35_ , in_50_ , in_32_ , in_30_ , in_33_ , in_17_ , in_31_ , in_44_ , in_1_ , in_23_ , in_52_ , in_20_ , in_46_ , in_13_ , in_63_ , in_47_ ;
  output out_1_ , out_3_ , out_6_ , out_2_ , out_0_ , out_4_ , out_5_ ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 ;
  assign n65 = in_15_ & in_14_ ;
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  assign n76 = in_12_ | in_13_ ;
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  assign n85 = in_4_ | in_5_ ;
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  assign n89 = in_0_ | in_1_ ;
  buffer buf_n90( .i (n89), .o (n90) );
  assign n91 = in_3_ & in_2_ ;
  buffer buf_n92( .i (n91), .o (n92) );
  assign n93 = ( n86 & n90 ) | ( n86 & n92 ) | ( n90 & n92 ) ;
  buffer buf_n94( .i (n93), .o (n94) );
  assign n100 = ( ~n86 & n90 ) | ( ~n86 & n92 ) | ( n90 & n92 ) ;
  buffer buf_n101( .i (n100), .o (n101) );
  assign n102 = ( n88 & ~n94 ) | ( n88 & n101 ) | ( ~n94 & n101 ) ;
  buffer buf_n103( .i (n102), .o (n103) );
  assign n104 = in_11_ & in_10_ ;
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  assign n108 = in_7_ & in_6_ ;
  buffer buf_n109( .i (n108), .o (n109) );
  assign n110 = in_9_ | in_8_ ;
  buffer buf_n111( .i (n110), .o (n111) );
  assign n112 = ( n105 & n109 ) | ( n105 & n111 ) | ( n109 & n111 ) ;
  buffer buf_n113( .i (n112), .o (n113) );
  assign n119 = ( ~n105 & n109 ) | ( ~n105 & n111 ) | ( n109 & n111 ) ;
  buffer buf_n120( .i (n119), .o (n120) );
  assign n121 = ( n107 & ~n113 ) | ( n107 & n120 ) | ( ~n113 & n120 ) ;
  buffer buf_n122( .i (n121), .o (n122) );
  assign n123 = ( n81 & n103 ) | ( n81 & n122 ) | ( n103 & n122 ) ;
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  assign n128 = ( ~n81 & n103 ) | ( ~n81 & n122 ) | ( n103 & n122 ) ;
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  assign n131 = ( n84 & ~n125 ) | ( n84 & n130 ) | ( ~n125 & n130 ) ;
  buffer buf_n132( .i (n131), .o (n132) );
  assign n133 = n75 & n132 ;
  buffer buf_n134( .i (n133), .o (n134) );
  assign n135 = n75 | n132 ;
  buffer buf_n136( .i (n135), .o (n136) );
  assign n137 = ~n134 & n136 ;
  buffer buf_n138( .i (n137), .o (n138) );
  assign n139 = in_30_ & in_31_ ;
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  assign n150 = in_29_ | in_28_ ;
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  assign n159 = in_21_ | in_20_ ;
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  assign n163 = in_16_ | in_17_ ;
  buffer buf_n164( .i (n163), .o (n164) );
  assign n165 = in_18_ & in_19_ ;
  buffer buf_n166( .i (n165), .o (n166) );
  assign n167 = ( n160 & n164 ) | ( n160 & n166 ) | ( n164 & n166 ) ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n174 = ( ~n160 & n164 ) | ( ~n160 & n166 ) | ( n164 & n166 ) ;
  buffer buf_n175( .i (n174), .o (n175) );
  assign n176 = ( n162 & ~n168 ) | ( n162 & n175 ) | ( ~n168 & n175 ) ;
  buffer buf_n177( .i (n176), .o (n177) );
  assign n178 = in_27_ & in_26_ ;
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  assign n182 = in_22_ & in_23_ ;
  buffer buf_n183( .i (n182), .o (n183) );
  assign n184 = in_25_ | in_24_ ;
  buffer buf_n185( .i (n184), .o (n185) );
  assign n186 = ( n179 & n183 ) | ( n179 & n185 ) | ( n183 & n185 ) ;
  buffer buf_n187( .i (n186), .o (n187) );
  assign n193 = ( ~n179 & n183 ) | ( ~n179 & n185 ) | ( n183 & n185 ) ;
  buffer buf_n194( .i (n193), .o (n194) );
  assign n195 = ( n181 & ~n187 ) | ( n181 & n194 ) | ( ~n187 & n194 ) ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n197 = ( n155 & n177 ) | ( n155 & n196 ) | ( n177 & n196 ) ;
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  assign n202 = ( ~n155 & n177 ) | ( ~n155 & n196 ) | ( n177 & n196 ) ;
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  assign n205 = ( n158 & ~n199 ) | ( n158 & n204 ) | ( ~n199 & n204 ) ;
  buffer buf_n206( .i (n205), .o (n206) );
  assign n207 = n149 & n206 ;
  buffer buf_n208( .i (n207), .o (n208) );
  assign n209 = n149 | n206 ;
  buffer buf_n210( .i (n209), .o (n210) );
  assign n211 = ~n208 & n210 ;
  buffer buf_n212( .i (n211), .o (n212) );
  assign n213 = n138 & n212 ;
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  assign n218 = n138 | n212 ;
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  assign n221 = ~n215 & n220 ;
  buffer buf_n222( .i (n221), .o (n222) );
  assign n223 = in_46_ & in_47_ ;
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  assign n234 = in_45_ | in_44_ ;
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  assign n243 = in_37_ | in_36_ ;
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  assign n247 = in_32_ | in_33_ ;
  buffer buf_n248( .i (n247), .o (n248) );
  assign n249 = in_34_ & in_35_ ;
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = ( n244 & n248 ) | ( n244 & n250 ) | ( n248 & n250 ) ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n258 = ( ~n244 & n248 ) | ( ~n244 & n250 ) | ( n248 & n250 ) ;
  buffer buf_n259( .i (n258), .o (n259) );
  assign n260 = ( n246 & ~n252 ) | ( n246 & n259 ) | ( ~n252 & n259 ) ;
  buffer buf_n261( .i (n260), .o (n261) );
  assign n262 = in_42_ & in_43_ ;
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  assign n266 = in_38_ & in_39_ ;
  buffer buf_n267( .i (n266), .o (n267) );
  assign n268 = in_40_ | in_41_ ;
  buffer buf_n269( .i (n268), .o (n269) );
  assign n270 = ( n263 & n267 ) | ( n263 & n269 ) | ( n267 & n269 ) ;
  buffer buf_n271( .i (n270), .o (n271) );
  assign n277 = ( ~n263 & n267 ) | ( ~n263 & n269 ) | ( n267 & n269 ) ;
  buffer buf_n278( .i (n277), .o (n278) );
  assign n279 = ( n265 & ~n271 ) | ( n265 & n278 ) | ( ~n271 & n278 ) ;
  buffer buf_n280( .i (n279), .o (n280) );
  assign n281 = ( n239 & n261 ) | ( n239 & n280 ) | ( n261 & n280 ) ;
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  assign n286 = ( ~n239 & n261 ) | ( ~n239 & n280 ) | ( n261 & n280 ) ;
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  assign n289 = ( n242 & ~n283 ) | ( n242 & n288 ) | ( ~n283 & n288 ) ;
  buffer buf_n290( .i (n289), .o (n290) );
  assign n291 = n233 & n290 ;
  buffer buf_n292( .i (n291), .o (n292) );
  assign n293 = n233 | n290 ;
  buffer buf_n294( .i (n293), .o (n294) );
  assign n295 = ~n292 & n294 ;
  buffer buf_n296( .i (n295), .o (n296) );
  assign n297 = in_62_ & in_63_ ;
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  assign n308 = in_61_ | in_60_ ;
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  assign n317 = in_53_ | in_52_ ;
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  assign n321 = in_48_ | in_49_ ;
  buffer buf_n322( .i (n321), .o (n322) );
  assign n323 = in_51_ & in_50_ ;
  buffer buf_n324( .i (n323), .o (n324) );
  assign n325 = ( n318 & n322 ) | ( n318 & n324 ) | ( n322 & n324 ) ;
  buffer buf_n326( .i (n325), .o (n326) );
  assign n332 = ( ~n318 & n322 ) | ( ~n318 & n324 ) | ( n322 & n324 ) ;
  buffer buf_n333( .i (n332), .o (n333) );
  assign n334 = ( n320 & ~n326 ) | ( n320 & n333 ) | ( ~n326 & n333 ) ;
  buffer buf_n335( .i (n334), .o (n335) );
  assign n336 = in_59_ & in_58_ ;
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  assign n340 = in_54_ & in_55_ ;
  buffer buf_n341( .i (n340), .o (n341) );
  assign n342 = in_57_ | in_56_ ;
  buffer buf_n343( .i (n342), .o (n343) );
  assign n344 = ( n337 & n341 ) | ( n337 & n343 ) | ( n341 & n343 ) ;
  buffer buf_n345( .i (n344), .o (n345) );
  assign n351 = ( ~n337 & n341 ) | ( ~n337 & n343 ) | ( n341 & n343 ) ;
  buffer buf_n352( .i (n351), .o (n352) );
  assign n353 = ( n339 & ~n345 ) | ( n339 & n352 ) | ( ~n345 & n352 ) ;
  buffer buf_n354( .i (n353), .o (n354) );
  assign n355 = ( n313 & n335 ) | ( n313 & n354 ) | ( n335 & n354 ) ;
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  assign n360 = ( ~n313 & n335 ) | ( ~n313 & n354 ) | ( n335 & n354 ) ;
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  assign n363 = ( n316 & ~n357 ) | ( n316 & n362 ) | ( ~n357 & n362 ) ;
  buffer buf_n364( .i (n363), .o (n364) );
  assign n365 = n307 | n364 ;
  buffer buf_n366( .i (n365), .o (n366) );
  assign n367 = n307 & n364 ;
  buffer buf_n368( .i (n367), .o (n368) );
  assign n369 = n366 & ~n368 ;
  buffer buf_n370( .i (n369), .o (n370) );
  assign n371 = n296 & n370 ;
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  assign n376 = n296 | n370 ;
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  assign n379 = ~n373 & n378 ;
  buffer buf_n380( .i (n379), .o (n380) );
  assign n381 = n222 & n380 ;
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  assign n387 = n222 | n380 ;
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  assign n390 = ~n383 & n389 ;
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  assign n399 = ( n99 & n118 ) | ( n99 & n125 ) | ( n118 & n125 ) ;
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n405( .i (n124), .o (n405) );
  assign n406 = ( n99 & n118 ) | ( n99 & ~n405 ) | ( n118 & ~n405 ) ;
  buffer buf_n407( .i (n406), .o (n407) );
  assign n408 = ( n127 & ~n400 ) | ( n127 & n407 ) | ( ~n400 & n407 ) ;
  buffer buf_n409( .i (n408), .o (n409) );
  assign n410 = n134 & n409 ;
  buffer buf_n411( .i (n410), .o (n411) );
  assign n412 = n404 & n411 ;
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  assign n419 = n404 | n411 ;
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  assign n422 = ~n414 & n421 ;
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  assign n424 = ( n173 & n192 ) | ( n173 & n199 ) | ( n192 & n199 ) ;
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n430( .i (n198), .o (n430) );
  assign n431 = ( n173 & n192 ) | ( n173 & ~n430 ) | ( n192 & ~n430 ) ;
  buffer buf_n432( .i (n431), .o (n432) );
  assign n433 = ( n201 & ~n425 ) | ( n201 & n432 ) | ( ~n425 & n432 ) ;
  buffer buf_n434( .i (n433), .o (n434) );
  assign n435 = n208 & n434 ;
  buffer buf_n436( .i (n435), .o (n436) );
  assign n437 = n429 & n436 ;
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  assign n444 = n429 | n436 ;
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  assign n447 = ~n439 & n446 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = n423 & n448 ;
  assign n450 = n423 | n448 ;
  assign n451 = ~n449 & n450 ;
  buffer buf_n452( .i (n451), .o (n452) );
  assign n453 = n134 | n409 ;
  buffer buf_n454( .i (n453), .o (n454) );
  assign n455 = ~n411 & n454 ;
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  assign n458 = n208 | n434 ;
  buffer buf_n459( .i (n458), .o (n459) );
  assign n460 = ~n436 & n459 ;
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  assign n463 = ( n215 & n457 ) | ( n215 & n462 ) | ( n457 & n462 ) ;
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  assign n468 = n452 & n467 ;
  assign n469 = n452 | n467 ;
  assign n470 = ~n468 & n469 ;
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  assign n472 = ( n257 & n276 ) | ( n257 & n283 ) | ( n276 & n283 ) ;
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n478( .i (n282), .o (n478) );
  assign n479 = ( n257 & n276 ) | ( n257 & ~n478 ) | ( n276 & ~n478 ) ;
  buffer buf_n480( .i (n479), .o (n480) );
  assign n481 = ( n285 & ~n473 ) | ( n285 & n480 ) | ( ~n473 & n480 ) ;
  buffer buf_n482( .i (n481), .o (n482) );
  assign n483 = n292 & n482 ;
  buffer buf_n484( .i (n483), .o (n484) );
  assign n485 = n477 & n484 ;
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  assign n492 = n477 | n484 ;
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  assign n495 = ~n487 & n494 ;
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  assign n497 = ( n331 & n350 ) | ( n331 & n357 ) | ( n350 & n357 ) ;
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n503( .i (n356), .o (n503) );
  assign n504 = ( n331 & n350 ) | ( n331 & ~n503 ) | ( n350 & ~n503 ) ;
  buffer buf_n505( .i (n504), .o (n505) );
  assign n506 = ( n359 & ~n498 ) | ( n359 & n505 ) | ( ~n498 & n505 ) ;
  buffer buf_n507( .i (n506), .o (n507) );
  assign n508 = n368 & n507 ;
  buffer buf_n509( .i (n508), .o (n509) );
  assign n510 = n502 & n509 ;
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  assign n517 = n502 | n509 ;
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  assign n520 = ~n512 & n519 ;
  buffer buf_n521( .i (n520), .o (n521) );
  assign n522 = n496 & n521 ;
  assign n523 = n496 | n521 ;
  assign n524 = ~n522 & n523 ;
  buffer buf_n525( .i (n524), .o (n525) );
  assign n526 = n292 | n482 ;
  buffer buf_n527( .i (n526), .o (n527) );
  assign n528 = ~n484 & n527 ;
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  assign n531 = n368 | n507 ;
  buffer buf_n532( .i (n531), .o (n532) );
  assign n533 = ~n509 & n532 ;
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  assign n536 = ( n373 & n530 ) | ( n373 & n535 ) | ( n530 & n535 ) ;
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  assign n541 = n525 & n540 ;
  assign n542 = n525 | n540 ;
  assign n543 = ~n541 & n542 ;
  buffer buf_n544( .i (n543), .o (n544) );
  assign n545 = n471 & n544 ;
  assign n546 = n471 | n544 ;
  assign n547 = ~n545 & n546 ;
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  assign n549 = n456 & n461 ;
  assign n550 = n456 | n461 ;
  assign n551 = ~n549 & n550 ;
  buffer buf_n552( .i (n551), .o (n552) );
  assign n553 = n217 & n552 ;
  assign n554 = n217 | n552 ;
  assign n555 = ~n553 & n554 ;
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  assign n557 = n529 & n534 ;
  assign n558 = n529 | n534 ;
  assign n559 = ~n557 & n558 ;
  buffer buf_n560( .i (n559), .o (n560) );
  assign n561 = n375 & n560 ;
  assign n562 = n375 | n560 ;
  assign n563 = ~n561 & n562 ;
  buffer buf_n564( .i (n563), .o (n564) );
  assign n565 = ( n383 & n556 ) | ( n383 & n564 ) | ( n556 & n564 ) ;
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  assign n571 = n548 & n570 ;
  assign n572 = n548 | n570 ;
  assign n573 = ~n571 & n572 ;
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  assign n575 = ( n423 & n448 ) | ( n423 & n464 ) | ( n448 & n464 ) ;
  buffer buf_n576( .i (n575), .o (n576) );
  assign n577 = ( n418 & n443 ) | ( n418 & n576 ) | ( n443 & n576 ) ;
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  assign n585 = ( n496 & n521 ) | ( n496 & n537 ) | ( n521 & n537 ) ;
  buffer buf_n586( .i (n585), .o (n586) );
  assign n587 = ( n491 & n516 ) | ( n491 & n586 ) | ( n516 & n586 ) ;
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  assign n595 = n415 & n440 ;
  assign n596 = n415 | n440 ;
  assign n597 = ~n595 & n596 ;
  buffer buf_n598( .i (n597), .o (n598) );
  assign n599 = n576 & n598 ;
  assign n600 = n576 | n598 ;
  assign n601 = ~n599 & n600 ;
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  assign n606 = n488 & n513 ;
  assign n607 = n488 | n513 ;
  assign n608 = ~n606 & n607 ;
  buffer buf_n609( .i (n608), .o (n609) );
  assign n610 = n586 & n609 ;
  assign n611 = n586 | n609 ;
  assign n612 = ~n610 & n611 ;
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  assign n617 = ( n471 & n544 ) | ( n471 & n567 ) | ( n544 & n567 ) ;
  buffer buf_n618( .i (n617), .o (n618) );
  assign n619 = ( n605 & n616 ) | ( n605 & n618 ) | ( n616 & n618 ) ;
  buffer buf_n620( .i (n619), .o (n620) );
  assign n621 = ( n584 & n594 ) | ( n584 & n620 ) | ( n594 & n620 ) ;
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  assign n623 = n556 & n564 ;
  assign n624 = n556 | n564 ;
  assign n625 = ~n623 & n624 ;
  buffer buf_n626( .i (n625), .o (n626) );
  assign n627 = n386 & n626 ;
  assign n628 = n386 | n626 ;
  assign n629 = ~n627 & n628 ;
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  assign n634 = n602 & n613 ;
  assign n635 = n602 | n613 ;
  assign n636 = ~n634 & n635 ;
  buffer buf_n637( .i (n636), .o (n637) );
  assign n638 = n618 & n637 ;
  assign n639 = n618 | n637 ;
  assign n640 = ~n638 & n639 ;
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  assign n643 = n578 & n588 ;
  assign n644 = n578 | n588 ;
  assign n645 = ~n643 & n644 ;
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  assign n650 = n620 & n649 ;
  assign n651 = n620 | n649 ;
  assign n652 = ~n650 & n651 ;
  assign out_1_ = n398 ;
  assign out_3_ = n574 ;
  assign out_6_ = n622 ;
  assign out_2_ = n633 ;
  assign out_0_ = 1'b0 ;
  assign out_4_ = n642 ;
  assign out_5_ = n652 ;
endmodule
