module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( b_4_ , a_6_ , a_7_ , a_1_ , a_0_ , a_2_ , c , b_7_ , a_5_ , b_3_ , b_2_ , b_1_ , b_6_ , a_3_ , b_5_ , a_4_ , b_0_ , cout , s_6_ , s_3_ , s_4_ , s_5_ , s_0_ , s_2_ , s_7_ , s_1_ );
  input b_4_ , a_6_ , a_7_ , a_1_ , a_0_ , a_2_ , c , b_7_ , a_5_ , b_3_ , b_2_ , b_1_ , b_6_ , a_3_ , b_5_ , a_4_ , b_0_ ;
  output cout , s_6_ , s_3_ , s_4_ , s_5_ , s_0_ , s_2_ , s_7_ , s_1_ ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 ;
  assign n18 = a_7_ & b_7_ ;
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  assign n24 = a_7_ | b_7_ ;
  assign n25 = ~n19 & n24 ;
  buffer buf_n26( .i (n25), .o (n26) );
  assign n27 = a_6_ & b_6_ ;
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  assign n33 = a_6_ | b_6_ ;
  assign n34 = ~n28 & n33 ;
  buffer buf_n35( .i (n34), .o (n35) );
  assign n36 = a_5_ & b_5_ ;
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  assign n42 = b_4_ & a_4_ ;
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  assign n48 = b_3_ & a_3_ ;
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  assign n54 = b_3_ | a_3_ ;
  assign n55 = ~n49 & n54 ;
  buffer buf_n56( .i (n55), .o (n56) );
  assign n57 = a_2_ & b_2_ ;
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  assign n63 = a_2_ | b_2_ ;
  assign n64 = ~n58 & n63 ;
  buffer buf_n65( .i (n64), .o (n65) );
  assign n66 = a_1_ & b_1_ ;
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  assign n69 = a_1_ | b_1_ ;
  buffer buf_n70( .i (n69), .o (n70) );
  assign n71 = a_0_ & b_0_ ;
  buffer buf_n72( .i (n71), .o (n72) );
  assign n77 = n70 & n72 ;
  assign n78 = n68 | n77 ;
  buffer buf_n79( .i (n78), .o (n79) );
  assign n80 = n65 & n79 ;
  buffer buf_n81( .i (n80), .o (n81) );
  assign n82 = n62 | n81 ;
  buffer buf_n83( .i (n82), .o (n83) );
  assign n84 = n56 & n83 ;
  buffer buf_n85( .i (n84), .o (n85) );
  assign n86 = n53 | n85 ;
  buffer buf_n87( .i (n86), .o (n87) );
  assign n88 = b_4_ | a_4_ ;
  assign n89 = ~n43 & n88 ;
  buffer buf_n90( .i (n89), .o (n90) );
  assign n91 = n87 & n90 ;
  buffer buf_n92( .i (n91), .o (n92) );
  assign n93 = n47 | n92 ;
  buffer buf_n94( .i (n93), .o (n94) );
  assign n95 = a_5_ | b_5_ ;
  assign n96 = ~n37 & n95 ;
  buffer buf_n97( .i (n96), .o (n97) );
  assign n98 = n94 & n97 ;
  buffer buf_n99( .i (n98), .o (n99) );
  assign n100 = n41 | n99 ;
  buffer buf_n101( .i (n100), .o (n101) );
  assign n102 = n35 & n101 ;
  buffer buf_n103( .i (n102), .o (n103) );
  assign n104 = n32 | n103 ;
  buffer buf_n105( .i (n104), .o (n105) );
  assign n106 = n26 & n105 ;
  buffer buf_n107( .i (n106), .o (n107) );
  assign n108 = n23 | n107 ;
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  assign n112 = n26 | n105 ;
  buffer buf_n113( .i (n112), .o (n113) );
  assign n114 = ~n107 & n113 ;
  buffer buf_n115( .i (n114), .o (n115) );
  assign n116 = n35 | n101 ;
  buffer buf_n117( .i (n116), .o (n117) );
  assign n118 = ~n103 & n117 ;
  buffer buf_n119( .i (n118), .o (n119) );
  assign n120 = n87 | n90 ;
  buffer buf_n121( .i (n120), .o (n121) );
  assign n122 = ~n92 & n121 ;
  buffer buf_n123( .i (n122), .o (n123) );
  assign n124 = n56 | n83 ;
  buffer buf_n125( .i (n124), .o (n125) );
  assign n126 = ~n85 & n125 ;
  buffer buf_n127( .i (n126), .o (n127) );
  assign n128 = n65 | n79 ;
  buffer buf_n129( .i (n128), .o (n129) );
  assign n130 = ~n81 & n129 ;
  buffer buf_n131( .i (n130), .o (n131) );
  assign n132 = ~n67 & n70 ;
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  assign n138 = a_0_ | b_0_ ;
  assign n139 = ~n72 & n138 ;
  buffer buf_n140( .i (n139), .o (n140) );
  assign n141 = c & n140 ;
  buffer buf_n142( .i (n141), .o (n142) );
  assign n143 = n135 & n142 ;
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  assign n146 = n131 & n145 ;
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  assign n150 = n127 & n149 ;
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  assign n154 = n123 & n153 ;
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  assign n158 = n94 | n97 ;
  buffer buf_n159( .i (n158), .o (n159) );
  assign n160 = ~n99 & n159 ;
  buffer buf_n161( .i (n160), .o (n161) );
  assign n162 = n157 & n161 ;
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  assign n166 = n119 & n165 ;
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  assign n170 = n115 & n169 ;
  buffer buf_n171( .i (n170), .o (n171) );
  assign n172 = n111 | n171 ;
  assign n173 = n119 | n165 ;
  buffer buf_n174( .i (n173), .o (n174) );
  assign n175 = ~n167 & n174 ;
  assign n176 = n127 | n149 ;
  buffer buf_n177( .i (n176), .o (n177) );
  assign n178 = ~n151 & n177 ;
  assign n179 = n123 | n153 ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = ~n155 & n180 ;
  assign n182 = n157 | n161 ;
  buffer buf_n183( .i (n182), .o (n183) );
  assign n184 = ~n163 & n183 ;
  assign n185 = c | n140 ;
  buffer buf_n186( .i (n185), .o (n186) );
  assign n187 = ~n142 & n186 ;
  assign n188 = n131 | n145 ;
  buffer buf_n189( .i (n188), .o (n189) );
  assign n190 = ~n147 & n189 ;
  assign n191 = n115 | n169 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = ~n171 & n192 ;
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  assign n194 = n76 | n142 ;
  buffer buf_n195( .i (n194), .o (n195) );
  assign n196 = n137 | n195 ;
  assign n197 = n137 & n195 ;
  assign n198 = n196 & ~n197 ;
  assign cout = n172 ;
  assign s_6_ = n175 ;
  assign s_3_ = n178 ;
  assign s_4_ = n181 ;
  assign s_5_ = n184 ;
  assign s_0_ = n187 ;
  assign s_2_ = n190 ;
  assign s_7_ = n193 ;
  assign s_1_ = n198 ;
endmodule
