module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 ;
  assign n65 = x0 & x15 ;
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  assign n75 = x33 | x61 ;
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  assign n83 = x2 | x19 ;
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  assign n87 = x1 | x56 ;
  buffer buf_n88( .i (n87), .o (n88) );
  assign n89 = x25 & x45 ;
  buffer buf_n90( .i (n89), .o (n90) );
  assign n91 = ( n84 & n88 ) | ( n84 & n90 ) | ( n88 & n90 ) ;
  buffer buf_n92( .i (n91), .o (n92) );
  assign n97 = ( ~n84 & n88 ) | ( ~n84 & n90 ) | ( n88 & n90 ) ;
  buffer buf_n98( .i (n97), .o (n98) );
  assign n99 = ( n86 & ~n92 ) | ( n86 & n98 ) | ( ~n92 & n98 ) ;
  buffer buf_n100( .i (n99), .o (n100) );
  assign n101 = x7 & x28 ;
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  assign n105 = x21 & x22 ;
  buffer buf_n106( .i (n105), .o (n106) );
  assign n107 = x38 | x42 ;
  buffer buf_n108( .i (n107), .o (n108) );
  assign n109 = ( n102 & n106 ) | ( n102 & n108 ) | ( n106 & n108 ) ;
  buffer buf_n110( .i (n109), .o (n110) );
  assign n115 = ( ~n102 & n106 ) | ( ~n102 & n108 ) | ( n106 & n108 ) ;
  buffer buf_n116( .i (n115), .o (n116) );
  assign n117 = ( n104 & ~n110 ) | ( n104 & n116 ) | ( ~n110 & n116 ) ;
  buffer buf_n118( .i (n117), .o (n118) );
  assign n119 = ( n80 & n100 ) | ( n80 & n118 ) | ( n100 & n118 ) ;
  buffer buf_n120( .i (n119), .o (n120) );
  assign n123 = ( ~n80 & n100 ) | ( ~n80 & n118 ) | ( n100 & n118 ) ;
  buffer buf_n124( .i (n123), .o (n124) );
  assign n125 = ( n82 & ~n120 ) | ( n82 & n124 ) | ( ~n120 & n124 ) ;
  buffer buf_n126( .i (n125), .o (n126) );
  assign n127 = n74 & n126 ;
  buffer buf_n128( .i (n127), .o (n128) );
  assign n129 = n74 | n126 ;
  buffer buf_n130( .i (n129), .o (n130) );
  assign n131 = ~n128 & n130 ;
  buffer buf_n132( .i (n131), .o (n132) );
  assign n133 = x51 & x54 ;
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  assign n143 = x3 | x20 ;
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  assign n151 = x30 | x59 ;
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  assign n155 = x11 | x53 ;
  buffer buf_n156( .i (n155), .o (n156) );
  assign n157 = x37 & x47 ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n159 = ( n152 & n156 ) | ( n152 & n158 ) | ( n156 & n158 ) ;
  buffer buf_n160( .i (n159), .o (n160) );
  assign n165 = ( ~n152 & n156 ) | ( ~n152 & n158 ) | ( n156 & n158 ) ;
  buffer buf_n166( .i (n165), .o (n166) );
  assign n167 = ( n154 & ~n160 ) | ( n154 & n166 ) | ( ~n160 & n166 ) ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = x29 & x41 ;
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  assign n173 = x32 & x57 ;
  buffer buf_n174( .i (n173), .o (n174) );
  assign n175 = x31 | x40 ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n177 = ( n170 & n174 ) | ( n170 & n176 ) | ( n174 & n176 ) ;
  buffer buf_n178( .i (n177), .o (n178) );
  assign n183 = ( ~n170 & n174 ) | ( ~n170 & n176 ) | ( n174 & n176 ) ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n185 = ( n172 & ~n178 ) | ( n172 & n184 ) | ( ~n178 & n184 ) ;
  buffer buf_n186( .i (n185), .o (n186) );
  assign n187 = ( n148 & n168 ) | ( n148 & n186 ) | ( n168 & n186 ) ;
  buffer buf_n188( .i (n187), .o (n188) );
  assign n191 = ( ~n148 & n168 ) | ( ~n148 & n186 ) | ( n168 & n186 ) ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = ( n150 & ~n188 ) | ( n150 & n192 ) | ( ~n188 & n192 ) ;
  buffer buf_n194( .i (n193), .o (n194) );
  assign n195 = n142 & n194 ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n197 = n142 | n194 ;
  buffer buf_n198( .i (n197), .o (n198) );
  assign n199 = ~n196 & n198 ;
  buffer buf_n200( .i (n199), .o (n200) );
  assign n201 = n132 & n200 ;
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  assign n206 = n132 | n200 ;
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  assign n209 = ~n203 & n208 ;
  buffer buf_n210( .i (n209), .o (n210) );
  assign n211 = x60 & x63 ;
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  assign n221 = x27 | x55 ;
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  assign n229 = x13 | x35 ;
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  assign n233 = x50 | x52 ;
  buffer buf_n234( .i (n233), .o (n234) );
  assign n235 = x23 & x48 ;
  buffer buf_n236( .i (n235), .o (n236) );
  assign n237 = ( n230 & n234 ) | ( n230 & n236 ) | ( n234 & n236 ) ;
  buffer buf_n238( .i (n237), .o (n238) );
  assign n243 = ( ~n230 & n234 ) | ( ~n230 & n236 ) | ( n234 & n236 ) ;
  buffer buf_n244( .i (n243), .o (n244) );
  assign n245 = ( n232 & ~n238 ) | ( n232 & n244 ) | ( ~n238 & n244 ) ;
  buffer buf_n246( .i (n245), .o (n246) );
  assign n247 = x6 & x12 ;
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = x4 & x39 ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n253 = x18 | x43 ;
  buffer buf_n254( .i (n253), .o (n254) );
  assign n255 = ( n248 & n252 ) | ( n248 & n254 ) | ( n252 & n254 ) ;
  buffer buf_n256( .i (n255), .o (n256) );
  assign n261 = ( ~n248 & n252 ) | ( ~n248 & n254 ) | ( n252 & n254 ) ;
  buffer buf_n262( .i (n261), .o (n262) );
  assign n263 = ( n250 & ~n256 ) | ( n250 & n262 ) | ( ~n256 & n262 ) ;
  buffer buf_n264( .i (n263), .o (n264) );
  assign n265 = ( n226 & n246 ) | ( n226 & n264 ) | ( n246 & n264 ) ;
  buffer buf_n266( .i (n265), .o (n266) );
  assign n269 = ( ~n226 & n246 ) | ( ~n226 & n264 ) | ( n246 & n264 ) ;
  buffer buf_n270( .i (n269), .o (n270) );
  assign n271 = ( n228 & ~n266 ) | ( n228 & n270 ) | ( ~n266 & n270 ) ;
  buffer buf_n272( .i (n271), .o (n272) );
  assign n273 = n220 & n272 ;
  buffer buf_n274( .i (n273), .o (n274) );
  assign n275 = n220 | n272 ;
  buffer buf_n276( .i (n275), .o (n276) );
  assign n277 = ~n274 & n276 ;
  buffer buf_n278( .i (n277), .o (n278) );
  assign n279 = x16 & x62 ;
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  assign n289 = x14 | x17 ;
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  assign n297 = x5 | x58 ;
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  assign n301 = x9 | x46 ;
  buffer buf_n302( .i (n301), .o (n302) );
  assign n303 = x36 & x49 ;
  buffer buf_n304( .i (n303), .o (n304) );
  assign n305 = ( n298 & n302 ) | ( n298 & n304 ) | ( n302 & n304 ) ;
  buffer buf_n306( .i (n305), .o (n306) );
  assign n311 = ( ~n298 & n302 ) | ( ~n298 & n304 ) | ( n302 & n304 ) ;
  buffer buf_n312( .i (n311), .o (n312) );
  assign n313 = ( n300 & ~n306 ) | ( n300 & n312 ) | ( ~n306 & n312 ) ;
  buffer buf_n314( .i (n313), .o (n314) );
  assign n315 = x8 & x34 ;
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  assign n319 = x10 & x44 ;
  buffer buf_n320( .i (n319), .o (n320) );
  assign n321 = x24 | x26 ;
  buffer buf_n322( .i (n321), .o (n322) );
  assign n323 = ( n316 & n320 ) | ( n316 & n322 ) | ( n320 & n322 ) ;
  buffer buf_n324( .i (n323), .o (n324) );
  assign n329 = ( ~n316 & n320 ) | ( ~n316 & n322 ) | ( n320 & n322 ) ;
  buffer buf_n330( .i (n329), .o (n330) );
  assign n331 = ( n318 & ~n324 ) | ( n318 & n330 ) | ( ~n324 & n330 ) ;
  buffer buf_n332( .i (n331), .o (n332) );
  assign n333 = ( n294 & n314 ) | ( n294 & n332 ) | ( n314 & n332 ) ;
  buffer buf_n334( .i (n333), .o (n334) );
  assign n337 = ( ~n294 & n314 ) | ( ~n294 & n332 ) | ( n314 & n332 ) ;
  buffer buf_n338( .i (n337), .o (n338) );
  assign n339 = ( n296 & ~n334 ) | ( n296 & n338 ) | ( ~n334 & n338 ) ;
  buffer buf_n340( .i (n339), .o (n340) );
  assign n341 = n288 | n340 ;
  buffer buf_n342( .i (n341), .o (n342) );
  assign n343 = n288 & n340 ;
  buffer buf_n344( .i (n343), .o (n344) );
  assign n345 = n342 & ~n344 ;
  buffer buf_n346( .i (n345), .o (n346) );
  assign n347 = n278 & n346 ;
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  assign n352 = n278 | n346 ;
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  assign n355 = ~n349 & n354 ;
  buffer buf_n356( .i (n355), .o (n356) );
  assign n357 = n210 & n356 ;
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  assign n363 = n210 | n356 ;
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  assign n366 = ~n359 & n365 ;
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  assign n374 = ( n96 & n114 ) | ( n96 & n120 ) | ( n114 & n120 ) ;
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  assign n380 = ( n96 & n114 ) | ( n96 & ~n120 ) | ( n114 & ~n120 ) ;
  buffer buf_n381( .i (n380), .o (n381) );
  assign n382 = ( n122 & ~n375 ) | ( n122 & n381 ) | ( ~n375 & n381 ) ;
  buffer buf_n383( .i (n382), .o (n383) );
  assign n384 = n128 & n383 ;
  buffer buf_n385( .i (n384), .o (n385) );
  assign n386 = n379 & n385 ;
  buffer buf_n387( .i (n386), .o (n387) );
  assign n392 = n379 | n385 ;
  buffer buf_n393( .i (n392), .o (n393) );
  assign n394 = ~n387 & n393 ;
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  assign n396 = ( n164 & n182 ) | ( n164 & n188 ) | ( n182 & n188 ) ;
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  assign n402 = ( n164 & n182 ) | ( n164 & ~n188 ) | ( n182 & ~n188 ) ;
  buffer buf_n403( .i (n402), .o (n403) );
  assign n404 = ( n190 & ~n397 ) | ( n190 & n403 ) | ( ~n397 & n403 ) ;
  buffer buf_n405( .i (n404), .o (n405) );
  assign n406 = n196 & n405 ;
  buffer buf_n407( .i (n406), .o (n407) );
  assign n408 = n401 & n407 ;
  buffer buf_n409( .i (n408), .o (n409) );
  assign n414 = n401 | n407 ;
  buffer buf_n415( .i (n414), .o (n415) );
  assign n416 = ~n409 & n415 ;
  buffer buf_n417( .i (n416), .o (n417) );
  assign n418 = n395 & n417 ;
  assign n419 = n395 | n417 ;
  assign n420 = ~n418 & n419 ;
  buffer buf_n421( .i (n420), .o (n421) );
  assign n422 = n128 | n383 ;
  buffer buf_n423( .i (n422), .o (n423) );
  assign n424 = ~n385 & n423 ;
  buffer buf_n425( .i (n424), .o (n425) );
  assign n426 = n196 | n405 ;
  buffer buf_n427( .i (n426), .o (n427) );
  assign n428 = ~n407 & n427 ;
  buffer buf_n429( .i (n428), .o (n429) );
  assign n430 = ( n202 & n425 ) | ( n202 & n429 ) | ( n425 & n429 ) ;
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  assign n435 = n421 & n434 ;
  assign n436 = n421 | n434 ;
  assign n437 = ~n435 & n436 ;
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  assign n439 = ( n242 & n260 ) | ( n242 & n266 ) | ( n260 & n266 ) ;
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  assign n445 = ( n242 & n260 ) | ( n242 & ~n266 ) | ( n260 & ~n266 ) ;
  buffer buf_n446( .i (n445), .o (n446) );
  assign n447 = ( n268 & ~n440 ) | ( n268 & n446 ) | ( ~n440 & n446 ) ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = n274 & n448 ;
  buffer buf_n450( .i (n449), .o (n450) );
  assign n451 = n444 & n450 ;
  buffer buf_n452( .i (n451), .o (n452) );
  assign n457 = n444 | n450 ;
  buffer buf_n458( .i (n457), .o (n458) );
  assign n459 = ~n452 & n458 ;
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  assign n461 = ( n310 & n328 ) | ( n310 & n334 ) | ( n328 & n334 ) ;
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  assign n467 = ( n310 & n328 ) | ( n310 & ~n334 ) | ( n328 & ~n334 ) ;
  buffer buf_n468( .i (n467), .o (n468) );
  assign n469 = ( n336 & ~n462 ) | ( n336 & n468 ) | ( ~n462 & n468 ) ;
  buffer buf_n470( .i (n469), .o (n470) );
  assign n471 = n344 & n470 ;
  buffer buf_n472( .i (n471), .o (n472) );
  assign n473 = n466 & n472 ;
  buffer buf_n474( .i (n473), .o (n474) );
  assign n479 = n466 | n472 ;
  buffer buf_n480( .i (n479), .o (n480) );
  assign n481 = ~n474 & n480 ;
  buffer buf_n482( .i (n481), .o (n482) );
  assign n483 = n460 & n482 ;
  assign n484 = n460 | n482 ;
  assign n485 = ~n483 & n484 ;
  buffer buf_n486( .i (n485), .o (n486) );
  assign n487 = n274 | n448 ;
  buffer buf_n488( .i (n487), .o (n488) );
  assign n489 = ~n450 & n488 ;
  buffer buf_n490( .i (n489), .o (n490) );
  assign n491 = n344 | n470 ;
  buffer buf_n492( .i (n491), .o (n492) );
  assign n493 = ~n472 & n492 ;
  buffer buf_n494( .i (n493), .o (n494) );
  assign n495 = ( n348 & n490 ) | ( n348 & n494 ) | ( n490 & n494 ) ;
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  assign n500 = n486 & n499 ;
  assign n501 = n486 | n499 ;
  assign n502 = ~n500 & n501 ;
  buffer buf_n503( .i (n502), .o (n503) );
  assign n504 = n438 & n503 ;
  assign n505 = n438 | n503 ;
  assign n506 = ~n504 & n505 ;
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  assign n508 = n425 & n429 ;
  assign n509 = n425 | n429 ;
  assign n510 = ~n508 & n509 ;
  buffer buf_n511( .i (n510), .o (n511) );
  assign n512 = n205 & n511 ;
  assign n513 = n205 | n511 ;
  assign n514 = ~n512 & n513 ;
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  assign n516 = n490 & n494 ;
  assign n517 = n490 | n494 ;
  assign n518 = ~n516 & n517 ;
  buffer buf_n519( .i (n518), .o (n519) );
  assign n520 = n351 & n519 ;
  assign n521 = n351 | n519 ;
  assign n522 = ~n520 & n521 ;
  buffer buf_n523( .i (n522), .o (n523) );
  assign n524 = ( n359 & n515 ) | ( n359 & n523 ) | ( n515 & n523 ) ;
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  assign n529 = n507 & n528 ;
  assign n530 = n507 | n528 ;
  assign n531 = ~n529 & n530 ;
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  assign n533 = ( n395 & n417 ) | ( n395 & n431 ) | ( n417 & n431 ) ;
  buffer buf_n534( .i (n533), .o (n534) );
  assign n536 = ( n391 & n413 ) | ( n391 & n534 ) | ( n413 & n534 ) ;
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  assign n544 = ( n460 & n482 ) | ( n460 & n496 ) | ( n482 & n496 ) ;
  buffer buf_n545( .i (n544), .o (n545) );
  assign n547 = ( n456 & n478 ) | ( n456 & n545 ) | ( n478 & n545 ) ;
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n535( .i (n534), .o (n535) );
  assign n555 = n389 & n411 ;
  assign n556 = n389 | n411 ;
  assign n557 = ~n555 & n556 ;
  buffer buf_n558( .i (n557), .o (n558) );
  assign n559 = n535 & n558 ;
  assign n560 = n535 | n558 ;
  assign n561 = ~n559 & n560 ;
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n546( .i (n545), .o (n546) );
  assign n565 = n454 & n476 ;
  assign n566 = n454 | n476 ;
  assign n567 = ~n565 & n566 ;
  buffer buf_n568( .i (n567), .o (n568) );
  assign n569 = n546 & n568 ;
  assign n570 = n546 | n568 ;
  assign n571 = ~n569 & n570 ;
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  assign n575 = ( n438 & n503 ) | ( n438 & n525 ) | ( n503 & n525 ) ;
  buffer buf_n576( .i (n575), .o (n576) );
  assign n578 = ( n564 & n574 ) | ( n564 & n576 ) | ( n574 & n576 ) ;
  buffer buf_n579( .i (n578), .o (n579) );
  assign n580 = ( n543 & n554 ) | ( n543 & n579 ) | ( n554 & n579 ) ;
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  assign n582 = n515 & n523 ;
  assign n583 = n515 | n523 ;
  assign n584 = ~n582 & n583 ;
  buffer buf_n585( .i (n584), .o (n585) );
  assign n586 = n362 & n585 ;
  assign n587 = n362 | n585 ;
  assign n588 = ~n586 & n587 ;
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n577( .i (n576), .o (n577) );
  assign n592 = n562 & n572 ;
  assign n593 = n562 | n572 ;
  assign n594 = ~n592 & n593 ;
  buffer buf_n595( .i (n594), .o (n595) );
  assign n596 = n577 & n595 ;
  assign n597 = n577 | n595 ;
  assign n598 = ~n596 & n597 ;
  buffer buf_n599( .i (n598), .o (n599) );
  assign n600 = n540 & n551 ;
  assign n601 = n540 | n551 ;
  assign n602 = ~n600 & n601 ;
  buffer buf_n603( .i (n602), .o (n603) );
  assign n604 = n579 & n603 ;
  assign n605 = n579 | n603 ;
  assign n606 = ~n604 & n605 ;
  assign y0 = n373 ;
  assign y1 = n532 ;
  assign y2 = n581 ;
  assign y3 = n591 ;
  assign y4 = 1'b0 ;
  assign y5 = n599 ;
  assign y6 = n606 ;
endmodule
