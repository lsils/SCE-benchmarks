module adder(b_4_,a_6_,a_7_,a_1_,a_0_,a_2_,c,b_7_,a_5_,b_3_,b_2_,b_1_,b_6_,a_3_,b_5_,a_4_,b_0_,cout,s_6_,s_3_,s_4_,s_5_,s_0_,s_2_,s_7_,s_1_);
    wire jinkela_wire_0;
    wire jinkela_wire_1;
    wire jinkela_wire_2;
    wire jinkela_wire_3;
    wire jinkela_wire_4;
    wire jinkela_wire_5;
    wire jinkela_wire_6;
    wire jinkela_wire_7;
    wire jinkela_wire_8;
    wire jinkela_wire_9;
    wire jinkela_wire_10;
    wire jinkela_wire_11;
    wire jinkela_wire_12;
    wire jinkela_wire_13;
    wire jinkela_wire_14;
    wire jinkela_wire_15;
    wire jinkela_wire_16;
    wire jinkela_wire_17;
    wire jinkela_wire_18;
    wire jinkela_wire_19;
    wire jinkela_wire_20;
    wire jinkela_wire_21;
    wire jinkela_wire_22;
    wire jinkela_wire_23;
    wire jinkela_wire_24;
    wire jinkela_wire_25;
    wire jinkela_wire_26;
    wire jinkela_wire_27;
    wire jinkela_wire_28;
    wire jinkela_wire_29;
    wire jinkela_wire_30;
    wire jinkela_wire_31;
    wire jinkela_wire_32;
    wire jinkela_wire_33;
    wire jinkela_wire_34;
    wire jinkela_wire_35;
    wire jinkela_wire_36;
    wire jinkela_wire_37;
    wire jinkela_wire_38;
    wire jinkela_wire_39;
    wire jinkela_wire_40;
    wire jinkela_wire_41;
    wire jinkela_wire_42;
    wire jinkela_wire_43;
    wire jinkela_wire_44;
    wire jinkela_wire_45;
    wire jinkela_wire_46;
    wire jinkela_wire_47;
    wire jinkela_wire_48;
    wire jinkela_wire_49;
    wire jinkela_wire_50;
    wire jinkela_wire_51;
    wire jinkela_wire_52;
    wire jinkela_wire_53;
    wire jinkela_wire_54;
    wire jinkela_wire_55;
    wire jinkela_wire_56;
    wire jinkela_wire_57;
    wire jinkela_wire_58;
    wire jinkela_wire_59;
    wire jinkela_wire_60;
    wire jinkela_wire_61;
    wire jinkela_wire_62;
    wire jinkela_wire_63;
    wire jinkela_wire_64;
    wire jinkela_wire_65;
    wire jinkela_wire_66;
    wire jinkela_wire_67;
    input b_4_;
    input a_6_;
    input a_7_;
    input a_1_;
    input a_0_;
    input a_2_;
    input c;
    input b_7_;
    input a_5_;
    input b_3_;
    input b_2_;
    input b_1_;
    input b_6_;
    input a_3_;
    input b_5_;
    input a_4_;
    input b_0_;
    output cout;
    output s_6_;
    output s_3_;
    output s_4_;
    output s_5_;
    output s_0_;
    output s_2_;
    output s_7_;
    output s_1_;

    or_bb n_116_ (
        .a(jinkela_wire_20),
        .b(jinkela_wire_40),
        .c(jinkela_wire_55)
    );

    and_ii n_117_ (
        .a(jinkela_wire_55),
        .b(jinkela_wire_63),
        .c(jinkela_wire_28)
    );

    and_bb n_118_ (
        .a(jinkela_wire_55),
        .b(jinkela_wire_63),
        .c(jinkela_wire_23)
    );

    or_bb n_119_ (
        .a(jinkela_wire_23),
        .b(jinkela_wire_28),
        .c(jinkela_wire_32)
    );

    or_bb n_120_ (
        .a(jinkela_wire_32),
        .b(jinkela_wire_13),
        .c(jinkela_wire_66)
    );

    and_bb n_121_ (
        .a(jinkela_wire_32),
        .b(jinkela_wire_13),
        .c(jinkela_wire_17)
    );

    and_bi n_122_ (
        .a(jinkela_wire_66),
        .b(jinkela_wire_17),
        .c(s_5_)
    );

    and_ii n_123_ (
        .a(jinkela_wire_28),
        .b(jinkela_wire_40),
        .c(jinkela_wire_57)
    );

    and_bb n_124_ (
        .a(b_6_),
        .b(a_6_),
        .c(jinkela_wire_54)
    );

    and_ii n_125_ (
        .a(b_6_),
        .b(a_6_),
        .c(jinkela_wire_22)
    );

    or_bb n_126_ (
        .a(jinkela_wire_22),
        .b(jinkela_wire_54),
        .c(jinkela_wire_3)
    );

    and_ii n_127_ (
        .a(jinkela_wire_3),
        .b(jinkela_wire_57),
        .c(jinkela_wire_21)
    );

    and_bb n_128_ (
        .a(jinkela_wire_3),
        .b(jinkela_wire_57),
        .c(jinkela_wire_18)
    );

    or_bb n_129_ (
        .a(jinkela_wire_18),
        .b(jinkela_wire_21),
        .c(jinkela_wire_7)
    );

    or_bb n_130_ (
        .a(jinkela_wire_7),
        .b(jinkela_wire_66),
        .c(jinkela_wire_0)
    );

    and_bb n_131_ (
        .a(jinkela_wire_7),
        .b(jinkela_wire_66),
        .c(jinkela_wire_10)
    );

    and_bi n_132_ (
        .a(jinkela_wire_0),
        .b(jinkela_wire_10),
        .c(s_6_)
    );

    and_ii n_133_ (
        .a(jinkela_wire_21),
        .b(jinkela_wire_54),
        .c(jinkela_wire_51)
    );

    and_bb n_134_ (
        .a(b_7_),
        .b(a_7_),
        .c(jinkela_wire_26)
    );

    and_ii n_135_ (
        .a(b_7_),
        .b(a_7_),
        .c(jinkela_wire_1)
    );

    or_bb n_136_ (
        .a(jinkela_wire_1),
        .b(jinkela_wire_26),
        .c(jinkela_wire_29)
    );

    and_ii n_137_ (
        .a(jinkela_wire_29),
        .b(jinkela_wire_51),
        .c(jinkela_wire_31)
    );

    and_bb n_138_ (
        .a(jinkela_wire_29),
        .b(jinkela_wire_51),
        .c(jinkela_wire_50)
    );

    or_bb n_139_ (
        .a(jinkela_wire_50),
        .b(jinkela_wire_31),
        .c(jinkela_wire_11)
    );

    and_ii n_140_ (
        .a(jinkela_wire_11),
        .b(jinkela_wire_0),
        .c(jinkela_wire_34)
    );

    or_ii n_141_ (
        .a(jinkela_wire_11),
        .b(jinkela_wire_0),
        .c(jinkela_wire_43)
    );

    and_bi n_142_ (
        .a(jinkela_wire_43),
        .b(jinkela_wire_34),
        .c(s_7_)
    );

    or_bb n_143_ (
        .a(jinkela_wire_31),
        .b(jinkela_wire_26),
        .c(jinkela_wire_49)
    );

    or_bb n_144_ (
        .a(jinkela_wire_49),
        .b(jinkela_wire_34),
        .c(cout)
    );

    or_ii n_074_ (
        .a(b_1_),
        .b(a_1_),
        .c(jinkela_wire_42)
    );

    and_ii n_075_ (
        .a(b_1_),
        .b(a_1_),
        .c(jinkela_wire_33)
    );

    and_bi n_076_ (
        .a(jinkela_wire_42),
        .b(jinkela_wire_33),
        .c(jinkela_wire_9)
    );

    and_ii n_077_ (
        .a(jinkela_wire_8),
        .b(jinkela_wire_6),
        .c(jinkela_wire_14)
    );

    or_bi n_078_ (
        .a(jinkela_wire_9),
        .b(jinkela_wire_14),
        .c(jinkela_wire_56)
    );

    and_bi n_079_ (
        .a(jinkela_wire_9),
        .b(jinkela_wire_14),
        .c(jinkela_wire_47)
    );

    and_bi n_080_ (
        .a(jinkela_wire_56),
        .b(jinkela_wire_47),
        .c(s_1_)
    );

    or_ii n_081_ (
        .a(jinkela_wire_9),
        .b(jinkela_wire_8),
        .c(jinkela_wire_46)
    );

    or_ii n_082_ (
        .a(b_2_),
        .b(a_2_),
        .c(jinkela_wire_2)
    );

    or_bb n_083_ (
        .a(b_2_),
        .b(a_2_),
        .c(jinkela_wire_37)
    );

    or_ii n_084_ (
        .a(jinkela_wire_37),
        .b(jinkela_wire_2),
        .c(jinkela_wire_41)
    );

    and_bi n_085_ (
        .a(jinkela_wire_6),
        .b(jinkela_wire_33),
        .c(jinkela_wire_65)
    );

    and_bi n_086_ (
        .a(jinkela_wire_42),
        .b(jinkela_wire_65),
        .c(jinkela_wire_38)
    );

    and_ii n_087_ (
        .a(jinkela_wire_38),
        .b(jinkela_wire_41),
        .c(jinkela_wire_27)
    );

    and_bb n_088_ (
        .a(jinkela_wire_38),
        .b(jinkela_wire_41),
        .c(jinkela_wire_53)
    );

    or_bb n_089_ (
        .a(jinkela_wire_53),
        .b(jinkela_wire_27),
        .c(jinkela_wire_25)
    );

    or_bb n_090_ (
        .a(jinkela_wire_25),
        .b(jinkela_wire_46),
        .c(jinkela_wire_16)
    );

    and_bb n_091_ (
        .a(jinkela_wire_25),
        .b(jinkela_wire_46),
        .c(jinkela_wire_58)
    );

    and_bi n_092_ (
        .a(jinkela_wire_16),
        .b(jinkela_wire_58),
        .c(s_2_)
    );

    and_bi n_093_ (
        .a(jinkela_wire_2),
        .b(jinkela_wire_27),
        .c(jinkela_wire_15)
    );

    and_bb n_094_ (
        .a(b_3_),
        .b(a_3_),
        .c(jinkela_wire_44)
    );

    and_ii n_095_ (
        .a(b_3_),
        .b(a_3_),
        .c(jinkela_wire_60)
    );

    or_bb n_096_ (
        .a(jinkela_wire_60),
        .b(jinkela_wire_44),
        .c(jinkela_wire_48)
    );

    and_ii n_097_ (
        .a(jinkela_wire_48),
        .b(jinkela_wire_15),
        .c(jinkela_wire_5)
    );

    and_bb n_098_ (
        .a(jinkela_wire_48),
        .b(jinkela_wire_15),
        .c(jinkela_wire_35)
    );

    or_bb n_099_ (
        .a(jinkela_wire_35),
        .b(jinkela_wire_5),
        .c(jinkela_wire_62)
    );

    or_bb n_100_ (
        .a(jinkela_wire_62),
        .b(jinkela_wire_16),
        .c(jinkela_wire_12)
    );

    and_bb n_101_ (
        .a(jinkela_wire_62),
        .b(jinkela_wire_16),
        .c(jinkela_wire_59)
    );

    and_bi n_102_ (
        .a(jinkela_wire_12),
        .b(jinkela_wire_59),
        .c(s_3_)
    );

    and_ii n_103_ (
        .a(jinkela_wire_5),
        .b(jinkela_wire_44),
        .c(jinkela_wire_24)
    );

    and_bb n_104_ (
        .a(b_4_),
        .b(a_4_),
        .c(jinkela_wire_30)
    );

    and_ii n_105_ (
        .a(b_4_),
        .b(a_4_),
        .c(jinkela_wire_45)
    );

    and_bb n_068_ (
        .a(b_0_),
        .b(a_0_),
        .c(jinkela_wire_6)
    );

    or_bb n_106_ (
        .a(jinkela_wire_45),
        .b(jinkela_wire_30),
        .c(jinkela_wire_19)
    );

    and_ii n_107_ (
        .a(jinkela_wire_19),
        .b(jinkela_wire_24),
        .c(jinkela_wire_52)
    );

    and_bb n_108_ (
        .a(jinkela_wire_19),
        .b(jinkela_wire_24),
        .c(jinkela_wire_36)
    );

    or_bb n_109_ (
        .a(jinkela_wire_36),
        .b(jinkela_wire_52),
        .c(jinkela_wire_61)
    );

    or_bb n_110_ (
        .a(jinkela_wire_61),
        .b(jinkela_wire_12),
        .c(jinkela_wire_13)
    );

    and_ii n_073_ (
        .a(jinkela_wire_64),
        .b(jinkela_wire_8),
        .c(s_0_)
    );

    and_bb n_111_ (
        .a(jinkela_wire_61),
        .b(jinkela_wire_12),
        .c(jinkela_wire_39)
    );

    and_bi n_071_ (
        .a(c),
        .b(jinkela_wire_4),
        .c(jinkela_wire_8)
    );

    and_ii n_069_ (
        .a(b_0_),
        .b(a_0_),
        .c(jinkela_wire_67)
    );

    and_bi n_112_ (
        .a(jinkela_wire_13),
        .b(jinkela_wire_39),
        .c(s_4_)
    );

    or_bb n_070_ (
        .a(jinkela_wire_67),
        .b(jinkela_wire_6),
        .c(jinkela_wire_4)
    );

    and_ii n_113_ (
        .a(jinkela_wire_52),
        .b(jinkela_wire_30),
        .c(jinkela_wire_63)
    );

    and_bb n_114_ (
        .a(b_5_),
        .b(a_5_),
        .c(jinkela_wire_40)
    );

    and_bi n_072_ (
        .a(jinkela_wire_4),
        .b(c),
        .c(jinkela_wire_64)
    );

    and_ii n_115_ (
        .a(b_5_),
        .b(a_5_),
        .c(jinkela_wire_20)
    );

endmodule
