module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( N1 , N102 , N105 , N108 , N11 , N112 , N115 , N14 , N17 , N21 , N24 , N27 , N30 , N34 , N37 , N4 , N40 , N43 , N47 , N50 , N53 , N56 , N60 , N63 , N66 , N69 , N73 , N76 , N79 , N8 , N82 , N86 , N89 , N92 , N95 , N99 , N223 , N329 , N370 , N421 , N430 , N431 , N432 );
  input N1 , N102 , N105 , N108 , N11 , N112 , N115 , N14 , N17 , N21 , N24 , N27 , N30 , N34 , N37 , N4 , N40 , N43 , N47 , N50 , N53 , N56 , N60 , N63 , N66 , N69 , N73 , N76 , N79 , N8 , N82 , N86 , N89 , N92 , N95 , N99 ;
  output N223 , N329 , N370 , N421 , N430 , N431 , N432 ;
  wire n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 ;
  buffer buf_n209( .i (N24), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n241( .i (N30), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  assign n615 = ~n211 & n243 ;
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n46( .i (N102), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n84( .i (N108), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  assign n622 = ~n49 & n87 ;
  assign n623 = n616 | n622 ;
  buffer buf_n37( .i (N1), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n278( .i (N4), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  assign n624 = ~n39 & n280 ;
  buffer buf_n548( .i (N89), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n586( .i (N95), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  assign n625 = ~n549 & n587 ;
  buffer buf_n462( .i (N76), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n519( .i (N82), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  assign n626 = ~n463 & n520 ;
  assign n627 = n625 | n626 ;
  assign n628 = n624 | n627 ;
  buffer buf_n412( .i (N63), .o (n412) );
  buffer buf_n434( .i (N69), .o (n434) );
  assign n629 = ~n412 & n434 ;
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n269( .i (N37), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n317( .i (N43), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  assign n638 = ~n270 & n318 ;
  assign n639 = n630 | n638 ;
  buffer buf_n346( .i (N50), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n384( .i (N56), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  assign n640 = ~n347 & n385 ;
  buffer buf_n94( .i (N11), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n180( .i (N17), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  assign n641 = ~n95 & n181 ;
  assign n642 = n640 | n641 ;
  assign n643 = n639 | n642 ;
  assign n644 = n628 | n643 ;
  assign n645 = n623 | n644 ;
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n103( .i (N112), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n647( .i (n646), .o (n647) );
  assign n648 = n54 & n647 ;
  assign n649 = n93 & ~n648 ;
  buffer buf_n650( .i (n649), .o (n650) );
  assign n659 = ~n114 & n650 ;
  buffer buf_n529( .i (N86), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  assign n660 = n470 & n647 ;
  assign n661 = n528 & ~n660 ;
  buffer buf_n662( .i (n661), .o (n662) );
  assign n671 = ~n540 & n662 ;
  assign n672 = n659 | n671 ;
  buffer buf_n250( .i (N34), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  assign n673 = n249 & ~n647 ;
  assign n674 = n621 | n673 ;
  buffer buf_n675( .i (n674), .o (n675) );
  assign n684 = ~n261 & n675 ;
  buffer buf_n190( .i (N21), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  assign n685 = n102 & n647 ;
  assign n686 = n189 & ~n685 ;
  buffer buf_n687( .i (n686), .o (n687) );
  assign n696 = ~n201 & n687 ;
  assign n697 = n684 | n696 ;
  assign n698 = n672 | n697 ;
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n500( .i (N8), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n700( .i (n646), .o (n700) );
  assign n701 = n45 & n700 ;
  assign n702 = n287 & ~n701 ;
  buffer buf_n703( .i (n702), .o (n703) );
  assign n712 = ~n511 & n703 ;
  buffer buf_n596( .i (N99), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  assign n713 = n556 & n700 ;
  assign n714 = n595 & ~n713 ;
  buffer buf_n715( .i (n714), .o (n715) );
  assign n724 = ~n607 & n715 ;
  assign n725 = n712 | n724 ;
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n394( .i (N60), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  assign n727 = n354 & n700 ;
  assign n728 = n393 & ~n727 ;
  buffer buf_n729( .i (n728), .o (n729) );
  assign n737 = ~n405 & n729 ;
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n443( .i (N73), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  assign n739 = n442 & ~n700 ;
  assign n740 = n637 | n739 ;
  buffer buf_n741( .i (n740), .o (n741) );
  assign n750 = ~n454 & n741 ;
  buffer buf_n327( .i (N47), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n751( .i (n646), .o (n751) );
  assign n752 = n277 & n751 ;
  assign n753 = n326 & ~n752 ;
  buffer buf_n754( .i (n753), .o (n754) );
  assign n763 = ~n338 & n754 ;
  assign n764 = n750 | n763 ;
  assign n765 = n738 | n764 ;
  assign n766 = n726 | n765 ;
  assign n767 = n699 | n766 ;
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n288( .i (N40), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n769( .i (n768), .o (n769) );
  assign n770 = n268 & n769 ;
  assign n771 = n683 & ~n770 ;
  buffer buf_n772( .i (n771), .o (n772) );
  assign n781 = ~n309 & n772 ;
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n55( .i (N105), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  assign n783 = n614 & n769 ;
  assign n784 = n723 & ~n783 ;
  buffer buf_n785( .i (n784), .o (n785) );
  assign n794 = ~n76 & n785 ;
  buffer buf_n212( .i (N27), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  assign n795 = n208 & n769 ;
  assign n796 = n695 & ~n795 ;
  buffer buf_n797( .i (n796), .o (n797) );
  assign n806 = ~n233 & n797 ;
  assign n807 = n794 | n806 ;
  assign n808 = n782 | n807 ;
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n152( .i (N14), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  assign n810 = n518 & n769 ;
  assign n811 = n711 & ~n810 ;
  buffer buf_n812( .i (n811), .o (n812) );
  assign n820 = ~n173 & n812 ;
  buffer buf_n557( .i (N92), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n821( .i (n768), .o (n821) );
  assign n822 = n547 & n821 ;
  assign n823 = n670 & ~n822 ;
  buffer buf_n824( .i (n823), .o (n824) );
  assign n833 = ~n578 & n824 ;
  assign n834 = n820 | n833 ;
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n471( .i (N79), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  assign n836 = n461 & n821 ;
  assign n837 = n749 & ~n836 ;
  buffer buf_n838( .i (n837), .o (n838) );
  assign n847 = ~n492 & n838 ;
  buffer buf_n413( .i (N66), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  assign n848 = n411 & n768 ;
  assign n849 = n736 & ~n848 ;
  buffer buf_n850( .i (n849), .o (n850) );
  assign n860 = ~n433 & n850 ;
  buffer buf_n861( .i (n860), .o (n861) );
  assign n870 = n847 | n861 ;
  buffer buf_n355( .i (N53), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  assign n871 = n345 & n821 ;
  assign n872 = n762 & ~n871 ;
  buffer buf_n873( .i (n872), .o (n873) );
  assign n882 = ~n376 & n873 ;
  buffer buf_n122( .i (N115), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  assign n883 = n121 & n821 ;
  assign n884 = n658 & ~n883 ;
  buffer buf_n885( .i (n884), .o (n885) );
  assign n895 = ~n143 & n885 ;
  assign n896 = n882 | n895 ;
  assign n897 = n870 | n896 ;
  assign n898 = n835 | n897 ;
  assign n899 = n809 | n898 ;
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n901( .i (n900), .o (n901) );
  assign n903 = n316 & n901 ;
  assign n904 = n780 & ~n903 ;
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  assign n910 = n240 & n901 ;
  assign n911 = n805 & ~n910 ;
  buffer buf_n912( .i (n911), .o (n912) );
  assign n918 = n905 | n912 ;
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  assign n921 = n383 & n901 ;
  assign n922 = n881 & ~n921 ;
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n902( .i (n901), .o (n902) );
  assign n925 = n859 & ~n902 ;
  assign n926 = n869 | n925 ;
  assign n927 = n923 | n926 ;
  buffer buf_n928( .i (n927), .o (n928) );
  assign n929 = n919 | n928 ;
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n931( .i (n900), .o (n931) );
  assign n932 = n585 & n931 ;
  assign n933 = n832 & ~n932 ;
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  assign n935 = n499 & n931 ;
  assign n936 = n846 & ~n935 ;
  buffer buf_n937( .i (n936), .o (n937) );
  assign n940 = n934 | n937 ;
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  assign n942 = n83 & n931 ;
  assign n943 = n793 & ~n942 ;
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  assign n945 = n151 & n902 ;
  assign n946 = n894 & ~n945 ;
  assign n947 = n944 | n946 ;
  buffer buf_n948( .i (n947), .o (n948) );
  assign n949 = n941 | n948 ;
  buffer buf_n950( .i (n949), .o (n950) );
  assign n951 = n930 | n950 ;
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  assign n952 = n179 & n900 ;
  assign n953 = n819 & ~n952 ;
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  assign n961 = n951 & ~n960 ;
  buffer buf_n920( .i (n919), .o (n920) );
  assign n962 = ~n928 & n941 ;
  assign n963 = n920 | n962 ;
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  assign n964 = ~n928 & n939 ;
  buffer buf_n924( .i (n923), .o (n924) );
  assign n965 = ~n934 & n944 ;
  assign n966 = n924 | n965 ;
  buffer buf_n967( .i (n966), .o (n967) );
  assign n968 = n964 | n967 ;
  assign n969 = ~n909 & n968 ;
  assign n970 = n917 | n969 ;
  assign N223 = n646 ;
  assign N329 = n768 ;
  assign N370 = n900 ;
  assign N421 = n961 ;
  assign N430 = n930 ;
  assign N431 = n963 ;
  assign N432 = n970 ;
endmodule
