module top( b_4_ , a_1_ , a_2_ , b_1_ , b_7_ , a_6_ , a_4_ , b_2_ , a_7_ , a_5_ , b_5_ , b_3_ , b_6_ , b_0_ , a_3_ , a_0_ , s_1_ , s_8_ , s_3_ , s_5_ , s_9_ , s_2_ , s_11_ , s_15_ , s_4_ , s_10_ , s_14_ , s_7_ , s_13_ , s_12_ , s_6_ , s_0_ );
  input b_4_ , a_1_ , a_2_ , b_1_ , b_7_ , a_6_ , a_4_ , b_2_ , a_7_ , a_5_ , b_5_ , b_3_ , b_6_ , b_0_ , a_3_ , a_0_ ;
  output s_1_ , s_8_ , s_3_ , s_5_ , s_9_ , s_2_ , s_11_ , s_15_ , s_4_ , s_10_ , s_14_ , s_7_ , s_13_ , s_12_ , s_6_ , s_0_ ;
  wire n53 , n55 , n57 , n65 , n67 , n132 , n142 , n144 , n146 , n152 , n158 , n160 , n162 , n164 , n166 , n172 , n186 , n188 , n190 , n192 , n207 , n221 , n231 , n233 , n235 , n241 , n243 , n245 , n251 , n253 , n255 , n261 , n263 , n265 , n267 , n269 , n276 , n282 , n284 , n286 , n292 , n294 , n296 , n298 , n300 , n307 , n310 , n313 , n319 , n326 , n328 , n330 , n332 , n334 , n335 , n336 , n340 , n343 , n352 , n358 , n364 , n366 , n368 , n370 , n372 , n374 , n376 , n378 , n381 , n387 , n394 , n395 , n396 , n400 , n402 , n404 , n406 , n412 , n414 , n421 , n423 , n425 , n427 , n429 , n435 , n437 , n439 , n441 , n443 , n445 , n447 , n449 , n451 , n454 , n456 , n463 , n469 , n471 , n473 , n475 , n478 , n484 , n486 , n493 , n495 , n497 , n499 , n501 , n507 , n509 , n516 , n518 , n520 , n522 , n524 , n530 , n532 , n534 , n536 , n538 , n540 , n542 , n544 , n546 , n548 , n550 , n554 , n557 , n559 , n565 , n571 , n573 , n575 , n577 , n579 , n585 , n592 , n595 , n597 , n599 , n605 , n607 , n609 , n611 , n617 , n619 , n621 , n623 , n626 , n632 , n642 , n644 , n665 , n667 , n678 , n680 , n682 , n684 , n686 , n692 , n694 , n696 , n698 , n700 , n702 , n712 , n718 , n720 , n722 , n724 , n726 , n728 , n730 , n732 , n734 , n736 , n738 , n744 , n750 , n752 , n754 , n756 , n758 , n765 , n768 , n769 , n772 , n786 , n806 , n816 , n818 , n820 , n822 , n824 , n830 , n832 , n834 , n836 , n839 , n847 , n853 , n855 , n857 , n859 , n861 , n863 , n865 , n867 , n869 , n871 , n873 , n879 , n885 , n887 , n889 , n891 , n893 , n895 , n897 , n903 , n905 , n907 , n909 , n911 , n919 , n924 , n930 , n932 , n934 , n936 , n938 , n940 , n942 , n944 , n946 , n954 , n956 , n958 , n962 , n970 , n975 , n977 , n979 , n981 , n983 , n985 , n987 , n1011 , n1013 , n1062 , n1064 , n1101 , n1103 , n1105 , n1120 , n1135 , n1145 , n1147 , n1153 , n1155 , n1157 , n1159 , n1161 , n1169 , n1176 , n1178 , n1180 , n1183 , n1185 , n1191 , n1193 , n1195 , n1197 , n1200 , n1207 , n1209 , n1211 , n1218 , n1220 , n1226 , n1228 , n1230 , n1232 , n1234 , n1236 , n1238 , n1244 , n1246 , n1248 , n1250 , n1252 , n1254 , n1266 , n1279 , n1289 , n1290 , n1291 , n1312 , n1314 , n1371 , n1373 , n1383 , n1389 , n1403 , n1405 , n1407 , n1409 , n1419 , n1431 , n1434 , n1436 , n1438 , n1440 , n1455 , n1469 , n1475 , n1481 , n1483 , n1485 , n1487 , n1489 , n1491 , n1501 , n1507 , n1509 , n1511 , n1513 , n1515 , n1517 , n1519 , n1521 , n1523 , n1525 , n1527 , n1533 , n1539 , n1541 , n1543 , n1545 , n1547 , n1549 , n1551 , n1557 , n1559 , n1561 , n1563 , n1565 , n1572 , n1574 , n1576 , n1583 , n1589 , n1604 , n1606 , n1608 , n1610 , n1612 , n1633 , n1635 , n1652 , n1654 , n1656 , n1658 , n1675 , n1676 , n1678 , n1680 , n1693 , n1695 , n1697 , n1699 , n1701 , n1714 , n1718 , n1720 , n1742 , n1763 , n1764 , n1765 , n1768 , n1778 , n1786 , n1792 , n1794 , n1796 , n1798 , n1800 , n1802 , n1804 , n1810 , n1818 , n1820 , n1822 , n1824 , n1826 , n1828 , n1872 , n1874 , n1916 , n1918 , n1926 , n1928 , n1934 , n1940 , n1948 , n1950 , n1952 , n1954 , n1956 , n1992 , n1994 , n2026 , n2028 , n2032 , n2034 , n2064 , n2066 , n2092 , n2094 , n2096 , n2098 , n2100 , n2102 , n2104 , n2105 , n2107 , n2152 , n2154 , n2171 , n2173 , n2174 , n2176 , n2204 , n2206 , n2211 , n2213 , n2222 , n2224 , n2256 ;
  buffer buf_n19( .i (a_1_), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n47( .i (b_0_), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  assign n53 = n20 & n48 ;
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n23( .i (b_1_), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n51( .i (a_0_), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  assign n55 = n24 & n52 ;
  buffer buf_n56( .i (n55), .o (n56) );
  assign n57 = n54 & n56 ;
  buffer buf_n58( .i (n57), .o (n58) );
  assign n65 = n54 | n56 ;
  buffer buf_n66( .i (n65), .o (n66) );
  assign n67 = ~n58 & n66 ;
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n41( .i (b_6_), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  assign n132 = n20 & n42 ;
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n17( .i (b_4_), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n21( .i (a_2_), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  assign n142 = n18 & n22 ;
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n39( .i (b_3_), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n49( .i (a_3_), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  assign n144 = n40 & n50 ;
  buffer buf_n145( .i (n144), .o (n145) );
  assign n146 = n143 & n145 ;
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n37( .i (b_5_), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  assign n152 = n20 & n38 ;
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  assign n158 = n143 | n145 ;
  buffer buf_n159( .i (n158), .o (n159) );
  assign n160 = ~n147 & n159 ;
  buffer buf_n161( .i (n160), .o (n161) );
  assign n162 = n157 & n161 ;
  buffer buf_n163( .i (n162), .o (n163) );
  assign n164 = n151 | n163 ;
  buffer buf_n165( .i (n164), .o (n165) );
  assign n166 = n141 & n165 ;
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n25( .i (b_7_), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  assign n172 = n26 & n52 ;
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  assign n186 = n141 | n165 ;
  buffer buf_n187( .i (n186), .o (n187) );
  assign n188 = ~n167 & n187 ;
  buffer buf_n189( .i (n188), .o (n189) );
  assign n190 = n185 & n189 ;
  buffer buf_n191( .i (n190), .o (n191) );
  assign n192 = n171 | n191 ;
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  assign n207 = n20 & n26 ;
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  assign n221 = n22 & n42 ;
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  assign n231 = n18 & n50 ;
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n29( .i (a_4_), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  assign n233 = n30 & n40 ;
  buffer buf_n234( .i (n233), .o (n234) );
  assign n235 = n232 & n234 ;
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  assign n241 = n232 | n234 ;
  buffer buf_n242( .i (n241), .o (n242) );
  assign n243 = ~n236 & n242 ;
  buffer buf_n244( .i (n243), .o (n244) );
  assign n245 = n22 & n38 ;
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = n244 & n250 ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n253 = n240 | n252 ;
  buffer buf_n254( .i (n253), .o (n254) );
  assign n255 = n230 & n254 ;
  buffer buf_n256( .i (n255), .o (n256) );
  assign n261 = n230 | n254 ;
  buffer buf_n262( .i (n261), .o (n262) );
  assign n263 = ~n256 & n262 ;
  buffer buf_n264( .i (n263), .o (n264) );
  assign n265 = n220 & n264 ;
  buffer buf_n266( .i (n265), .o (n266) );
  assign n267 = n220 | n264 ;
  buffer buf_n268( .i (n267), .o (n268) );
  assign n269 = ~n266 & n268 ;
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  assign n276 = n38 & n50 ;
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  assign n282 = n18 & n30 ;
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n35( .i (a_5_), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  assign n284 = n36 & n40 ;
  buffer buf_n285( .i (n284), .o (n285) );
  assign n286 = n283 & n285 ;
  buffer buf_n287( .i (n286), .o (n287) );
  assign n292 = n283 | n285 ;
  buffer buf_n293( .i (n292), .o (n293) );
  assign n294 = ~n287 & n293 ;
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = n281 & n295 ;
  buffer buf_n297( .i (n296), .o (n297) );
  assign n298 = n281 | n295 ;
  buffer buf_n299( .i (n298), .o (n299) );
  assign n300 = ~n297 & n299 ;
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n27( .i (a_6_), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  assign n307 = n24 & n28 ;
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n33( .i (a_7_), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  assign n310 = n34 & n48 ;
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  assign n313 = n309 & n312 ;
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n31( .i (b_2_), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  assign n319 = n32 & n36 ;
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  assign n326 = n309 | n312 ;
  buffer buf_n327( .i (n326), .o (n327) );
  assign n328 = ~n314 & n327 ;
  buffer buf_n329( .i (n328), .o (n329) );
  assign n330 = n325 & n329 ;
  buffer buf_n331( .i (n330), .o (n331) );
  assign n332 = n318 | n331 ;
  buffer buf_n333( .i (n332), .o (n333) );
  assign n334 = n24 & n34 ;
  assign n335 = n28 & n32 ;
  assign n336 = n334 | n335 ;
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  assign n340 = n32 & n34 ;
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  assign n343 = n309 & n342 ;
  buffer buf_n344( .i (n343), .o (n344) );
  assign n352 = n339 & ~n344 ;
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  assign n358 = n333 & n357 ;
  buffer buf_n359( .i (n358), .o (n359) );
  assign n364 = n333 | n357 ;
  buffer buf_n365( .i (n364), .o (n365) );
  assign n366 = ~n359 & n365 ;
  buffer buf_n367( .i (n366), .o (n367) );
  assign n368 = n306 & n367 ;
  buffer buf_n369( .i (n368), .o (n369) );
  assign n370 = n306 | n367 ;
  buffer buf_n371( .i (n370), .o (n371) );
  assign n372 = ~n369 & n371 ;
  buffer buf_n373( .i (n372), .o (n373) );
  assign n374 = n325 | n329 ;
  buffer buf_n375( .i (n374), .o (n375) );
  assign n376 = ~n331 & n375 ;
  buffer buf_n377( .i (n376), .o (n377) );
  assign n378 = n36 & n48 ;
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  assign n381 = n309 & n380 ;
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  assign n387 = n30 & n32 ;
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  assign n394 = n24 & n36 ;
  assign n395 = n28 & n48 ;
  assign n396 = n394 | n395 ;
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  assign n400 = ~n382 & n399 ;
  buffer buf_n401( .i (n400), .o (n401) );
  assign n402 = n393 & n401 ;
  buffer buf_n403( .i (n402), .o (n403) );
  assign n404 = n386 | n403 ;
  buffer buf_n405( .i (n404), .o (n405) );
  assign n406 = n377 & n405 ;
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  assign n412 = n244 | n250 ;
  buffer buf_n413( .i (n412), .o (n413) );
  assign n414 = ~n252 & n413 ;
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  assign n421 = n377 | n405 ;
  buffer buf_n422( .i (n421), .o (n422) );
  assign n423 = ~n407 & n422 ;
  buffer buf_n424( .i (n423), .o (n424) );
  assign n425 = n420 & n424 ;
  buffer buf_n426( .i (n425), .o (n426) );
  assign n427 = n411 | n426 ;
  buffer buf_n428( .i (n427), .o (n428) );
  assign n429 = n373 & n428 ;
  buffer buf_n430( .i (n429), .o (n430) );
  assign n435 = n373 | n428 ;
  buffer buf_n436( .i (n435), .o (n436) );
  assign n437 = ~n430 & n436 ;
  buffer buf_n438( .i (n437), .o (n438) );
  assign n439 = n275 & n438 ;
  buffer buf_n440( .i (n439), .o (n440) );
  assign n441 = n275 | n438 ;
  buffer buf_n442( .i (n441), .o (n442) );
  assign n443 = ~n440 & n442 ;
  buffer buf_n444( .i (n443), .o (n444) );
  assign n445 = n420 | n424 ;
  buffer buf_n446( .i (n445), .o (n446) );
  assign n447 = ~n426 & n446 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = n393 | n401 ;
  buffer buf_n450( .i (n449), .o (n450) );
  assign n451 = ~n403 & n450 ;
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n23), .o (n453) );
  assign n454 = n30 & n453 ;
  buffer buf_n455( .i (n454), .o (n455) );
  assign n456 = n379 & n455 ;
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n31), .o (n462) );
  assign n463 = n50 & n462 ;
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  assign n469 = n379 | n455 ;
  buffer buf_n470( .i (n469), .o (n470) );
  assign n471 = ~n457 & n470 ;
  buffer buf_n472( .i (n471), .o (n472) );
  assign n473 = n468 & n472 ;
  buffer buf_n474( .i (n473), .o (n474) );
  assign n475 = n461 | n474 ;
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  assign n478 = n452 & n477 ;
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  assign n484 = n157 | n161 ;
  buffer buf_n485( .i (n484), .o (n485) );
  assign n486 = ~n163 & n485 ;
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  assign n493 = n452 | n477 ;
  buffer buf_n494( .i (n493), .o (n494) );
  assign n495 = ~n479 & n494 ;
  buffer buf_n496( .i (n495), .o (n496) );
  assign n497 = n492 & n496 ;
  buffer buf_n498( .i (n497), .o (n498) );
  assign n499 = n483 | n498 ;
  buffer buf_n500( .i (n499), .o (n500) );
  assign n501 = n448 & n500 ;
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  assign n507 = n185 | n189 ;
  buffer buf_n508( .i (n507), .o (n508) );
  assign n509 = ~n191 & n508 ;
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  assign n516 = n448 | n500 ;
  buffer buf_n517( .i (n516), .o (n517) );
  assign n518 = ~n502 & n517 ;
  buffer buf_n519( .i (n518), .o (n519) );
  assign n520 = n515 & n519 ;
  buffer buf_n521( .i (n520), .o (n521) );
  assign n522 = n506 | n521 ;
  buffer buf_n523( .i (n522), .o (n523) );
  assign n524 = n444 & n523 ;
  buffer buf_n525( .i (n524), .o (n525) );
  assign n530 = n444 | n523 ;
  buffer buf_n531( .i (n530), .o (n531) );
  assign n532 = ~n525 & n531 ;
  buffer buf_n533( .i (n532), .o (n533) );
  assign n534 = n206 & n533 ;
  buffer buf_n535( .i (n534), .o (n535) );
  assign n536 = n206 | n533 ;
  buffer buf_n537( .i (n536), .o (n537) );
  assign n538 = ~n535 & n537 ;
  buffer buf_n539( .i (n538), .o (n539) );
  assign n540 = n515 | n519 ;
  buffer buf_n541( .i (n540), .o (n541) );
  assign n542 = ~n521 & n541 ;
  buffer buf_n543( .i (n542), .o (n543) );
  assign n544 = n492 | n496 ;
  buffer buf_n545( .i (n544), .o (n545) );
  assign n546 = ~n498 & n545 ;
  buffer buf_n547( .i (n546), .o (n547) );
  assign n548 = n468 | n472 ;
  buffer buf_n549( .i (n548), .o (n549) );
  assign n550 = ~n474 & n549 ;
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n29), .o (n552) );
  buffer buf_n553( .i (n47), .o (n553) );
  assign n554 = n552 & n553 ;
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n49), .o (n556) );
  assign n557 = n453 & n556 ;
  buffer buf_n558( .i (n557), .o (n558) );
  assign n559 = n555 & n558 ;
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  assign n565 = n22 & n462 ;
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  assign n571 = n555 | n558 ;
  buffer buf_n572( .i (n571), .o (n572) );
  assign n573 = ~n560 & n572 ;
  buffer buf_n574( .i (n573), .o (n574) );
  assign n575 = n570 & n574 ;
  buffer buf_n576( .i (n575), .o (n576) );
  assign n577 = n564 | n576 ;
  buffer buf_n578( .i (n577), .o (n578) );
  assign n579 = n551 & n578 ;
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  assign n585 = n38 & n52 ;
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n19), .o (n591) );
  assign n592 = n18 & n591 ;
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n21), .o (n594) );
  assign n595 = n40 & n594 ;
  buffer buf_n596( .i (n595), .o (n596) );
  assign n597 = n593 | n596 ;
  buffer buf_n598( .i (n597), .o (n598) );
  assign n599 = n593 & n596 ;
  buffer buf_n600( .i (n599), .o (n600) );
  assign n605 = n598 & ~n600 ;
  buffer buf_n606( .i (n605), .o (n606) );
  assign n607 = n590 & n606 ;
  buffer buf_n608( .i (n607), .o (n608) );
  assign n609 = n590 | n606 ;
  buffer buf_n610( .i (n609), .o (n610) );
  assign n611 = ~n608 & n610 ;
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  assign n617 = n551 | n578 ;
  buffer buf_n618( .i (n617), .o (n618) );
  assign n619 = ~n580 & n618 ;
  buffer buf_n620( .i (n619), .o (n620) );
  assign n621 = n616 & n620 ;
  buffer buf_n622( .i (n621), .o (n622) );
  assign n623 = n584 | n622 ;
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  assign n626 = n547 & n625 ;
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  assign n632 = n42 & n52 ;
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  assign n642 = n604 | n608 ;
  buffer buf_n643( .i (n642), .o (n643) );
  assign n644 = n641 & n643 ;
  buffer buf_n645( .i (n644), .o (n645) );
  assign n665 = n641 | n643 ;
  buffer buf_n666( .i (n665), .o (n666) );
  assign n667 = ~n645 & n666 ;
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  assign n678 = n547 | n625 ;
  buffer buf_n679( .i (n678), .o (n679) );
  assign n680 = ~n627 & n679 ;
  buffer buf_n681( .i (n680), .o (n681) );
  assign n682 = n677 & n681 ;
  buffer buf_n683( .i (n682), .o (n683) );
  assign n684 = n631 | n683 ;
  buffer buf_n685( .i (n684), .o (n685) );
  assign n686 = n543 & n685 ;
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  assign n692 = n543 | n685 ;
  buffer buf_n693( .i (n692), .o (n693) );
  assign n694 = ~n687 & n693 ;
  buffer buf_n695( .i (n694), .o (n695) );
  assign n696 = n664 & n695 ;
  buffer buf_n697( .i (n696), .o (n697) );
  assign n698 = n691 | n697 ;
  buffer buf_n699( .i (n698), .o (n699) );
  assign n700 = n539 | n699 ;
  buffer buf_n701( .i (n700), .o (n701) );
  assign n702 = n539 & n699 ;
  buffer buf_n703( .i (n702), .o (n703) );
  assign n712 = n701 & ~n703 ;
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  assign n718 = n664 | n695 ;
  buffer buf_n719( .i (n718), .o (n719) );
  assign n720 = ~n697 & n719 ;
  buffer buf_n721( .i (n720), .o (n721) );
  assign n722 = n677 | n681 ;
  buffer buf_n723( .i (n722), .o (n723) );
  assign n724 = ~n683 & n723 ;
  buffer buf_n725( .i (n724), .o (n725) );
  assign n726 = n616 | n620 ;
  buffer buf_n727( .i (n726), .o (n727) );
  assign n728 = ~n622 & n727 ;
  buffer buf_n729( .i (n728), .o (n729) );
  assign n730 = n570 | n574 ;
  buffer buf_n731( .i (n730), .o (n731) );
  assign n732 = ~n576 & n731 ;
  buffer buf_n733( .i (n732), .o (n733) );
  assign n734 = n453 & n594 ;
  buffer buf_n735( .i (n734), .o (n735) );
  assign n736 = n553 & n556 ;
  buffer buf_n737( .i (n736), .o (n737) );
  assign n738 = n735 & n737 ;
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  assign n744 = n462 & n591 ;
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  assign n750 = n735 | n737 ;
  buffer buf_n751( .i (n750), .o (n751) );
  assign n752 = ~n739 & n751 ;
  buffer buf_n753( .i (n752), .o (n753) );
  assign n754 = n749 & n753 ;
  buffer buf_n755( .i (n754), .o (n755) );
  assign n756 = n743 | n755 ;
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = n733 & n757 ;
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n39), .o (n764) );
  assign n765 = n591 & n764 ;
  buffer buf_n766( .i (n17), .o (n766) );
  buffer buf_n767( .i (n51), .o (n767) );
  assign n768 = n766 & n767 ;
  assign n769 = n765 | n768 ;
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  assign n772 = n764 & n767 ;
  buffer buf_n773( .i (n772), .o (n773) );
  assign n786 = n593 & n773 ;
  buffer buf_n787( .i (n786), .o (n787) );
  assign n806 = n771 & ~n787 ;
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  assign n816 = n733 | n757 ;
  buffer buf_n817( .i (n816), .o (n817) );
  assign n818 = ~n759 & n817 ;
  buffer buf_n819( .i (n818), .o (n819) );
  assign n820 = n815 & n819 ;
  buffer buf_n821( .i (n820), .o (n821) );
  assign n822 = n763 | n821 ;
  buffer buf_n823( .i (n822), .o (n823) );
  assign n824 = n729 & n823 ;
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  assign n830 = n729 | n823 ;
  buffer buf_n831( .i (n830), .o (n831) );
  assign n832 = ~n825 & n831 ;
  buffer buf_n833( .i (n832), .o (n833) );
  assign n834 = n805 & n833 ;
  buffer buf_n835( .i (n834), .o (n835) );
  assign n836 = n829 | n835 ;
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  assign n839 = n725 & n838 ;
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  assign n847 = n721 & n846 ;
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  assign n853 = n721 | n846 ;
  buffer buf_n854( .i (n853), .o (n854) );
  assign n855 = ~n848 & n854 ;
  buffer buf_n856( .i (n855), .o (n856) );
  assign n857 = n725 | n838 ;
  buffer buf_n858( .i (n857), .o (n858) );
  assign n859 = ~n840 & n858 ;
  buffer buf_n860( .i (n859), .o (n860) );
  assign n861 = n805 | n833 ;
  buffer buf_n862( .i (n861), .o (n862) );
  assign n863 = ~n835 & n862 ;
  buffer buf_n864( .i (n863), .o (n864) );
  assign n865 = n815 | n819 ;
  buffer buf_n866( .i (n865), .o (n866) );
  assign n867 = ~n821 & n866 ;
  buffer buf_n868( .i (n867), .o (n868) );
  assign n869 = n453 & n591 ;
  buffer buf_n870( .i (n869), .o (n870) );
  assign n871 = n553 & n594 ;
  buffer buf_n872( .i (n871), .o (n872) );
  assign n873 = n870 & n872 ;
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  assign n879 = n462 & n767 ;
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  assign n885 = n870 | n872 ;
  buffer buf_n886( .i (n885), .o (n886) );
  assign n887 = ~n874 & n886 ;
  buffer buf_n888( .i (n887), .o (n888) );
  assign n889 = n884 & n888 ;
  buffer buf_n890( .i (n889), .o (n890) );
  assign n891 = n878 | n890 ;
  buffer buf_n892( .i (n891), .o (n892) );
  assign n893 = n749 | n753 ;
  buffer buf_n894( .i (n893), .o (n894) );
  assign n895 = ~n755 & n894 ;
  buffer buf_n896( .i (n895), .o (n896) );
  assign n897 = n892 & n896 ;
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  assign n903 = n892 | n896 ;
  buffer buf_n904( .i (n903), .o (n904) );
  assign n905 = ~n898 & n904 ;
  buffer buf_n906( .i (n905), .o (n906) );
  assign n907 = n785 & n906 ;
  buffer buf_n908( .i (n907), .o (n908) );
  assign n909 = n902 | n908 ;
  buffer buf_n910( .i (n909), .o (n910) );
  assign n911 = n868 & n910 ;
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  assign n919 = n864 & n918 ;
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  assign n924 = n860 & n923 ;
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  assign n930 = n860 | n923 ;
  buffer buf_n931( .i (n930), .o (n931) );
  assign n932 = ~n925 & n931 ;
  buffer buf_n933( .i (n932), .o (n933) );
  assign n934 = n864 | n918 ;
  buffer buf_n935( .i (n934), .o (n935) );
  assign n936 = ~n920 & n935 ;
  buffer buf_n937( .i (n936), .o (n937) );
  assign n938 = n868 | n910 ;
  buffer buf_n939( .i (n938), .o (n939) );
  assign n940 = ~n912 & n939 ;
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  assign n942 = n884 | n888 ;
  buffer buf_n943( .i (n942), .o (n943) );
  assign n944 = ~n890 & n943 ;
  buffer buf_n945( .i (n944), .o (n945) );
  assign n946 = n64 & n945 ;
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  assign n954 = n785 | n906 ;
  buffer buf_n955( .i (n954), .o (n955) );
  assign n956 = ~n908 & n955 ;
  buffer buf_n957( .i (n956), .o (n957) );
  assign n958 = n953 & n957 ;
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  assign n962 = n941 & n961 ;
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  assign n970 = n937 & n969 ;
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  assign n975 = n933 & n974 ;
  buffer buf_n976( .i (n975), .o (n976) );
  assign n977 = n929 | n976 ;
  buffer buf_n978( .i (n977), .o (n978) );
  assign n979 = n856 & n978 ;
  buffer buf_n980( .i (n979), .o (n980) );
  assign n981 = n852 | n980 ;
  buffer buf_n982( .i (n981), .o (n982) );
  assign n983 = n717 & n982 ;
  buffer buf_n984( .i (n983), .o (n984) );
  assign n985 = n717 | n982 ;
  buffer buf_n986( .i (n985), .o (n986) );
  assign n987 = ~n984 & n986 ;
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  assign n1011 = n953 | n957 ;
  buffer buf_n1012( .i (n1011), .o (n1012) );
  assign n1013 = ~n959 & n1012 ;
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  assign n1062 = n937 | n969 ;
  buffer buf_n1063( .i (n1062), .o (n1063) );
  assign n1064 = ~n971 & n1063 ;
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  assign n1101 = n711 | n984 ;
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  assign n1103 = n529 | n535 ;
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  assign n1105 = n260 | n266 ;
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  assign n1120 = n26 & n594 ;
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n41), .o (n1134) );
  assign n1135 = n556 & n1134 ;
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  assign n1145 = n291 | n297 ;
  buffer buf_n1146( .i (n1145), .o (n1146) );
  assign n1147 = n1144 & n1146 ;
  buffer buf_n1148( .i (n1147), .o (n1148) );
  assign n1153 = n1144 | n1146 ;
  buffer buf_n1154( .i (n1153), .o (n1154) );
  assign n1155 = ~n1148 & n1154 ;
  buffer buf_n1156( .i (n1155), .o (n1156) );
  assign n1157 = n1133 & n1156 ;
  buffer buf_n1158( .i (n1157), .o (n1158) );
  assign n1159 = n1133 | n1156 ;
  buffer buf_n1160( .i (n1159), .o (n1160) );
  assign n1161 = ~n1158 & n1160 ;
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n37), .o (n1168) );
  assign n1169 = n552 & n1168 ;
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n35), .o (n1175) );
  assign n1176 = n766 & n1175 ;
  buffer buf_n1177( .i (n1176), .o (n1177) );
  assign n1178 = n28 & n764 ;
  buffer buf_n1179( .i (n1178), .o (n1179) );
  assign n1180 = n1177 | n1179 ;
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n27), .o (n1182) );
  assign n1183 = n766 & n1182 ;
  buffer buf_n1184( .i (n1183), .o (n1184) );
  assign n1185 = n285 & n1184 ;
  buffer buf_n1186( .i (n1185), .o (n1186) );
  assign n1191 = n1181 & ~n1186 ;
  buffer buf_n1192( .i (n1191), .o (n1192) );
  assign n1193 = n1174 & n1192 ;
  buffer buf_n1194( .i (n1193), .o (n1194) );
  assign n1195 = n1174 | n1192 ;
  buffer buf_n1196( .i (n1195), .o (n1196) );
  assign n1197 = ~n1194 & n1196 ;
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n308), .o (n1199) );
  assign n1200 = n342 & ~n1199 ;
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  assign n1207 = n1198 & n1206 ;
  buffer buf_n1208( .i (n1207), .o (n1208) );
  assign n1209 = n1198 | n1206 ;
  buffer buf_n1210( .i (n1209), .o (n1210) );
  assign n1211 = ~n1208 & n1210 ;
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  assign n1218 = n363 | n369 ;
  buffer buf_n1219( .i (n1218), .o (n1219) );
  assign n1220 = n1217 & n1219 ;
  buffer buf_n1221( .i (n1220), .o (n1221) );
  assign n1226 = n1217 | n1219 ;
  buffer buf_n1227( .i (n1226), .o (n1227) );
  assign n1228 = ~n1221 & n1227 ;
  buffer buf_n1229( .i (n1228), .o (n1229) );
  assign n1230 = n1167 & n1229 ;
  buffer buf_n1231( .i (n1230), .o (n1231) );
  assign n1232 = n1167 | n1229 ;
  buffer buf_n1233( .i (n1232), .o (n1233) );
  assign n1234 = ~n1231 & n1233 ;
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  assign n1236 = n434 | n440 ;
  buffer buf_n1237( .i (n1236), .o (n1237) );
  assign n1238 = n1235 & n1237 ;
  buffer buf_n1239( .i (n1238), .o (n1239) );
  assign n1244 = n1235 | n1237 ;
  buffer buf_n1245( .i (n1244), .o (n1245) );
  assign n1246 = ~n1239 & n1245 ;
  buffer buf_n1247( .i (n1246), .o (n1247) );
  assign n1248 = n1119 & n1247 ;
  buffer buf_n1249( .i (n1248), .o (n1249) );
  assign n1250 = n1119 | n1247 ;
  buffer buf_n1251( .i (n1250), .o (n1251) );
  assign n1252 = ~n1249 & n1251 ;
  buffer buf_n1253( .i (n1252), .o (n1253) );
  assign n1254 = n1104 & n1253 ;
  buffer buf_n1255( .i (n1254), .o (n1255) );
  assign n1266 = n1104 | n1253 ;
  buffer buf_n1267( .i (n1266), .o (n1267) );
  assign n1279 = ~n1255 & n1267 ;
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  assign n1289 = n1102 | n1288 ;
  assign n1290 = n1102 & n1288 ;
  assign n1291 = n1289 & ~n1290 ;
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  assign n1312 = n64 | n945 ;
  buffer buf_n1313( .i (n1312), .o (n1313) );
  assign n1314 = ~n947 & n1313 ;
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  assign n1371 = n1190 | n1194 ;
  buffer buf_n1372( .i (n1371), .o (n1372) );
  assign n1373 = n552 & n1134 ;
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  assign n1383 = n1372 & n1382 ;
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  assign n1389 = n26 & n556 ;
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  assign n1403 = n1372 | n1382 ;
  buffer buf_n1404( .i (n1403), .o (n1404) );
  assign n1405 = ~n1384 & n1404 ;
  buffer buf_n1406( .i (n1405), .o (n1406) );
  assign n1407 = n1402 & n1406 ;
  buffer buf_n1408( .i (n1407), .o (n1408) );
  assign n1409 = n1388 | n1408 ;
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  assign n1419 = n34 & n1168 ;
  buffer buf_n1420( .i (n1419), .o (n1420) );
  assign n1431 = n1184 & n1420 ;
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n33), .o (n1433) );
  assign n1434 = n766 & n1433 ;
  buffer buf_n1435( .i (n1434), .o (n1435) );
  assign n1436 = n1168 & n1182 ;
  buffer buf_n1437( .i (n1436), .o (n1437) );
  assign n1438 = n1435 | n1437 ;
  buffer buf_n1439( .i (n1438), .o (n1439) );
  assign n1440 = ~n1432 & n1439 ;
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n25), .o (n1454) );
  assign n1455 = n552 & n1454 ;
  buffer buf_n1456( .i (n1455), .o (n1456) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  assign n1469 = n1179 & n1435 ;
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  assign n1475 = n1168 & n1175 ;
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  assign n1481 = n764 & n1433 ;
  buffer buf_n1482( .i (n1481), .o (n1482) );
  assign n1483 = n1184 | n1482 ;
  buffer buf_n1484( .i (n1483), .o (n1484) );
  assign n1485 = ~n1470 & n1484 ;
  buffer buf_n1486( .i (n1485), .o (n1486) );
  assign n1487 = n1480 & n1486 ;
  buffer buf_n1488( .i (n1487), .o (n1488) );
  assign n1489 = n1474 | n1488 ;
  buffer buf_n1490( .i (n1489), .o (n1490) );
  assign n1491 = n1134 & n1175 ;
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  assign n1501 = n1490 & n1500 ;
  buffer buf_n1502( .i (n1501), .o (n1502) );
  assign n1507 = n1490 | n1500 ;
  buffer buf_n1508( .i (n1507), .o (n1508) );
  assign n1509 = ~n1502 & n1508 ;
  buffer buf_n1510( .i (n1509), .o (n1510) );
  assign n1511 = n1468 & n1510 ;
  buffer buf_n1512( .i (n1511), .o (n1512) );
  assign n1513 = n1468 | n1510 ;
  buffer buf_n1514( .i (n1513), .o (n1514) );
  assign n1515 = ~n1512 & n1514 ;
  buffer buf_n1516( .i (n1515), .o (n1516) );
  assign n1517 = n1453 & n1516 ;
  buffer buf_n1518( .i (n1517), .o (n1518) );
  assign n1519 = n1453 | n1516 ;
  buffer buf_n1520( .i (n1519), .o (n1520) );
  assign n1521 = ~n1518 & n1520 ;
  buffer buf_n1522( .i (n1521), .o (n1522) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  assign n1523 = n351 | n1208 ;
  buffer buf_n1524( .i (n1523), .o (n1524) );
  assign n1525 = n1480 | n1486 ;
  buffer buf_n1526( .i (n1525), .o (n1526) );
  assign n1527 = ~n1488 & n1526 ;
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  assign n1533 = n1524 & n1532 ;
  buffer buf_n1534( .i (n1533), .o (n1534) );
  buffer buf_n1535( .i (n1534), .o (n1535) );
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  assign n1539 = n1524 | n1532 ;
  buffer buf_n1540( .i (n1539), .o (n1540) );
  assign n1541 = ~n1534 & n1540 ;
  buffer buf_n1542( .i (n1541), .o (n1542) );
  assign n1543 = n1402 | n1406 ;
  buffer buf_n1544( .i (n1543), .o (n1544) );
  assign n1545 = ~n1408 & n1544 ;
  buffer buf_n1546( .i (n1545), .o (n1546) );
  assign n1547 = n1542 & n1546 ;
  buffer buf_n1548( .i (n1547), .o (n1548) );
  assign n1549 = n1538 | n1548 ;
  buffer buf_n1550( .i (n1549), .o (n1550) );
  assign n1551 = n1522 & n1550 ;
  buffer buf_n1552( .i (n1551), .o (n1552) );
  assign n1557 = n1522 | n1550 ;
  buffer buf_n1558( .i (n1557), .o (n1558) );
  assign n1559 = ~n1552 & n1558 ;
  buffer buf_n1560( .i (n1559), .o (n1560) );
  assign n1561 = n1418 & n1560 ;
  buffer buf_n1562( .i (n1561), .o (n1562) );
  assign n1563 = n1418 | n1560 ;
  buffer buf_n1564( .i (n1563), .o (n1564) );
  assign n1565 = ~n1562 & n1564 ;
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  assign n1572 = n1225 | n1231 ;
  buffer buf_n1573( .i (n1572), .o (n1573) );
  assign n1574 = n1542 | n1546 ;
  buffer buf_n1575( .i (n1574), .o (n1575) );
  assign n1576 = ~n1548 & n1575 ;
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  assign n1583 = n1573 & n1582 ;
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  assign n1589 = n1152 | n1158 ;
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  assign n1604 = n1573 | n1582 ;
  buffer buf_n1605( .i (n1604), .o (n1605) );
  assign n1606 = ~n1584 & n1605 ;
  buffer buf_n1607( .i (n1606), .o (n1607) );
  assign n1608 = n1603 & n1607 ;
  buffer buf_n1609( .i (n1608), .o (n1609) );
  assign n1610 = n1588 | n1609 ;
  buffer buf_n1611( .i (n1610), .o (n1611) );
  assign n1612 = n1571 & n1611 ;
  buffer buf_n1613( .i (n1612), .o (n1613) );
  assign n1633 = n1571 | n1611 ;
  buffer buf_n1634( .i (n1633), .o (n1634) );
  assign n1635 = ~n1613 & n1634 ;
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n1637( .i (n1636), .o (n1637) );
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  assign n1652 = n1243 | n1249 ;
  buffer buf_n1653( .i (n1652), .o (n1653) );
  assign n1654 = n1603 | n1607 ;
  buffer buf_n1655( .i (n1654), .o (n1655) );
  assign n1656 = ~n1609 & n1655 ;
  buffer buf_n1657( .i (n1656), .o (n1657) );
  assign n1658 = n1653 & n1657 ;
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  assign n1675 = n1102 | n1265 ;
  assign n1676 = n1278 & n1675 ;
  buffer buf_n1677( .i (n1676), .o (n1677) );
  assign n1678 = n1653 | n1657 ;
  buffer buf_n1679( .i (n1678), .o (n1679) );
  assign n1680 = ~n1659 & n1679 ;
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  assign n1693 = n1677 & n1692 ;
  buffer buf_n1694( .i (n1693), .o (n1694) );
  assign n1695 = n1674 | n1694 ;
  buffer buf_n1696( .i (n1695), .o (n1696) );
  assign n1697 = n1651 | n1696 ;
  buffer buf_n1698( .i (n1697), .o (n1698) );
  assign n1699 = n1651 & n1696 ;
  buffer buf_n1700( .i (n1699), .o (n1700) );
  assign n1701 = n1698 & ~n1700 ;
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  assign n1714 = n1134 & n1182 ;
  buffer buf_n1715( .i (n1714), .o (n1715) );
  assign n1718 = n1433 & n1454 ;
  buffer buf_n1719( .i (n1718), .o (n1719) );
  assign n1720 = n1715 & n1719 ;
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  assign n1742 = ~n1715 & n1719 ;
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n41), .o (n1762) );
  assign n1763 = n1433 & n1762 ;
  assign n1764 = n1182 & n1454 ;
  assign n1765 = n1763 | n1764 ;
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  assign n1768 = ~n1721 & n1767 ;
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  assign n1778 = n1175 & n1454 ;
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  assign n1786 = n46 & n1432 ;
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  assign n1792 = n1432 | n1717 ;
  buffer buf_n1793( .i (n1792), .o (n1793) );
  assign n1794 = ~n1787 & n1793 ;
  buffer buf_n1795( .i (n1794), .o (n1795) );
  assign n1796 = n1785 & n1795 ;
  buffer buf_n1797( .i (n1796), .o (n1797) );
  assign n1798 = n1785 | n1795 ;
  buffer buf_n1799( .i (n1798), .o (n1799) );
  assign n1800 = ~n1797 & n1799 ;
  buffer buf_n1801( .i (n1800), .o (n1801) );
  assign n1802 = n1430 & n1801 ;
  buffer buf_n1803( .i (n1802), .o (n1803) );
  assign n1804 = n1777 & n1803 ;
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  assign n1810 = n1791 | n1797 ;
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  buffer buf_n1813( .i (n1812), .o (n1813) );
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  assign n1818 = n1777 | n1803 ;
  buffer buf_n1819( .i (n1818), .o (n1819) );
  assign n1820 = ~n1805 & n1819 ;
  buffer buf_n1821( .i (n1820), .o (n1821) );
  assign n1822 = n1817 & n1821 ;
  buffer buf_n1823( .i (n1822), .o (n1823) );
  assign n1824 = n1809 | n1823 ;
  buffer buf_n1825( .i (n1824), .o (n1825) );
  assign n1826 = n1761 & n1825 ;
  buffer buf_n1827( .i (n1826), .o (n1827) );
  assign n1828 = n1741 | n1827 ;
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  buffer buf_n1846( .i (n1845), .o (n1846) );
  buffer buf_n1847( .i (n1846), .o (n1847) );
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  assign n1872 = n1761 | n1825 ;
  buffer buf_n1873( .i (n1872), .o (n1873) );
  assign n1874 = ~n1827 & n1873 ;
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  buffer buf_n1879( .i (n1878), .o (n1879) );
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n1888( .i (n1887), .o (n1888) );
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1907( .i (n1906), .o (n1907) );
  buffer buf_n1908( .i (n1907), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n1915( .i (n1914), .o (n1915) );
  assign n1916 = n1817 | n1821 ;
  buffer buf_n1917( .i (n1916), .o (n1917) );
  assign n1918 = ~n1823 & n1917 ;
  buffer buf_n1919( .i (n1918), .o (n1919) );
  buffer buf_n1920( .i (n1919), .o (n1920) );
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  assign n1926 = n1430 | n1801 ;
  buffer buf_n1927( .i (n1926), .o (n1927) );
  assign n1928 = ~n1803 & n1927 ;
  buffer buf_n1929( .i (n1928), .o (n1929) );
  buffer buf_n1930( .i (n1929), .o (n1930) );
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  assign n1934 = n1518 & n1933 ;
  buffer buf_n1935( .i (n1934), .o (n1935) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  assign n1940 = n1506 | n1512 ;
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  assign n1948 = n1518 | n1933 ;
  buffer buf_n1949( .i (n1948), .o (n1949) );
  assign n1950 = ~n1935 & n1949 ;
  buffer buf_n1951( .i (n1950), .o (n1951) );
  assign n1952 = n1947 & n1951 ;
  buffer buf_n1953( .i (n1952), .o (n1953) );
  assign n1954 = n1939 | n1953 ;
  buffer buf_n1955( .i (n1954), .o (n1955) );
  assign n1956 = n1925 & n1955 ;
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  buffer buf_n1960( .i (n1959), .o (n1960) );
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n1967( .i (n1966), .o (n1967) );
  buffer buf_n1968( .i (n1967), .o (n1968) );
  buffer buf_n1969( .i (n1968), .o (n1969) );
  buffer buf_n1970( .i (n1969), .o (n1970) );
  buffer buf_n1971( .i (n1970), .o (n1971) );
  buffer buf_n1972( .i (n1971), .o (n1972) );
  buffer buf_n1973( .i (n1972), .o (n1973) );
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  buffer buf_n1983( .i (n1982), .o (n1983) );
  buffer buf_n1984( .i (n1983), .o (n1984) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n1986( .i (n1985), .o (n1986) );
  buffer buf_n1987( .i (n1986), .o (n1987) );
  buffer buf_n1988( .i (n1987), .o (n1988) );
  buffer buf_n1989( .i (n1988), .o (n1989) );
  buffer buf_n1990( .i (n1989), .o (n1990) );
  buffer buf_n1991( .i (n1990), .o (n1991) );
  assign n1992 = n1925 | n1955 ;
  buffer buf_n1993( .i (n1992), .o (n1993) );
  assign n1994 = ~n1957 & n1993 ;
  buffer buf_n1995( .i (n1994), .o (n1995) );
  buffer buf_n1996( .i (n1995), .o (n1996) );
  buffer buf_n1997( .i (n1996), .o (n1997) );
  buffer buf_n1998( .i (n1997), .o (n1998) );
  buffer buf_n1999( .i (n1998), .o (n1999) );
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n2001( .i (n2000), .o (n2001) );
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n2003), .o (n2004) );
  buffer buf_n2005( .i (n2004), .o (n2005) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n2007( .i (n2006), .o (n2007) );
  buffer buf_n2008( .i (n2007), .o (n2008) );
  buffer buf_n2009( .i (n2008), .o (n2009) );
  buffer buf_n2010( .i (n2009), .o (n2010) );
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n2012( .i (n2011), .o (n2012) );
  buffer buf_n2013( .i (n2012), .o (n2013) );
  buffer buf_n2014( .i (n2013), .o (n2014) );
  buffer buf_n2015( .i (n2014), .o (n2015) );
  buffer buf_n2016( .i (n2015), .o (n2016) );
  buffer buf_n2017( .i (n2016), .o (n2017) );
  buffer buf_n2018( .i (n2017), .o (n2018) );
  buffer buf_n2019( .i (n2018), .o (n2019) );
  buffer buf_n2020( .i (n2019), .o (n2020) );
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2025( .i (n2024), .o (n2025) );
  assign n2026 = n1947 | n1951 ;
  buffer buf_n2027( .i (n2026), .o (n2027) );
  assign n2028 = ~n1953 & n2027 ;
  buffer buf_n2029( .i (n2028), .o (n2029) );
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n2031( .i (n2030), .o (n2031) );
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n1556( .i (n1555), .o (n1556) );
  assign n2032 = n1556 | n1562 ;
  buffer buf_n2033( .i (n2032), .o (n2033) );
  assign n2034 = n2031 & n2033 ;
  buffer buf_n2035( .i (n2034), .o (n2035) );
  buffer buf_n2036( .i (n2035), .o (n2036) );
  buffer buf_n2037( .i (n2036), .o (n2037) );
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  buffer buf_n2055( .i (n2054), .o (n2055) );
  buffer buf_n2056( .i (n2055), .o (n2056) );
  buffer buf_n2057( .i (n2056), .o (n2057) );
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  assign n2064 = n2031 | n2033 ;
  buffer buf_n2065( .i (n2064), .o (n2065) );
  assign n2066 = ~n2035 & n2065 ;
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n2073( .i (n2072), .o (n2073) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n2075( .i (n2074), .o (n2075) );
  buffer buf_n2076( .i (n2075), .o (n2076) );
  buffer buf_n2077( .i (n2076), .o (n2077) );
  buffer buf_n2078( .i (n2077), .o (n2078) );
  buffer buf_n2079( .i (n2078), .o (n2079) );
  buffer buf_n2080( .i (n2079), .o (n2080) );
  buffer buf_n2081( .i (n2080), .o (n2081) );
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2089( .i (n2088), .o (n2089) );
  buffer buf_n2090( .i (n2089), .o (n2090) );
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  assign n2092 = n1632 | n1700 ;
  buffer buf_n2093( .i (n2092), .o (n2093) );
  assign n2094 = n2091 & n2093 ;
  buffer buf_n2095( .i (n2094), .o (n2095) );
  assign n2096 = n2063 | n2095 ;
  buffer buf_n2097( .i (n2096), .o (n2097) );
  assign n2098 = n2025 & n2097 ;
  buffer buf_n2099( .i (n2098), .o (n2099) );
  assign n2100 = n1991 | n2099 ;
  buffer buf_n2101( .i (n2100), .o (n2101) );
  assign n2102 = n1915 & n2101 ;
  buffer buf_n2103( .i (n2102), .o (n2103) );
  assign n2104 = n1871 | n2103 ;
  assign n2105 = n941 | n961 ;
  buffer buf_n2106( .i (n2105), .o (n2106) );
  assign n2107 = ~n963 & n2106 ;
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n2111( .i (n2110), .o (n2111) );
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  buffer buf_n2119( .i (n2118), .o (n2119) );
  buffer buf_n2120( .i (n2119), .o (n2120) );
  buffer buf_n2121( .i (n2120), .o (n2121) );
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  buffer buf_n2129( .i (n2128), .o (n2129) );
  buffer buf_n2130( .i (n2129), .o (n2130) );
  buffer buf_n2131( .i (n2130), .o (n2131) );
  buffer buf_n2132( .i (n2131), .o (n2132) );
  buffer buf_n2133( .i (n2132), .o (n2133) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  buffer buf_n2137( .i (n2136), .o (n2137) );
  buffer buf_n2138( .i (n2137), .o (n2138) );
  buffer buf_n2139( .i (n2138), .o (n2139) );
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n2143( .i (n2142), .o (n2143) );
  buffer buf_n2144( .i (n2143), .o (n2144) );
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  assign n2152 = n1677 | n1692 ;
  buffer buf_n2153( .i (n2152), .o (n2153) );
  assign n2154 = ~n1694 & n2153 ;
  buffer buf_n2155( .i (n2154), .o (n2155) );
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n2158( .i (n2157), .o (n2158) );
  buffer buf_n2159( .i (n2158), .o (n2159) );
  buffer buf_n2160( .i (n2159), .o (n2160) );
  buffer buf_n2161( .i (n2160), .o (n2161) );
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n2163( .i (n2162), .o (n2163) );
  buffer buf_n2164( .i (n2163), .o (n2164) );
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n2166( .i (n2165), .o (n2166) );
  buffer buf_n2167( .i (n2166), .o (n2167) );
  buffer buf_n2168( .i (n2167), .o (n2168) );
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  assign n2171 = n1915 | n2101 ;
  buffer buf_n2172( .i (n2171), .o (n2172) );
  assign n2173 = ~n2103 & n2172 ;
  assign n2174 = n856 | n978 ;
  buffer buf_n2175( .i (n2174), .o (n2175) );
  assign n2176 = ~n980 & n2175 ;
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n2177), .o (n2178) );
  buffer buf_n2179( .i (n2178), .o (n2179) );
  buffer buf_n2180( .i (n2179), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  buffer buf_n2182( .i (n2181), .o (n2182) );
  buffer buf_n2183( .i (n2182), .o (n2183) );
  buffer buf_n2184( .i (n2183), .o (n2184) );
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  buffer buf_n2187( .i (n2186), .o (n2187) );
  buffer buf_n2188( .i (n2187), .o (n2188) );
  buffer buf_n2189( .i (n2188), .o (n2189) );
  buffer buf_n2190( .i (n2189), .o (n2190) );
  buffer buf_n2191( .i (n2190), .o (n2191) );
  buffer buf_n2192( .i (n2191), .o (n2192) );
  buffer buf_n2193( .i (n2192), .o (n2193) );
  buffer buf_n2194( .i (n2193), .o (n2194) );
  buffer buf_n2195( .i (n2194), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  buffer buf_n2197( .i (n2196), .o (n2197) );
  buffer buf_n2198( .i (n2197), .o (n2198) );
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n2200( .i (n2199), .o (n2200) );
  buffer buf_n2201( .i (n2200), .o (n2201) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  buffer buf_n2203( .i (n2202), .o (n2203) );
  assign n2204 = n2025 | n2097 ;
  buffer buf_n2205( .i (n2204), .o (n2205) );
  assign n2206 = ~n2099 & n2205 ;
  buffer buf_n2207( .i (n2206), .o (n2207) );
  buffer buf_n2208( .i (n2207), .o (n2208) );
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  assign n2211 = n2091 | n2093 ;
  buffer buf_n2212( .i (n2211), .o (n2212) );
  assign n2213 = ~n2095 & n2212 ;
  buffer buf_n2214( .i (n2213), .o (n2214) );
  buffer buf_n2215( .i (n2214), .o (n2215) );
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n2221( .i (n2220), .o (n2221) );
  assign n2222 = n933 | n974 ;
  buffer buf_n2223( .i (n2222), .o (n2223) );
  assign n2224 = ~n976 & n2223 ;
  buffer buf_n2225( .i (n2224), .o (n2225) );
  buffer buf_n2226( .i (n2225), .o (n2226) );
  buffer buf_n2227( .i (n2226), .o (n2227) );
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  buffer buf_n2231( .i (n2230), .o (n2231) );
  buffer buf_n2232( .i (n2231), .o (n2232) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  buffer buf_n2235( .i (n2234), .o (n2235) );
  buffer buf_n2236( .i (n2235), .o (n2236) );
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  buffer buf_n2250( .i (n2249), .o (n2250) );
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  assign n2256 = n553 & n767 ;
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  buffer buf_n2265( .i (n2264), .o (n2265) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  buffer buf_n2269( .i (n2268), .o (n2269) );
  buffer buf_n2270( .i (n2269), .o (n2270) );
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2273( .i (n2272), .o (n2273) );
  buffer buf_n2274( .i (n2273), .o (n2274) );
  buffer buf_n2275( .i (n2274), .o (n2275) );
  buffer buf_n2276( .i (n2275), .o (n2276) );
  buffer buf_n2277( .i (n2276), .o (n2277) );
  buffer buf_n2278( .i (n2277), .o (n2278) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  buffer buf_n2280( .i (n2279), .o (n2280) );
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n2289( .i (n2288), .o (n2289) );
  buffer buf_n2290( .i (n2289), .o (n2290) );
  buffer buf_n2291( .i (n2290), .o (n2291) );
  buffer buf_n2292( .i (n2291), .o (n2292) );
  buffer buf_n2293( .i (n2292), .o (n2293) );
  buffer buf_n2294( .i (n2293), .o (n2294) );
  buffer buf_n2295( .i (n2294), .o (n2295) );
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n2297( .i (n2296), .o (n2297) );
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  buffer buf_n2307( .i (n2306), .o (n2307) );
  buffer buf_n2308( .i (n2307), .o (n2308) );
  buffer buf_n2309( .i (n2308), .o (n2309) );
  buffer buf_n2310( .i (n2309), .o (n2310) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n2321( .i (n2320), .o (n2321) );
  buffer buf_n2322( .i (n2321), .o (n2322) );
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  assign s_1_ = n131 ;
  assign s_8_ = n1010 ;
  assign s_3_ = n1061 ;
  assign s_5_ = n1100 ;
  assign s_9_ = n1311 ;
  assign s_2_ = n1370 ;
  assign s_11_ = n1713 ;
  assign s_15_ = n2104 ;
  assign s_4_ = n2151 ;
  assign s_10_ = n2170 ;
  assign s_14_ = n2173 ;
  assign s_7_ = n2203 ;
  assign s_13_ = n2210 ;
  assign s_12_ = n2221 ;
  assign s_6_ = n2255 ;
  assign s_0_ = n2324 ;
endmodule
