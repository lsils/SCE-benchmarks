module sorter48(a_44_,a_5_,a_38_,a_43_,a_20_,a_27_,a_8_,a_40_,a_47_,a_11_,a_0_,a_6_,a_16_,a_9_,a_31_,a_4_,a_30_,a_35_,a_26_,a_19_,a_7_,a_13_,a_45_,a_34_,a_42_,a_14_,a_41_,a_17_,a_37_,a_18_,a_29_,a_21_,a_32_,a_22_,a_36_,a_3_,a_28_,a_46_,a_25_,a_10_,a_12_,a_33_,a_24_,a_1_,a_15_,a_2_,a_39_,a_23_,b_47_,b_43_,b_40_,b_11_,b_7_,b_5_,b_32_,b_17_,b_29_,b_25_,b_12_,b_16_,b_1_,b_42_,b_0_,b_28_,b_9_,b_36_,b_2_,b_20_,b_41_,b_33_,b_31_,b_34_,b_13_,b_21_,b_35_,b_39_,b_27_,b_46_,b_4_,b_14_,b_37_,b_22_,b_6_,b_38_,b_18_,b_15_,b_30_,b_8_,b_26_,b_24_,b_19_,b_23_,b_10_,b_3_,b_45_,b_44_);
    wire jinkela_wire_0;
    wire jinkela_wire_1;
    wire jinkela_wire_2;
    wire jinkela_wire_3;
    wire jinkela_wire_4;
    wire jinkela_wire_5;
    wire jinkela_wire_6;
    wire jinkela_wire_7;
    wire jinkela_wire_8;
    wire jinkela_wire_9;
    wire jinkela_wire_10;
    wire jinkela_wire_11;
    wire jinkela_wire_12;
    wire jinkela_wire_13;
    wire jinkela_wire_14;
    wire jinkela_wire_15;
    wire jinkela_wire_16;
    wire jinkela_wire_17;
    wire jinkela_wire_18;
    wire jinkela_wire_19;
    wire jinkela_wire_20;
    wire jinkela_wire_21;
    wire jinkela_wire_22;
    wire jinkela_wire_23;
    wire jinkela_wire_24;
    wire jinkela_wire_25;
    wire jinkela_wire_26;
    wire jinkela_wire_27;
    wire jinkela_wire_28;
    wire jinkela_wire_29;
    wire jinkela_wire_30;
    wire jinkela_wire_31;
    wire jinkela_wire_32;
    wire jinkela_wire_33;
    wire jinkela_wire_34;
    wire jinkela_wire_35;
    wire jinkela_wire_36;
    wire jinkela_wire_37;
    wire jinkela_wire_38;
    wire jinkela_wire_39;
    wire jinkela_wire_40;
    wire jinkela_wire_41;
    wire jinkela_wire_42;
    wire jinkela_wire_43;
    wire jinkela_wire_44;
    wire jinkela_wire_45;
    wire jinkela_wire_46;
    wire jinkela_wire_47;
    wire jinkela_wire_48;
    wire jinkela_wire_49;
    wire jinkela_wire_50;
    wire jinkela_wire_51;
    wire jinkela_wire_52;
    wire jinkela_wire_53;
    wire jinkela_wire_54;
    wire jinkela_wire_55;
    wire jinkela_wire_56;
    wire jinkela_wire_57;
    wire jinkela_wire_58;
    wire jinkela_wire_59;
    wire jinkela_wire_60;
    wire jinkela_wire_61;
    wire jinkela_wire_62;
    wire jinkela_wire_63;
    wire jinkela_wire_64;
    wire jinkela_wire_65;
    wire jinkela_wire_66;
    wire jinkela_wire_67;
    wire jinkela_wire_68;
    wire jinkela_wire_69;
    wire jinkela_wire_70;
    wire jinkela_wire_71;
    wire jinkela_wire_72;
    wire jinkela_wire_73;
    wire jinkela_wire_74;
    wire jinkela_wire_75;
    wire jinkela_wire_76;
    wire jinkela_wire_77;
    wire jinkela_wire_78;
    wire jinkela_wire_79;
    wire jinkela_wire_80;
    wire jinkela_wire_81;
    wire jinkela_wire_82;
    wire jinkela_wire_83;
    wire jinkela_wire_84;
    wire jinkela_wire_85;
    wire jinkela_wire_86;
    wire jinkela_wire_87;
    wire jinkela_wire_88;
    wire jinkela_wire_89;
    wire jinkela_wire_90;
    wire jinkela_wire_91;
    wire jinkela_wire_92;
    wire jinkela_wire_93;
    wire jinkela_wire_94;
    wire jinkela_wire_95;
    wire jinkela_wire_96;
    wire jinkela_wire_97;
    wire jinkela_wire_98;
    wire jinkela_wire_99;
    wire jinkela_wire_100;
    wire jinkela_wire_101;
    wire jinkela_wire_102;
    wire jinkela_wire_103;
    wire jinkela_wire_104;
    wire jinkela_wire_105;
    wire jinkela_wire_106;
    wire jinkela_wire_107;
    wire jinkela_wire_108;
    wire jinkela_wire_109;
    wire jinkela_wire_110;
    wire jinkela_wire_111;
    wire jinkela_wire_112;
    wire jinkela_wire_113;
    wire jinkela_wire_114;
    wire jinkela_wire_115;
    wire jinkela_wire_116;
    wire jinkela_wire_117;
    wire jinkela_wire_118;
    wire jinkela_wire_119;
    wire jinkela_wire_120;
    wire jinkela_wire_121;
    wire jinkela_wire_122;
    wire jinkela_wire_123;
    wire jinkela_wire_124;
    wire jinkela_wire_125;
    wire jinkela_wire_126;
    wire jinkela_wire_127;
    wire jinkela_wire_128;
    wire jinkela_wire_129;
    wire jinkela_wire_130;
    wire jinkela_wire_131;
    wire jinkela_wire_132;
    wire jinkela_wire_133;
    wire jinkela_wire_134;
    wire jinkela_wire_135;
    wire jinkela_wire_136;
    wire jinkela_wire_137;
    wire jinkela_wire_138;
    wire jinkela_wire_139;
    wire jinkela_wire_140;
    wire jinkela_wire_141;
    wire jinkela_wire_142;
    wire jinkela_wire_143;
    wire jinkela_wire_144;
    wire jinkela_wire_145;
    wire jinkela_wire_146;
    wire jinkela_wire_147;
    wire jinkela_wire_148;
    wire jinkela_wire_149;
    wire jinkela_wire_150;
    wire jinkela_wire_151;
    wire jinkela_wire_152;
    wire jinkela_wire_153;
    wire jinkela_wire_154;
    wire jinkela_wire_155;
    wire jinkela_wire_156;
    wire jinkela_wire_157;
    wire jinkela_wire_158;
    wire jinkela_wire_159;
    wire jinkela_wire_160;
    wire jinkela_wire_161;
    wire jinkela_wire_162;
    wire jinkela_wire_163;
    wire jinkela_wire_164;
    wire jinkela_wire_165;
    wire jinkela_wire_166;
    wire jinkela_wire_167;
    wire jinkela_wire_168;
    wire jinkela_wire_169;
    wire jinkela_wire_170;
    wire jinkela_wire_171;
    wire jinkela_wire_172;
    wire jinkela_wire_173;
    wire jinkela_wire_174;
    wire jinkela_wire_175;
    wire jinkela_wire_176;
    wire jinkela_wire_177;
    wire jinkela_wire_178;
    wire jinkela_wire_179;
    wire jinkela_wire_180;
    wire jinkela_wire_181;
    wire jinkela_wire_182;
    wire jinkela_wire_183;
    wire jinkela_wire_184;
    wire jinkela_wire_185;
    wire jinkela_wire_186;
    wire jinkela_wire_187;
    wire jinkela_wire_188;
    wire jinkela_wire_189;
    wire jinkela_wire_190;
    wire jinkela_wire_191;
    wire jinkela_wire_192;
    wire jinkela_wire_193;
    wire jinkela_wire_194;
    wire jinkela_wire_195;
    wire jinkela_wire_196;
    wire jinkela_wire_197;
    wire jinkela_wire_198;
    wire jinkela_wire_199;
    wire jinkela_wire_200;
    wire jinkela_wire_201;
    wire jinkela_wire_202;
    wire jinkela_wire_203;
    wire jinkela_wire_204;
    wire jinkela_wire_205;
    wire jinkela_wire_206;
    wire jinkela_wire_207;
    wire jinkela_wire_208;
    wire jinkela_wire_209;
    wire jinkela_wire_210;
    wire jinkela_wire_211;
    wire jinkela_wire_212;
    wire jinkela_wire_213;
    wire jinkela_wire_214;
    wire jinkela_wire_215;
    wire jinkela_wire_216;
    wire jinkela_wire_217;
    wire jinkela_wire_218;
    wire jinkela_wire_219;
    wire jinkela_wire_220;
    wire jinkela_wire_221;
    wire jinkela_wire_222;
    wire jinkela_wire_223;
    wire jinkela_wire_224;
    wire jinkela_wire_225;
    wire jinkela_wire_226;
    wire jinkela_wire_227;
    wire jinkela_wire_228;
    wire jinkela_wire_229;
    wire jinkela_wire_230;
    wire jinkela_wire_231;
    wire jinkela_wire_232;
    wire jinkela_wire_233;
    wire jinkela_wire_234;
    wire jinkela_wire_235;
    wire jinkela_wire_236;
    wire jinkela_wire_237;
    wire jinkela_wire_238;
    wire jinkela_wire_239;
    wire jinkela_wire_240;
    wire jinkela_wire_241;
    wire jinkela_wire_242;
    wire jinkela_wire_243;
    wire jinkela_wire_244;
    wire jinkela_wire_245;
    wire jinkela_wire_246;
    wire jinkela_wire_247;
    wire jinkela_wire_248;
    wire jinkela_wire_249;
    wire jinkela_wire_250;
    wire jinkela_wire_251;
    wire jinkela_wire_252;
    wire jinkela_wire_253;
    wire jinkela_wire_254;
    wire jinkela_wire_255;
    wire jinkela_wire_256;
    wire jinkela_wire_257;
    wire jinkela_wire_258;
    wire jinkela_wire_259;
    wire jinkela_wire_260;
    wire jinkela_wire_261;
    wire jinkela_wire_262;
    wire jinkela_wire_263;
    wire jinkela_wire_264;
    wire jinkela_wire_265;
    wire jinkela_wire_266;
    wire jinkela_wire_267;
    wire jinkela_wire_268;
    wire jinkela_wire_269;
    wire jinkela_wire_270;
    wire jinkela_wire_271;
    wire jinkela_wire_272;
    wire jinkela_wire_273;
    wire jinkela_wire_274;
    wire jinkela_wire_275;
    wire jinkela_wire_276;
    wire jinkela_wire_277;
    wire jinkela_wire_278;
    wire jinkela_wire_279;
    wire jinkela_wire_280;
    wire jinkela_wire_281;
    wire jinkela_wire_282;
    wire jinkela_wire_283;
    wire jinkela_wire_284;
    wire jinkela_wire_285;
    wire jinkela_wire_286;
    wire jinkela_wire_287;
    wire jinkela_wire_288;
    wire jinkela_wire_289;
    wire jinkela_wire_290;
    wire jinkela_wire_291;
    wire jinkela_wire_292;
    wire jinkela_wire_293;
    wire jinkela_wire_294;
    wire jinkela_wire_295;
    wire jinkela_wire_296;
    wire jinkela_wire_297;
    wire jinkela_wire_298;
    wire jinkela_wire_299;
    wire jinkela_wire_300;
    wire jinkela_wire_301;
    wire jinkela_wire_302;
    wire jinkela_wire_303;
    wire jinkela_wire_304;
    wire jinkela_wire_305;
    wire jinkela_wire_306;
    wire jinkela_wire_307;
    wire jinkela_wire_308;
    wire jinkela_wire_309;
    wire jinkela_wire_310;
    wire jinkela_wire_311;
    wire jinkela_wire_312;
    wire jinkela_wire_313;
    wire jinkela_wire_314;
    wire jinkela_wire_315;
    wire jinkela_wire_316;
    wire jinkela_wire_317;
    wire jinkela_wire_318;
    wire jinkela_wire_319;
    wire jinkela_wire_320;
    wire jinkela_wire_321;
    wire jinkela_wire_322;
    wire jinkela_wire_323;
    wire jinkela_wire_324;
    wire jinkela_wire_325;
    wire jinkela_wire_326;
    wire jinkela_wire_327;
    wire jinkela_wire_328;
    wire jinkela_wire_329;
    wire jinkela_wire_330;
    wire jinkela_wire_331;
    wire jinkela_wire_332;
    wire jinkela_wire_333;
    wire jinkela_wire_334;
    wire jinkela_wire_335;
    wire jinkela_wire_336;
    wire jinkela_wire_337;
    wire jinkela_wire_338;
    wire jinkela_wire_339;
    wire jinkela_wire_340;
    wire jinkela_wire_341;
    wire jinkela_wire_342;
    wire jinkela_wire_343;
    wire jinkela_wire_344;
    wire jinkela_wire_345;
    wire jinkela_wire_346;
    wire jinkela_wire_347;
    wire jinkela_wire_348;
    wire jinkela_wire_349;
    wire jinkela_wire_350;
    wire jinkela_wire_351;
    wire jinkela_wire_352;
    wire jinkela_wire_353;
    wire jinkela_wire_354;
    wire jinkela_wire_355;
    wire jinkela_wire_356;
    wire jinkela_wire_357;
    wire jinkela_wire_358;
    wire jinkela_wire_359;
    wire jinkela_wire_360;
    wire jinkela_wire_361;
    wire jinkela_wire_362;
    wire jinkela_wire_363;
    wire jinkela_wire_364;
    wire jinkela_wire_365;
    wire jinkela_wire_366;
    wire jinkela_wire_367;
    wire jinkela_wire_368;
    wire jinkela_wire_369;
    wire jinkela_wire_370;
    wire jinkela_wire_371;
    wire jinkela_wire_372;
    wire jinkela_wire_373;
    wire jinkela_wire_374;
    wire jinkela_wire_375;
    wire jinkela_wire_376;
    wire jinkela_wire_377;
    wire jinkela_wire_378;
    wire jinkela_wire_379;
    wire jinkela_wire_380;
    wire jinkela_wire_381;
    wire jinkela_wire_382;
    wire jinkela_wire_383;
    wire jinkela_wire_384;
    wire jinkela_wire_385;
    wire jinkela_wire_386;
    wire jinkela_wire_387;
    wire jinkela_wire_388;
    wire jinkela_wire_389;
    wire jinkela_wire_390;
    wire jinkela_wire_391;
    wire jinkela_wire_392;
    wire jinkela_wire_393;
    wire jinkela_wire_394;
    wire jinkela_wire_395;
    wire jinkela_wire_396;
    wire jinkela_wire_397;
    wire jinkela_wire_398;
    wire jinkela_wire_399;
    wire jinkela_wire_400;
    wire jinkela_wire_401;
    wire jinkela_wire_402;
    wire jinkela_wire_403;
    wire jinkela_wire_404;
    wire jinkela_wire_405;
    wire jinkela_wire_406;
    wire jinkela_wire_407;
    wire jinkela_wire_408;
    wire jinkela_wire_409;
    wire jinkela_wire_410;
    wire jinkela_wire_411;
    wire jinkela_wire_412;
    wire jinkela_wire_413;
    wire jinkela_wire_414;
    wire jinkela_wire_415;
    wire jinkela_wire_416;
    wire jinkela_wire_417;
    wire jinkela_wire_418;
    wire jinkela_wire_419;
    wire jinkela_wire_420;
    wire jinkela_wire_421;
    wire jinkela_wire_422;
    wire jinkela_wire_423;
    wire jinkela_wire_424;
    wire jinkela_wire_425;
    wire jinkela_wire_426;
    wire jinkela_wire_427;
    wire jinkela_wire_428;
    wire jinkela_wire_429;
    wire jinkela_wire_430;
    wire jinkela_wire_431;
    wire jinkela_wire_432;
    wire jinkela_wire_433;
    wire jinkela_wire_434;
    wire jinkela_wire_435;
    wire jinkela_wire_436;
    wire jinkela_wire_437;
    wire jinkela_wire_438;
    wire jinkela_wire_439;
    wire jinkela_wire_440;
    wire jinkela_wire_441;
    wire jinkela_wire_442;
    wire jinkela_wire_443;
    wire jinkela_wire_444;
    wire jinkela_wire_445;
    wire jinkela_wire_446;
    wire jinkela_wire_447;
    wire jinkela_wire_448;
    wire jinkela_wire_449;
    wire jinkela_wire_450;
    wire jinkela_wire_451;
    wire jinkela_wire_452;
    wire jinkela_wire_453;
    wire jinkela_wire_454;
    wire jinkela_wire_455;
    wire jinkela_wire_456;
    wire jinkela_wire_457;
    wire jinkela_wire_458;
    wire jinkela_wire_459;
    wire jinkela_wire_460;
    wire jinkela_wire_461;
    wire jinkela_wire_462;
    wire jinkela_wire_463;
    wire jinkela_wire_464;
    wire jinkela_wire_465;
    wire jinkela_wire_466;
    wire jinkela_wire_467;
    wire jinkela_wire_468;
    wire jinkela_wire_469;
    wire jinkela_wire_470;
    wire jinkela_wire_471;
    wire jinkela_wire_472;
    wire jinkela_wire_473;
    wire jinkela_wire_474;
    wire jinkela_wire_475;
    wire jinkela_wire_476;
    wire jinkela_wire_477;
    wire jinkela_wire_478;
    wire jinkela_wire_479;
    wire jinkela_wire_480;
    wire jinkela_wire_481;
    wire jinkela_wire_482;
    wire jinkela_wire_483;
    wire jinkela_wire_484;
    wire jinkela_wire_485;
    wire jinkela_wire_486;
    wire jinkela_wire_487;
    wire jinkela_wire_488;
    wire jinkela_wire_489;
    wire jinkela_wire_490;
    wire jinkela_wire_491;
    wire jinkela_wire_492;
    wire jinkela_wire_493;
    wire jinkela_wire_494;
    wire jinkela_wire_495;
    wire jinkela_wire_496;
    wire jinkela_wire_497;
    wire jinkela_wire_498;
    wire jinkela_wire_499;
    wire jinkela_wire_500;
    wire jinkela_wire_501;
    wire jinkela_wire_502;
    wire jinkela_wire_503;
    wire jinkela_wire_504;
    wire jinkela_wire_505;
    wire jinkela_wire_506;
    wire jinkela_wire_507;
    wire jinkela_wire_508;
    wire jinkela_wire_509;
    wire jinkela_wire_510;
    wire jinkela_wire_511;
    wire jinkela_wire_512;
    wire jinkela_wire_513;
    wire jinkela_wire_514;
    wire jinkela_wire_515;
    wire jinkela_wire_516;
    wire jinkela_wire_517;
    wire jinkela_wire_518;
    wire jinkela_wire_519;
    wire jinkela_wire_520;
    wire jinkela_wire_521;
    wire jinkela_wire_522;
    wire jinkela_wire_523;
    wire jinkela_wire_524;
    wire jinkela_wire_525;
    wire jinkela_wire_526;
    wire jinkela_wire_527;
    wire jinkela_wire_528;
    wire jinkela_wire_529;
    wire jinkela_wire_530;
    wire jinkela_wire_531;
    wire jinkela_wire_532;
    wire jinkela_wire_533;
    wire jinkela_wire_534;
    wire jinkela_wire_535;
    wire jinkela_wire_536;
    wire jinkela_wire_537;
    wire jinkela_wire_538;
    wire jinkela_wire_539;
    wire jinkela_wire_540;
    wire jinkela_wire_541;
    wire jinkela_wire_542;
    wire jinkela_wire_543;
    wire jinkela_wire_544;
    wire jinkela_wire_545;
    wire jinkela_wire_546;
    wire jinkela_wire_547;
    wire jinkela_wire_548;
    wire jinkela_wire_549;
    wire jinkela_wire_550;
    wire jinkela_wire_551;
    wire jinkela_wire_552;
    wire jinkela_wire_553;
    wire jinkela_wire_554;
    wire jinkela_wire_555;
    wire jinkela_wire_556;
    wire jinkela_wire_557;
    wire jinkela_wire_558;
    wire jinkela_wire_559;
    wire jinkela_wire_560;
    wire jinkela_wire_561;
    wire jinkela_wire_562;
    wire jinkela_wire_563;
    wire jinkela_wire_564;
    wire jinkela_wire_565;
    wire jinkela_wire_566;
    wire jinkela_wire_567;
    wire jinkela_wire_568;
    wire jinkela_wire_569;
    wire jinkela_wire_570;
    wire jinkela_wire_571;
    wire jinkela_wire_572;
    wire jinkela_wire_573;
    wire jinkela_wire_574;
    wire jinkela_wire_575;
    wire jinkela_wire_576;
    wire jinkela_wire_577;
    wire jinkela_wire_578;
    wire jinkela_wire_579;
    wire jinkela_wire_580;
    wire jinkela_wire_581;
    wire jinkela_wire_582;
    wire jinkela_wire_583;
    wire jinkela_wire_584;
    wire jinkela_wire_585;
    wire jinkela_wire_586;
    wire jinkela_wire_587;
    wire jinkela_wire_588;
    wire jinkela_wire_589;
    wire jinkela_wire_590;
    wire jinkela_wire_591;
    wire jinkela_wire_592;
    wire jinkela_wire_593;
    wire jinkela_wire_594;
    wire jinkela_wire_595;
    wire jinkela_wire_596;
    wire jinkela_wire_597;
    wire jinkela_wire_598;
    wire jinkela_wire_599;
    wire jinkela_wire_600;
    wire jinkela_wire_601;
    wire jinkela_wire_602;
    wire jinkela_wire_603;
    wire jinkela_wire_604;
    wire jinkela_wire_605;
    wire jinkela_wire_606;
    wire jinkela_wire_607;
    wire jinkela_wire_608;
    wire jinkela_wire_609;
    wire jinkela_wire_610;
    wire jinkela_wire_611;
    wire jinkela_wire_612;
    wire jinkela_wire_613;
    wire jinkela_wire_614;
    wire jinkela_wire_615;
    wire jinkela_wire_616;
    wire jinkela_wire_617;
    wire jinkela_wire_618;
    wire jinkela_wire_619;
    wire jinkela_wire_620;
    wire jinkela_wire_621;
    wire jinkela_wire_622;
    wire jinkela_wire_623;
    wire jinkela_wire_624;
    wire jinkela_wire_625;
    wire jinkela_wire_626;
    wire jinkela_wire_627;
    wire jinkela_wire_628;
    wire jinkela_wire_629;
    wire jinkela_wire_630;
    wire jinkela_wire_631;
    wire jinkela_wire_632;
    wire jinkela_wire_633;
    wire jinkela_wire_634;
    wire jinkela_wire_635;
    wire jinkela_wire_636;
    wire jinkela_wire_637;
    wire jinkela_wire_638;
    wire jinkela_wire_639;
    wire jinkela_wire_640;
    wire jinkela_wire_641;
    wire jinkela_wire_642;
    wire jinkela_wire_643;
    wire jinkela_wire_644;
    wire jinkela_wire_645;
    wire jinkela_wire_646;
    wire jinkela_wire_647;
    wire jinkela_wire_648;
    wire jinkela_wire_649;
    wire jinkela_wire_650;
    wire jinkela_wire_651;
    wire jinkela_wire_652;
    wire jinkela_wire_653;
    wire jinkela_wire_654;
    wire jinkela_wire_655;
    wire jinkela_wire_656;
    wire jinkela_wire_657;
    wire jinkela_wire_658;
    wire jinkela_wire_659;
    wire jinkela_wire_660;
    wire jinkela_wire_661;
    wire jinkela_wire_662;
    wire jinkela_wire_663;
    wire jinkela_wire_664;
    wire jinkela_wire_665;
    wire jinkela_wire_666;
    wire jinkela_wire_667;
    wire jinkela_wire_668;
    wire jinkela_wire_669;
    wire jinkela_wire_670;
    wire jinkela_wire_671;
    wire jinkela_wire_672;
    wire jinkela_wire_673;
    wire jinkela_wire_674;
    wire jinkela_wire_675;
    wire jinkela_wire_676;
    wire jinkela_wire_677;
    wire jinkela_wire_678;
    wire jinkela_wire_679;
    wire jinkela_wire_680;
    wire jinkela_wire_681;
    wire jinkela_wire_682;
    wire jinkela_wire_683;
    wire jinkela_wire_684;
    wire jinkela_wire_685;
    wire jinkela_wire_686;
    wire jinkela_wire_687;
    wire jinkela_wire_688;
    wire jinkela_wire_689;
    wire jinkela_wire_690;
    wire jinkela_wire_691;
    wire jinkela_wire_692;
    wire jinkela_wire_693;
    wire jinkela_wire_694;
    wire jinkela_wire_695;
    wire jinkela_wire_696;
    wire jinkela_wire_697;
    wire jinkela_wire_698;
    wire jinkela_wire_699;
    wire jinkela_wire_700;
    wire jinkela_wire_701;
    wire jinkela_wire_702;
    wire jinkela_wire_703;
    wire jinkela_wire_704;
    wire jinkela_wire_705;
    wire jinkela_wire_706;
    wire jinkela_wire_707;
    wire jinkela_wire_708;
    wire jinkela_wire_709;
    wire jinkela_wire_710;
    wire jinkela_wire_711;
    wire jinkela_wire_712;
    wire jinkela_wire_713;
    wire jinkela_wire_714;
    wire jinkela_wire_715;
    wire jinkela_wire_716;
    wire jinkela_wire_717;
    wire jinkela_wire_718;
    wire jinkela_wire_719;
    wire jinkela_wire_720;
    wire jinkela_wire_721;
    wire jinkela_wire_722;
    wire jinkela_wire_723;
    wire jinkela_wire_724;
    wire jinkela_wire_725;
    wire jinkela_wire_726;
    wire jinkela_wire_727;
    wire jinkela_wire_728;
    wire jinkela_wire_729;
    wire jinkela_wire_730;
    wire jinkela_wire_731;
    wire jinkela_wire_732;
    wire jinkela_wire_733;
    wire jinkela_wire_734;
    wire jinkela_wire_735;
    wire jinkela_wire_736;
    wire jinkela_wire_737;
    wire jinkela_wire_738;
    wire jinkela_wire_739;
    wire jinkela_wire_740;
    wire jinkela_wire_741;
    wire jinkela_wire_742;
    wire jinkela_wire_743;
    wire jinkela_wire_744;
    wire jinkela_wire_745;
    wire jinkela_wire_746;
    wire jinkela_wire_747;
    wire jinkela_wire_748;
    wire jinkela_wire_749;
    wire jinkela_wire_750;
    wire jinkela_wire_751;
    wire jinkela_wire_752;
    wire jinkela_wire_753;
    wire jinkela_wire_754;
    wire jinkela_wire_755;
    wire jinkela_wire_756;
    wire jinkela_wire_757;
    wire jinkela_wire_758;
    wire jinkela_wire_759;
    wire jinkela_wire_760;
    wire jinkela_wire_761;
    wire jinkela_wire_762;
    wire jinkela_wire_763;
    wire jinkela_wire_764;
    wire jinkela_wire_765;
    wire jinkela_wire_766;
    wire jinkela_wire_767;
    wire jinkela_wire_768;
    wire jinkela_wire_769;
    wire jinkela_wire_770;
    wire jinkela_wire_771;
    wire jinkela_wire_772;
    wire jinkela_wire_773;
    wire jinkela_wire_774;
    wire jinkela_wire_775;
    wire jinkela_wire_776;
    wire jinkela_wire_777;
    wire jinkela_wire_778;
    wire jinkela_wire_779;
    wire jinkela_wire_780;
    wire jinkela_wire_781;
    wire jinkela_wire_782;
    wire jinkela_wire_783;
    wire jinkela_wire_784;
    wire jinkela_wire_785;
    wire jinkela_wire_786;
    wire jinkela_wire_787;
    wire jinkela_wire_788;
    wire jinkela_wire_789;
    wire jinkela_wire_790;
    wire jinkela_wire_791;
    wire jinkela_wire_792;
    wire jinkela_wire_793;
    wire jinkela_wire_794;
    wire jinkela_wire_795;
    wire jinkela_wire_796;
    wire jinkela_wire_797;
    wire jinkela_wire_798;
    wire jinkela_wire_799;
    wire jinkela_wire_800;
    wire jinkela_wire_801;
    wire jinkela_wire_802;
    wire jinkela_wire_803;
    wire jinkela_wire_804;
    wire jinkela_wire_805;
    wire jinkela_wire_806;
    wire jinkela_wire_807;
    wire jinkela_wire_808;
    wire jinkela_wire_809;
    wire jinkela_wire_810;
    wire jinkela_wire_811;
    wire jinkela_wire_812;
    wire jinkela_wire_813;
    wire jinkela_wire_814;
    wire jinkela_wire_815;
    wire jinkela_wire_816;
    wire jinkela_wire_817;
    wire jinkela_wire_818;
    wire jinkela_wire_819;
    wire jinkela_wire_820;
    wire jinkela_wire_821;
    wire jinkela_wire_822;
    wire jinkela_wire_823;
    wire jinkela_wire_824;
    wire jinkela_wire_825;
    wire jinkela_wire_826;
    wire jinkela_wire_827;
    wire jinkela_wire_828;
    wire jinkela_wire_829;
    wire jinkela_wire_830;
    wire jinkela_wire_831;
    input a_44_;
    input a_5_;
    input a_38_;
    input a_43_;
    input a_20_;
    input a_27_;
    input a_8_;
    input a_40_;
    input a_47_;
    input a_11_;
    input a_0_;
    input a_6_;
    input a_16_;
    input a_9_;
    input a_31_;
    input a_4_;
    input a_30_;
    input a_35_;
    input a_26_;
    input a_19_;
    input a_7_;
    input a_13_;
    input a_45_;
    input a_34_;
    input a_42_;
    input a_14_;
    input a_41_;
    input a_17_;
    input a_37_;
    input a_18_;
    input a_29_;
    input a_21_;
    input a_32_;
    input a_22_;
    input a_36_;
    input a_3_;
    input a_28_;
    input a_46_;
    input a_25_;
    input a_10_;
    input a_12_;
    input a_33_;
    input a_24_;
    input a_1_;
    input a_15_;
    input a_2_;
    input a_39_;
    input a_23_;
    output b_47_;
    output b_43_;
    output b_40_;
    output b_11_;
    output b_7_;
    output b_5_;
    output b_32_;
    output b_17_;
    output b_29_;
    output b_25_;
    output b_12_;
    output b_16_;
    output b_1_;
    output b_42_;
    output b_0_;
    output b_28_;
    output b_9_;
    output b_36_;
    output b_2_;
    output b_20_;
    output b_41_;
    output b_33_;
    output b_31_;
    output b_34_;
    output b_13_;
    output b_21_;
    output b_35_;
    output b_39_;
    output b_27_;
    output b_46_;
    output b_4_;
    output b_14_;
    output b_37_;
    output b_22_;
    output b_6_;
    output b_38_;
    output b_18_;
    output b_15_;
    output b_30_;
    output b_8_;
    output b_26_;
    output b_24_;
    output b_19_;
    output b_23_;
    output b_10_;
    output b_3_;
    output b_45_;
    output b_44_;

    or_bb _0631_ (
        .b(jinkela_wire_410),
        .a(jinkela_wire_57),
        .c(jinkela_wire_563)
    );

    maj_bbb _0632_ (
        .c(jinkela_wire_356),
        .b(jinkela_wire_816),
        .a(jinkela_wire_410),
        .d(jinkela_wire_663)
    );

    and_bb _0633_ (
        .b(jinkela_wire_356),
        .a(jinkela_wire_816),
        .c(jinkela_wire_142)
    );

    and_bb _0634_ (
        .b(jinkela_wire_410),
        .a(jinkela_wire_142),
        .c(jinkela_wire_723)
    );

    or_bb _0635_ (
        .b(jinkela_wire_649),
        .a(jinkela_wire_542),
        .c(jinkela_wire_200)
    );

    or_bb _0636_ (
        .b(jinkela_wire_76),
        .a(jinkela_wire_200),
        .c(jinkela_wire_419)
    );

    maj_bbb _0637_ (
        .c(jinkela_wire_649),
        .b(jinkela_wire_542),
        .a(jinkela_wire_76),
        .d(jinkela_wire_334)
    );

    and_bb _0638_ (
        .b(jinkela_wire_649),
        .a(jinkela_wire_542),
        .c(jinkela_wire_22)
    );

    and_bb _0639_ (
        .b(jinkela_wire_76),
        .a(jinkela_wire_22),
        .c(jinkela_wire_381)
    );

    or_bb _0640_ (
        .b(jinkela_wire_817),
        .a(jinkela_wire_239),
        .c(jinkela_wire_425)
    );

    and_bb _0641_ (
        .b(jinkela_wire_817),
        .a(jinkela_wire_239),
        .c(jinkela_wire_794)
    );

    or_bb _0642_ (
        .b(jinkela_wire_226),
        .a(jinkela_wire_829),
        .c(jinkela_wire_583)
    );

    and_bb _0643_ (
        .b(jinkela_wire_226),
        .a(jinkela_wire_829),
        .c(jinkela_wire_557)
    );

    or_bb _0644_ (
        .b(jinkela_wire_70),
        .a(jinkela_wire_543),
        .c(jinkela_wire_367)
    );

    and_bb _0645_ (
        .b(jinkela_wire_70),
        .a(jinkela_wire_543),
        .c(jinkela_wire_83)
    );

    or_bb _0646_ (
        .b(jinkela_wire_425),
        .a(jinkela_wire_583),
        .c(jinkela_wire_647)
    );

    or_bb _0647_ (
        .b(jinkela_wire_367),
        .a(jinkela_wire_647),
        .c(jinkela_wire_429)
    );

    maj_bbb _0648_ (
        .c(jinkela_wire_425),
        .b(jinkela_wire_583),
        .a(jinkela_wire_367),
        .d(jinkela_wire_819)
    );

    and_bb _0649_ (
        .b(jinkela_wire_425),
        .a(jinkela_wire_583),
        .c(jinkela_wire_360)
    );

    and_bb _0650_ (
        .b(jinkela_wire_367),
        .a(jinkela_wire_360),
        .c(jinkela_wire_290)
    );

    or_bb _0651_ (
        .b(jinkela_wire_794),
        .a(jinkela_wire_557),
        .c(jinkela_wire_62)
    );

    or_bb _0652_ (
        .b(jinkela_wire_83),
        .a(jinkela_wire_62),
        .c(jinkela_wire_291)
    );

    maj_bbb _0653_ (
        .c(jinkela_wire_794),
        .b(jinkela_wire_557),
        .a(jinkela_wire_83),
        .d(jinkela_wire_638)
    );

    and_bb _0654_ (
        .b(jinkela_wire_794),
        .a(jinkela_wire_557),
        .c(jinkela_wire_336)
    );

    and_bb _0655_ (
        .b(jinkela_wire_83),
        .a(jinkela_wire_336),
        .c(jinkela_wire_330)
    );

    or_bb _0656_ (
        .b(jinkela_wire_691),
        .a(jinkela_wire_819),
        .c(jinkela_wire_377)
    );

    and_bb _0657_ (
        .b(jinkela_wire_691),
        .a(jinkela_wire_819),
        .c(jinkela_wire_637)
    );

    or_bb _0658_ (
        .b(jinkela_wire_711),
        .a(jinkela_wire_290),
        .c(jinkela_wire_323)
    );

    and_bb _0659_ (
        .b(jinkela_wire_711),
        .a(jinkela_wire_290),
        .c(jinkela_wire_814)
    );

    or_bb _0660_ (
        .b(jinkela_wire_580),
        .a(jinkela_wire_291),
        .c(jinkela_wire_703)
    );

    and_bb _0661_ (
        .b(jinkela_wire_580),
        .a(jinkela_wire_291),
        .c(jinkela_wire_221)
    );

    or_bb _0662_ (
        .b(jinkela_wire_156),
        .a(jinkela_wire_638),
        .c(jinkela_wire_240)
    );

    and_bb _0663_ (
        .b(jinkela_wire_156),
        .a(jinkela_wire_638),
        .c(jinkela_wire_500)
    );

    or_bb _0664_ (
        .b(jinkela_wire_401),
        .a(jinkela_wire_330),
        .c(jinkela_wire_781)
    );

    and_bb _0665_ (
        .b(jinkela_wire_401),
        .a(jinkela_wire_330),
        .c(jinkela_wire_112)
    );

    or_bb _0666_ (
        .b(jinkela_wire_459),
        .a(jinkela_wire_563),
        .c(jinkela_wire_287)
    );

    and_bb _0667_ (
        .b(jinkela_wire_459),
        .a(jinkela_wire_563),
        .c(jinkela_wire_434)
    );

    or_bb _0668_ (
        .b(jinkela_wire_395),
        .a(jinkela_wire_663),
        .c(jinkela_wire_90)
    );

    and_bb _0669_ (
        .b(jinkela_wire_395),
        .a(jinkela_wire_663),
        .c(jinkela_wire_585)
    );

    or_bb _0670_ (
        .b(jinkela_wire_92),
        .a(jinkela_wire_723),
        .c(jinkela_wire_759)
    );

    and_bb _0671_ (
        .b(jinkela_wire_92),
        .a(jinkela_wire_723),
        .c(jinkela_wire_78)
    );

    or_bb _0672_ (
        .b(jinkela_wire_278),
        .a(jinkela_wire_419),
        .c(jinkela_wire_549)
    );

    or_bb _0208_ (
        .b(jinkela_wire_466),
        .a(jinkela_wire_241),
        .c(jinkela_wire_173)
    );

    or_bb _0715_ (
        .b(jinkela_wire_734),
        .a(jinkela_wire_138),
        .c(jinkela_wire_575)
    );

    maj_bbb _0925_ (
        .c(jinkela_wire_246),
        .b(jinkela_wire_123),
        .a(jinkela_wire_565),
        .d(b_19_)
    );

    maj_bbb _0209_ (
        .c(jinkela_wire_212),
        .b(jinkela_wire_146),
        .a(jinkela_wire_466),
        .d(jinkela_wire_207)
    );

    maj_bbb _0716_ (
        .c(jinkela_wire_63),
        .b(jinkela_wire_704),
        .a(jinkela_wire_734),
        .d(jinkela_wire_642)
    );

    and_bb _0926_ (
        .b(jinkela_wire_246),
        .a(jinkela_wire_123),
        .c(jinkela_wire_665)
    );

    and_bb _0210_ (
        .b(jinkela_wire_212),
        .a(jinkela_wire_146),
        .c(jinkela_wire_99)
    );

    and_bb _0717_ (
        .b(jinkela_wire_63),
        .a(jinkela_wire_704),
        .c(jinkela_wire_779)
    );

    and_bb _0927_ (
        .b(jinkela_wire_565),
        .a(jinkela_wire_665),
        .c(b_18_)
    );

    and_bb _0211_ (
        .b(jinkela_wire_466),
        .a(jinkela_wire_99),
        .c(jinkela_wire_117)
    );

    and_bb _0718_ (
        .b(jinkela_wire_734),
        .a(jinkela_wire_779),
        .c(jinkela_wire_113)
    );

    or_bb _0928_ (
        .b(jinkela_wire_431),
        .a(jinkela_wire_368),
        .c(jinkela_wire_338)
    );

    or_bb _0212_ (
        .b(jinkela_wire_18),
        .a(jinkela_wire_570),
        .c(jinkela_wire_536)
    );

    or_bb _0719_ (
        .b(jinkela_wire_599),
        .a(jinkela_wire_351),
        .c(jinkela_wire_311)
    );

    and_bb _0929_ (
        .b(jinkela_wire_431),
        .a(jinkela_wire_368),
        .c(jinkela_wire_825)
    );

    and_bb _0213_ (
        .b(jinkela_wire_18),
        .a(jinkela_wire_570),
        .c(jinkela_wire_608)
    );

    or_bb _0720_ (
        .b(jinkela_wire_47),
        .a(jinkela_wire_311),
        .c(jinkela_wire_307)
    );

    or_bb _0930_ (
        .b(jinkela_wire_380),
        .a(jinkela_wire_295),
        .c(jinkela_wire_150)
    );

    or_bb _0214_ (
        .b(jinkela_wire_765),
        .a(jinkela_wire_327),
        .c(jinkela_wire_133)
    );

    maj_bbb _0721_ (
        .c(jinkela_wire_599),
        .b(jinkela_wire_351),
        .a(jinkela_wire_47),
        .d(jinkela_wire_732)
    );

    and_bb _0931_ (
        .b(jinkela_wire_380),
        .a(jinkela_wire_295),
        .c(jinkela_wire_172)
    );

    and_bb _0215_ (
        .b(jinkela_wire_765),
        .a(jinkela_wire_327),
        .c(jinkela_wire_483)
    );

    and_bb _0722_ (
        .b(jinkela_wire_599),
        .a(jinkela_wire_351),
        .c(jinkela_wire_506)
    );

    or_bb _0932_ (
        .b(jinkela_wire_784),
        .a(jinkela_wire_679),
        .c(jinkela_wire_668)
    );

    or_bb _0216_ (
        .b(jinkela_wire_445),
        .a(jinkela_wire_292),
        .c(jinkela_wire_91)
    );

    and_bb _0723_ (
        .b(jinkela_wire_47),
        .a(jinkela_wire_506),
        .c(jinkela_wire_514)
    );

    and_bb _0933_ (
        .b(jinkela_wire_784),
        .a(jinkela_wire_679),
        .c(jinkela_wire_680)
    );

    and_bb _0217_ (
        .b(jinkela_wire_445),
        .a(jinkela_wire_292),
        .c(jinkela_wire_693)
    );

    or_bb _0724_ (
        .b(jinkela_wire_287),
        .a(jinkela_wire_489),
        .c(jinkela_wire_498)
    );

    or_bb _0934_ (
        .b(jinkela_wire_204),
        .a(jinkela_wire_664),
        .c(jinkela_wire_443)
    );

    or_bb _0218_ (
        .b(jinkela_wire_708),
        .a(jinkela_wire_173),
        .c(jinkela_wire_329)
    );

    and_bb _0725_ (
        .b(jinkela_wire_287),
        .a(jinkela_wire_489),
        .c(jinkela_wire_454)
    );

    and_bb _0935_ (
        .b(jinkela_wire_204),
        .a(jinkela_wire_664),
        .c(jinkela_wire_403)
    );

    and_bb _0219_ (
        .b(jinkela_wire_708),
        .a(jinkela_wire_173),
        .c(jinkela_wire_176)
    );

    or_bb _0726_ (
        .b(jinkela_wire_90),
        .a(jinkela_wire_377),
        .c(jinkela_wire_48)
    );

    or_bb _0936_ (
        .b(jinkela_wire_52),
        .a(jinkela_wire_277),
        .c(jinkela_wire_120)
    );

    or_bb _0220_ (
        .b(jinkela_wire_624),
        .a(jinkela_wire_207),
        .c(jinkela_wire_251)
    );

    and_bb _0727_ (
        .b(jinkela_wire_90),
        .a(jinkela_wire_377),
        .c(jinkela_wire_331)
    );

    and_bb _0937_ (
        .b(jinkela_wire_52),
        .a(jinkela_wire_277),
        .c(jinkela_wire_526)
    );

    and_bb _0221_ (
        .b(jinkela_wire_624),
        .a(jinkela_wire_207),
        .c(jinkela_wire_619)
    );

    or_bb _0728_ (
        .b(jinkela_wire_759),
        .a(jinkela_wire_323),
        .c(jinkela_wire_522)
    );

    or_bb _0938_ (
        .b(jinkela_wire_137),
        .a(jinkela_wire_447),
        .c(jinkela_wire_300)
    );

    or_bb _0222_ (
        .b(jinkela_wire_699),
        .a(jinkela_wire_117),
        .c(jinkela_wire_27)
    );

    and_bb _0729_ (
        .b(jinkela_wire_759),
        .a(jinkela_wire_323),
        .c(jinkela_wire_738)
    );

    and_bb _0939_ (
        .b(jinkela_wire_137),
        .a(jinkela_wire_447),
        .c(jinkela_wire_108)
    );

    and_bb _0223_ (
        .b(jinkela_wire_699),
        .a(jinkela_wire_117),
        .c(jinkela_wire_94)
    );

    or_bb _0730_ (
        .b(jinkela_wire_549),
        .a(jinkela_wire_703),
        .c(jinkela_wire_705)
    );

    or_bb _0940_ (
        .b(jinkela_wire_250),
        .a(jinkela_wire_96),
        .c(jinkela_wire_276)
    );

    or_bb _0224_ (
        .b(jinkela_wire_94),
        .a(jinkela_wire_693),
        .c(jinkela_wire_768)
    );

    and_bb _0731_ (
        .b(jinkela_wire_549),
        .a(jinkela_wire_703),
        .c(jinkela_wire_310)
    );

    and_bb _0941_ (
        .b(jinkela_wire_250),
        .a(jinkela_wire_96),
        .c(jinkela_wire_795)
    );

    and_bb _0225_ (
        .b(jinkela_wire_94),
        .a(jinkela_wire_693),
        .c(jinkela_wire_216)
    );

    or_bb _0732_ (
        .b(jinkela_wire_325),
        .a(jinkela_wire_240),
        .c(jinkela_wire_66)
    );

    or_bb _0942_ (
        .b(jinkela_wire_525),
        .a(jinkela_wire_211),
        .c(jinkela_wire_160)
    );

    or_bb _0226_ (
        .b(jinkela_wire_619),
        .a(jinkela_wire_483),
        .c(jinkela_wire_26)
    );

    and_bb _0733_ (
        .b(jinkela_wire_325),
        .a(jinkela_wire_240),
        .c(jinkela_wire_630)
    );

    and_bb _0943_ (
        .b(jinkela_wire_525),
        .a(jinkela_wire_211),
        .c(jinkela_wire_265)
    );

    and_bb _0227_ (
        .b(jinkela_wire_619),
        .a(jinkela_wire_483),
        .c(jinkela_wire_363)
    );

    or_bb _0734_ (
        .b(jinkela_wire_761),
        .a(jinkela_wire_781),
        .c(jinkela_wire_464)
    );

    or_bb _0944_ (
        .b(jinkela_wire_474),
        .a(jinkela_wire_564),
        .c(jinkela_wire_214)
    );

    or_bb _0228_ (
        .b(jinkela_wire_176),
        .a(jinkela_wire_608),
        .c(jinkela_wire_726)
    );

    and_bb _0735_ (
        .b(jinkela_wire_761),
        .a(jinkela_wire_781),
        .c(jinkela_wire_587)
    );

    and_bb _0945_ (
        .b(jinkela_wire_474),
        .a(jinkela_wire_564),
        .c(jinkela_wire_428)
    );

    and_bb _0229_ (
        .b(jinkela_wire_176),
        .a(jinkela_wire_608),
        .c(jinkela_wire_423)
    );

    or_bb _0736_ (
        .b(jinkela_wire_587),
        .a(jinkela_wire_738),
        .c(jinkela_wire_771)
    );

    or_bb _0946_ (
        .b(jinkela_wire_164),
        .a(jinkela_wire_590),
        .c(jinkela_wire_597)
    );

    or_bb _0230_ (
        .b(jinkela_wire_768),
        .a(jinkela_wire_26),
        .c(jinkela_wire_326)
    );

    and_bb _0737_ (
        .b(jinkela_wire_587),
        .a(jinkela_wire_738),
        .c(jinkela_wire_191)
    );

    and_bb _0947_ (
        .b(jinkela_wire_164),
        .a(jinkela_wire_590),
        .c(jinkela_wire_554)
    );

    or_bb _0231_ (
        .b(jinkela_wire_726),
        .a(jinkela_wire_326),
        .c(jinkela_wire_584)
    );

    or_bb _0738_ (
        .b(jinkela_wire_630),
        .a(jinkela_wire_331),
        .c(jinkela_wire_724)
    );

    or_bb _0948_ (
        .b(jinkela_wire_609),
        .a(jinkela_wire_353),
        .c(jinkela_wire_252)
    );

    maj_bbb _0232_ (
        .c(jinkela_wire_768),
        .b(jinkela_wire_26),
        .a(jinkela_wire_726),
        .d(jinkela_wire_249)
    );

    and_bb _0739_ (
        .b(jinkela_wire_630),
        .a(jinkela_wire_331),
        .c(jinkela_wire_567)
    );

    and_bb _0949_ (
        .b(jinkela_wire_609),
        .a(jinkela_wire_353),
        .c(jinkela_wire_774)
    );

    and_bb _0233_ (
        .b(jinkela_wire_768),
        .a(jinkela_wire_26),
        .c(jinkela_wire_548)
    );

    or_bb _0740_ (
        .b(jinkela_wire_310),
        .a(jinkela_wire_454),
        .c(jinkela_wire_102)
    );

    or_bb _0950_ (
        .b(jinkela_wire_206),
        .a(jinkela_wire_695),
        .c(jinkela_wire_387)
    );

    and_bb _0234_ (
        .b(jinkela_wire_726),
        .a(jinkela_wire_548),
        .c(jinkela_wire_769)
    );

    and_bb _0741_ (
        .b(jinkela_wire_310),
        .a(jinkela_wire_454),
        .c(jinkela_wire_65)
    );

    and_bb _0951_ (
        .b(jinkela_wire_206),
        .a(jinkela_wire_695),
        .c(jinkela_wire_129)
    );

    or_bb _0235_ (
        .b(jinkela_wire_216),
        .a(jinkela_wire_363),
        .c(jinkela_wire_477)
    );

    or_bb _0742_ (
        .b(jinkela_wire_771),
        .a(jinkela_wire_724),
        .c(jinkela_wire_254)
    );

    or_bb _0952_ (
        .b(jinkela_wire_108),
        .a(jinkela_wire_129),
        .c(jinkela_wire_139)
    );

    or_bb _0236_ (
        .b(jinkela_wire_423),
        .a(jinkela_wire_477),
        .c(jinkela_wire_382)
    );

    or_bb _0743_ (
        .b(jinkela_wire_102),
        .a(jinkela_wire_254),
        .c(jinkela_wire_165)
    );

    and_bb _0953_ (
        .b(jinkela_wire_108),
        .a(jinkela_wire_129),
        .c(jinkela_wire_553)
    );

    maj_bbb _0237_ (
        .c(jinkela_wire_216),
        .b(jinkela_wire_363),
        .a(jinkela_wire_423),
        .d(jinkela_wire_107)
    );

    maj_bbb _0744_ (
        .c(jinkela_wire_771),
        .b(jinkela_wire_724),
        .a(jinkela_wire_102),
        .d(jinkela_wire_725)
    );

    or_bb _0954_ (
        .b(jinkela_wire_795),
        .a(jinkela_wire_825),
        .c(jinkela_wire_430)
    );

    and_bb _0238_ (
        .b(jinkela_wire_216),
        .a(jinkela_wire_363),
        .c(jinkela_wire_280)
    );

    and_bb _0745_ (
        .b(jinkela_wire_771),
        .a(jinkela_wire_724),
        .c(jinkela_wire_742)
    );

    and_bb _0955_ (
        .b(jinkela_wire_795),
        .a(jinkela_wire_825),
        .c(jinkela_wire_375)
    );

    and_bb _0239_ (
        .b(jinkela_wire_423),
        .a(jinkela_wire_280),
        .c(jinkela_wire_39)
    );

    and_bb _0746_ (
        .b(jinkela_wire_102),
        .a(jinkela_wire_742),
        .c(jinkela_wire_15)
    );

    or_bb _0956_ (
        .b(jinkela_wire_265),
        .a(jinkela_wire_172),
        .c(jinkela_wire_68)
    );

    or_bb _0240_ (
        .b(jinkela_wire_27),
        .a(jinkela_wire_91),
        .c(jinkela_wire_376)
    );

    or_bb _0747_ (
        .b(jinkela_wire_191),
        .a(jinkela_wire_567),
        .c(jinkela_wire_722)
    );

    and_bb _0957_ (
        .b(jinkela_wire_265),
        .a(jinkela_wire_172),
        .c(jinkela_wire_332)
    );

    and_bb _0241_ (
        .b(jinkela_wire_27),
        .a(jinkela_wire_91),
        .c(jinkela_wire_195)
    );

    or_bb _0748_ (
        .b(jinkela_wire_65),
        .a(jinkela_wire_722),
        .c(jinkela_wire_255)
    );

    or_bb _0958_ (
        .b(jinkela_wire_428),
        .a(jinkela_wire_680),
        .c(jinkela_wire_248)
    );

    or_bb _0242_ (
        .b(jinkela_wire_251),
        .a(jinkela_wire_133),
        .c(jinkela_wire_818)
    );

    maj_bbb _0749_ (
        .c(jinkela_wire_191),
        .b(jinkela_wire_567),
        .a(jinkela_wire_65),
        .d(jinkela_wire_710)
    );

    and_bb _0959_ (
        .b(jinkela_wire_428),
        .a(jinkela_wire_680),
        .c(jinkela_wire_217)
    );

    and_bb _0243_ (
        .b(jinkela_wire_251),
        .a(jinkela_wire_133),
        .c(jinkela_wire_515)
    );

    and_bb _0750_ (
        .b(jinkela_wire_191),
        .a(jinkela_wire_567),
        .c(jinkela_wire_313)
    );

    or_bb _0960_ (
        .b(jinkela_wire_554),
        .a(jinkela_wire_403),
        .c(jinkela_wire_23)
    );

    or_bb _0244_ (
        .b(jinkela_wire_329),
        .a(jinkela_wire_536),
        .c(jinkela_wire_222)
    );

    and_bb _0751_ (
        .b(jinkela_wire_65),
        .a(jinkela_wire_313),
        .c(jinkela_wire_651)
    );

    and_bb _0961_ (
        .b(jinkela_wire_554),
        .a(jinkela_wire_403),
        .c(jinkela_wire_625)
    );

    and_bb _0245_ (
        .b(jinkela_wire_329),
        .a(jinkela_wire_536),
        .c(jinkela_wire_757)
    );

    or_bb _0752_ (
        .b(jinkela_wire_464),
        .a(jinkela_wire_522),
        .c(jinkela_wire_256)
    );

    or_bb _0962_ (
        .b(jinkela_wire_774),
        .a(jinkela_wire_526),
        .c(jinkela_wire_116)
    );

    or_bb _0246_ (
        .b(jinkela_wire_376),
        .a(jinkela_wire_818),
        .c(jinkela_wire_754)
    );

    and_bb _0753_ (
        .b(jinkela_wire_464),
        .a(jinkela_wire_522),
        .c(jinkela_wire_24)
    );

    and_bb _0963_ (
        .b(jinkela_wire_774),
        .a(jinkela_wire_526),
        .c(jinkela_wire_149)
    );

    or_bb _0247_ (
        .b(jinkela_wire_222),
        .a(jinkela_wire_754),
        .c(jinkela_wire_468)
    );

    or_bb _0754_ (
        .b(jinkela_wire_66),
        .a(jinkela_wire_48),
        .c(jinkela_wire_537)
    );

    or_bb _0964_ (
        .b(jinkela_wire_149),
        .a(jinkela_wire_332),
        .c(jinkela_wire_535)
    );

    maj_bbb _0248_ (
        .c(jinkela_wire_376),
        .b(jinkela_wire_818),
        .a(jinkela_wire_222),
        .d(jinkela_wire_208)
    );

    and_bb _0755_ (
        .b(jinkela_wire_66),
        .a(jinkela_wire_48),
        .c(jinkela_wire_413)
    );

    and_bb _0965_ (
        .b(jinkela_wire_149),
        .a(jinkela_wire_332),
        .c(jinkela_wire_260)
    );

    and_bb _0249_ (
        .b(jinkela_wire_376),
        .a(jinkela_wire_818),
        .c(jinkela_wire_242)
    );

    or_bb _0756_ (
        .b(jinkela_wire_705),
        .a(jinkela_wire_498),
        .c(jinkela_wire_352)
    );

    or_bb _0966_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_375),
        .c(jinkela_wire_369)
    );

    or_bb _0166_ (
        .b(a_42_),
        .a(jinkela_wire_787),
        .c(jinkela_wire_263)
    );

    and_bb _0250_ (
        .b(jinkela_wire_222),
        .a(jinkela_wire_242),
        .c(jinkela_wire_547)
    );

    or_bb _0292_ (
        .b(jinkela_wire_452),
        .a(jinkela_wire_203),
        .c(jinkela_wire_778)
    );

    maj_bbb _0167_ (
        .c(a_44_),
        .b(a_43_),
        .a(a_42_),
        .d(jinkela_wire_154)
    );

    or_bb _0251_ (
        .b(jinkela_wire_195),
        .a(jinkela_wire_515),
        .c(jinkela_wire_415)
    );

    and_bb _0293_ (
        .b(jinkela_wire_452),
        .a(jinkela_wire_203),
        .c(jinkela_wire_197)
    );

    and_bb _0168_ (
        .b(a_44_),
        .a(a_43_),
        .c(jinkela_wire_79)
    );

    or_bb _0252_ (
        .b(jinkela_wire_757),
        .a(jinkela_wire_415),
        .c(jinkela_wire_50)
    );

    or_bb _0294_ (
        .b(jinkela_wire_683),
        .a(jinkela_wire_675),
        .c(jinkela_wire_682)
    );

    and_bb _0169_ (
        .b(a_42_),
        .a(jinkela_wire_79),
        .c(jinkela_wire_613)
    );

    maj_bbb _0253_ (
        .c(jinkela_wire_195),
        .b(jinkela_wire_515),
        .a(jinkela_wire_757),
        .d(jinkela_wire_821)
    );

    and_bb _0295_ (
        .b(jinkela_wire_683),
        .a(jinkela_wire_675),
        .c(jinkela_wire_366)
    );

    or_bb _0170_ (
        .b(jinkela_wire_436),
        .a(jinkela_wire_613),
        .c(jinkela_wire_807)
    );

    and_bb _0254_ (
        .b(jinkela_wire_195),
        .a(jinkela_wire_515),
        .c(jinkela_wire_460)
    );

    or_bb _0296_ (
        .b(jinkela_wire_576),
        .a(jinkela_wire_418),
        .c(jinkela_wire_550)
    );

    and_bb _0171_ (
        .b(jinkela_wire_436),
        .a(jinkela_wire_613),
        .c(jinkela_wire_261)
    );

    and_bb _0255_ (
        .b(jinkela_wire_757),
        .a(jinkela_wire_460),
        .c(jinkela_wire_394)
    );

    and_bb _0297_ (
        .b(jinkela_wire_576),
        .a(jinkela_wire_418),
        .c(jinkela_wire_741)
    );

    or_bb _0172_ (
        .b(jinkela_wire_293),
        .a(jinkela_wire_154),
        .c(jinkela_wire_645)
    );

    or_bb _0256_ (
        .b(a_35_),
        .a(a_34_),
        .c(jinkela_wire_361)
    );

    or_bb _0298_ (
        .b(jinkela_wire_778),
        .a(jinkela_wire_682),
        .c(jinkela_wire_469)
    );

    and_bb _0173_ (
        .b(jinkela_wire_293),
        .a(jinkela_wire_154),
        .c(jinkela_wire_672)
    );

    or_bb _0257_ (
        .b(a_33_),
        .a(jinkela_wire_361),
        .c(jinkela_wire_114)
    );

    or_bb _0299_ (
        .b(jinkela_wire_550),
        .a(jinkela_wire_469),
        .c(jinkela_wire_7)
    );

    or_bb _0174_ (
        .b(jinkela_wire_616),
        .a(jinkela_wire_263),
        .c(jinkela_wire_450)
    );

    maj_bbb _0258_ (
        .c(a_35_),
        .b(a_34_),
        .a(a_33_),
        .d(jinkela_wire_45)
    );

    maj_bbb _0300_ (
        .c(jinkela_wire_778),
        .b(jinkela_wire_682),
        .a(jinkela_wire_550),
        .d(jinkela_wire_688)
    );

    or_bb _0312_ (
        .b(jinkela_wire_471),
        .a(jinkela_wire_541),
        .c(jinkela_wire_601)
    );

    and_bb _0175_ (
        .b(jinkela_wire_616),
        .a(jinkela_wire_263),
        .c(jinkela_wire_698)
    );

    and_bb _0259_ (
        .b(a_35_),
        .a(a_34_),
        .c(jinkela_wire_100)
    );

    and_bb _0301_ (
        .b(jinkela_wire_778),
        .a(jinkela_wire_682),
        .c(jinkela_wire_588)
    );

    or_bb _0176_ (
        .b(jinkela_wire_807),
        .a(jinkela_wire_645),
        .c(jinkela_wire_720)
    );

    and_bb _0260_ (
        .b(a_33_),
        .a(jinkela_wire_100),
        .c(jinkela_wire_41)
    );

    and_bb _0302_ (
        .b(jinkela_wire_550),
        .a(jinkela_wire_588),
        .c(jinkela_wire_541)
    );

    and_bb _0313_ (
        .b(jinkela_wire_471),
        .a(jinkela_wire_541),
        .c(jinkela_wire_81)
    );

    or_bb _0177_ (
        .b(jinkela_wire_450),
        .a(jinkela_wire_720),
        .c(jinkela_wire_699)
    );

    or_bb _0261_ (
        .b(a_32_),
        .a(a_31_),
        .c(jinkela_wire_220)
    );

    or_bb _0303_ (
        .b(jinkela_wire_197),
        .a(jinkela_wire_366),
        .c(jinkela_wire_125)
    );

    and_bb _0311_ (
        .b(jinkela_wire_626),
        .a(jinkela_wire_688),
        .c(jinkela_wire_215)
    );

    maj_bbb _0178_ (
        .c(jinkela_wire_807),
        .b(jinkela_wire_645),
        .a(jinkela_wire_450),
        .d(jinkela_wire_624)
    );

    or_bb _0262_ (
        .b(a_30_),
        .a(jinkela_wire_220),
        .c(jinkela_wire_11)
    );

    or_bb _0304_ (
        .b(jinkela_wire_741),
        .a(jinkela_wire_125),
        .c(jinkela_wire_648)
    );

    and_bb _0179_ (
        .b(jinkela_wire_807),
        .a(jinkela_wire_645),
        .c(jinkela_wire_294)
    );

    maj_bbb _0263_ (
        .c(a_32_),
        .b(a_31_),
        .a(a_30_),
        .d(jinkela_wire_632)
    );

    maj_bbb _0305_ (
        .c(jinkela_wire_197),
        .b(jinkela_wire_366),
        .a(jinkela_wire_741),
        .d(jinkela_wire_730)
    );

    and_bb _0180_ (
        .b(jinkela_wire_450),
        .a(jinkela_wire_294),
        .c(jinkela_wire_708)
    );

    and_bb _0264_ (
        .b(a_32_),
        .a(a_31_),
        .c(jinkela_wire_247)
    );

    and_bb _0306_ (
        .b(jinkela_wire_197),
        .a(jinkela_wire_366),
        .c(jinkela_wire_101)
    );

    or_bb _0181_ (
        .b(jinkela_wire_261),
        .a(jinkela_wire_672),
        .c(jinkela_wire_772)
    );

    and_bb _0265_ (
        .b(a_30_),
        .a(jinkela_wire_247),
        .c(jinkela_wire_43)
    );

    and_bb _0307_ (
        .b(jinkela_wire_741),
        .a(jinkela_wire_101),
        .c(jinkela_wire_752)
    );

    or_bb _0182_ (
        .b(jinkela_wire_698),
        .a(jinkela_wire_772),
        .c(jinkela_wire_445)
    );

    or_bb _0266_ (
        .b(jinkela_wire_114),
        .a(jinkela_wire_43),
        .c(jinkela_wire_731)
    );

    or_bb _0308_ (
        .b(jinkela_wire_457),
        .a(jinkela_wire_7),
        .c(jinkela_wire_364)
    );

    maj_bbb _0183_ (
        .c(jinkela_wire_261),
        .b(jinkela_wire_672),
        .a(jinkela_wire_698),
        .d(jinkela_wire_765)
    );

    and_bb _0267_ (
        .b(jinkela_wire_114),
        .a(jinkela_wire_43),
        .c(jinkela_wire_14)
    );

    and_bb _0309_ (
        .b(jinkela_wire_457),
        .a(jinkela_wire_7),
        .c(jinkela_wire_422)
    );

    and_bb _0184_ (
        .b(jinkela_wire_261),
        .a(jinkela_wire_672),
        .c(jinkela_wire_1)
    );

    or_bb _0268_ (
        .b(jinkela_wire_45),
        .a(jinkela_wire_632),
        .c(jinkela_wire_718)
    );

    or_bb _0310_ (
        .b(jinkela_wire_626),
        .a(jinkela_wire_688),
        .c(jinkela_wire_491)
    );

    and_bb _0185_ (
        .b(jinkela_wire_698),
        .a(jinkela_wire_1),
        .c(jinkela_wire_18)
    );

    and_bb _0269_ (
        .b(jinkela_wire_45),
        .a(jinkela_wire_632),
        .c(jinkela_wire_350)
    );

    or_bb _0314_ (
        .b(jinkela_wire_692),
        .a(jinkela_wire_648),
        .c(jinkela_wire_13)
    );

    or_bb _0186_ (
        .b(a_41_),
        .a(a_40_),
        .c(jinkela_wire_767)
    );

    or_bb _0270_ (
        .b(jinkela_wire_41),
        .a(jinkela_wire_11),
        .c(jinkela_wire_21)
    );

    and_bb _0315_ (
        .b(jinkela_wire_692),
        .a(jinkela_wire_648),
        .c(jinkela_wire_780)
    );

    or_bb _0187_ (
        .b(a_39_),
        .a(jinkela_wire_767),
        .c(jinkela_wire_777)
    );

    and_bb _0271_ (
        .b(jinkela_wire_41),
        .a(jinkela_wire_11),
        .c(jinkela_wire_272)
    );

    or_bb _0316_ (
        .b(jinkela_wire_797),
        .a(jinkela_wire_730),
        .c(jinkela_wire_275)
    );

    maj_bbb _1021_ (
        .c(jinkela_wire_620),
        .b(jinkela_wire_530),
        .a(jinkela_wire_73),
        .d(b_37_)
    );

    maj_bbb _0188_ (
        .c(a_41_),
        .b(a_40_),
        .a(a_39_),
        .d(jinkela_wire_507)
    );

    or_bb _0272_ (
        .b(jinkela_wire_731),
        .a(jinkela_wire_718),
        .c(jinkela_wire_155)
    );

    and_bb _0317_ (
        .b(jinkela_wire_797),
        .a(jinkela_wire_730),
        .c(jinkela_wire_465)
    );

    and_bb _0189_ (
        .b(a_41_),
        .a(a_40_),
        .c(jinkela_wire_159)
    );

    or_bb _0273_ (
        .b(jinkela_wire_21),
        .a(jinkela_wire_155),
        .c(jinkela_wire_739)
    );

    or_bb _0318_ (
        .b(jinkela_wire_739),
        .a(jinkela_wire_752),
        .c(jinkela_wire_582)
    );

    and_bb _0190_ (
        .b(a_39_),
        .a(jinkela_wire_159),
        .c(jinkela_wire_389)
    );

    maj_bbb _0274_ (
        .c(jinkela_wire_731),
        .b(jinkela_wire_718),
        .a(jinkela_wire_21),
        .d(jinkela_wire_797)
    );

    and_bb _0319_ (
        .b(jinkela_wire_739),
        .a(jinkela_wire_752),
        .c(jinkela_wire_745)
    );

    or_bb _0191_ (
        .b(a_38_),
        .a(a_37_),
        .c(jinkela_wire_827)
    );

    and_bb _0275_ (
        .b(jinkela_wire_731),
        .a(jinkela_wire_718),
        .c(jinkela_wire_158)
    );

    or_bb _0320_ (
        .b(jinkela_wire_745),
        .a(jinkela_wire_81),
        .c(jinkela_wire_618)
    );

    or_bb _0192_ (
        .b(a_36_),
        .a(jinkela_wire_827),
        .c(jinkela_wire_56)
    );

    and_bb _0276_ (
        .b(jinkela_wire_21),
        .a(jinkela_wire_158),
        .c(jinkela_wire_692)
    );

    and_bb _0321_ (
        .b(jinkela_wire_745),
        .a(jinkela_wire_81),
        .c(jinkela_wire_88)
    );

    maj_bbb _0193_ (
        .c(a_38_),
        .b(a_37_),
        .a(a_36_),
        .d(jinkela_wire_122)
    );

    or_bb _0277_ (
        .b(jinkela_wire_14),
        .a(jinkela_wire_350),
        .c(jinkela_wire_659)
    );

    or_bb _0322_ (
        .b(jinkela_wire_465),
        .a(jinkela_wire_215),
        .c(jinkela_wire_451)
    );

    and_bb _0194_ (
        .b(a_38_),
        .a(a_37_),
        .c(jinkela_wire_432)
    );

    or_bb _0278_ (
        .b(jinkela_wire_272),
        .a(jinkela_wire_659),
        .c(jinkela_wire_471)
    );

    and_bb _0323_ (
        .b(jinkela_wire_465),
        .a(jinkela_wire_215),
        .c(jinkela_wire_286)
    );

    and_bb _0195_ (
        .b(a_36_),
        .a(jinkela_wire_432),
        .c(jinkela_wire_444)
    );

    maj_bbb _0279_ (
        .c(jinkela_wire_14),
        .b(jinkela_wire_350),
        .a(jinkela_wire_272),
        .d(jinkela_wire_626)
    );

    or_bb _0324_ (
        .b(jinkela_wire_780),
        .a(jinkela_wire_422),
        .c(jinkela_wire_385)
    );

    or_bb _0196_ (
        .b(jinkela_wire_777),
        .a(jinkela_wire_444),
        .c(jinkela_wire_341)
    );

    and_bb _0280_ (
        .b(jinkela_wire_14),
        .a(jinkela_wire_350),
        .c(jinkela_wire_747)
    );

    and_bb _0325_ (
        .b(jinkela_wire_780),
        .a(jinkela_wire_422),
        .c(jinkela_wire_764)
    );

    and_bb _0197_ (
        .b(jinkela_wire_777),
        .a(jinkela_wire_444),
        .c(jinkela_wire_212)
    );

    and_bb _0281_ (
        .b(jinkela_wire_272),
        .a(jinkela_wire_747),
        .c(jinkela_wire_457)
    );

    or_bb _0326_ (
        .b(jinkela_wire_618),
        .a(jinkela_wire_451),
        .c(jinkela_wire_37)
    );

    or_bb _0198_ (
        .b(jinkela_wire_507),
        .a(jinkela_wire_122),
        .c(jinkela_wire_521)
    );

    or_bb _0282_ (
        .b(a_29_),
        .a(a_28_),
        .c(jinkela_wire_233)
    );

    or_bb _0327_ (
        .b(jinkela_wire_385),
        .a(jinkela_wire_37),
        .c(jinkela_wire_805)
    );

    and_bb _0199_ (
        .b(jinkela_wire_507),
        .a(jinkela_wire_122),
        .c(jinkela_wire_146)
    );

    or_bb _0283_ (
        .b(a_27_),
        .a(jinkela_wire_233),
        .c(jinkela_wire_452)
    );

    maj_bbb _0328_ (
        .c(jinkela_wire_618),
        .b(jinkela_wire_451),
        .a(jinkela_wire_385),
        .d(jinkela_wire_28)
    );

    or_bb _0200_ (
        .b(jinkela_wire_389),
        .a(jinkela_wire_56),
        .c(jinkela_wire_671)
    );

    maj_bbb _0284_ (
        .c(a_29_),
        .b(a_28_),
        .a(a_27_),
        .d(jinkela_wire_683)
    );

    and_bb _0329_ (
        .b(jinkela_wire_618),
        .a(jinkela_wire_451),
        .c(jinkela_wire_560)
    );

    and_bb _0201_ (
        .b(jinkela_wire_389),
        .a(jinkela_wire_56),
        .c(jinkela_wire_466)
    );

    and_bb _0285_ (
        .b(a_29_),
        .a(a_28_),
        .c(jinkela_wire_494)
    );

    and_bb _0330_ (
        .b(jinkela_wire_385),
        .a(jinkela_wire_560),
        .c(jinkela_wire_762)
    );

    or_bb _0202_ (
        .b(jinkela_wire_341),
        .a(jinkela_wire_521),
        .c(jinkela_wire_496)
    );

    and_bb _0286_ (
        .b(a_27_),
        .a(jinkela_wire_494),
        .c(jinkela_wire_576)
    );

    or_bb _0331_ (
        .b(jinkela_wire_88),
        .a(jinkela_wire_286),
        .c(jinkela_wire_527)
    );

    or_bb _0203_ (
        .b(jinkela_wire_671),
        .a(jinkela_wire_496),
        .c(jinkela_wire_570)
    );

    or_bb _0287_ (
        .b(a_26_),
        .a(a_25_),
        .c(jinkela_wire_744)
    );

    or_bb _0332_ (
        .b(jinkela_wire_764),
        .a(jinkela_wire_527),
        .c(jinkela_wire_80)
    );

    maj_bbb _0204_ (
        .c(jinkela_wire_341),
        .b(jinkela_wire_521),
        .a(jinkela_wire_671),
        .d(jinkela_wire_327)
    );

    or_bb _0288_ (
        .b(a_24_),
        .a(jinkela_wire_744),
        .c(jinkela_wire_418)
    );

    maj_bbb _0333_ (
        .c(jinkela_wire_88),
        .b(jinkela_wire_286),
        .a(jinkela_wire_764),
        .d(jinkela_wire_820)
    );

    and_bb _0205_ (
        .b(jinkela_wire_341),
        .a(jinkela_wire_521),
        .c(jinkela_wire_449)
    );

    maj_bbb _0289_ (
        .c(a_26_),
        .b(a_25_),
        .a(a_24_),
        .d(jinkela_wire_675)
    );

    and_bb _0334_ (
        .b(jinkela_wire_88),
        .a(jinkela_wire_286),
        .c(jinkela_wire_266)
    );

    and_bb _0206_ (
        .b(jinkela_wire_671),
        .a(jinkela_wire_449),
        .c(jinkela_wire_292)
    );

    and_bb _0290_ (
        .b(a_26_),
        .a(a_25_),
        .c(jinkela_wire_355)
    );

    and_bb _0335_ (
        .b(jinkela_wire_764),
        .a(jinkela_wire_266),
        .c(jinkela_wire_441)
    );

    or_bb _0207_ (
        .b(jinkela_wire_212),
        .a(jinkela_wire_146),
        .c(jinkela_wire_241)
    );

    and_bb _0291_ (
        .b(a_24_),
        .a(jinkela_wire_355),
        .c(jinkela_wire_203)
    );

    or_bb _0336_ (
        .b(jinkela_wire_582),
        .a(jinkela_wire_601),
        .c(jinkela_wire_193)
    );

    and_bb _0337_ (
        .b(jinkela_wire_582),
        .a(jinkela_wire_601),
        .c(jinkela_wire_166)
    );

    and_bb _0757_ (
        .b(jinkela_wire_705),
        .a(jinkela_wire_498),
        .c(jinkela_wire_676)
    );

    and_bb _0799_ (
        .b(jinkela_wire_77),
        .a(jinkela_wire_307),
        .c(jinkela_wire_0)
    );

    and_bb _0967_ (
        .b(jinkela_wire_625),
        .a(jinkela_wire_375),
        .c(jinkela_wire_25)
    );

    or_bb _0338_ (
        .b(jinkela_wire_275),
        .a(jinkela_wire_491),
        .c(jinkela_wire_437)
    );

    or_bb _0758_ (
        .b(jinkela_wire_256),
        .a(jinkela_wire_537),
        .c(jinkela_wire_830)
    );

    or_bb _0800_ (
        .b(jinkela_wire_442),
        .a(jinkela_wire_732),
        .c(jinkela_wire_204)
    );

    or_bb _0968_ (
        .b(jinkela_wire_217),
        .a(jinkela_wire_553),
        .c(jinkela_wire_593)
    );

    and_bb _0339_ (
        .b(jinkela_wire_275),
        .a(jinkela_wire_491),
        .c(jinkela_wire_162)
    );

    or_bb _0759_ (
        .b(jinkela_wire_352),
        .a(jinkela_wire_830),
        .c(jinkela_wire_480)
    );

    and_bb _0801_ (
        .b(jinkela_wire_442),
        .a(jinkela_wire_732),
        .c(jinkela_wire_269)
    );

    and_bb _0969_ (
        .b(jinkela_wire_217),
        .a(jinkela_wire_553),
        .c(jinkela_wire_740)
    );

    or_bb _0340_ (
        .b(jinkela_wire_13),
        .a(jinkela_wire_364),
        .c(jinkela_wire_808)
    );

    maj_bbb _0760_ (
        .c(jinkela_wire_256),
        .b(jinkela_wire_537),
        .a(jinkela_wire_352),
        .d(jinkela_wire_533)
    );

    or_bb _0802_ (
        .b(jinkela_wire_509),
        .a(jinkela_wire_514),
        .c(jinkela_wire_52)
    );

    or_bb _0970_ (
        .b(jinkela_wire_535),
        .a(jinkela_wire_369),
        .c(jinkela_wire_511)
    );

    or_bb _1026_ (
        .b(jinkela_wire_231),
        .a(jinkela_wire_273),
        .c(jinkela_wire_237)
    );

    and_bb _0341_ (
        .b(jinkela_wire_13),
        .a(jinkela_wire_364),
        .c(jinkela_wire_677)
    );

    and_bb _0761_ (
        .b(jinkela_wire_256),
        .a(jinkela_wire_537),
        .c(jinkela_wire_391)
    );

    and_bb _0803_ (
        .b(jinkela_wire_509),
        .a(jinkela_wire_514),
        .c(jinkela_wire_472)
    );

    or_bb _0971_ (
        .b(jinkela_wire_593),
        .a(jinkela_wire_511),
        .c(b_29_)
    );

    or_bb _0342_ (
        .b(jinkela_wire_193),
        .a(jinkela_wire_437),
        .c(jinkela_wire_831)
    );

    and_bb _0762_ (
        .b(jinkela_wire_352),
        .a(jinkela_wire_391),
        .c(jinkela_wire_411)
    );

    or_bb _0804_ (
        .b(jinkela_wire_595),
        .a(jinkela_wire_2),
        .c(jinkela_wire_137)
    );

    maj_bbb _0972_ (
        .c(jinkela_wire_535),
        .b(jinkela_wire_369),
        .a(jinkela_wire_593),
        .d(b_28_)
    );

    or_bb _0343_ (
        .b(jinkela_wire_808),
        .a(jinkela_wire_831),
        .c(jinkela_wire_349)
    );

    or_bb _0763_ (
        .b(jinkela_wire_24),
        .a(jinkela_wire_413),
        .c(jinkela_wire_60)
    );

    and_bb _0805_ (
        .b(jinkela_wire_595),
        .a(jinkela_wire_2),
        .c(jinkela_wire_229)
    );

    and_bb _0973_ (
        .b(jinkela_wire_535),
        .a(jinkela_wire_369),
        .c(jinkela_wire_402)
    );

    maj_bbb _0344_ (
        .c(jinkela_wire_193),
        .b(jinkela_wire_437),
        .a(jinkela_wire_808),
        .d(jinkela_wire_170)
    );

    or_bb _0764_ (
        .b(jinkela_wire_676),
        .a(jinkela_wire_60),
        .c(jinkela_wire_333)
    );

    or_bb _0806_ (
        .b(jinkela_wire_715),
        .a(jinkela_wire_103),
        .c(jinkela_wire_250)
    );

    and_bb _0974_ (
        .b(jinkela_wire_593),
        .a(jinkela_wire_402),
        .c(b_27_)
    );

    and_bb _0345_ (
        .b(jinkela_wire_193),
        .a(jinkela_wire_437),
        .c(jinkela_wire_304)
    );

    maj_bbb _0765_ (
        .c(jinkela_wire_24),
        .b(jinkela_wire_413),
        .a(jinkela_wire_676),
        .d(jinkela_wire_315)
    );

    and_bb _0807_ (
        .b(jinkela_wire_715),
        .a(jinkela_wire_103),
        .c(jinkela_wire_610)
    );

    or_bb _0975_ (
        .b(jinkela_wire_260),
        .a(jinkela_wire_25),
        .c(jinkela_wire_187)
    );

    and_bb _0346_ (
        .b(jinkela_wire_808),
        .a(jinkela_wire_304),
        .c(jinkela_wire_728)
    );

    and_bb _0766_ (
        .b(jinkela_wire_24),
        .a(jinkela_wire_413),
        .c(jinkela_wire_735)
    );

    or_bb _0808_ (
        .b(jinkela_wire_416),
        .a(jinkela_wire_144),
        .c(jinkela_wire_525)
    );

    or_bb _0976_ (
        .b(jinkela_wire_740),
        .a(jinkela_wire_187),
        .c(b_26_)
    );

    or_bb _0347_ (
        .b(jinkela_wire_166),
        .a(jinkela_wire_162),
        .c(jinkela_wire_343)
    );

    and_bb _0767_ (
        .b(jinkela_wire_676),
        .a(jinkela_wire_735),
        .c(jinkela_wire_760)
    );

    and_bb _0809_ (
        .b(jinkela_wire_416),
        .a(jinkela_wire_144),
        .c(jinkela_wire_312)
    );

    maj_bbb _0977_ (
        .c(jinkela_wire_260),
        .b(jinkela_wire_25),
        .a(jinkela_wire_740),
        .d(b_25_)
    );

    or_bb _0348_ (
        .b(jinkela_wire_677),
        .a(jinkela_wire_343),
        .c(jinkela_wire_815)
    );

    or_bb _0768_ (
        .b(jinkela_wire_119),
        .a(jinkela_wire_480),
        .c(jinkela_wire_695)
    );

    or_bb _0810_ (
        .b(jinkela_wire_179),
        .a(jinkela_wire_362),
        .c(jinkela_wire_474)
    );

    and_bb _0978_ (
        .b(jinkela_wire_260),
        .a(jinkela_wire_25),
        .c(jinkela_wire_186)
    );

    maj_bbb _0349_ (
        .c(jinkela_wire_166),
        .b(jinkela_wire_162),
        .a(jinkela_wire_677),
        .d(jinkela_wire_479)
    );

    and_bb _0769_ (
        .b(jinkela_wire_119),
        .a(jinkela_wire_480),
        .c(jinkela_wire_678)
    );

    and_bb _0811_ (
        .b(jinkela_wire_179),
        .a(jinkela_wire_362),
        .c(jinkela_wire_426)
    );

    and_bb _0979_ (
        .b(jinkela_wire_740),
        .a(jinkela_wire_186),
        .c(b_24_)
    );

    and_bb _0350_ (
        .b(jinkela_wire_166),
        .a(jinkela_wire_162),
        .c(jinkela_wire_46)
    );

    or_bb _0770_ (
        .b(jinkela_wire_285),
        .a(jinkela_wire_533),
        .c(jinkela_wire_368)
    );

    or_bb _0812_ (
        .b(jinkela_wire_298),
        .a(jinkela_wire_478),
        .c(jinkela_wire_164)
    );

    or_bb _0980_ (
        .b(jinkela_wire_116),
        .a(jinkela_wire_68),
        .c(jinkela_wire_532)
    );

    and_bb _0351_ (
        .b(jinkela_wire_677),
        .a(jinkela_wire_46),
        .c(jinkela_wire_497)
    );

    and_bb _0771_ (
        .b(jinkela_wire_285),
        .a(jinkela_wire_533),
        .c(jinkela_wire_631)
    );

    and_bb _0813_ (
        .b(jinkela_wire_298),
        .a(jinkela_wire_478),
        .c(jinkela_wire_458)
    );

    and_bb _0981_ (
        .b(jinkela_wire_116),
        .a(jinkela_wire_68),
        .c(jinkela_wire_793)
    );

    or_bb _0352_ (
        .b(jinkela_wire_107),
        .a(jinkela_wire_170),
        .c(jinkela_wire_520)
    );

    or_bb _0772_ (
        .b(jinkela_wire_461),
        .a(jinkela_wire_411),
        .c(jinkela_wire_295)
    );

    or_bb _0814_ (
        .b(jinkela_wire_199),
        .a(jinkela_wire_51),
        .c(jinkela_wire_609)
    );

    or_bb _0982_ (
        .b(jinkela_wire_23),
        .a(jinkela_wire_430),
        .c(jinkela_wire_789)
    );

    and_bb _0353_ (
        .b(jinkela_wire_107),
        .a(jinkela_wire_170),
        .c(jinkela_wire_357)
    );

    and_bb _0773_ (
        .b(jinkela_wire_461),
        .a(jinkela_wire_411),
        .c(jinkela_wire_89)
    );

    and_bb _0815_ (
        .b(jinkela_wire_199),
        .a(jinkela_wire_51),
        .c(jinkela_wire_174)
    );

    and_bb _0983_ (
        .b(jinkela_wire_23),
        .a(jinkela_wire_430),
        .c(jinkela_wire_345)
    );

    or_bb _0354_ (
        .b(jinkela_wire_382),
        .a(jinkela_wire_728),
        .c(jinkela_wire_85)
    );

    or_bb _0774_ (
        .b(jinkela_wire_596),
        .a(jinkela_wire_333),
        .c(jinkela_wire_679)
    );

    or_bb _0816_ (
        .b(jinkela_wire_335),
        .a(jinkela_wire_631),
        .c(jinkela_wire_34)
    );

    or_bb _0984_ (
        .b(jinkela_wire_248),
        .a(jinkela_wire_139),
        .c(jinkela_wire_5)
    );

    and_bb _0355_ (
        .b(jinkela_wire_382),
        .a(jinkela_wire_728),
        .c(jinkela_wire_244)
    );

    and_bb _0775_ (
        .b(jinkela_wire_596),
        .a(jinkela_wire_333),
        .c(jinkela_wire_228)
    );

    and_bb _0817_ (
        .b(jinkela_wire_335),
        .a(jinkela_wire_631),
        .c(jinkela_wire_185)
    );

    and_bb _0985_ (
        .b(jinkela_wire_248),
        .a(jinkela_wire_139),
        .c(jinkela_wire_503)
    );

    or_bb _0356_ (
        .b(jinkela_wire_769),
        .a(jinkela_wire_815),
        .c(jinkela_wire_299)
    );

    or_bb _0776_ (
        .b(jinkela_wire_510),
        .a(jinkela_wire_315),
        .c(jinkela_wire_664)
    );

    or_bb _0818_ (
        .b(jinkela_wire_669),
        .a(jinkela_wire_89),
        .c(jinkela_wire_354)
    );

    or_bb _0986_ (
        .b(jinkela_wire_532),
        .a(jinkela_wire_789),
        .c(jinkela_wire_393)
    );

    and_bb _0357_ (
        .b(jinkela_wire_769),
        .a(jinkela_wire_815),
        .c(jinkela_wire_259)
    );

    and_bb _0777_ (
        .b(jinkela_wire_510),
        .a(jinkela_wire_315),
        .c(jinkela_wire_455)
    );

    and_bb _0819_ (
        .b(jinkela_wire_669),
        .a(jinkela_wire_89),
        .c(jinkela_wire_798)
    );

    or_bb _0987_ (
        .b(jinkela_wire_5),
        .a(jinkela_wire_393),
        .c(b_35_)
    );

    or_bb _0358_ (
        .b(jinkela_wire_249),
        .a(jinkela_wire_479),
        .c(jinkela_wire_810)
    );

    or_bb _0778_ (
        .b(jinkela_wire_670),
        .a(jinkela_wire_760),
        .c(jinkela_wire_277)
    );

    or_bb _0820_ (
        .b(jinkela_wire_0),
        .a(jinkela_wire_228),
        .c(jinkela_wire_486)
    );

    maj_bbb _0988_ (
        .c(jinkela_wire_532),
        .b(jinkela_wire_789),
        .a(jinkela_wire_5),
        .d(b_34_)
    );

    and_bb _0359_ (
        .b(jinkela_wire_249),
        .a(jinkela_wire_479),
        .c(jinkela_wire_636)
    );

    and_bb _0779_ (
        .b(jinkela_wire_670),
        .a(jinkela_wire_760),
        .c(jinkela_wire_538)
    );

    and_bb _0821_ (
        .b(jinkela_wire_0),
        .a(jinkela_wire_228),
        .c(jinkela_wire_592)
    );

    and_bb _0989_ (
        .b(jinkela_wire_532),
        .a(jinkela_wire_789),
        .c(jinkela_wire_386)
    );

    or_bb _0360_ (
        .b(jinkela_wire_584),
        .a(jinkela_wire_497),
        .c(jinkela_wire_614)
    );

    or_bb _0780_ (
        .b(jinkela_wire_783),
        .a(jinkela_wire_165),
        .c(jinkela_wire_447)
    );

    or_bb _0822_ (
        .b(jinkela_wire_269),
        .a(jinkela_wire_455),
        .c(jinkela_wire_650)
    );

    and_bb _0990_ (
        .b(jinkela_wire_5),
        .a(jinkela_wire_386),
        .c(b_33_)
    );

    and_bb _0361_ (
        .b(jinkela_wire_584),
        .a(jinkela_wire_497),
        .c(jinkela_wire_36)
    );

    and_bb _0781_ (
        .b(jinkela_wire_783),
        .a(jinkela_wire_165),
        .c(jinkela_wire_667)
    );

    and_bb _0823_ (
        .b(jinkela_wire_269),
        .a(jinkela_wire_455),
        .c(jinkela_wire_316)
    );

    or_bb _0991_ (
        .b(jinkela_wire_793),
        .a(jinkela_wire_345),
        .c(jinkela_wire_143)
    );

    or_bb _0362_ (
        .b(jinkela_wire_394),
        .a(jinkela_wire_805),
        .c(jinkela_wire_337)
    );

    or_bb _0782_ (
        .b(jinkela_wire_574),
        .a(jinkela_wire_725),
        .c(jinkela_wire_96)
    );

    or_bb _0824_ (
        .b(jinkela_wire_472),
        .a(jinkela_wire_538),
        .c(jinkela_wire_685)
    );

    or_bb _0992_ (
        .b(jinkela_wire_503),
        .a(jinkela_wire_143),
        .c(b_32_)
    );

    and_bb _0363_ (
        .b(jinkela_wire_394),
        .a(jinkela_wire_805),
        .c(jinkela_wire_558)
    );

    and_bb _0783_ (
        .b(jinkela_wire_574),
        .a(jinkela_wire_725),
        .c(jinkela_wire_392)
    );

    and_bb _0825_ (
        .b(jinkela_wire_472),
        .a(jinkela_wire_538),
        .c(jinkela_wire_135)
    );

    maj_bbb _0993_ (
        .c(jinkela_wire_793),
        .b(jinkela_wire_345),
        .a(jinkela_wire_503),
        .d(b_31_)
    );

    or_bb _0364_ (
        .b(jinkela_wire_821),
        .a(jinkela_wire_28),
        .c(jinkela_wire_98)
    );

    or_bb _0784_ (
        .b(jinkela_wire_607),
        .a(jinkela_wire_15),
        .c(jinkela_wire_211)
    );

    or_bb _0826_ (
        .b(jinkela_wire_229),
        .a(jinkela_wire_667),
        .c(jinkela_wire_38)
    );

    and_bb _0994_ (
        .b(jinkela_wire_793),
        .a(jinkela_wire_345),
        .c(jinkela_wire_775)
    );

    and_bb _0365_ (
        .b(jinkela_wire_821),
        .a(jinkela_wire_28),
        .c(jinkela_wire_201)
    );

    and_bb _0785_ (
        .b(jinkela_wire_607),
        .a(jinkela_wire_15),
        .c(jinkela_wire_182)
    );

    and_bb _0827_ (
        .b(jinkela_wire_229),
        .a(jinkela_wire_667),
        .c(jinkela_wire_405)
    );

    and_bb _0995_ (
        .b(jinkela_wire_503),
        .a(jinkela_wire_775),
        .c(b_30_)
    );

    or_bb _0366_ (
        .b(jinkela_wire_50),
        .a(jinkela_wire_762),
        .c(jinkela_wire_33)
    );

    or_bb _0786_ (
        .b(jinkela_wire_435),
        .a(jinkela_wire_255),
        .c(jinkela_wire_564)
    );

    or_bb _0828_ (
        .b(jinkela_wire_610),
        .a(jinkela_wire_392),
        .c(jinkela_wire_64)
    );

    or_bb _0996_ (
        .b(jinkela_wire_300),
        .a(jinkela_wire_387),
        .c(jinkela_wire_652)
    );

    and_bb _0367_ (
        .b(jinkela_wire_50),
        .a(jinkela_wire_762),
        .c(jinkela_wire_106)
    );

    and_bb _0787_ (
        .b(jinkela_wire_435),
        .a(jinkela_wire_255),
        .c(jinkela_wire_72)
    );

    and_bb _0829_ (
        .b(jinkela_wire_610),
        .a(jinkela_wire_392),
        .c(jinkela_wire_267)
    );

    and_bb _0997_ (
        .b(jinkela_wire_300),
        .a(jinkela_wire_387),
        .c(jinkela_wire_324)
    );

    or_bb _0368_ (
        .b(jinkela_wire_547),
        .a(jinkela_wire_80),
        .c(jinkela_wire_681)
    );

    or_bb _0788_ (
        .b(jinkela_wire_439),
        .a(jinkela_wire_710),
        .c(jinkela_wire_590)
    );

    or_bb _0830_ (
        .b(jinkela_wire_312),
        .a(jinkela_wire_182),
        .c(jinkela_wire_598)
    );

    or_bb _0998_ (
        .b(jinkela_wire_276),
        .a(jinkela_wire_338),
        .c(jinkela_wire_273)
    );

    and_bb _0369_ (
        .b(jinkela_wire_547),
        .a(jinkela_wire_80),
        .c(jinkela_wire_790)
    );

    and_bb _0789_ (
        .b(jinkela_wire_439),
        .a(jinkela_wire_710),
        .c(jinkela_wire_53)
    );

    and_bb _0831_ (
        .b(jinkela_wire_312),
        .a(jinkela_wire_182),
        .c(jinkela_wire_314)
    );

    and_bb _0999_ (
        .b(jinkela_wire_276),
        .a(jinkela_wire_338),
        .c(jinkela_wire_223)
    );

    or_bb _0370_ (
        .b(jinkela_wire_208),
        .a(jinkela_wire_820),
        .c(jinkela_wire_721)
    );

    or_bb _0790_ (
        .b(jinkela_wire_238),
        .a(jinkela_wire_651),
        .c(jinkela_wire_353)
    );

    or_bb _0832_ (
        .b(jinkela_wire_426),
        .a(jinkela_wire_72),
        .c(jinkela_wire_782)
    );

    or_bb _1000_ (
        .b(jinkela_wire_160),
        .a(jinkela_wire_150),
        .c(jinkela_wire_579)
    );

    and_bb _0371_ (
        .b(jinkela_wire_208),
        .a(jinkela_wire_820),
        .c(jinkela_wire_397)
    );

    and_bb _0791_ (
        .b(jinkela_wire_238),
        .a(jinkela_wire_651),
        .c(jinkela_wire_225)
    );

    and_bb _0833_ (
        .b(jinkela_wire_426),
        .a(jinkela_wire_72),
        .c(jinkela_wire_157)
    );

    and_bb _1001_ (
        .b(jinkela_wire_160),
        .a(jinkela_wire_150),
        .c(jinkela_wire_502)
    );

    or_bb _0372_ (
        .b(jinkela_wire_468),
        .a(jinkela_wire_441),
        .c(jinkela_wire_534)
    );

    or_bb _0792_ (
        .b(jinkela_wire_82),
        .a(jinkela_wire_575),
        .c(jinkela_wire_206)
    );

    or_bb _0834_ (
        .b(jinkela_wire_458),
        .a(jinkela_wire_53),
        .c(jinkela_wire_271)
    );

    or_bb _1002_ (
        .b(jinkela_wire_214),
        .a(jinkela_wire_668),
        .c(jinkela_wire_339)
    );

    and_bb _0373_ (
        .b(jinkela_wire_468),
        .a(jinkela_wire_441),
        .c(jinkela_wire_568)
    );

    and_bb _0793_ (
        .b(jinkela_wire_82),
        .a(jinkela_wire_575),
        .c(jinkela_wire_342)
    );

    and_bb _0835_ (
        .b(jinkela_wire_458),
        .a(jinkela_wire_53),
        .c(jinkela_wire_749)
    );

    and_bb _1003_ (
        .b(jinkela_wire_214),
        .a(jinkela_wire_668),
        .c(jinkela_wire_198)
    );

    or_bb _0374_ (
        .b(jinkela_wire_39),
        .a(jinkela_wire_349),
        .c(jinkela_wire_513)
    );

    or_bb _0794_ (
        .b(jinkela_wire_205),
        .a(jinkela_wire_642),
        .c(jinkela_wire_431)
    );

    or_bb _0836_ (
        .b(jinkela_wire_174),
        .a(jinkela_wire_225),
        .c(jinkela_wire_417)
    );

    or_bb _1004_ (
        .b(jinkela_wire_597),
        .a(jinkela_wire_443),
        .c(jinkela_wire_231)
    );

    and_bb _0375_ (
        .b(jinkela_wire_39),
        .a(jinkela_wire_349),
        .c(jinkela_wire_617)
    );

    and_bb _0795_ (
        .b(jinkela_wire_205),
        .a(jinkela_wire_642),
        .c(jinkela_wire_335)
    );

    and_bb _0837_ (
        .b(jinkela_wire_174),
        .a(jinkela_wire_225),
        .c(jinkela_wire_512)
    );

    and_bb _1005_ (
        .b(jinkela_wire_597),
        .a(jinkela_wire_443),
        .c(jinkela_wire_194)
    );

    or_bb _0376_ (
        .b(jinkela_wire_558),
        .a(jinkela_wire_617),
        .c(jinkela_wire_136)
    );

    or_bb _0796_ (
        .b(jinkela_wire_727),
        .a(jinkela_wire_113),
        .c(jinkela_wire_380)
    );

    or_bb _0838_ (
        .b(jinkela_wire_342),
        .a(jinkela_wire_678),
        .c(jinkela_wire_97)
    );

    or_bb _1006_ (
        .b(jinkela_wire_252),
        .a(jinkela_wire_120),
        .c(jinkela_wire_105)
    );

    and_bb _0377_ (
        .b(jinkela_wire_558),
        .a(jinkela_wire_617),
        .c(jinkela_wire_71)
    );

    and_bb _0797_ (
        .b(jinkela_wire_727),
        .a(jinkela_wire_113),
        .c(jinkela_wire_669)
    );

    and_bb _0839_ (
        .b(jinkela_wire_342),
        .a(jinkela_wire_678),
        .c(jinkela_wire_684)
    );

    and_bb _1007_ (
        .b(jinkela_wire_252),
        .a(jinkela_wire_120),
        .c(jinkela_wire_646)
    );

    or_bb _0378_ (
        .b(jinkela_wire_201),
        .a(jinkela_wire_357),
        .c(jinkela_wire_87)
    );

    or_bb _0798_ (
        .b(jinkela_wire_77),
        .a(jinkela_wire_307),
        .c(jinkela_wire_784)
    );

    or_bb _0840_ (
        .b(jinkela_wire_405),
        .a(jinkela_wire_684),
        .c(jinkela_wire_8)
    );

    or_bb _1008_ (
        .b(jinkela_wire_646),
        .a(jinkela_wire_502),
        .c(jinkela_wire_571)
    );

    and_bb _0379_ (
        .b(jinkela_wire_201),
        .a(jinkela_wire_357),
        .c(jinkela_wire_210)
    );

    or_bb _0380_ (
        .b(jinkela_wire_106),
        .a(jinkela_wire_244),
        .c(jinkela_wire_482)
    );

    and_bb _0381_ (
        .b(jinkela_wire_106),
        .a(jinkela_wire_244),
        .c(jinkela_wire_183)
    );

    or_bb _0382_ (
        .b(jinkela_wire_790),
        .a(jinkela_wire_259),
        .c(jinkela_wire_58)
    );

    and_bb _0383_ (
        .b(jinkela_wire_790),
        .a(jinkela_wire_259),
        .c(jinkela_wire_358)
    );

    or_bb _0384_ (
        .b(jinkela_wire_397),
        .a(jinkela_wire_636),
        .c(jinkela_wire_140)
    );

    and_bb _0385_ (
        .b(jinkela_wire_397),
        .a(jinkela_wire_636),
        .c(jinkela_wire_346)
    );

    or_bb _0386_ (
        .b(jinkela_wire_568),
        .a(jinkela_wire_36),
        .c(jinkela_wire_95)
    );

    and_bb _0387_ (
        .b(jinkela_wire_568),
        .a(jinkela_wire_36),
        .c(jinkela_wire_202)
    );

    or_bb _0388_ (
        .b(jinkela_wire_202),
        .a(jinkela_wire_183),
        .c(jinkela_wire_627)
    );

    and_bb _0389_ (
        .b(jinkela_wire_202),
        .a(jinkela_wire_183),
        .c(jinkela_wire_49)
    );

    or_bb _0390_ (
        .b(jinkela_wire_346),
        .a(jinkela_wire_210),
        .c(jinkela_wire_308)
    );

    and_bb _0391_ (
        .b(jinkela_wire_346),
        .a(jinkela_wire_210),
        .c(jinkela_wire_641)
    );

    or_bb _0392_ (
        .b(jinkela_wire_358),
        .a(jinkela_wire_71),
        .c(jinkela_wire_192)
    );

    and_bb _0393_ (
        .b(jinkela_wire_358),
        .a(jinkela_wire_71),
        .c(jinkela_wire_414)
    );

    or_bb _0394_ (
        .b(jinkela_wire_627),
        .a(jinkela_wire_308),
        .c(jinkela_wire_6)
    );

    or_bb _0395_ (
        .b(jinkela_wire_192),
        .a(jinkela_wire_6),
        .c(jinkela_wire_670)
    );

    maj_bbb _0396_ (
        .c(jinkela_wire_627),
        .b(jinkela_wire_308),
        .a(jinkela_wire_192),
        .d(jinkela_wire_510)
    );

    and_bb _0397_ (
        .b(jinkela_wire_627),
        .a(jinkela_wire_308),
        .c(jinkela_wire_523)
    );

    and_bb _0398_ (
        .b(jinkela_wire_192),
        .a(jinkela_wire_523),
        .c(jinkela_wire_596)
    );

    or_bb _0399_ (
        .b(jinkela_wire_49),
        .a(jinkela_wire_641),
        .c(jinkela_wire_602)
    );

    or_bb _0400_ (
        .b(jinkela_wire_414),
        .a(jinkela_wire_602),
        .c(jinkela_wire_461)
    );

    maj_bbb _0401_ (
        .c(jinkela_wire_49),
        .b(jinkela_wire_641),
        .a(jinkela_wire_414),
        .d(jinkela_wire_285)
    );

    and_bb _0402_ (
        .b(jinkela_wire_49),
        .a(jinkela_wire_641),
        .c(jinkela_wire_218)
    );

    and_bb _0403_ (
        .b(jinkela_wire_414),
        .a(jinkela_wire_218),
        .c(jinkela_wire_119)
    );

    or_bb _0404_ (
        .b(jinkela_wire_95),
        .a(jinkela_wire_482),
        .c(jinkela_wire_127)
    );

    and_bb _0405_ (
        .b(jinkela_wire_95),
        .a(jinkela_wire_482),
        .c(jinkela_wire_751)
    );

    or_bb _0406_ (
        .b(jinkela_wire_140),
        .a(jinkela_wire_87),
        .c(jinkela_wire_303)
    );

    and_bb _0407_ (
        .b(jinkela_wire_140),
        .a(jinkela_wire_87),
        .c(jinkela_wire_566)
    );

    or_bb _0408_ (
        .b(jinkela_wire_58),
        .a(jinkela_wire_136),
        .c(jinkela_wire_378)
    );

    and_bb _0409_ (
        .b(jinkela_wire_58),
        .a(jinkela_wire_136),
        .c(jinkela_wire_268)
    );

    or_bb _0410_ (
        .b(jinkela_wire_127),
        .a(jinkela_wire_303),
        .c(jinkela_wire_687)
    );

    or_bb _0411_ (
        .b(jinkela_wire_378),
        .a(jinkela_wire_687),
        .c(jinkela_wire_238)
    );

    maj_bbb _0412_ (
        .c(jinkela_wire_127),
        .b(jinkela_wire_303),
        .a(jinkela_wire_378),
        .d(jinkela_wire_439)
    );

    and_bb _0413_ (
        .b(jinkela_wire_127),
        .a(jinkela_wire_303),
        .c(jinkela_wire_9)
    );

    or_bb _0923_ (
        .b(jinkela_wire_246),
        .a(jinkela_wire_123),
        .c(jinkela_wire_453)
    );

    and_bb _0414_ (
        .b(jinkela_wire_378),
        .a(jinkela_wire_9),
        .c(jinkela_wire_435)
    );

    or_bb _0415_ (
        .b(jinkela_wire_751),
        .a(jinkela_wire_566),
        .c(jinkela_wire_493)
    );

    or_bb _0416_ (
        .b(jinkela_wire_268),
        .a(jinkela_wire_493),
        .c(jinkela_wire_607)
    );

    maj_bbb _0417_ (
        .c(jinkela_wire_751),
        .b(jinkela_wire_566),
        .a(jinkela_wire_268),
        .d(jinkela_wire_574)
    );

    and_bb _0418_ (
        .b(jinkela_wire_751),
        .a(jinkela_wire_566),
        .c(jinkela_wire_600)
    );

    or_bb _0924_ (
        .b(jinkela_wire_565),
        .a(jinkela_wire_453),
        .c(b_20_)
    );

    and_bb _0419_ (
        .b(jinkela_wire_268),
        .a(jinkela_wire_600),
        .c(jinkela_wire_783)
    );

    or_bb _0420_ (
        .b(jinkela_wire_337),
        .a(jinkela_wire_513),
        .c(jinkela_wire_17)
    );

    and_bb _0421_ (
        .b(jinkela_wire_337),
        .a(jinkela_wire_513),
        .c(jinkela_wire_412)
    );

    and_bb _0841_ (
        .b(jinkela_wire_405),
        .a(jinkela_wire_684),
        .c(jinkela_wire_750)
    );

    or_bb _0422_ (
        .b(jinkela_wire_98),
        .a(jinkela_wire_520),
        .c(jinkela_wire_44)
    );

    or_bb _0842_ (
        .b(jinkela_wire_267),
        .a(jinkela_wire_185),
        .c(jinkela_wire_67)
    );

    and_bb _0423_ (
        .b(jinkela_wire_98),
        .a(jinkela_wire_520),
        .c(jinkela_wire_188)
    );

    and_bb _0843_ (
        .b(jinkela_wire_267),
        .a(jinkela_wire_185),
        .c(jinkela_wire_803)
    );

    or_bb _0424_ (
        .b(jinkela_wire_33),
        .a(jinkela_wire_85),
        .c(jinkela_wire_756)
    );

    or_bb _0844_ (
        .b(jinkela_wire_314),
        .a(jinkela_wire_798),
        .c(jinkela_wire_406)
    );

    and_bb _0425_ (
        .b(jinkela_wire_33),
        .a(jinkela_wire_85),
        .c(jinkela_wire_562)
    );

    and_bb _0845_ (
        .b(jinkela_wire_314),
        .a(jinkela_wire_798),
        .c(jinkela_wire_788)
    );

    or_bb _0426_ (
        .b(jinkela_wire_681),
        .a(jinkela_wire_299),
        .c(jinkela_wire_501)
    );

    or_bb _0846_ (
        .b(jinkela_wire_157),
        .a(jinkela_wire_592),
        .c(jinkela_wire_686)
    );

    and_bb _0427_ (
        .b(jinkela_wire_681),
        .a(jinkela_wire_299),
        .c(jinkela_wire_690)
    );

    and_bb _0847_ (
        .b(jinkela_wire_157),
        .a(jinkela_wire_592),
        .c(jinkela_wire_622)
    );

    or_bb _0428_ (
        .b(jinkela_wire_721),
        .a(jinkela_wire_810),
        .c(jinkela_wire_635)
    );

    or_bb _0848_ (
        .b(jinkela_wire_749),
        .a(jinkela_wire_316),
        .c(jinkela_wire_492)
    );

    and_bb _0429_ (
        .b(jinkela_wire_721),
        .a(jinkela_wire_810),
        .c(jinkela_wire_706)
    );

    and_bb _0849_ (
        .b(jinkela_wire_749),
        .a(jinkela_wire_316),
        .c(jinkela_wire_623)
    );

    or_bb _0430_ (
        .b(jinkela_wire_534),
        .a(jinkela_wire_614),
        .c(jinkela_wire_440)
    );

    or_bb _0850_ (
        .b(jinkela_wire_512),
        .a(jinkela_wire_135),
        .c(jinkela_wire_785)
    );

    and_bb _0431_ (
        .b(jinkela_wire_534),
        .a(jinkela_wire_614),
        .c(jinkela_wire_446)
    );

    and_bb _0851_ (
        .b(jinkela_wire_512),
        .a(jinkela_wire_135),
        .c(jinkela_wire_408)
    );

    or_bb _0432_ (
        .b(jinkela_wire_446),
        .a(jinkela_wire_562),
        .c(jinkela_wire_578)
    );

    or_bb _0852_ (
        .b(jinkela_wire_408),
        .a(jinkela_wire_788),
        .c(jinkela_wire_490)
    );

    and_bb _0433_ (
        .b(jinkela_wire_446),
        .a(jinkela_wire_562),
        .c(jinkela_wire_322)
    );

    and_bb _0853_ (
        .b(jinkela_wire_408),
        .a(jinkela_wire_788),
        .c(jinkela_wire_812)
    );

    or_bb _0434_ (
        .b(jinkela_wire_706),
        .a(jinkela_wire_188),
        .c(jinkela_wire_145)
    );

    or_bb _0854_ (
        .b(jinkela_wire_623),
        .a(jinkela_wire_803),
        .c(jinkela_wire_111)
    );

    and_bb _0435_ (
        .b(jinkela_wire_706),
        .a(jinkela_wire_188),
        .c(jinkela_wire_826)
    );

    and_bb _0855_ (
        .b(jinkela_wire_623),
        .a(jinkela_wire_803),
        .c(jinkela_wire_743)
    );

    or_bb _0436_ (
        .b(jinkela_wire_690),
        .a(jinkela_wire_412),
        .c(jinkela_wire_702)
    );

    or_bb _0856_ (
        .b(jinkela_wire_622),
        .a(jinkela_wire_750),
        .c(jinkela_wire_657)
    );

    and_bb _0437_ (
        .b(jinkela_wire_690),
        .a(jinkela_wire_412),
        .c(jinkela_wire_40)
    );

    and_bb _0857_ (
        .b(jinkela_wire_622),
        .a(jinkela_wire_750),
        .c(jinkela_wire_499)
    );

    or_bb _0438_ (
        .b(jinkela_wire_578),
        .a(jinkela_wire_145),
        .c(jinkela_wire_232)
    );

    or_bb _0858_ (
        .b(jinkela_wire_490),
        .a(jinkela_wire_111),
        .c(jinkela_wire_180)
    );

    or_bb _0439_ (
        .b(jinkela_wire_702),
        .a(jinkela_wire_232),
        .c(jinkela_wire_509)
    );

    or_bb _0859_ (
        .b(jinkela_wire_657),
        .a(jinkela_wire_180),
        .c(b_5_)
    );

    maj_bbb _0440_ (
        .c(jinkela_wire_578),
        .b(jinkela_wire_145),
        .a(jinkela_wire_702),
        .d(jinkela_wire_442)
    );

    maj_bbb _0860_ (
        .c(jinkela_wire_490),
        .b(jinkela_wire_111),
        .a(jinkela_wire_657),
        .d(b_4_)
    );

    and_bb _0441_ (
        .b(jinkela_wire_578),
        .a(jinkela_wire_145),
        .c(jinkela_wire_713)
    );

    and_bb _0861_ (
        .b(jinkela_wire_490),
        .a(jinkela_wire_111),
        .c(jinkela_wire_733)
    );

    and_bb _0442_ (
        .b(jinkela_wire_702),
        .a(jinkela_wire_713),
        .c(jinkela_wire_77)
    );

    and_bb _0862_ (
        .b(jinkela_wire_657),
        .a(jinkela_wire_733),
        .c(b_3_)
    );

    or_bb _0443_ (
        .b(jinkela_wire_322),
        .a(jinkela_wire_826),
        .c(jinkela_wire_556)
    );

    or_bb _0863_ (
        .b(jinkela_wire_812),
        .a(jinkela_wire_743),
        .c(jinkela_wire_110)
    );

    or_bb _0444_ (
        .b(jinkela_wire_40),
        .a(jinkela_wire_556),
        .c(jinkela_wire_727)
    );

    or_bb _0864_ (
        .b(jinkela_wire_499),
        .a(jinkela_wire_110),
        .c(b_2_)
    );

    maj_bbb _0445_ (
        .c(jinkela_wire_322),
        .b(jinkela_wire_826),
        .a(jinkela_wire_40),
        .d(jinkela_wire_205)
    );

    maj_bbb _0865_ (
        .c(jinkela_wire_812),
        .b(jinkela_wire_743),
        .a(jinkela_wire_499),
        .d(b_1_)
    );

    and_bb _0446_ (
        .b(jinkela_wire_322),
        .a(jinkela_wire_826),
        .c(jinkela_wire_209)
    );

    and_bb _0866_ (
        .b(jinkela_wire_812),
        .a(jinkela_wire_743),
        .c(jinkela_wire_224)
    );

    and_bb _0447_ (
        .b(jinkela_wire_40),
        .a(jinkela_wire_209),
        .c(jinkela_wire_82)
    );

    and_bb _0867_ (
        .b(jinkela_wire_499),
        .a(jinkela_wire_224),
        .c(b_0_)
    );

    or_bb _0448_ (
        .b(jinkela_wire_440),
        .a(jinkela_wire_756),
        .c(jinkela_wire_163)
    );

    or_bb _0868_ (
        .b(jinkela_wire_785),
        .a(jinkela_wire_406),
        .c(jinkela_wire_3)
    );

    and_bb _0449_ (
        .b(jinkela_wire_440),
        .a(jinkela_wire_756),
        .c(jinkela_wire_181)
    );

    and_bb _0869_ (
        .b(jinkela_wire_785),
        .a(jinkela_wire_406),
        .c(jinkela_wire_4)
    );

    or_bb _0450_ (
        .b(jinkela_wire_635),
        .a(jinkela_wire_44),
        .c(jinkela_wire_700)
    );

    or_bb _0870_ (
        .b(jinkela_wire_492),
        .a(jinkela_wire_67),
        .c(jinkela_wire_786)
    );

    and_bb _0451_ (
        .b(jinkela_wire_635),
        .a(jinkela_wire_44),
        .c(jinkela_wire_551)
    );

    and_bb _0871_ (
        .b(jinkela_wire_492),
        .a(jinkela_wire_67),
        .c(jinkela_wire_141)
    );

    or_bb _0452_ (
        .b(jinkela_wire_501),
        .a(jinkela_wire_17),
        .c(jinkela_wire_124)
    );

    or_bb _0872_ (
        .b(jinkela_wire_686),
        .a(jinkela_wire_8),
        .c(jinkela_wire_656)
    );

    and_bb _0453_ (
        .b(jinkela_wire_501),
        .a(jinkela_wire_17),
        .c(jinkela_wire_569)
    );

    and_bb _0873_ (
        .b(jinkela_wire_686),
        .a(jinkela_wire_8),
        .c(jinkela_wire_258)
    );

    or_bb _0454_ (
        .b(jinkela_wire_163),
        .a(jinkela_wire_700),
        .c(jinkela_wire_344)
    );

    or_bb _0874_ (
        .b(jinkela_wire_3),
        .a(jinkela_wire_786),
        .c(jinkela_wire_561)
    );

    or_bb _0455_ (
        .b(jinkela_wire_124),
        .a(jinkela_wire_344),
        .c(jinkela_wire_199)
    );

    or_bb _0875_ (
        .b(jinkela_wire_656),
        .a(jinkela_wire_561),
        .c(b_11_)
    );

    maj_bbb _0456_ (
        .c(jinkela_wire_163),
        .b(jinkela_wire_700),
        .a(jinkela_wire_124),
        .d(jinkela_wire_298)
    );

    maj_bbb _0876_ (
        .c(jinkela_wire_3),
        .b(jinkela_wire_786),
        .a(jinkela_wire_656),
        .d(b_10_)
    );

    and_bb _0457_ (
        .b(jinkela_wire_163),
        .a(jinkela_wire_700),
        .c(jinkela_wire_577)
    );

    and_bb _0877_ (
        .b(jinkela_wire_3),
        .a(jinkela_wire_786),
        .c(jinkela_wire_581)
    );

    and_bb _0458_ (
        .b(jinkela_wire_124),
        .a(jinkela_wire_577),
        .c(jinkela_wire_179)
    );

    and_bb _0878_ (
        .b(jinkela_wire_656),
        .a(jinkela_wire_581),
        .c(b_9_)
    );

    and_bb _0163_ (
        .b(a_47_),
        .a(a_46_),
        .c(jinkela_wire_399)
    );

    or_bb _0161_ (
        .b(a_45_),
        .a(jinkela_wire_806),
        .c(jinkela_wire_436)
    );

    or_bb _0459_ (
        .b(jinkela_wire_181),
        .a(jinkela_wire_551),
        .c(jinkela_wire_653)
    );

    or_bb _0879_ (
        .b(jinkela_wire_4),
        .a(jinkela_wire_141),
        .c(jinkela_wire_20)
    );

    maj_bbb _0162_ (
        .c(a_47_),
        .b(a_46_),
        .a(a_45_),
        .d(jinkela_wire_293)
    );

    or_bb _0460_ (
        .b(jinkela_wire_569),
        .a(jinkela_wire_653),
        .c(jinkela_wire_416)
    );

    or_bb _0880_ (
        .b(jinkela_wire_258),
        .a(jinkela_wire_20),
        .c(b_8_)
    );

    maj_bbb _0461_ (
        .c(jinkela_wire_181),
        .b(jinkela_wire_551),
        .a(jinkela_wire_569),
        .d(jinkela_wire_715)
    );

    or_bb _0160_ (
        .b(a_47_),
        .a(a_46_),
        .c(jinkela_wire_806)
    );

    maj_bbb _0881_ (
        .c(jinkela_wire_4),
        .b(jinkela_wire_141),
        .a(jinkela_wire_258),
        .d(b_7_)
    );

    and_bb _0164_ (
        .b(a_45_),
        .a(jinkela_wire_399),
        .c(jinkela_wire_616)
    );

    and_bb _0462_ (
        .b(jinkela_wire_181),
        .a(jinkela_wire_551),
        .c(jinkela_wire_388)
    );

    or_bb _0165_ (
        .b(a_44_),
        .a(a_43_),
        .c(jinkela_wire_787)
    );

    and_bb _0882_ (
        .b(jinkela_wire_4),
        .a(jinkela_wire_141),
        .c(jinkela_wire_318)
    );

    and_bb _0547_ (
        .b(jinkela_wire_694),
        .a(jinkela_wire_404),
        .c(jinkela_wire_605)
    );

    or_bb _0548_ (
        .b(jinkela_wire_707),
        .a(jinkela_wire_282),
        .c(jinkela_wire_169)
    );

    and_bb _0549_ (
        .b(jinkela_wire_707),
        .a(jinkela_wire_282),
        .c(jinkela_wire_384)
    );

    or_bb _0550_ (
        .b(jinkela_wire_488),
        .a(jinkela_wire_270),
        .c(jinkela_wire_758)
    );

    or_bb _0551_ (
        .b(jinkela_wire_169),
        .a(jinkela_wire_758),
        .c(jinkela_wire_128)
    );

    maj_bbb _0552_ (
        .c(jinkela_wire_488),
        .b(jinkela_wire_270),
        .a(jinkela_wire_169),
        .d(jinkela_wire_365)
    );

    and_bb _0553_ (
        .b(jinkela_wire_488),
        .a(jinkela_wire_270),
        .c(jinkela_wire_347)
    );

    and_bb _0554_ (
        .b(jinkela_wire_169),
        .a(jinkela_wire_347),
        .c(jinkela_wire_278)
    );

    or_bb _0555_ (
        .b(jinkela_wire_660),
        .a(jinkela_wire_605),
        .c(jinkela_wire_586)
    );

    or_bb _0556_ (
        .b(jinkela_wire_384),
        .a(jinkela_wire_586),
        .c(jinkela_wire_92)
    );

    maj_bbb _0557_ (
        .c(jinkela_wire_660),
        .b(jinkela_wire_605),
        .a(jinkela_wire_384),
        .d(jinkela_wire_395)
    );

    and_bb _0558_ (
        .b(jinkela_wire_660),
        .a(jinkela_wire_605),
        .c(jinkela_wire_709)
    );

    and_bb _0559_ (
        .b(jinkela_wire_384),
        .a(jinkela_wire_709),
        .c(jinkela_wire_459)
    );

    and_bb _0545_ (
        .b(jinkela_wire_190),
        .a(jinkela_wire_604),
        .c(jinkela_wire_660)
    );

    or_bb _0560_ (
        .b(a_11_),
        .a(a_10_),
        .c(jinkela_wire_572)
    );

    or_bb _0561_ (
        .b(a_9_),
        .a(jinkela_wire_572),
        .c(jinkela_wire_485)
    );

    maj_bbb _0562_ (
        .c(a_11_),
        .b(a_10_),
        .a(a_9_),
        .d(jinkela_wire_516)
    );

    and_bb _0563_ (
        .b(a_11_),
        .a(a_10_),
        .c(jinkela_wire_153)
    );

    and_bb _0564_ (
        .b(a_9_),
        .a(jinkela_wire_153),
        .c(jinkela_wire_438)
    );

    or_bb _0546_ (
        .b(jinkela_wire_694),
        .a(jinkela_wire_404),
        .c(jinkela_wire_270)
    );

    or_bb _0565_ (
        .b(a_8_),
        .a(a_7_),
        .c(jinkela_wire_433)
    );

    or_bb _0566_ (
        .b(a_6_),
        .a(jinkela_wire_433),
        .c(jinkela_wire_309)
    );

    maj_bbb _0567_ (
        .c(a_8_),
        .b(a_7_),
        .a(a_6_),
        .d(jinkela_wire_227)
    );

    and_bb _0568_ (
        .b(a_8_),
        .a(a_7_),
        .c(jinkela_wire_383)
    );

    and_bb _0569_ (
        .b(a_6_),
        .a(jinkela_wire_383),
        .c(jinkela_wire_130)
    );

    or_bb _0570_ (
        .b(jinkela_wire_485),
        .a(jinkela_wire_130),
        .c(jinkela_wire_161)
    );

    and_bb _0571_ (
        .b(jinkela_wire_485),
        .a(jinkela_wire_130),
        .c(jinkela_wire_148)
    );

    or_bb _0572_ (
        .b(jinkela_wire_516),
        .a(jinkela_wire_227),
        .c(jinkela_wire_372)
    );

    and_bb _0573_ (
        .b(jinkela_wire_516),
        .a(jinkela_wire_227),
        .c(jinkela_wire_115)
    );

    or_bb _0574_ (
        .b(jinkela_wire_438),
        .a(jinkela_wire_309),
        .c(jinkela_wire_802)
    );

    and_bb _0575_ (
        .b(jinkela_wire_438),
        .a(jinkela_wire_309),
        .c(jinkela_wire_545)
    );

    or_bb _0576_ (
        .b(jinkela_wire_161),
        .a(jinkela_wire_372),
        .c(jinkela_wire_629)
    );

    or_bb _0577_ (
        .b(jinkela_wire_802),
        .a(jinkela_wire_629),
        .c(jinkela_wire_178)
    );

    maj_bbb _0578_ (
        .c(jinkela_wire_161),
        .b(jinkela_wire_372),
        .a(jinkela_wire_802),
        .d(jinkela_wire_84)
    );

    and_bb _0579_ (
        .b(jinkela_wire_161),
        .a(jinkela_wire_372),
        .c(jinkela_wire_628)
    );

    and_bb _0580_ (
        .b(jinkela_wire_802),
        .a(jinkela_wire_628),
        .c(jinkela_wire_74)
    );

    or_bb _0581_ (
        .b(jinkela_wire_148),
        .a(jinkela_wire_115),
        .c(jinkela_wire_606)
    );

    and_bb _0629_ (
        .b(jinkela_wire_35),
        .a(jinkela_wire_398),
        .c(jinkela_wire_76)
    );

    or_bb _0582_ (
        .b(jinkela_wire_545),
        .a(jinkela_wire_606),
        .c(jinkela_wire_823)
    );

    maj_bbb _0583_ (
        .c(jinkela_wire_148),
        .b(jinkela_wire_115),
        .a(jinkela_wire_545),
        .d(jinkela_wire_712)
    );

    and_bb _0584_ (
        .b(jinkela_wire_148),
        .a(jinkela_wire_115),
        .c(jinkela_wire_719)
    );

    and_bb _0585_ (
        .b(jinkela_wire_545),
        .a(jinkela_wire_719),
        .c(jinkela_wire_603)
    );

    or_bb _0586_ (
        .b(a_5_),
        .a(a_4_),
        .c(jinkela_wire_540)
    );

    or_bb _0630_ (
        .b(jinkela_wire_356),
        .a(jinkela_wire_816),
        .c(jinkela_wire_57)
    );

    or_bb _0587_ (
        .b(a_3_),
        .a(jinkela_wire_540),
        .c(jinkela_wire_539)
    );

    maj_bbb _0588_ (
        .c(a_5_),
        .b(a_4_),
        .a(a_3_),
        .d(jinkela_wire_456)
    );

    and_bb _0463_ (
        .b(jinkela_wire_569),
        .a(jinkela_wire_388),
        .c(jinkela_wire_595)
    );

    and_bb _0505_ (
        .b(jinkela_wire_495),
        .a(jinkela_wire_30),
        .c(jinkela_wire_409)
    );

    and_bb _0589_ (
        .b(a_5_),
        .a(a_4_),
        .c(jinkela_wire_177)
    );

    and_bb _0673_ (
        .b(jinkela_wire_278),
        .a(jinkela_wire_419),
        .c(jinkela_wire_264)
    );

    and_bb _0883_ (
        .b(jinkela_wire_258),
        .a(jinkela_wire_318),
        .c(b_6_)
    );

    and_bb _1009_ (
        .b(jinkela_wire_646),
        .a(jinkela_wire_502),
        .c(jinkela_wire_620)
    );

    or_bb _0464_ (
        .b(a_23_),
        .a(a_22_),
        .c(jinkela_wire_19)
    );

    or_bb _0506_ (
        .b(jinkela_wire_390),
        .a(jinkela_wire_289),
        .c(jinkela_wire_716)
    );

    and_bb _0590_ (
        .b(a_3_),
        .a(jinkela_wire_177),
        .c(jinkela_wire_59)
    );

    or_bb _0674_ (
        .b(jinkela_wire_365),
        .a(jinkela_wire_334),
        .c(jinkela_wire_325)
    );

    or_bb _0884_ (
        .b(jinkela_wire_38),
        .a(jinkela_wire_97),
        .c(jinkela_wire_301)
    );

    or_bb _1010_ (
        .b(jinkela_wire_194),
        .a(jinkela_wire_223),
        .c(jinkela_wire_644)
    );

    or_bb _0465_ (
        .b(a_21_),
        .a(jinkela_wire_19),
        .c(jinkela_wire_467)
    );

    or_bb _0507_ (
        .b(jinkela_wire_10),
        .a(jinkela_wire_716),
        .c(jinkela_wire_196)
    );

    or_bb _0591_ (
        .b(a_2_),
        .a(a_1_),
        .c(jinkela_wire_773)
    );

    and_bb _0675_ (
        .b(jinkela_wire_365),
        .a(jinkela_wire_334),
        .c(jinkela_wire_528)
    );

    and_bb _0885_ (
        .b(jinkela_wire_38),
        .a(jinkela_wire_97),
        .c(jinkela_wire_697)
    );

    and_bb _1011_ (
        .b(jinkela_wire_194),
        .a(jinkela_wire_223),
        .c(jinkela_wire_530)
    );

    maj_bbb _0466_ (
        .c(a_23_),
        .b(a_22_),
        .a(a_21_),
        .d(jinkela_wire_175)
    );

    maj_bbb _0508_ (
        .c(jinkela_wire_390),
        .b(jinkela_wire_289),
        .a(jinkela_wire_10),
        .d(jinkela_wire_147)
    );

    or_bb _0592_ (
        .b(a_0_),
        .a(jinkela_wire_773),
        .c(jinkela_wire_640)
    );

    or_bb _0676_ (
        .b(jinkela_wire_128),
        .a(jinkela_wire_381),
        .c(jinkela_wire_761)
    );

    or_bb _0886_ (
        .b(jinkela_wire_64),
        .a(jinkela_wire_34),
        .c(jinkela_wire_219)
    );

    or_bb _1012_ (
        .b(jinkela_wire_198),
        .a(jinkela_wire_324),
        .c(jinkela_wire_320)
    );

    and_bb _0467_ (
        .b(a_23_),
        .a(a_22_),
        .c(jinkela_wire_639)
    );

    and_bb _0509_ (
        .b(jinkela_wire_390),
        .a(jinkela_wire_289),
        .c(jinkela_wire_770)
    );

    maj_bbb _0593_ (
        .c(a_2_),
        .b(a_1_),
        .a(a_0_),
        .d(jinkela_wire_151)
    );

    and_bb _0677_ (
        .b(jinkela_wire_128),
        .a(jinkela_wire_381),
        .c(jinkela_wire_666)
    );

    and_bb _0887_ (
        .b(jinkela_wire_64),
        .a(jinkela_wire_34),
        .c(jinkela_wire_189)
    );

    and_bb _1013_ (
        .b(jinkela_wire_198),
        .a(jinkela_wire_324),
        .c(jinkela_wire_73)
    );

    and_bb _0468_ (
        .b(a_21_),
        .a(jinkela_wire_639),
        .c(jinkela_wire_257)
    );

    and_bb _0510_ (
        .b(jinkela_wire_10),
        .a(jinkela_wire_770),
        .c(jinkela_wire_591)
    );

    and_bb _0594_ (
        .b(a_2_),
        .a(a_1_),
        .c(jinkela_wire_396)
    );

    or_bb _0678_ (
        .b(jinkela_wire_531),
        .a(jinkela_wire_429),
        .c(jinkela_wire_489)
    );

    or_bb _0888_ (
        .b(jinkela_wire_598),
        .a(jinkela_wire_354),
        .c(jinkela_wire_109)
    );

    or_bb _1014_ (
        .b(jinkela_wire_571),
        .a(jinkela_wire_644),
        .c(jinkela_wire_370)
    );

    or_bb _0469_ (
        .b(a_20_),
        .a(a_19_),
        .c(jinkela_wire_615)
    );

    or_bb _0511_ (
        .b(jinkela_wire_371),
        .a(jinkela_wire_546),
        .c(jinkela_wire_611)
    );

    and_bb _0595_ (
        .b(a_0_),
        .a(jinkela_wire_396),
        .c(jinkela_wire_281)
    );

    and_bb _0679_ (
        .b(jinkela_wire_531),
        .a(jinkela_wire_429),
        .c(jinkela_wire_655)
    );

    and_bb _0889_ (
        .b(jinkela_wire_598),
        .a(jinkela_wire_354),
        .c(jinkela_wire_519)
    );

    or_bb _1015_ (
        .b(jinkela_wire_320),
        .a(jinkela_wire_370),
        .c(b_41_)
    );

    or_bb _0470_ (
        .b(a_18_),
        .a(jinkela_wire_615),
        .c(jinkela_wire_16)
    );

    or_bb _0512_ (
        .b(jinkela_wire_409),
        .a(jinkela_wire_611),
        .c(jinkela_wire_420)
    );

    or_bb _0596_ (
        .b(jinkela_wire_539),
        .a(jinkela_wire_281),
        .c(jinkela_wire_243)
    );

    or_bb _0680_ (
        .b(jinkela_wire_434),
        .a(jinkela_wire_655),
        .c(jinkela_wire_813)
    );

    or_bb _0890_ (
        .b(jinkela_wire_782),
        .a(jinkela_wire_486),
        .c(jinkela_wire_508)
    );

    maj_bbb _1016_ (
        .c(jinkela_wire_571),
        .b(jinkela_wire_644),
        .a(jinkela_wire_320),
        .d(b_40_)
    );

    maj_bbb _0471_ (
        .c(a_20_),
        .b(a_19_),
        .a(a_18_),
        .d(jinkela_wire_171)
    );

    maj_bbb _0513_ (
        .c(jinkela_wire_371),
        .b(jinkela_wire_546),
        .a(jinkela_wire_409),
        .d(jinkela_wire_236)
    );

    and_bb _0597_ (
        .b(jinkela_wire_539),
        .a(jinkela_wire_281),
        .c(jinkela_wire_32)
    );

    and_bb _0681_ (
        .b(jinkela_wire_434),
        .a(jinkela_wire_655),
        .c(jinkela_wire_69)
    );

    and_bb _0891_ (
        .b(jinkela_wire_782),
        .a(jinkela_wire_486),
        .c(jinkela_wire_279)
    );

    and_bb _1017_ (
        .b(jinkela_wire_571),
        .a(jinkela_wire_644),
        .c(jinkela_wire_633)
    );

    and_bb _0472_ (
        .b(a_20_),
        .a(a_19_),
        .c(jinkela_wire_400)
    );

    and_bb _0514_ (
        .b(jinkela_wire_371),
        .a(jinkela_wire_546),
        .c(jinkela_wire_504)
    );

    or_bb _0598_ (
        .b(jinkela_wire_456),
        .a(jinkela_wire_151),
        .c(jinkela_wire_755)
    );

    or_bb _0682_ (
        .b(jinkela_wire_585),
        .a(jinkela_wire_637),
        .c(jinkela_wire_589)
    );

    or_bb _0892_ (
        .b(jinkela_wire_271),
        .a(jinkela_wire_650),
        .c(jinkela_wire_544)
    );

    and_bb _1018_ (
        .b(jinkela_wire_320),
        .a(jinkela_wire_633),
        .c(b_39_)
    );

    and_bb _0473_ (
        .b(a_18_),
        .a(jinkela_wire_400),
        .c(jinkela_wire_729)
    );

    and_bb _0515_ (
        .b(jinkela_wire_409),
        .a(jinkela_wire_504),
        .c(jinkela_wire_167)
    );

    and_bb _0599_ (
        .b(jinkela_wire_456),
        .a(jinkela_wire_151),
        .c(jinkela_wire_828)
    );

    and_bb _0683_ (
        .b(jinkela_wire_585),
        .a(jinkela_wire_637),
        .c(jinkela_wire_470)
    );

    and_bb _0893_ (
        .b(jinkela_wire_271),
        .a(jinkela_wire_650),
        .c(jinkela_wire_75)
    );

    or_bb _1019_ (
        .b(jinkela_wire_620),
        .a(jinkela_wire_530),
        .c(jinkela_wire_766)
    );

    or_bb _0474_ (
        .b(jinkela_wire_467),
        .a(jinkela_wire_729),
        .c(jinkela_wire_643)
    );

    or_bb _0516_ (
        .b(jinkela_wire_213),
        .a(jinkela_wire_196),
        .c(jinkela_wire_282)
    );

    or_bb _0600_ (
        .b(jinkela_wire_59),
        .a(jinkela_wire_640),
        .c(jinkela_wire_302)
    );

    or_bb _0684_ (
        .b(jinkela_wire_78),
        .a(jinkela_wire_814),
        .c(jinkela_wire_126)
    );

    or_bb _0894_ (
        .b(jinkela_wire_417),
        .a(jinkela_wire_685),
        .c(jinkela_wire_612)
    );

    or_bb _1020_ (
        .b(jinkela_wire_73),
        .a(jinkela_wire_766),
        .c(b_38_)
    );

    and_bb _0475_ (
        .b(jinkela_wire_467),
        .a(jinkela_wire_729),
        .c(jinkela_wire_184)
    );

    and_bb _0517_ (
        .b(jinkela_wire_213),
        .a(jinkela_wire_196),
        .c(jinkela_wire_689)
    );

    and_bb _0601_ (
        .b(jinkela_wire_59),
        .a(jinkela_wire_640),
        .c(jinkela_wire_374)
    );

    and_bb _0685_ (
        .b(jinkela_wire_78),
        .a(jinkela_wire_814),
        .c(jinkela_wire_317)
    );

    and_bb _0713_ (
        .b(jinkela_wire_746),
        .a(jinkela_wire_813),
        .c(jinkela_wire_47)
    );

    and_bb _0895_ (
        .b(jinkela_wire_417),
        .a(jinkela_wire_685),
        .c(jinkela_wire_737)
    );

    or_bb _0476_ (
        .b(jinkela_wire_175),
        .a(jinkela_wire_171),
        .c(jinkela_wire_31)
    );

    or_bb _0518_ (
        .b(jinkela_wire_505),
        .a(jinkela_wire_147),
        .c(jinkela_wire_404)
    );

    or_bb _0602_ (
        .b(jinkela_wire_243),
        .a(jinkela_wire_755),
        .c(jinkela_wire_634)
    );

    or_bb _0686_ (
        .b(jinkela_wire_264),
        .a(jinkela_wire_221),
        .c(jinkela_wire_746)
    );

    or_bb _0896_ (
        .b(jinkela_wire_737),
        .a(jinkela_wire_519),
        .c(jinkela_wire_559)
    );

    and_bb _1022_ (
        .b(jinkela_wire_620),
        .a(jinkela_wire_530),
        .c(jinkela_wire_696)
    );

    and_bb _0477_ (
        .b(jinkela_wire_175),
        .a(jinkela_wire_171),
        .c(jinkela_wire_29)
    );

    and_bb _0519_ (
        .b(jinkela_wire_505),
        .a(jinkela_wire_147),
        .c(jinkela_wire_340)
    );

    or_bb _0603_ (
        .b(jinkela_wire_302),
        .a(jinkela_wire_634),
        .c(jinkela_wire_168)
    );

    and_bb _0687_ (
        .b(jinkela_wire_264),
        .a(jinkela_wire_221),
        .c(jinkela_wire_824)
    );

    and_bb _0897_ (
        .b(jinkela_wire_737),
        .a(jinkela_wire_519),
        .c(jinkela_wire_763)
    );

    and_bb _1023_ (
        .b(jinkela_wire_73),
        .a(jinkela_wire_696),
        .c(b_36_)
    );

    or_bb _0478_ (
        .b(jinkela_wire_257),
        .a(jinkela_wire_16),
        .c(jinkela_wire_359)
    );

    or_bb _0520_ (
        .b(jinkela_wire_296),
        .a(jinkela_wire_591),
        .c(jinkela_wire_604)
    );

    maj_bbb _0604_ (
        .c(jinkela_wire_243),
        .b(jinkela_wire_755),
        .a(jinkela_wire_302),
        .d(jinkela_wire_594)
    );

    or_bb _0688_ (
        .b(jinkela_wire_528),
        .a(jinkela_wire_500),
        .c(jinkela_wire_245)
    );

    or_bb _0898_ (
        .b(jinkela_wire_75),
        .a(jinkela_wire_189),
        .c(jinkela_wire_230)
    );

    or_bb _1024_ (
        .b(jinkela_wire_105),
        .a(jinkela_wire_579),
        .c(jinkela_wire_463)
    );

    and_bb _0479_ (
        .b(jinkela_wire_257),
        .a(jinkela_wire_16),
        .c(jinkela_wire_809)
    );

    and_bb _0521_ (
        .b(jinkela_wire_296),
        .a(jinkela_wire_591),
        .c(jinkela_wire_822)
    );

    and_bb _0605_ (
        .b(jinkela_wire_243),
        .a(jinkela_wire_755),
        .c(jinkela_wire_673)
    );

    and_bb _0689_ (
        .b(jinkela_wire_528),
        .a(jinkela_wire_500),
        .c(jinkela_wire_811)
    );

    and_bb _0899_ (
        .b(jinkela_wire_75),
        .a(jinkela_wire_189),
        .c(jinkela_wire_792)
    );

    and_bb _1025_ (
        .b(jinkela_wire_105),
        .a(jinkela_wire_579),
        .c(jinkela_wire_714)
    );

    or_bb _0480_ (
        .b(jinkela_wire_643),
        .a(jinkela_wire_31),
        .c(jinkela_wire_621)
    );

    or_bb _0522_ (
        .b(jinkela_wire_552),
        .a(jinkela_wire_420),
        .c(jinkela_wire_707)
    );

    and_bb _0606_ (
        .b(jinkela_wire_302),
        .a(jinkela_wire_673),
        .c(jinkela_wire_121)
    );

    or_bb _0690_ (
        .b(jinkela_wire_666),
        .a(jinkela_wire_112),
        .c(jinkela_wire_658)
    );

    or_bb _0714_ (
        .b(jinkela_wire_63),
        .a(jinkela_wire_704),
        .c(jinkela_wire_138)
    );

    or_bb _0900_ (
        .b(jinkela_wire_279),
        .a(jinkela_wire_697),
        .c(jinkela_wire_484)
    );

    or_bb _0481_ (
        .b(jinkela_wire_359),
        .a(jinkela_wire_621),
        .c(jinkela_wire_288)
    );

    and_bb _0523_ (
        .b(jinkela_wire_552),
        .a(jinkela_wire_420),
        .c(jinkela_wire_118)
    );

    or_bb _0607_ (
        .b(jinkela_wire_32),
        .a(jinkela_wire_828),
        .c(jinkela_wire_555)
    );

    and_bb _0691_ (
        .b(jinkela_wire_666),
        .a(jinkela_wire_112),
        .c(jinkela_wire_800)
    );

    and_bb _0901_ (
        .b(jinkela_wire_279),
        .a(jinkela_wire_697),
        .c(jinkela_wire_573)
    );

    and_bb _1027_ (
        .b(jinkela_wire_231),
        .a(jinkela_wire_273),
        .c(jinkela_wire_473)
    );

    maj_bbb _0482_ (
        .c(jinkela_wire_643),
        .b(jinkela_wire_31),
        .a(jinkela_wire_359),
        .d(jinkela_wire_55)
    );

    or_bb _0524_ (
        .b(jinkela_wire_55),
        .a(jinkela_wire_236),
        .c(jinkela_wire_694)
    );

    or_bb _0608_ (
        .b(jinkela_wire_374),
        .a(jinkela_wire_555),
        .c(jinkela_wire_319)
    );

    or_bb _0692_ (
        .b(jinkela_wire_800),
        .a(jinkela_wire_317),
        .c(jinkela_wire_379)
    );

    or_bb _0902_ (
        .b(jinkela_wire_559),
        .a(jinkela_wire_230),
        .c(jinkela_wire_42)
    );

    or_bb _1028_ (
        .b(jinkela_wire_339),
        .a(jinkela_wire_652),
        .c(jinkela_wire_132)
    );

    and_bb _0483_ (
        .b(jinkela_wire_643),
        .a(jinkela_wire_31),
        .c(jinkela_wire_54)
    );

    and_bb _0525_ (
        .b(jinkela_wire_55),
        .a(jinkela_wire_236),
        .c(jinkela_wire_448)
    );

    maj_bbb _0609_ (
        .c(jinkela_wire_32),
        .b(jinkela_wire_828),
        .a(jinkela_wire_374),
        .d(jinkela_wire_253)
    );

    and_bb _0693_ (
        .b(jinkela_wire_800),
        .a(jinkela_wire_317),
        .c(jinkela_wire_328)
    );

    or_bb _0903_ (
        .b(jinkela_wire_484),
        .a(jinkela_wire_42),
        .c(b_17_)
    );

    and_bb _1029_ (
        .b(jinkela_wire_339),
        .a(jinkela_wire_652),
        .c(jinkela_wire_86)
    );

    and_bb _0484_ (
        .b(jinkela_wire_359),
        .a(jinkela_wire_54),
        .c(jinkela_wire_552)
    );

    or_bb _0526_ (
        .b(jinkela_wire_288),
        .a(jinkela_wire_167),
        .c(jinkela_wire_190)
    );

    and_bb _0610_ (
        .b(jinkela_wire_32),
        .a(jinkela_wire_828),
        .c(jinkela_wire_776)
    );

    or_bb _0694_ (
        .b(jinkela_wire_811),
        .a(jinkela_wire_470),
        .c(jinkela_wire_321)
    );

    maj_bbb _0904_ (
        .c(jinkela_wire_559),
        .b(jinkela_wire_230),
        .a(jinkela_wire_484),
        .d(b_16_)
    );

    or_bb _1030_ (
        .b(jinkela_wire_463),
        .a(jinkela_wire_237),
        .c(jinkela_wire_104)
    );

    or_bb _0485_ (
        .b(jinkela_wire_184),
        .a(jinkela_wire_29),
        .c(jinkela_wire_674)
    );

    and_bb _0527_ (
        .b(jinkela_wire_288),
        .a(jinkela_wire_167),
        .c(jinkela_wire_654)
    );

    and_bb _0611_ (
        .b(jinkela_wire_374),
        .a(jinkela_wire_776),
        .c(jinkela_wire_348)
    );

    and_bb _0695_ (
        .b(jinkela_wire_811),
        .a(jinkela_wire_470),
        .c(jinkela_wire_93)
    );

    and_bb _0905_ (
        .b(jinkela_wire_559),
        .a(jinkela_wire_230),
        .c(jinkela_wire_306)
    );

    or_bb _1031_ (
        .b(jinkela_wire_132),
        .a(jinkela_wire_104),
        .c(b_47_)
    );

    or_bb _0486_ (
        .b(jinkela_wire_809),
        .a(jinkela_wire_674),
        .c(jinkela_wire_296)
    );

    or_bb _0528_ (
        .b(jinkela_wire_654),
        .a(jinkela_wire_822),
        .c(jinkela_wire_518)
    );

    or_bb _0612_ (
        .b(jinkela_wire_603),
        .a(jinkela_wire_168),
        .c(jinkela_wire_543)
    );

    or_bb _0696_ (
        .b(jinkela_wire_824),
        .a(jinkela_wire_69),
        .c(jinkela_wire_234)
    );

    and_bb _0906_ (
        .b(jinkela_wire_484),
        .a(jinkela_wire_306),
        .c(b_15_)
    );

    maj_bbb _1032_ (
        .c(jinkela_wire_463),
        .b(jinkela_wire_237),
        .a(jinkela_wire_132),
        .d(b_46_)
    );

    maj_bbb _0487_ (
        .c(jinkela_wire_184),
        .b(jinkela_wire_29),
        .a(jinkela_wire_809),
        .d(jinkela_wire_505)
    );

    and_bb _0529_ (
        .b(jinkela_wire_654),
        .a(jinkela_wire_822),
        .c(jinkela_wire_487)
    );

    and_bb _0613_ (
        .b(jinkela_wire_603),
        .a(jinkela_wire_168),
        .c(jinkela_wire_398)
    );

    and_bb _0697_ (
        .b(jinkela_wire_824),
        .a(jinkela_wire_69),
        .c(jinkela_wire_131)
    );

    or_bb _0907_ (
        .b(jinkela_wire_763),
        .a(jinkela_wire_792),
        .c(jinkela_wire_736)
    );

    and_bb _1033_ (
        .b(jinkela_wire_463),
        .a(jinkela_wire_237),
        .c(jinkela_wire_791)
    );

    and_bb _0488_ (
        .b(jinkela_wire_184),
        .a(jinkela_wire_29),
        .c(jinkela_wire_274)
    );

    or_bb _0530_ (
        .b(jinkela_wire_448),
        .a(jinkela_wire_340),
        .c(jinkela_wire_424)
    );

    or_bb _0614_ (
        .b(jinkela_wire_712),
        .a(jinkela_wire_594),
        .c(jinkela_wire_829)
    );

    or_bb _0698_ (
        .b(jinkela_wire_379),
        .a(jinkela_wire_321),
        .c(jinkela_wire_804)
    );

    or_bb _0908_ (
        .b(jinkela_wire_573),
        .a(jinkela_wire_736),
        .c(b_14_)
    );

    and_bb _1034_ (
        .b(jinkela_wire_132),
        .a(jinkela_wire_791),
        .c(b_45_)
    );

    and_bb _0489_ (
        .b(jinkela_wire_809),
        .a(jinkela_wire_274),
        .c(jinkela_wire_213)
    );

    and_bb _0531_ (
        .b(jinkela_wire_448),
        .a(jinkela_wire_340),
        .c(jinkela_wire_305)
    );

    and_bb _0615_ (
        .b(jinkela_wire_712),
        .a(jinkela_wire_594),
        .c(jinkela_wire_799)
    );

    or_bb _0699_ (
        .b(jinkela_wire_234),
        .a(jinkela_wire_804),
        .c(jinkela_wire_2)
    );

    maj_bbb _0909_ (
        .c(jinkela_wire_763),
        .b(jinkela_wire_792),
        .a(jinkela_wire_573),
        .d(b_13_)
    );

    or_bb _1035_ (
        .b(jinkela_wire_714),
        .a(jinkela_wire_473),
        .c(jinkela_wire_152)
    );

    or_bb _0490_ (
        .b(a_17_),
        .a(a_16_),
        .c(jinkela_wire_476)
    );

    or_bb _0532_ (
        .b(jinkela_wire_118),
        .a(jinkela_wire_689),
        .c(jinkela_wire_701)
    );

    or_bb _0616_ (
        .b(jinkela_wire_823),
        .a(jinkela_wire_121),
        .c(jinkela_wire_239)
    );

    maj_bbb _0700_ (
        .c(jinkela_wire_379),
        .b(jinkela_wire_321),
        .a(jinkela_wire_234),
        .d(jinkela_wire_103)
    );

    and_bb _0910_ (
        .b(jinkela_wire_763),
        .a(jinkela_wire_792),
        .c(jinkela_wire_475)
    );

    or_bb _1036_ (
        .b(jinkela_wire_86),
        .a(jinkela_wire_152),
        .c(b_44_)
    );

    or_bb _0491_ (
        .b(a_15_),
        .a(jinkela_wire_476),
        .c(jinkela_wire_61)
    );

    and_bb _0533_ (
        .b(jinkela_wire_118),
        .a(jinkela_wire_689),
        .c(jinkela_wire_529)
    );

    and_bb _0617_ (
        .b(jinkela_wire_823),
        .a(jinkela_wire_121),
        .c(jinkela_wire_373)
    );

    and_bb _0701_ (
        .b(jinkela_wire_379),
        .a(jinkela_wire_321),
        .c(jinkela_wire_407)
    );

    and_bb _0911_ (
        .b(jinkela_wire_573),
        .a(jinkela_wire_475),
        .c(b_12_)
    );

    maj_bbb _1037_ (
        .c(jinkela_wire_714),
        .b(jinkela_wire_473),
        .a(jinkela_wire_86),
        .d(b_43_)
    );

    maj_bbb _0492_ (
        .c(a_17_),
        .b(a_16_),
        .a(a_15_),
        .d(jinkela_wire_134)
    );

    or_bb _0534_ (
        .b(jinkela_wire_518),
        .a(jinkela_wire_424),
        .c(jinkela_wire_753)
    );

    or_bb _0618_ (
        .b(jinkela_wire_74),
        .a(jinkela_wire_319),
        .c(jinkela_wire_70)
    );

    and_bb _0702_ (
        .b(jinkela_wire_234),
        .a(jinkela_wire_407),
        .c(jinkela_wire_144)
    );

    or_bb _0912_ (
        .b(jinkela_wire_612),
        .a(jinkela_wire_109),
        .c(jinkela_wire_284)
    );

    and_bb _1038_ (
        .b(jinkela_wire_714),
        .a(jinkela_wire_473),
        .c(jinkela_wire_462)
    );

    and_bb _0493_ (
        .b(a_17_),
        .a(a_16_),
        .c(jinkela_wire_481)
    );

    or_bb _0535_ (
        .b(jinkela_wire_701),
        .a(jinkela_wire_753),
        .c(jinkela_wire_401)
    );

    and_bb _0619_ (
        .b(jinkela_wire_74),
        .a(jinkela_wire_319),
        .c(jinkela_wire_35)
    );

    or_bb _0703_ (
        .b(jinkela_wire_328),
        .a(jinkela_wire_93),
        .c(jinkela_wire_283)
    );

    and_bb _0913_ (
        .b(jinkela_wire_612),
        .a(jinkela_wire_109),
        .c(jinkela_wire_246)
    );

    and_bb _1039_ (
        .b(jinkela_wire_86),
        .a(jinkela_wire_462),
        .c(b_42_)
    );

    and_bb _0494_ (
        .b(a_15_),
        .a(jinkela_wire_481),
        .c(jinkela_wire_495)
    );

    maj_bbb _0536_ (
        .c(jinkela_wire_518),
        .b(jinkela_wire_424),
        .a(jinkela_wire_701),
        .d(jinkela_wire_156)
    );

    or_bb _0620_ (
        .b(jinkela_wire_84),
        .a(jinkela_wire_253),
        .c(jinkela_wire_226)
    );

    or_bb _0704_ (
        .b(jinkela_wire_131),
        .a(jinkela_wire_283),
        .c(jinkela_wire_362)
    );

    or_bb _0914_ (
        .b(jinkela_wire_544),
        .a(jinkela_wire_219),
        .c(jinkela_wire_796)
    );

    or_bb _0495_ (
        .b(a_14_),
        .a(a_13_),
        .c(jinkela_wire_12)
    );

    and_bb _0537_ (
        .b(jinkela_wire_518),
        .a(jinkela_wire_424),
        .c(jinkela_wire_662)
    );

    and_bb _0621_ (
        .b(jinkela_wire_84),
        .a(jinkela_wire_253),
        .c(jinkela_wire_517)
    );

    maj_bbb _0705_ (
        .c(jinkela_wire_328),
        .b(jinkela_wire_93),
        .a(jinkela_wire_131),
        .d(jinkela_wire_478)
    );

    and_bb _0915_ (
        .b(jinkela_wire_544),
        .a(jinkela_wire_219),
        .c(jinkela_wire_123)
    );

    or_bb _0496_ (
        .b(a_12_),
        .a(jinkela_wire_12),
        .c(jinkela_wire_30)
    );

    and_bb _0538_ (
        .b(jinkela_wire_701),
        .a(jinkela_wire_662),
        .c(jinkela_wire_580)
    );

    or_bb _0622_ (
        .b(jinkela_wire_178),
        .a(jinkela_wire_348),
        .c(jinkela_wire_817)
    );

    and_bb _0706_ (
        .b(jinkela_wire_328),
        .a(jinkela_wire_93),
        .c(jinkela_wire_235)
    );

    or_bb _0916_ (
        .b(jinkela_wire_508),
        .a(jinkela_wire_301),
        .c(jinkela_wire_262)
    );

    maj_bbb _0497_ (
        .c(a_14_),
        .b(a_13_),
        .a(a_12_),
        .d(jinkela_wire_661)
    );

    or_bb _0539_ (
        .b(jinkela_wire_487),
        .a(jinkela_wire_305),
        .c(jinkela_wire_421)
    );

    and_bb _0623_ (
        .b(jinkela_wire_178),
        .a(jinkela_wire_348),
        .c(jinkela_wire_717)
    );

    and_bb _0707_ (
        .b(jinkela_wire_131),
        .a(jinkela_wire_235),
        .c(jinkela_wire_51)
    );

    and_bb _0917_ (
        .b(jinkela_wire_508),
        .a(jinkela_wire_301),
        .c(jinkela_wire_565)
    );

    and_bb _0498_ (
        .b(a_14_),
        .a(a_13_),
        .c(jinkela_wire_748)
    );

    or_bb _0540_ (
        .b(jinkela_wire_529),
        .a(jinkela_wire_421),
        .c(jinkela_wire_711)
    );

    or_bb _0624_ (
        .b(jinkela_wire_717),
        .a(jinkela_wire_373),
        .c(jinkela_wire_356)
    );

    or_bb _0708_ (
        .b(jinkela_wire_658),
        .a(jinkela_wire_126),
        .c(jinkela_wire_63)
    );

    or_bb _0918_ (
        .b(jinkela_wire_284),
        .a(jinkela_wire_796),
        .c(jinkela_wire_427)
    );

    and_bb _0499_ (
        .b(a_12_),
        .a(jinkela_wire_748),
        .c(jinkela_wire_297)
    );

    maj_bbb _0541_ (
        .c(jinkela_wire_487),
        .b(jinkela_wire_305),
        .a(jinkela_wire_529),
        .d(jinkela_wire_691)
    );

    and_bb _0625_ (
        .b(jinkela_wire_717),
        .a(jinkela_wire_373),
        .c(jinkela_wire_649)
    );

    and_bb _0709_ (
        .b(jinkela_wire_658),
        .a(jinkela_wire_126),
        .c(jinkela_wire_599)
    );

    or_bb _0919_ (
        .b(jinkela_wire_262),
        .a(jinkela_wire_427),
        .c(b_23_)
    );

    or_bb _0500_ (
        .b(jinkela_wire_61),
        .a(jinkela_wire_297),
        .c(jinkela_wire_390)
    );

    and_bb _0542_ (
        .b(jinkela_wire_487),
        .a(jinkela_wire_305),
        .c(jinkela_wire_801)
    );

    or_bb _0626_ (
        .b(jinkela_wire_517),
        .a(jinkela_wire_799),
        .c(jinkela_wire_816)
    );

    or_bb _0710_ (
        .b(jinkela_wire_245),
        .a(jinkela_wire_589),
        .c(jinkela_wire_704)
    );

    maj_bbb _0920_ (
        .c(jinkela_wire_284),
        .b(jinkela_wire_796),
        .a(jinkela_wire_262),
        .d(b_22_)
    );

    and_bb _0501_ (
        .b(jinkela_wire_61),
        .a(jinkela_wire_297),
        .c(jinkela_wire_371)
    );

    and_bb _0543_ (
        .b(jinkela_wire_529),
        .a(jinkela_wire_801),
        .c(jinkela_wire_531)
    );

    and_bb _0627_ (
        .b(jinkela_wire_517),
        .a(jinkela_wire_799),
        .c(jinkela_wire_542)
    );

    and_bb _0711_ (
        .b(jinkela_wire_245),
        .a(jinkela_wire_589),
        .c(jinkela_wire_351)
    );

    and_bb _0921_ (
        .b(jinkela_wire_284),
        .a(jinkela_wire_796),
        .c(jinkela_wire_524)
    );

    or_bb _0502_ (
        .b(jinkela_wire_134),
        .a(jinkela_wire_661),
        .c(jinkela_wire_289)
    );

    or_bb _0544_ (
        .b(jinkela_wire_190),
        .a(jinkela_wire_604),
        .c(jinkela_wire_488)
    );

    or_bb _0628_ (
        .b(jinkela_wire_35),
        .a(jinkela_wire_398),
        .c(jinkela_wire_410)
    );

    or_bb _0712_ (
        .b(jinkela_wire_746),
        .a(jinkela_wire_813),
        .c(jinkela_wire_734)
    );

    and_bb _0922_ (
        .b(jinkela_wire_262),
        .a(jinkela_wire_524),
        .c(b_21_)
    );

    and_bb _0503_ (
        .b(jinkela_wire_134),
        .a(jinkela_wire_661),
        .c(jinkela_wire_546)
    );

    or_bb _0504_ (
        .b(jinkela_wire_495),
        .a(jinkela_wire_30),
        .c(jinkela_wire_10)
    );

endmodule
