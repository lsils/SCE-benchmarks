module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( in_15_ , in_0_ , in_4_ , in_29_ , in_38_ , in_53_ , in_42_ , in_11_ , in_59_ , in_48_ , in_54_ , in_16_ , in_43_ , in_37_ , in_61_ , in_14_ , in_62_ , in_60_ , in_40_ , in_5_ , in_28_ , in_7_ , in_6_ , in_34_ , in_57_ , in_3_ , in_56_ , in_45_ , in_10_ , in_27_ , in_21_ , in_25_ , in_22_ , in_12_ , in_58_ , in_36_ , in_51_ , in_18_ , in_9_ , in_39_ , in_24_ , in_26_ , in_8_ , in_41_ , in_55_ , in_2_ , in_49_ , in_19_ , in_35_ , in_50_ , in_32_ , in_30_ , in_33_ , in_17_ , in_31_ , in_44_ , in_1_ , in_23_ , in_52_ , in_20_ , in_46_ , in_13_ , in_63_ , in_47_ , out_1_ , out_3_ , out_6_ , out_2_ , out_0_ , out_4_ , out_5_ );
  input in_15_ , in_0_ , in_4_ , in_29_ , in_38_ , in_53_ , in_42_ , in_11_ , in_59_ , in_48_ , in_54_ , in_16_ , in_43_ , in_37_ , in_61_ , in_14_ , in_62_ , in_60_ , in_40_ , in_5_ , in_28_ , in_7_ , in_6_ , in_34_ , in_57_ , in_3_ , in_56_ , in_45_ , in_10_ , in_27_ , in_21_ , in_25_ , in_22_ , in_12_ , in_58_ , in_36_ , in_51_ , in_18_ , in_9_ , in_39_ , in_24_ , in_26_ , in_8_ , in_41_ , in_55_ , in_2_ , in_49_ , in_19_ , in_35_ , in_50_ , in_32_ , in_30_ , in_33_ , in_17_ , in_31_ , in_44_ , in_1_ , in_23_ , in_52_ , in_20_ , in_46_ , in_13_ , in_63_ , in_47_ ;
  output out_1_ , out_3_ , out_6_ , out_2_ , out_0_ , out_4_ , out_5_ ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 ;
  assign n65 = in_15_ & in_14_ ;
  buffer buf_n66( .i (n65), .o (n66) );
  assign n67 = in_12_ | in_13_ ;
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  assign n71 = in_4_ | in_5_ ;
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  assign n75 = in_0_ | in_1_ ;
  buffer buf_n76( .i (n75), .o (n76) );
  assign n77 = in_3_ & in_2_ ;
  buffer buf_n78( .i (n77), .o (n78) );
  assign n79 = ( n72 & n76 ) | ( n72 & n78 ) | ( n76 & n78 ) ;
  buffer buf_n80( .i (n79), .o (n80) );
  assign n85 = ( ~n72 & n76 ) | ( ~n72 & n78 ) | ( n76 & n78 ) ;
  buffer buf_n86( .i (n85), .o (n86) );
  assign n87 = ( n74 & ~n80 ) | ( n74 & n86 ) | ( ~n80 & n86 ) ;
  buffer buf_n88( .i (n87), .o (n88) );
  assign n89 = in_11_ & in_10_ ;
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  assign n93 = in_7_ & in_6_ ;
  buffer buf_n94( .i (n93), .o (n94) );
  assign n95 = in_9_ | in_8_ ;
  buffer buf_n96( .i (n95), .o (n96) );
  assign n97 = ( n90 & n94 ) | ( n90 & n96 ) | ( n94 & n96 ) ;
  buffer buf_n98( .i (n97), .o (n98) );
  assign n103 = ( ~n90 & n94 ) | ( ~n90 & n96 ) | ( n94 & n96 ) ;
  buffer buf_n104( .i (n103), .o (n104) );
  assign n105 = ( n92 & ~n98 ) | ( n92 & n104 ) | ( ~n98 & n104 ) ;
  buffer buf_n106( .i (n105), .o (n106) );
  assign n107 = ( n68 & n88 ) | ( n68 & n106 ) | ( n88 & n106 ) ;
  buffer buf_n108( .i (n107), .o (n108) );
  assign n111 = ( ~n68 & n88 ) | ( ~n68 & n106 ) | ( n88 & n106 ) ;
  buffer buf_n112( .i (n111), .o (n112) );
  assign n113 = ( n70 & ~n108 ) | ( n70 & n112 ) | ( ~n108 & n112 ) ;
  buffer buf_n114( .i (n113), .o (n114) );
  assign n115 = n66 & n114 ;
  buffer buf_n116( .i (n115), .o (n116) );
  assign n117 = n66 | n114 ;
  buffer buf_n118( .i (n117), .o (n118) );
  assign n119 = ~n116 & n118 ;
  buffer buf_n120( .i (n119), .o (n120) );
  assign n121 = in_30_ & in_31_ ;
  buffer buf_n122( .i (n121), .o (n122) );
  assign n123 = in_29_ | in_28_ ;
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  assign n127 = in_21_ | in_20_ ;
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  assign n131 = in_16_ | in_17_ ;
  buffer buf_n132( .i (n131), .o (n132) );
  assign n133 = in_18_ & in_19_ ;
  buffer buf_n134( .i (n133), .o (n134) );
  assign n135 = ( n128 & n132 ) | ( n128 & n134 ) | ( n132 & n134 ) ;
  buffer buf_n136( .i (n135), .o (n136) );
  assign n141 = ( ~n128 & n132 ) | ( ~n128 & n134 ) | ( n132 & n134 ) ;
  buffer buf_n142( .i (n141), .o (n142) );
  assign n143 = ( n130 & ~n136 ) | ( n130 & n142 ) | ( ~n136 & n142 ) ;
  buffer buf_n144( .i (n143), .o (n144) );
  assign n145 = in_27_ & in_26_ ;
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  assign n149 = in_22_ & in_23_ ;
  buffer buf_n150( .i (n149), .o (n150) );
  assign n151 = in_25_ | in_24_ ;
  buffer buf_n152( .i (n151), .o (n152) );
  assign n153 = ( n146 & n150 ) | ( n146 & n152 ) | ( n150 & n152 ) ;
  buffer buf_n154( .i (n153), .o (n154) );
  assign n159 = ( ~n146 & n150 ) | ( ~n146 & n152 ) | ( n150 & n152 ) ;
  buffer buf_n160( .i (n159), .o (n160) );
  assign n161 = ( n148 & ~n154 ) | ( n148 & n160 ) | ( ~n154 & n160 ) ;
  buffer buf_n162( .i (n161), .o (n162) );
  assign n163 = ( n124 & n144 ) | ( n124 & n162 ) | ( n144 & n162 ) ;
  buffer buf_n164( .i (n163), .o (n164) );
  assign n167 = ( ~n124 & n144 ) | ( ~n124 & n162 ) | ( n144 & n162 ) ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = ( n126 & ~n164 ) | ( n126 & n168 ) | ( ~n164 & n168 ) ;
  buffer buf_n170( .i (n169), .o (n170) );
  assign n171 = n122 & n170 ;
  buffer buf_n172( .i (n171), .o (n172) );
  assign n173 = n122 | n170 ;
  buffer buf_n174( .i (n173), .o (n174) );
  assign n175 = ~n172 & n174 ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n177 = n120 & n176 ;
  buffer buf_n178( .i (n177), .o (n178) );
  assign n182 = n120 | n176 ;
  buffer buf_n183( .i (n182), .o (n183) );
  assign n184 = ~n178 & n183 ;
  buffer buf_n185( .i (n184), .o (n185) );
  assign n186 = in_46_ & in_47_ ;
  buffer buf_n187( .i (n186), .o (n187) );
  assign n188 = in_45_ | in_44_ ;
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  assign n192 = in_37_ | in_36_ ;
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  assign n196 = in_32_ | in_33_ ;
  buffer buf_n197( .i (n196), .o (n197) );
  assign n198 = in_34_ & in_35_ ;
  buffer buf_n199( .i (n198), .o (n199) );
  assign n200 = ( n193 & n197 ) | ( n193 & n199 ) | ( n197 & n199 ) ;
  buffer buf_n201( .i (n200), .o (n201) );
  assign n206 = ( ~n193 & n197 ) | ( ~n193 & n199 ) | ( n197 & n199 ) ;
  buffer buf_n207( .i (n206), .o (n207) );
  assign n208 = ( n195 & ~n201 ) | ( n195 & n207 ) | ( ~n201 & n207 ) ;
  buffer buf_n209( .i (n208), .o (n209) );
  assign n210 = in_42_ & in_43_ ;
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  assign n214 = in_38_ & in_39_ ;
  buffer buf_n215( .i (n214), .o (n215) );
  assign n216 = in_40_ | in_41_ ;
  buffer buf_n217( .i (n216), .o (n217) );
  assign n218 = ( n211 & n215 ) | ( n211 & n217 ) | ( n215 & n217 ) ;
  buffer buf_n219( .i (n218), .o (n219) );
  assign n224 = ( ~n211 & n215 ) | ( ~n211 & n217 ) | ( n215 & n217 ) ;
  buffer buf_n225( .i (n224), .o (n225) );
  assign n226 = ( n213 & ~n219 ) | ( n213 & n225 ) | ( ~n219 & n225 ) ;
  buffer buf_n227( .i (n226), .o (n227) );
  assign n228 = ( n189 & n209 ) | ( n189 & n227 ) | ( n209 & n227 ) ;
  buffer buf_n229( .i (n228), .o (n229) );
  assign n232 = ( ~n189 & n209 ) | ( ~n189 & n227 ) | ( n209 & n227 ) ;
  buffer buf_n233( .i (n232), .o (n233) );
  assign n234 = ( n191 & ~n229 ) | ( n191 & n233 ) | ( ~n229 & n233 ) ;
  buffer buf_n235( .i (n234), .o (n235) );
  assign n236 = n187 & n235 ;
  buffer buf_n237( .i (n236), .o (n237) );
  assign n238 = n187 | n235 ;
  buffer buf_n239( .i (n238), .o (n239) );
  assign n240 = ~n237 & n239 ;
  buffer buf_n241( .i (n240), .o (n241) );
  assign n242 = in_62_ & in_63_ ;
  buffer buf_n243( .i (n242), .o (n243) );
  assign n244 = in_61_ | in_60_ ;
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  assign n248 = in_53_ | in_52_ ;
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  assign n252 = in_48_ | in_49_ ;
  buffer buf_n253( .i (n252), .o (n253) );
  assign n254 = in_51_ & in_50_ ;
  buffer buf_n255( .i (n254), .o (n255) );
  assign n256 = ( n249 & n253 ) | ( n249 & n255 ) | ( n253 & n255 ) ;
  buffer buf_n257( .i (n256), .o (n257) );
  assign n262 = ( ~n249 & n253 ) | ( ~n249 & n255 ) | ( n253 & n255 ) ;
  buffer buf_n263( .i (n262), .o (n263) );
  assign n264 = ( n251 & ~n257 ) | ( n251 & n263 ) | ( ~n257 & n263 ) ;
  buffer buf_n265( .i (n264), .o (n265) );
  assign n266 = in_59_ & in_58_ ;
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  assign n270 = in_54_ & in_55_ ;
  buffer buf_n271( .i (n270), .o (n271) );
  assign n272 = in_57_ | in_56_ ;
  buffer buf_n273( .i (n272), .o (n273) );
  assign n274 = ( n267 & n271 ) | ( n267 & n273 ) | ( n271 & n273 ) ;
  buffer buf_n275( .i (n274), .o (n275) );
  assign n280 = ( ~n267 & n271 ) | ( ~n267 & n273 ) | ( n271 & n273 ) ;
  buffer buf_n281( .i (n280), .o (n281) );
  assign n282 = ( n269 & ~n275 ) | ( n269 & n281 ) | ( ~n275 & n281 ) ;
  buffer buf_n283( .i (n282), .o (n283) );
  assign n284 = ( n245 & n265 ) | ( n245 & n283 ) | ( n265 & n283 ) ;
  buffer buf_n285( .i (n284), .o (n285) );
  assign n288 = ( ~n245 & n265 ) | ( ~n245 & n283 ) | ( n265 & n283 ) ;
  buffer buf_n289( .i (n288), .o (n289) );
  assign n290 = ( n247 & ~n285 ) | ( n247 & n289 ) | ( ~n285 & n289 ) ;
  buffer buf_n291( .i (n290), .o (n291) );
  assign n292 = n243 | n291 ;
  buffer buf_n293( .i (n292), .o (n293) );
  assign n294 = n243 & n291 ;
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = n293 & ~n295 ;
  buffer buf_n297( .i (n296), .o (n297) );
  assign n298 = n241 & n297 ;
  buffer buf_n299( .i (n298), .o (n299) );
  assign n303 = n241 | n297 ;
  buffer buf_n304( .i (n303), .o (n304) );
  assign n305 = ~n299 & n304 ;
  buffer buf_n306( .i (n305), .o (n306) );
  assign n307 = n185 & n306 ;
  buffer buf_n308( .i (n307), .o (n308) );
  assign n314 = n185 | n306 ;
  buffer buf_n315( .i (n314), .o (n315) );
  assign n316 = ~n308 & n315 ;
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  assign n317 = ( n84 & n102 ) | ( n84 & n108 ) | ( n102 & n108 ) ;
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  assign n323 = ( n84 & n102 ) | ( n84 & ~n108 ) | ( n102 & ~n108 ) ;
  buffer buf_n324( .i (n323), .o (n324) );
  assign n325 = ( n110 & ~n318 ) | ( n110 & n324 ) | ( ~n318 & n324 ) ;
  buffer buf_n326( .i (n325), .o (n326) );
  assign n327 = n116 & n326 ;
  buffer buf_n328( .i (n327), .o (n328) );
  assign n329 = n322 & n328 ;
  buffer buf_n330( .i (n329), .o (n330) );
  assign n335 = n322 | n328 ;
  buffer buf_n336( .i (n335), .o (n336) );
  assign n337 = ~n330 & n336 ;
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  assign n339 = ( n140 & n158 ) | ( n140 & n164 ) | ( n158 & n164 ) ;
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  assign n345 = ( n140 & n158 ) | ( n140 & ~n164 ) | ( n158 & ~n164 ) ;
  buffer buf_n346( .i (n345), .o (n346) );
  assign n347 = ( n166 & ~n340 ) | ( n166 & n346 ) | ( ~n340 & n346 ) ;
  buffer buf_n348( .i (n347), .o (n348) );
  assign n349 = n172 & n348 ;
  buffer buf_n350( .i (n349), .o (n350) );
  assign n351 = n344 & n350 ;
  buffer buf_n352( .i (n351), .o (n352) );
  assign n357 = n344 | n350 ;
  buffer buf_n358( .i (n357), .o (n358) );
  assign n359 = ~n352 & n358 ;
  buffer buf_n360( .i (n359), .o (n360) );
  assign n361 = n338 & n360 ;
  assign n362 = n338 | n360 ;
  assign n363 = ~n361 & n362 ;
  buffer buf_n364( .i (n363), .o (n364) );
  assign n365 = n116 | n326 ;
  buffer buf_n366( .i (n365), .o (n366) );
  assign n367 = ~n328 & n366 ;
  buffer buf_n368( .i (n367), .o (n368) );
  assign n369 = n172 | n348 ;
  buffer buf_n370( .i (n369), .o (n370) );
  assign n371 = ~n350 & n370 ;
  buffer buf_n372( .i (n371), .o (n372) );
  assign n373 = ( n178 & n368 ) | ( n178 & n372 ) | ( n368 & n372 ) ;
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  assign n378 = n364 & n377 ;
  assign n379 = n364 | n377 ;
  assign n380 = ~n378 & n379 ;
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  assign n382 = ( n205 & n223 ) | ( n205 & n229 ) | ( n223 & n229 ) ;
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  assign n388 = ( n205 & n223 ) | ( n205 & ~n229 ) | ( n223 & ~n229 ) ;
  buffer buf_n389( .i (n388), .o (n389) );
  assign n390 = ( n231 & ~n383 ) | ( n231 & n389 ) | ( ~n383 & n389 ) ;
  buffer buf_n391( .i (n390), .o (n391) );
  assign n392 = n237 & n391 ;
  buffer buf_n393( .i (n392), .o (n393) );
  assign n394 = n387 & n393 ;
  buffer buf_n395( .i (n394), .o (n395) );
  assign n400 = n387 | n393 ;
  buffer buf_n401( .i (n400), .o (n401) );
  assign n402 = ~n395 & n401 ;
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  assign n404 = ( n261 & n279 ) | ( n261 & n285 ) | ( n279 & n285 ) ;
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  assign n410 = ( n261 & n279 ) | ( n261 & ~n285 ) | ( n279 & ~n285 ) ;
  buffer buf_n411( .i (n410), .o (n411) );
  assign n412 = ( n287 & ~n405 ) | ( n287 & n411 ) | ( ~n405 & n411 ) ;
  buffer buf_n413( .i (n412), .o (n413) );
  assign n414 = n295 & n413 ;
  buffer buf_n415( .i (n414), .o (n415) );
  assign n416 = n409 & n415 ;
  buffer buf_n417( .i (n416), .o (n417) );
  assign n422 = n409 | n415 ;
  buffer buf_n423( .i (n422), .o (n423) );
  assign n424 = ~n417 & n423 ;
  buffer buf_n425( .i (n424), .o (n425) );
  assign n426 = n403 & n425 ;
  assign n427 = n403 | n425 ;
  assign n428 = ~n426 & n427 ;
  buffer buf_n429( .i (n428), .o (n429) );
  assign n430 = n237 | n391 ;
  buffer buf_n431( .i (n430), .o (n431) );
  assign n432 = ~n393 & n431 ;
  buffer buf_n433( .i (n432), .o (n433) );
  assign n434 = n295 | n413 ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n436 = ~n415 & n435 ;
  buffer buf_n437( .i (n436), .o (n437) );
  assign n438 = ( n299 & n433 ) | ( n299 & n437 ) | ( n433 & n437 ) ;
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  assign n443 = n429 & n442 ;
  assign n444 = n429 | n442 ;
  assign n445 = ~n443 & n444 ;
  buffer buf_n446( .i (n445), .o (n446) );
  assign n447 = n381 & n446 ;
  assign n448 = n381 | n446 ;
  assign n449 = ~n447 & n448 ;
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  assign n451 = n368 & n372 ;
  assign n452 = n368 | n372 ;
  assign n453 = ~n451 & n452 ;
  buffer buf_n454( .i (n453), .o (n454) );
  assign n455 = n181 & n454 ;
  assign n456 = n181 | n454 ;
  assign n457 = ~n455 & n456 ;
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  assign n459 = n433 & n437 ;
  assign n460 = n433 | n437 ;
  assign n461 = ~n459 & n460 ;
  buffer buf_n462( .i (n461), .o (n462) );
  assign n463 = n302 & n462 ;
  assign n464 = n302 | n462 ;
  assign n465 = ~n463 & n464 ;
  buffer buf_n466( .i (n465), .o (n466) );
  assign n467 = ( n310 & n458 ) | ( n310 & n466 ) | ( n458 & n466 ) ;
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  assign n472 = n450 & n471 ;
  assign n473 = n450 | n471 ;
  assign n474 = ~n472 & n473 ;
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  assign n475 = ( n338 & n360 ) | ( n338 & n374 ) | ( n360 & n374 ) ;
  buffer buf_n476( .i (n475), .o (n476) );
  assign n477 = ( n334 & n356 ) | ( n334 & n476 ) | ( n356 & n476 ) ;
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  assign n485 = ( n403 & n425 ) | ( n403 & n439 ) | ( n425 & n439 ) ;
  buffer buf_n486( .i (n485), .o (n486) );
  assign n487 = ( n399 & n421 ) | ( n399 & n486 ) | ( n421 & n486 ) ;
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  assign n495 = n330 & n352 ;
  assign n496 = n330 | n352 ;
  assign n497 = ~n495 & n496 ;
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  assign n500 = n476 & n499 ;
  assign n501 = n476 | n499 ;
  assign n502 = ~n500 & n501 ;
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  assign n507 = n395 & n417 ;
  assign n508 = n395 | n417 ;
  assign n509 = ~n507 & n508 ;
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  assign n512 = n486 & n511 ;
  assign n513 = n486 | n511 ;
  assign n514 = ~n512 & n513 ;
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  assign n519 = ( n381 & n446 ) | ( n381 & n468 ) | ( n446 & n468 ) ;
  buffer buf_n520( .i (n519), .o (n520) );
  assign n521 = ( n506 & n518 ) | ( n506 & n520 ) | ( n518 & n520 ) ;
  buffer buf_n522( .i (n521), .o (n522) );
  assign n523 = ( n484 & n494 ) | ( n484 & n522 ) | ( n494 & n522 ) ;
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  assign n524 = n458 & n466 ;
  assign n525 = n458 | n466 ;
  assign n526 = ~n524 & n525 ;
  buffer buf_n527( .i (n526), .o (n527) );
  assign n528 = n313 & n527 ;
  assign n529 = n313 | n527 ;
  assign n530 = ~n528 & n529 ;
  assign n531 = n503 & n515 ;
  assign n532 = n503 | n515 ;
  assign n533 = ~n531 & n532 ;
  buffer buf_n534( .i (n533), .o (n534) );
  assign n535 = n520 & n534 ;
  assign n536 = n520 | n534 ;
  assign n537 = ~n535 & n536 ;
  assign n538 = n478 & n488 ;
  assign n539 = n478 | n488 ;
  assign n540 = ~n538 & n539 ;
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  assign n545 = n522 & n544 ;
  assign n546 = n522 | n544 ;
  assign n547 = ~n545 & n546 ;
  assign out_1_ = n316 ;
  assign out_3_ = n474 ;
  assign out_6_ = n523 ;
  assign out_2_ = n530 ;
  assign out_0_ = 1'b0 ;
  assign out_4_ = n537 ;
  assign out_5_ = n547 ;
endmodule
