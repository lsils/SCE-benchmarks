module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G158 , G159 , G16 , G160 , G161 , G162 , G163 , G164 , G165 , G166 , G167 , G168 , G169 , G17 , G170 , G171 , G172 , G173 , G174 , G175 , G176 , G177 , G178 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 , G5193 , G5194 , G5195 , G5196 , G5197 , G5198 , G5199 , G5200 , G5201 , G5202 , G5203 , G5204 , G5205 , G5206 , G5207 , G5208 , G5209 , G5210 , G5211 , G5212 , G5213 , G5214 , G5215 , G5216 , G5217 , G5218 , G5219 , G5220 , G5221 , G5222 , G5223 , G5224 , G5225 , G5226 , G5227 , G5228 , G5229 , G5230 , G5231 , G5232 , G5233 , G5234 , G5235 , G5236 , G5237 , G5238 , G5239 , G5240 , G5241 , G5242 , G5243 , G5244 , G5245 , G5246 , G5247 , G5248 , G5249 , G5250 , G5251 , G5252 , G5253 , G5254 , G5255 , G5256 , G5257 , G5258 , G5259 , G5260 , G5261 , G5262 , G5263 , G5264 , G5265 , G5266 , G5267 , G5268 , G5269 , G5270 , G5271 , G5272 , G5273 , G5274 , G5275 , G5276 , G5277 , G5278 , G5279 , G5280 , G5281 , G5282 , G5283 , G5284 , G5285 , G5286 , G5287 , G5288 , G5289 , G5290 , G5291 , G5292 , G5293 , G5294 , G5295 , G5296 , G5297 , G5298 , G5299 , G5300 , G5301 , G5302 , G5303 , G5304 , G5305 , G5306 , G5307 , G5308 , G5309 , G5310 , G5311 , G5312 , G5313 , G5314 , G5315 );
  input G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G158 , G159 , G16 , G160 , G161 , G162 , G163 , G164 , G165 , G166 , G167 , G168 , G169 , G17 , G170 , G171 , G172 , G173 , G174 , G175 , G176 , G177 , G178 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 ;
  output G5193 , G5194 , G5195 , G5196 , G5197 , G5198 , G5199 , G5200 , G5201 , G5202 , G5203 , G5204 , G5205 , G5206 , G5207 , G5208 , G5209 , G5210 , G5211 , G5212 , G5213 , G5214 , G5215 , G5216 , G5217 , G5218 , G5219 , G5220 , G5221 , G5222 , G5223 , G5224 , G5225 , G5226 , G5227 , G5228 , G5229 , G5230 , G5231 , G5232 , G5233 , G5234 , G5235 , G5236 , G5237 , G5238 , G5239 , G5240 , G5241 , G5242 , G5243 , G5244 , G5245 , G5246 , G5247 , G5248 , G5249 , G5250 , G5251 , G5252 , G5253 , G5254 , G5255 , G5256 , G5257 , G5258 , G5259 , G5260 , G5261 , G5262 , G5263 , G5264 , G5265 , G5266 , G5267 , G5268 , G5269 , G5270 , G5271 , G5272 , G5273 , G5274 , G5275 , G5276 , G5277 , G5278 , G5279 , G5280 , G5281 , G5282 , G5283 , G5284 , G5285 , G5286 , G5287 , G5288 , G5289 , G5290 , G5291 , G5292 , G5293 , G5294 , G5295 , G5296 , G5297 , G5298 , G5299 , G5300 , G5301 , G5302 , G5303 , G5304 , G5305 , G5306 , G5307 , G5308 , G5309 , G5310 , G5311 , G5312 , G5313 , G5314 , G5315 ;
  wire n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 ;
  buffer buf_n847( .i (G66), .o (n847) );
  inverter inv_n3898( .i (n847), .o (n3898) );
  buffer buf_n287( .i (G113), .o (n287) );
  inverter inv_n3899( .i (n287), .o (n3899) );
  buffer buf_n766( .i (G165), .o (n766) );
  inverter inv_n3900( .i (n766), .o (n3900) );
  inverter inv_n736( .i (G151), .o (n736) );
  buffer buf_n444( .i (G127), .o (n444) );
  inverter inv_n3901( .i (n444), .o (n3901) );
  buffer buf_n487( .i (G131), .o (n487) );
  inverter inv_n3902( .i (n487), .o (n3902) );
  buffer buf_n738( .i (G153), .o (n738) );
  buffer buf_n740( .i (G156), .o (n740) );
  assign n998 = n738 & n740 ;
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n737( .i (G152), .o (n737) );
  inverter inv_n3903( .i (n737), .o (n3903) );
  buffer buf_n406( .i (G125), .o (n406) );
  inverter inv_n3904( .i (n406), .o (n3904) );
  buffer buf_n468( .i (G129), .o (n468) );
  inverter inv_n3905( .i (n468), .o (n3905) );
  buffer buf_n848( .i (n847), .o (n848) );
  assign n1000 = G67 & n848 ;
  buffer buf_n997( .i (G99), .o (n997) );
  inverter inv_n3906( .i (n997), .o (n3906) );
  inverter inv_n3907( .i (n738), .o (n3907) );
  inverter inv_n3908( .i (n740), .o (n3908) );
  buffer buf_n739( .i (G155), .o (n739) );
  inverter inv_n3909( .i (n739), .o (n3909) );
  buffer buf_n179( .i (G1), .o (n179) );
  assign n1001 = G134 & n179 ;
  assign n1002 = G63 & ~n766 ;
  buffer buf_n279( .i (G11), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  assign n1003 = G164 | ~n284 ;
  assign n1004 = G136 & G154 ;
  buffer buf_n1005( .i (n1004), .o (n1005) );
  inverter inv_n3910( .i (n1005), .o (n3910) );
  buffer buf_n844( .i (G64), .o (n844) );
  buffer buf_n299( .i (G114), .o (n299) );
  assign n1006 = G12 & n279 ;
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  assign n1011 = ~G65 | ~n1010 ;
  inverter inv_n3913( .i (n1007), .o (n3913) );
  inverter inv_n3911( .i (n179), .o (n3911) );
  inverter inv_n3912( .i (n299), .o (n3912) );
  buffer buf_n763( .i (G163), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  assign n1012 = G34 & n765 ;
  assign n1013 = G33 & ~n765 ;
  assign n1014 = n1012 | n1013 ;
  assign n1015 = ~n1010 | ~n1014 ;
  assign n1016 = G13 & n764 ;
  assign n1017 = G35 & ~n764 ;
  assign n1018 = n1016 | n1017 ;
  assign n1019 = n1009 & n1018 ;
  inverter inv_n1020( .i (n1019), .o (n1020) );
  assign n1021 = ~G32 | ~n1010 ;
  assign n1022 = G9 & ~n765 ;
  assign n1023 = G8 & n764 ;
  assign n1024 = n1008 & ~n1023 ;
  assign n1025 = ~n1022 & n1024 ;
  assign n1026 = n848 & ~n1025 ;
  assign n1027 = G30 & ~n765 ;
  buffer buf_n1028( .i (n763), .o (n1028) );
  assign n1029 = G10 & n1028 ;
  assign n1030 = n1008 & ~n1029 ;
  assign n1031 = ~n1027 & n1030 ;
  assign n1032 = n848 & ~n1031 ;
  buffer buf_n1033( .i (n1028), .o (n1033) );
  assign n1034 = G7 & ~n1033 ;
  assign n1035 = G28 & n1028 ;
  assign n1036 = n1008 & ~n1035 ;
  assign n1037 = ~n1034 & n1036 ;
  assign n1038 = n848 & ~n1037 ;
  assign n1039 = G29 & ~n1033 ;
  assign n1040 = G31 & n1028 ;
  buffer buf_n1041( .i (n1007), .o (n1041) );
  assign n1042 = ~n1040 & n1041 ;
  assign n1043 = ~n1039 & n1042 ;
  buffer buf_n1044( .i (n847), .o (n1044) );
  assign n1045 = ~n1043 & n1044 ;
  buffer buf_n665( .i (G145), .o (n665) );
  buffer buf_n180( .i (G100), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n311( .i (G117), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  assign n1046 = n181 | n312 ;
  buffer buf_n184( .i (G101), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  assign n1047 = ~n185 & n312 ;
  assign n1048 = n1046 & ~n1047 ;
  assign n1049 = n665 & ~n1048 ;
  buffer buf_n188( .i (G102), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  assign n1050 = n189 & n312 ;
  buffer buf_n993( .i (G98), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n1051( .i (n311), .o (n1051) );
  assign n1052 = n994 & ~n1051 ;
  assign n1053 = n1050 | n1052 ;
  assign n1054 = ~n665 & n1053 ;
  assign n1055 = n1049 | n1054 ;
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n668( .i (G146), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n325( .i (G119), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  assign n1066 = n181 | n328 ;
  assign n1067 = ~n185 & n328 ;
  assign n1068 = n1066 & ~n1067 ;
  assign n1069 = n670 & ~n1068 ;
  assign n1070 = n189 & n328 ;
  buffer buf_n1071( .i (n327), .o (n1071) );
  assign n1072 = n994 & ~n1071 ;
  assign n1073 = n1070 | n1072 ;
  assign n1074 = ~n670 & n1073 ;
  assign n1075 = n1069 | n1074 ;
  buffer buf_n1076( .i (n1075), .o (n1076) );
  assign n1086 = n1056 & n1076 ;
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n717( .i (G150), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n445( .i (G128), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n776( .i (G169), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  assign n1097 = n464 | n777 ;
  buffer buf_n773( .i (G168), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  assign n1098 = n464 & ~n774 ;
  assign n1099 = n1097 & ~n1098 ;
  assign n1100 = n735 & ~n1099 ;
  buffer buf_n770( .i (G167), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  assign n1101 = n464 & n771 ;
  buffer buf_n767( .i (G166), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n1102( .i (n463), .o (n1102) );
  assign n1103 = n768 & ~n1102 ;
  assign n1104 = n1101 | n1103 ;
  assign n1105 = ~n735 & n1104 ;
  assign n1106 = n1100 | n1105 ;
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  assign n1108 = n288 | n996 ;
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  assign n1109 = ~n191 & n288 ;
  assign n1110 = n1108 & ~n1109 ;
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n300( .i (G115), .o (n300) );
  assign n1127 = n183 | n300 ;
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  assign n1128 = ~n187 & n300 ;
  assign n1129 = n1127 & ~n1128 ;
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n1141 = n1111 & ~n1130 ;
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n469( .i (G130), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  assign n1149 = n181 | n477 ;
  assign n1150 = ~n185 & n477 ;
  assign n1151 = n1149 & ~n1150 ;
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n686( .i (G148), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  assign n1165 = ~n698 & n768 ;
  assign n1166 = n698 & ~n777 ;
  assign n1167 = n1165 | n1166 ;
  buffer buf_n1168( .i (n1167), .o (n1168) );
  assign n1169 = ~n1161 & n1168 ;
  assign n1170 = n1148 & n1169 ;
  assign n1171 = n1107 & n1170 ;
  buffer buf_n671( .i (G147), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n341( .i (G121), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  assign n1172 = n356 | n777 ;
  assign n1173 = n356 & ~n774 ;
  assign n1174 = n1172 & ~n1173 ;
  assign n1175 = n685 & ~n1174 ;
  assign n1176 = n356 & n771 ;
  buffer buf_n1177( .i (n355), .o (n1177) );
  assign n1178 = n768 & ~n1177 ;
  assign n1179 = n1176 | n1178 ;
  assign n1180 = ~n685 & n1179 ;
  assign n1181 = n1175 | n1180 ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n699( .i (G149), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n423( .i (G126), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n1183( .i (n776), .o (n1183) );
  assign n1184 = n440 | n1183 ;
  assign n1185 = n440 & ~n774 ;
  assign n1186 = n1184 & ~n1185 ;
  assign n1187 = n715 & ~n1186 ;
  assign n1188 = n440 & n771 ;
  buffer buf_n1189( .i (n439), .o (n1189) );
  buffer buf_n1190( .i (n767), .o (n1190) );
  assign n1191 = ~n1189 & n1190 ;
  assign n1192 = n1188 | n1191 ;
  assign n1193 = ~n715 & n1192 ;
  assign n1194 = n1187 | n1193 ;
  buffer buf_n1195( .i (n1194), .o (n1195) );
  assign n1196 = n1182 & n1195 ;
  assign n1197 = n1171 & n1196 ;
  assign n1198 = n1096 & n1197 ;
  buffer buf_n569( .i (G140), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n947( .i (G94), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  assign n1199 = n969 | n1183 ;
  buffer buf_n1200( .i (n773), .o (n1200) );
  assign n1201 = n969 & ~n1200 ;
  assign n1202 = n1199 & ~n1201 ;
  assign n1203 = n590 & ~n1202 ;
  buffer buf_n1204( .i (n770), .o (n1204) );
  assign n1205 = n969 & n1204 ;
  buffer buf_n1206( .i (n968), .o (n1206) );
  assign n1207 = n1190 & ~n1206 ;
  assign n1208 = n1205 | n1207 ;
  assign n1209 = ~n590 & n1208 ;
  assign n1210 = n1203 | n1209 ;
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n622( .i (G143), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n894( .i (G90), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  assign n1215 = n914 | n1183 ;
  assign n1216 = n914 & ~n1200 ;
  assign n1217 = n1215 & ~n1216 ;
  assign n1218 = n641 & ~n1217 ;
  assign n1219 = n914 & n1204 ;
  buffer buf_n1220( .i (n913), .o (n1220) );
  assign n1221 = n1190 & ~n1220 ;
  assign n1222 = n1219 | n1221 ;
  assign n1223 = ~n641 & n1222 ;
  assign n1224 = n1218 | n1223 ;
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n642( .i (G144), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n919( .i (G92), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  assign n1228 = n942 | n1183 ;
  assign n1229 = n942 & ~n1200 ;
  assign n1230 = n1228 & ~n1229 ;
  assign n1231 = n664 & ~n1230 ;
  assign n1232 = n942 & n1204 ;
  buffer buf_n1233( .i (n941), .o (n1233) );
  assign n1234 = n1190 & ~n1233 ;
  assign n1235 = n1232 | n1234 ;
  assign n1236 = ~n664 & n1235 ;
  assign n1237 = n1231 | n1236 ;
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  assign n1241 = n1227 & n1240 ;
  assign n1242 = n1214 & n1241 ;
  buffer buf_n491( .i (G135), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n258( .i (G109), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n778( .i (n777), .o (n778) );
  assign n1243 = n278 | n778 ;
  buffer buf_n775( .i (n774), .o (n775) );
  assign n1244 = n278 & ~n775 ;
  assign n1245 = n1243 & ~n1244 ;
  assign n1246 = n510 & ~n1245 ;
  buffer buf_n772( .i (n771), .o (n772) );
  assign n1247 = n278 & n772 ;
  buffer buf_n769( .i (n768), .o (n769) );
  assign n1248 = ~n278 & n769 ;
  assign n1249 = n1247 | n1248 ;
  assign n1250 = ~n510 & n1249 ;
  assign n1251 = n1246 | n1250 ;
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n591( .i (G141), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n974( .i (G96), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  assign n1254 = n778 | n992 ;
  assign n1255 = ~n775 & n992 ;
  assign n1256 = n1254 & ~n1255 ;
  assign n1257 = n608 & ~n1256 ;
  assign n1258 = n772 & n992 ;
  assign n1259 = n769 & ~n992 ;
  assign n1260 = n1258 | n1259 ;
  assign n1261 = ~n608 & n1260 ;
  assign n1262 = n1257 | n1261 ;
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  assign n1265 = n1253 & n1264 ;
  buffer buf_n548( .i (G139), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n234( .i (G107), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  assign n1266 = n254 | n778 ;
  assign n1267 = n254 & ~n775 ;
  assign n1268 = n1266 & ~n1267 ;
  assign n1269 = n567 & ~n1268 ;
  assign n1270 = n254 & n772 ;
  buffer buf_n1271( .i (n253), .o (n1271) );
  assign n1272 = n769 & ~n1271 ;
  assign n1273 = n1270 | n1272 ;
  assign n1274 = ~n567 & n1273 ;
  assign n1275 = n1269 | n1274 ;
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n609( .i (G142), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n869( .i (G88), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  assign n1277 = n187 | n882 ;
  assign n1278 = ~n183 & n882 ;
  assign n1279 = n1277 & ~n1278 ;
  assign n1280 = n621 & ~n1279 ;
  assign n1281 = n882 & n996 ;
  buffer buf_n1282( .i (n881), .o (n1282) );
  assign n1283 = n191 & ~n1282 ;
  assign n1284 = n1281 | n1283 ;
  assign n1285 = ~n621 & n1284 ;
  assign n1286 = n1280 | n1285 ;
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  assign n1297 = n1276 & n1295 ;
  buffer buf_n511( .i (G137), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n192( .i (G103), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  assign n1298 = n210 | n778 ;
  assign n1299 = n210 & ~n775 ;
  assign n1300 = n1298 & ~n1299 ;
  assign n1301 = n528 & ~n1300 ;
  assign n1302 = n210 & n772 ;
  assign n1303 = ~n210 & n769 ;
  assign n1304 = n1302 | n1303 ;
  assign n1305 = ~n528 & n1304 ;
  assign n1306 = n1301 | n1305 ;
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n529( .i (G138), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n211( .i (G105), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n1308( .i (n776), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  assign n1310 = n230 | n1309 ;
  buffer buf_n1311( .i (n1200), .o (n1311) );
  assign n1312 = n230 & ~n1311 ;
  assign n1313 = n1310 & ~n1312 ;
  assign n1314 = n547 & ~n1313 ;
  buffer buf_n1315( .i (n1204), .o (n1315) );
  assign n1316 = n230 & n1315 ;
  buffer buf_n1317( .i (n229), .o (n1317) );
  buffer buf_n1318( .i (n767), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  assign n1320 = ~n1317 & n1319 ;
  assign n1321 = n1316 | n1320 ;
  assign n1322 = ~n547 & n1321 ;
  assign n1323 = n1314 | n1322 ;
  buffer buf_n1324( .i (n1323), .o (n1324) );
  assign n1325 = n1307 & n1324 ;
  assign n1326 = n1297 & n1325 ;
  assign n1327 = n1265 & n1326 ;
  assign n1328 = n1242 & n1327 ;
  buffer buf_n382( .i (G124), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  assign n1329 = n388 & n974 ;
  assign n1330 = G97 & ~n388 ;
  assign n1331 = n1329 | n1330 ;
  buffer buf_n1332( .i (n1331), .o (n1332) );
  assign n1350 = n591 & n1332 ;
  buffer buf_n1351( .i (n1350), .o (n1351) );
  assign n1355 = n591 | n1332 ;
  buffer buf_n1356( .i (n1355), .o (n1356) );
  assign n1359 = ~n1351 & n1356 ;
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  assign n1368 = n258 & n386 ;
  assign n1369 = G110 & ~n386 ;
  assign n1370 = n1368 | n1369 ;
  buffer buf_n1371( .i (n1370), .o (n1371) );
  assign n1394 = n491 & n1371 ;
  buffer buf_n1395( .i (n1394), .o (n1395) );
  assign n1408 = n491 | n1371 ;
  buffer buf_n1409( .i (n1408), .o (n1409) );
  assign n1418 = ~n1395 & n1409 ;
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  assign n1436 = n234 & n386 ;
  buffer buf_n1437( .i (n385), .o (n1437) );
  assign n1438 = G108 & ~n1437 ;
  assign n1439 = n1436 | n1438 ;
  buffer buf_n1440( .i (n1439), .o (n1440) );
  assign n1463 = n548 | n1440 ;
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  assign n1473 = n548 & n1440 ;
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  assign n1491 = n1466 & ~n1476 ;
  buffer buf_n1492( .i (n1491), .o (n1492) );
  assign n1507 = n1421 & n1492 ;
  buffer buf_n1508( .i (n1507), .o (n1508) );
  assign n1511 = n211 & n387 ;
  assign n1512 = G106 & ~n387 ;
  assign n1513 = n1511 | n1512 ;
  buffer buf_n1514( .i (n1513), .o (n1514) );
  assign n1536 = n529 & n1514 ;
  buffer buf_n1537( .i (n1536), .o (n1537) );
  assign n1538 = n529 | n1514 ;
  buffer buf_n1539( .i (n1538), .o (n1539) );
  assign n1542 = ~n1537 & n1539 ;
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  assign n1559 = n192 & n388 ;
  buffer buf_n1560( .i (n387), .o (n1560) );
  assign n1561 = G104 & ~n1560 ;
  assign n1562 = n1559 | n1561 ;
  buffer buf_n1563( .i (n1562), .o (n1563) );
  assign n1584 = n511 | n1563 ;
  buffer buf_n1585( .i (n1584), .o (n1585) );
  assign n1590 = n511 & n1563 ;
  buffer buf_n1591( .i (n1590), .o (n1591) );
  assign n1597 = n1585 & ~n1591 ;
  buffer buf_n1598( .i (n1597), .o (n1598) );
  assign n1613 = n1544 & n1598 ;
  buffer buf_n1614( .i (n1613), .o (n1614) );
  assign n1623 = n1508 & n1614 ;
  buffer buf_n1624( .i (n1623), .o (n1624) );
  assign n1634 = n1364 & n1624 ;
  buffer buf_n1635( .i (n1634), .o (n1635) );
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n1637( .i (n1636), .o (n1637) );
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  assign n1644 = n385 & n869 ;
  assign n1645 = G89 & ~n385 ;
  assign n1646 = n1644 | n1645 ;
  buffer buf_n1647( .i (n1646), .o (n1647) );
  assign n1668 = n609 & n1647 ;
  buffer buf_n1669( .i (n1668), .o (n1669) );
  assign n1689 = n609 | n1647 ;
  buffer buf_n1690( .i (n1689), .o (n1690) );
  assign n1709 = ~n1669 & n1690 ;
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1729( .i (n384), .o (n1729) );
  assign n1730 = n894 & n1729 ;
  assign n1731 = G91 & ~n1729 ;
  assign n1732 = n1730 | n1731 ;
  buffer buf_n1733( .i (n1732), .o (n1733) );
  assign n1757 = n622 & n1733 ;
  buffer buf_n1758( .i (n1757), .o (n1758) );
  assign n1775 = n622 | n1733 ;
  buffer buf_n1776( .i (n1775), .o (n1776) );
  assign n1785 = ~n1758 & n1776 ;
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  assign n1803 = n382 & n919 ;
  assign n1804 = G93 & ~n382 ;
  assign n1805 = n1803 | n1804 ;
  buffer buf_n1806( .i (n1805), .o (n1806) );
  assign n1833 = n642 & n1806 ;
  buffer buf_n1834( .i (n1833), .o (n1834) );
  assign n1838 = n642 | n1806 ;
  buffer buf_n1839( .i (n1838), .o (n1839) );
  assign n1841 = ~n1834 & n1839 ;
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  assign n1862 = n383 & n947 ;
  assign n1863 = G95 & ~n383 ;
  assign n1864 = n1862 | n1863 ;
  buffer buf_n1865( .i (n1864), .o (n1865) );
  assign n1888 = n569 & n1865 ;
  buffer buf_n1889( .i (n1888), .o (n1889) );
  assign n1907 = n569 | n1865 ;
  buffer buf_n1908( .i (n1907), .o (n1908) );
  assign n1926 = ~n1889 & n1908 ;
  buffer buf_n1927( .i (n1926), .o (n1927) );
  assign n1946 = n1843 & n1927 ;
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  buffer buf_n1954( .i (n1953), .o (n1954) );
  buffer buf_n1955( .i (n1954), .o (n1955) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  buffer buf_n1960( .i (n1959), .o (n1960) );
  assign n1961 = n1799 & n1960 ;
  buffer buf_n1962( .i (n1961), .o (n1962) );
  assign n1963 = n1725 & n1962 ;
  buffer buf_n1964( .i (n1963), .o (n1964) );
  assign n1965 = n1643 & n1964 ;
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n360( .i (G123), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  assign n1967 = n365 | n406 ;
  buffer buf_n1968( .i (n1967), .o (n1968) );
  assign n1983 = n686 & n1968 ;
  buffer buf_n1984( .i (n1983), .o (n1984) );
  assign n1993 = n686 | n1968 ;
  buffer buf_n1994( .i (n1993), .o (n1994) );
  assign n2003 = ~n1984 & n1994 ;
  buffer buf_n2004( .i (n2003), .o (n2004) );
  assign n2014 = n360 & n445 ;
  assign n2015 = ~n360 & n468 ;
  assign n2016 = n2014 | n2015 ;
  buffer buf_n2017( .i (n2016), .o (n2017) );
  buffer buf_n2018( .i (n2017), .o (n2018) );
  buffer buf_n2019( .i (n2018), .o (n2019) );
  assign n2036 = n719 | n2019 ;
  buffer buf_n2037( .i (n2036), .o (n2037) );
  assign n2052 = n362 & n469 ;
  assign n2053 = ~n362 & n487 ;
  assign n2054 = n2052 | n2053 ;
  buffer buf_n2055( .i (n2054), .o (n2055) );
  assign n2075 = n717 & n2017 ;
  buffer buf_n2076( .i (n2075), .o (n2076) );
  assign n2093 = n2055 | n2076 ;
  buffer buf_n2094( .i (n2093), .o (n2094) );
  assign n2099 = n2037 & ~n2094 ;
  buffer buf_n2100( .i (n2099), .o (n2100) );
  assign n2115 = n362 & n423 ;
  buffer buf_n2116( .i (n361), .o (n2116) );
  assign n2117 = n444 & ~n2116 ;
  assign n2118 = n2115 | n2117 ;
  buffer buf_n2119( .i (n2118), .o (n2119) );
  assign n2136 = n699 & n2119 ;
  buffer buf_n2137( .i (n2136), .o (n2137) );
  assign n2140 = n699 | n2119 ;
  buffer buf_n2141( .i (n2140), .o (n2141) );
  assign n2143 = ~n2137 & n2141 ;
  buffer buf_n2144( .i (n2143), .o (n2144) );
  assign n2158 = n2100 & n2144 ;
  buffer buf_n2159( .i (n2158), .o (n2159) );
  assign n2164 = n2004 & n2159 ;
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n2166( .i (n2165), .o (n2166) );
  buffer buf_n2167( .i (n2166), .o (n2167) );
  buffer buf_n2168( .i (n2167), .o (n2168) );
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  buffer buf_n2171( .i (n2170), .o (n2171) );
  buffer buf_n2172( .i (n2171), .o (n2172) );
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n2175( .i (n2174), .o (n2175) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n2177), .o (n2178) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  assign n2179 = n311 & n369 ;
  assign n2180 = G118 & ~n369 ;
  assign n2181 = n2179 | n2180 ;
  buffer buf_n2182( .i (n2181), .o (n2182) );
  buffer buf_n2183( .i (n2182), .o (n2183) );
  assign n2186 = n666 & n2183 ;
  buffer buf_n2187( .i (n2186), .o (n2187) );
  buffer buf_n2188( .i (n2187), .o (n2188) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n2184( .i (n2183), .o (n2184) );
  assign n2193 = n667 | n2184 ;
  buffer buf_n2194( .i (n2193), .o (n2194) );
  assign n2198 = ~n2188 & n2194 ;
  buffer buf_n2199( .i (n2198), .o (n2199) );
  assign n2204 = n325 & n367 ;
  assign n2205 = G120 & ~n367 ;
  assign n2206 = n2204 | n2205 ;
  buffer buf_n2207( .i (n2206), .o (n2207) );
  assign n2222 = n668 & n2207 ;
  buffer buf_n2223( .i (n2222), .o (n2223) );
  assign n2231 = n668 | n2207 ;
  buffer buf_n2232( .i (n2231), .o (n2232) );
  assign n2240 = ~n2223 & n2232 ;
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  assign n2250 = n2199 & n2245 ;
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  assign n2257 = n287 & n371 ;
  assign n2258 = n299 & ~n371 ;
  assign n2259 = n2257 | n2258 ;
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  buffer buf_n2265( .i (n2264), .o (n2265) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  assign n2275 = n307 & n379 ;
  assign n2276 = G116 & ~n379 ;
  assign n2277 = n2275 | n2276 ;
  buffer buf_n2278( .i (n2277), .o (n2278) );
  assign n2281 = n2268 | n2278 ;
  buffer buf_n2282( .i (n2281), .o (n2282) );
  assign n2283 = G122 | n363 ;
  buffer buf_n2284( .i (n2283), .o (n2284) );
  assign n2301 = ~n341 & n364 ;
  assign n2302 = n2284 & ~n2301 ;
  buffer buf_n2303( .i (n2302), .o (n2303) );
  assign n2318 = n671 & n2303 ;
  buffer buf_n2319( .i (n2318), .o (n2319) );
  assign n2327 = n671 | n2303 ;
  buffer buf_n2328( .i (n2327), .o (n2328) );
  assign n2335 = ~n2319 & n2328 ;
  buffer buf_n2336( .i (n2335), .o (n2336) );
  buffer buf_n2337( .i (n2336), .o (n2337) );
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  buffer buf_n2340( .i (n2339), .o (n2340) );
  buffer buf_n2341( .i (n2340), .o (n2341) );
  buffer buf_n2342( .i (n2341), .o (n2342) );
  buffer buf_n2343( .i (n2342), .o (n2343) );
  buffer buf_n2344( .i (n2343), .o (n2344) );
  buffer buf_n2345( .i (n2344), .o (n2345) );
  buffer buf_n2346( .i (n2345), .o (n2346) );
  buffer buf_n2347( .i (n2346), .o (n2347) );
  buffer buf_n2348( .i (n2347), .o (n2348) );
  buffer buf_n2349( .i (n2348), .o (n2349) );
  assign n2350 = ~n2282 & n2349 ;
  assign n2351 = n2256 & n2350 ;
  assign n2352 = n2178 & n2351 ;
  buffer buf_n2353( .i (n2352), .o (n2353) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  assign n2354 = n298 | n310 ;
  assign n2355 = n298 & n310 ;
  assign n2356 = n2354 & ~n2355 ;
  buffer buf_n2357( .i (n2356), .o (n2357) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  assign n2358 = n324 & ~n340 ;
  assign n2359 = ~n324 & n340 ;
  assign n2360 = n2358 | n2359 ;
  buffer buf_n2361( .i (n2360), .o (n2361) );
  assign n2362 = ~n2357 & n2361 ;
  assign n2363 = n2357 & ~n2361 ;
  assign n2364 = n2362 | n2363 ;
  buffer buf_n2365( .i (n2364), .o (n2365) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n488( .i (G132), .o (n488) );
  assign n2366 = n486 & ~n488 ;
  assign n2367 = ~n486 & n488 ;
  assign n2368 = n2366 | n2367 ;
  buffer buf_n2369( .i (n2368), .o (n2369) );
  assign n2370 = n359 & ~n2369 ;
  assign n2371 = ~n359 & n2369 ;
  assign n2372 = n2370 | n2371 ;
  buffer buf_n2373( .i (n2372), .o (n2373) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  assign n2374 = n443 & ~n467 ;
  assign n2375 = ~n443 & n467 ;
  assign n2376 = n2374 | n2375 ;
  buffer buf_n2377( .i (n2376), .o (n2377) );
  assign n2378 = n2373 & ~n2377 ;
  assign n2379 = ~n2373 & n2377 ;
  assign n2380 = n2378 | n2379 ;
  buffer buf_n2381( .i (n2380), .o (n2381) );
  assign n2382 = n2365 | n2381 ;
  assign n2383 = n2365 & n2381 ;
  assign n2384 = n2382 & ~n2383 ;
  buffer buf_n2385( .i (n2384), .o (n2385) );
  inverter inv_n3914( .i (n2385), .o (n3914) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  assign n2386 = n893 | n918 ;
  assign n2387 = n893 & n918 ;
  assign n2388 = n2386 & ~n2387 ;
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  assign n2390 = n946 & ~n973 ;
  assign n2391 = ~n946 & n973 ;
  assign n2392 = n2390 | n2391 ;
  buffer buf_n2393( .i (n2392), .o (n2393) );
  assign n2394 = ~n2389 & n2393 ;
  assign n2395 = n2389 & ~n2393 ;
  assign n2396 = n2394 | n2395 ;
  buffer buf_n2397( .i (n2396), .o (n2397) );
  buffer buf_n2398( .i (n209), .o (n2398) );
  buffer buf_n2399( .i (n991), .o (n2399) );
  assign n2400 = n2398 | n2399 ;
  assign n2401 = n2398 & n2399 ;
  assign n2402 = n2400 & ~n2401 ;
  buffer buf_n2403( .i (n2402), .o (n2403) );
  buffer buf_n285( .i (G111), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n2404( .i (n277), .o (n2404) );
  assign n2405 = ~n286 & n2404 ;
  assign n2406 = n286 & ~n2404 ;
  assign n2407 = n2405 | n2406 ;
  buffer buf_n2408( .i (n2407), .o (n2408) );
  assign n2409 = n2403 | n2408 ;
  assign n2410 = n2403 & n2408 ;
  assign n2411 = n2409 & ~n2410 ;
  buffer buf_n2412( .i (n2411), .o (n2412) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  assign n2413 = n233 & ~n257 ;
  assign n2414 = ~n233 & n257 ;
  assign n2415 = n2413 | n2414 ;
  buffer buf_n2416( .i (n2415), .o (n2416) );
  assign n2417 = n2412 & ~n2416 ;
  assign n2418 = ~n2412 & n2416 ;
  assign n2419 = n2417 | n2418 ;
  buffer buf_n2420( .i (n2419), .o (n2420) );
  assign n2421 = n2397 & n2420 ;
  assign n2422 = n2397 | n2420 ;
  assign n2423 = ~n2421 & n2422 ;
  buffer buf_n2424( .i (n2423), .o (n2424) );
  inverter inv_n3915( .i (n2424), .o (n3915) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  assign n2425 = n1395 & n1464 ;
  buffer buf_n2426( .i (n2425), .o (n2426) );
  assign n2432 = n1475 | n1537 ;
  assign n2433 = n2426 | n2432 ;
  assign n2434 = n1541 & n2433 ;
  buffer buf_n2435( .i (n2434), .o (n2435) );
  assign n2446 = n1360 & n1598 ;
  assign n2447 = n2435 & n2446 ;
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  assign n2448 = n1358 & n1593 ;
  assign n2449 = n1354 | n2448 ;
  assign n2450 = n2447 | n2449 ;
  buffer buf_n2451( .i (n2450), .o (n2451) );
  buffer buf_n2452( .i (n2451), .o (n2452) );
  buffer buf_n2453( .i (n2452), .o (n2453) );
  buffer buf_n2454( .i (n2453), .o (n2454) );
  buffer buf_n2455( .i (n2454), .o (n2455) );
  buffer buf_n2456( .i (n2455), .o (n2456) );
  buffer buf_n2457( .i (n2456), .o (n2457) );
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n2460( .i (n2459), .o (n2460) );
  buffer buf_n2461( .i (n2460), .o (n2461) );
  assign n2462 = n1964 & n2461 ;
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  assign n2463 = n1840 & n1889 ;
  buffer buf_n2464( .i (n2463), .o (n2464) );
  assign n2470 = n1837 | n2464 ;
  buffer buf_n2471( .i (n2470), .o (n2471) );
  buffer buf_n2472( .i (n2471), .o (n2472) );
  buffer buf_n2473( .i (n2472), .o (n2473) );
  assign n2486 = n1780 & n2473 ;
  buffer buf_n2487( .i (n2486), .o (n2487) );
  buffer buf_n2488( .i (n2487), .o (n2488) );
  buffer buf_n2489( .i (n2488), .o (n2489) );
  buffer buf_n2490( .i (n2489), .o (n2490) );
  buffer buf_n2491( .i (n2490), .o (n2491) );
  buffer buf_n2492( .i (n2491), .o (n2492) );
  buffer buf_n2493( .i (n2492), .o (n2493) );
  buffer buf_n2494( .i (n2493), .o (n2494) );
  buffer buf_n2495( .i (n2494), .o (n2495) );
  buffer buf_n2496( .i (n2495), .o (n2496) );
  buffer buf_n2497( .i (n2496), .o (n2497) );
  assign n2498 = n1774 | n2497 ;
  buffer buf_n2499( .i (n2498), .o (n2499) );
  assign n2500 = n1708 & n2499 ;
  assign n2501 = n1688 | n2500 ;
  assign n2502 = n2462 | n2501 ;
  buffer buf_n2503( .i (n2502), .o (n2503) );
  assign n2504 = ~n2268 & n2278 ;
  inverter inv_n2505( .i (n2504), .o (n2505) );
  buffer buf_n800( .i (G176), .o (n800) );
  buffer buf_n806( .i (G177), .o (n806) );
  assign n2506 = n800 & ~n806 ;
  buffer buf_n2507( .i (n2506), .o (n2507) );
  buffer buf_n2508( .i (n2507), .o (n2508) );
  buffer buf_n2509( .i (n2508), .o (n2509) );
  buffer buf_n2510( .i (n2509), .o (n2510) );
  assign n2517 = G60 & n2510 ;
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n823( .i (G21), .o (n823) );
  buffer buf_n2056( .i (n2055), .o (n2056) );
  buffer buf_n2057( .i (n2056), .o (n2057) );
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  buffer buf_n2064( .i (n2063), .o (n2064) );
  buffer buf_n2065( .i (n2064), .o (n2065) );
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n2073( .i (n2072), .o (n2073) );
  assign n2518 = ~n823 & n2073 ;
  assign n2519 = n823 & ~n2073 ;
  assign n2520 = n2518 | n2519 ;
  buffer buf_n2521( .i (n2520), .o (n2521) );
  assign n2522 = ~n804 & n2521 ;
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  assign n2523 = n803 & ~n1164 ;
  assign n2524 = n810 & ~n2523 ;
  assign n2525 = ~n2522 & n2524 ;
  assign n2526 = n2517 | n2525 ;
  buffer buf_n2527( .i (n2526), .o (n2527) );
  inverter inv_n3916( .i (n2527), .o (n3916) );
  assign n2529 = G58 & n2509 ;
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n2102( .i (n2101), .o (n2102) );
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n2111( .i (n2110), .o (n2111) );
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2077( .i (n2076), .o (n2077) );
  buffer buf_n2078( .i (n2077), .o (n2078) );
  buffer buf_n2079( .i (n2078), .o (n2079) );
  buffer buf_n2080( .i (n2079), .o (n2080) );
  buffer buf_n2081( .i (n2080), .o (n2081) );
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2089( .i (n2088), .o (n2089) );
  buffer buf_n2090( .i (n2089), .o (n2090) );
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  assign n2530 = n2051 & ~n2092 ;
  assign n2531 = n2072 & ~n2530 ;
  assign n2532 = n2114 | n2531 ;
  buffer buf_n2533( .i (n2532), .o (n2533) );
  assign n2536 = n803 | n2533 ;
  assign n2537 = n802 & n1107 ;
  assign n2538 = n809 & ~n2537 ;
  assign n2539 = n2536 & n2538 ;
  assign n2540 = n2529 | n2539 ;
  buffer buf_n2541( .i (n2540), .o (n2541) );
  inverter inv_n3917( .i (n2541), .o (n3917) );
  assign n2544 = G48 & n2510 ;
  buffer buf_n814( .i (G2), .o (n814) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  assign n2545 = n814 & n1427 ;
  buffer buf_n2546( .i (n2545), .o (n2546) );
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  buffer buf_n2551( .i (n2550), .o (n2551) );
  buffer buf_n2552( .i (n2551), .o (n2552) );
  buffer buf_n2553( .i (n2552), .o (n2553) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  assign n2554 = n822 | n1435 ;
  assign n2555 = ~n2553 & n2554 ;
  buffer buf_n2556( .i (n2555), .o (n2556) );
  assign n2557 = n804 | n2556 ;
  assign n2558 = n803 & n1252 ;
  assign n2559 = n810 & ~n2558 ;
  assign n2560 = n2557 & n2559 ;
  assign n2561 = n2544 | n2560 ;
  buffer buf_n2562( .i (n2561), .o (n2562) );
  inverter inv_n3918( .i (n2562), .o (n3918) );
  buffer buf_n2269( .i (n2268), .o (n2269) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  assign n2565 = n2269 & n2279 ;
  assign n2566 = n2282 & ~n2565 ;
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n788( .i (G173), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n2563( .i (n2562), .o (n2563) );
  buffer buf_n2564( .i (n2563), .o (n2564) );
  assign n2575 = n791 | n2564 ;
  buffer buf_n784( .i (G172), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n2528( .i (n2527), .o (n2528) );
  assign n2576 = n790 & ~n2528 ;
  assign n2577 = n787 & ~n2576 ;
  assign n2578 = n2575 & n2577 ;
  buffer buf_n830( .i (G3), .o (n830) );
  assign n2579 = ~n784 & n788 ;
  buffer buf_n2580( .i (n2579), .o (n2580) );
  buffer buf_n2581( .i (n2580), .o (n2581) );
  assign n2582 = n830 & n2581 ;
  buffer buf_n824( .i (G22), .o (n824) );
  assign n2583 = n784 | n788 ;
  buffer buf_n2584( .i (n2583), .o (n2584) );
  buffer buf_n2585( .i (n2584), .o (n2585) );
  assign n2586 = n824 & ~n2585 ;
  assign n2587 = n2582 | n2586 ;
  assign n2588 = n2578 | n2587 ;
  assign n2589 = G19 & n2509 ;
  buffer buf_n1995( .i (n1994), .o (n1995) );
  buffer buf_n1996( .i (n1995), .o (n1996) );
  buffer buf_n1997( .i (n1996), .o (n1997) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n1986( .i (n1985), .o (n1986) );
  buffer buf_n2138( .i (n2137), .o (n2138) );
  buffer buf_n2139( .i (n2138), .o (n2139) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  assign n2590 = n2079 & n2142 ;
  assign n2591 = n2139 | n2590 ;
  buffer buf_n2592( .i (n2591), .o (n2592) );
  assign n2597 = n1986 | n2592 ;
  assign n2598 = n1997 & n2597 ;
  assign n2599 = n2165 | n2598 ;
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  buffer buf_n2602( .i (n2601), .o (n2602) );
  buffer buf_n2603( .i (n2602), .o (n2603) );
  buffer buf_n2604( .i (n2603), .o (n2604) );
  buffer buf_n2605( .i (n2604), .o (n2605) );
  buffer buf_n2606( .i (n2605), .o (n2606) );
  buffer buf_n2607( .i (n2606), .o (n2607) );
  assign n2608 = n2347 | n2607 ;
  assign n2609 = n2347 & n2607 ;
  assign n2610 = n2608 & ~n2609 ;
  buffer buf_n2611( .i (n2610), .o (n2611) );
  buffer buf_n2617( .i (n802), .o (n2617) );
  assign n2618 = n2611 & ~n2617 ;
  assign n2619 = n802 & n1182 ;
  assign n2620 = n809 & ~n2619 ;
  assign n2621 = ~n2618 & n2620 ;
  assign n2622 = n2589 | n2621 ;
  buffer buf_n2623( .i (n2622), .o (n2623) );
  inverter inv_n3919( .i (n2623), .o (n3919) );
  assign n2626 = G59 & n2507 ;
  buffer buf_n2005( .i (n2004), .o (n2005) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n2007( .i (n2006), .o (n2007) );
  buffer buf_n2008( .i (n2007), .o (n2008) );
  buffer buf_n2009( .i (n2008), .o (n2009) );
  buffer buf_n2010( .i (n2009), .o (n2010) );
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n2012( .i (n2011), .o (n2012) );
  buffer buf_n2013( .i (n2012), .o (n2013) );
  buffer buf_n2160( .i (n2159), .o (n2160) );
  buffer buf_n2161( .i (n2160), .o (n2161) );
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n2163( .i (n2162), .o (n2163) );
  buffer buf_n2593( .i (n2592), .o (n2593) );
  buffer buf_n2594( .i (n2593), .o (n2594) );
  buffer buf_n2595( .i (n2594), .o (n2595) );
  buffer buf_n2596( .i (n2595), .o (n2596) );
  assign n2627 = n2163 | n2596 ;
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  buffer buf_n2631( .i (n2630), .o (n2631) );
  assign n2632 = ~n2013 & n2631 ;
  assign n2633 = n2013 & ~n2631 ;
  assign n2634 = n2632 | n2633 ;
  buffer buf_n2635( .i (n2634), .o (n2635) );
  assign n2642 = ~n801 & n2635 ;
  assign n2643 = n800 & n1168 ;
  assign n2644 = n807 & ~n2643 ;
  assign n2645 = ~n2642 & n2644 ;
  assign n2646 = n2626 | n2645 ;
  buffer buf_n2647( .i (n2646), .o (n2647) );
  inverter inv_n3920( .i (n2647), .o (n3920) );
  assign n2652 = G50 & n2509 ;
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  buffer buf_n2152( .i (n2151), .o (n2152) );
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n2155( .i (n2154), .o (n2155) );
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  assign n2653 = n2091 | n2111 ;
  buffer buf_n2654( .i (n2653), .o (n2654) );
  assign n2655 = n2157 | n2654 ;
  assign n2656 = n2157 & n2654 ;
  assign n2657 = n2655 & ~n2656 ;
  buffer buf_n2658( .i (n2657), .o (n2658) );
  assign n2662 = ~n2617 & n2658 ;
  buffer buf_n2663( .i (n801), .o (n2663) );
  assign n2664 = n1195 & n2663 ;
  assign n2665 = n809 & ~n2664 ;
  assign n2666 = ~n2662 & n2665 ;
  assign n2667 = n2652 | n2666 ;
  buffer buf_n2668( .i (n2667), .o (n2668) );
  inverter inv_n3921( .i (n2668), .o (n3921) );
  buffer buf_n792( .i (G174), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  assign n2671 = n795 | n2564 ;
  buffer buf_n796( .i (G175), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  assign n2672 = n794 & ~n2528 ;
  assign n2673 = n799 & ~n2672 ;
  assign n2674 = n2671 & n2673 ;
  assign n2675 = n792 & ~n796 ;
  buffer buf_n2676( .i (n2675), .o (n2676) );
  buffer buf_n2677( .i (n2676), .o (n2677) );
  assign n2678 = n830 & n2677 ;
  assign n2679 = n792 | n796 ;
  buffer buf_n2680( .i (n2679), .o (n2680) );
  buffer buf_n2681( .i (n2680), .o (n2681) );
  assign n2682 = n824 & ~n2681 ;
  assign n2683 = n2678 | n2682 ;
  assign n2684 = n2674 | n2683 ;
  assign n2685 = G53 & n2510 ;
  assign n2686 = n814 & n1635 ;
  buffer buf_n2687( .i (n2686), .o (n2687) );
  buffer buf_n2688( .i (n2687), .o (n2688) );
  buffer buf_n2689( .i (n2688), .o (n2689) );
  buffer buf_n2690( .i (n2689), .o (n2690) );
  buffer buf_n2691( .i (n2690), .o (n2691) );
  buffer buf_n2692( .i (n2691), .o (n2692) );
  buffer buf_n2693( .i (n2692), .o (n2693) );
  buffer buf_n2694( .i (n2693), .o (n2694) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n1633( .i (n1632), .o (n1633) );
  assign n2695 = n821 & n1633 ;
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n2436( .i (n2435), .o (n2436) );
  assign n2696 = n1589 & n2436 ;
  assign n2697 = n1596 | n2696 ;
  buffer buf_n2698( .i (n2697), .o (n2698) );
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n2700( .i (n2699), .o (n2700) );
  assign n2701 = ~n1367 & n2700 ;
  assign n2702 = n1367 & ~n2700 ;
  assign n2703 = n2701 | n2702 ;
  buffer buf_n2704( .i (n2703), .o (n2704) );
  buffer buf_n2705( .i (n2704), .o (n2705) );
  buffer buf_n2706( .i (n2705), .o (n2706) );
  buffer buf_n2707( .i (n2706), .o (n2707) );
  buffer buf_n2708( .i (n2707), .o (n2708) );
  assign n2709 = n2695 | n2708 ;
  assign n2710 = ~n2694 & n2709 ;
  buffer buf_n2711( .i (n2710), .o (n2711) );
  assign n2715 = ~n804 & n2711 ;
  assign n2716 = n1263 & n2617 ;
  assign n2717 = n810 & ~n2716 ;
  assign n2718 = ~n2715 & n2717 ;
  assign n2719 = n2685 | n2718 ;
  buffer buf_n2720( .i (n2719), .o (n2720) );
  inverter inv_n3922( .i (n2720), .o (n3922) );
  buffer buf_n2723( .i (n2508), .o (n2723) );
  buffer buf_n2724( .i (n2723), .o (n2724) );
  assign n2725 = G57 & n2724 ;
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n2437( .i (n2436), .o (n2437) );
  buffer buf_n2438( .i (n2437), .o (n2438) );
  buffer buf_n2439( .i (n2438), .o (n2439) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  assign n2726 = n1510 & n1548 ;
  assign n2727 = n2439 | n2726 ;
  buffer buf_n2728( .i (n2727), .o (n2728) );
  buffer buf_n2729( .i (n2728), .o (n2729) );
  buffer buf_n2730( .i (n2729), .o (n2730) );
  buffer buf_n2731( .i (n2730), .o (n2731) );
  buffer buf_n2732( .i (n2731), .o (n2732) );
  buffer buf_n2733( .i (n2732), .o (n2733) );
  buffer buf_n2440( .i (n2439), .o (n2440) );
  buffer buf_n2441( .i (n2440), .o (n2441) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  buffer buf_n2443( .i (n2442), .o (n2443) );
  buffer buf_n2444( .i (n2443), .o (n2444) );
  buffer buf_n2445( .i (n2444), .o (n2445) );
  assign n2734 = n819 | n2445 ;
  assign n2735 = n2733 & n2734 ;
  buffer buf_n2736( .i (n2735), .o (n2736) );
  assign n2737 = ~n1612 & n2736 ;
  assign n2738 = n1612 & ~n2736 ;
  assign n2739 = n2737 | n2738 ;
  buffer buf_n2740( .i (n2739), .o (n2740) );
  buffer buf_n2742( .i (n2617), .o (n2742) );
  assign n2743 = n2740 & ~n2742 ;
  buffer buf_n2744( .i (n2663), .o (n2744) );
  assign n2745 = n1307 & n2744 ;
  buffer buf_n2746( .i (n808), .o (n2746) );
  buffer buf_n2747( .i (n2746), .o (n2747) );
  assign n2748 = ~n2745 & n2747 ;
  assign n2749 = ~n2743 & n2748 ;
  assign n2750 = n2725 | n2749 ;
  buffer buf_n2751( .i (n2750), .o (n2751) );
  inverter inv_n3923( .i (n2751), .o (n3923) );
  assign n2754 = G56 & n2724 ;
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n1556( .i (n1555), .o (n1556) );
  buffer buf_n1557( .i (n1556), .o (n1557) );
  buffer buf_n1558( .i (n1557), .o (n1558) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n1488( .i (n1487), .o (n1488) );
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  assign n2755 = n1407 | n2546 ;
  buffer buf_n2756( .i (n2755), .o (n2756) );
  assign n2761 = n1502 & n2756 ;
  buffer buf_n2762( .i (n2761), .o (n2762) );
  assign n2766 = n1490 | n2762 ;
  buffer buf_n2767( .i (n2766), .o (n2767) );
  assign n2768 = n1558 | n2767 ;
  assign n2769 = n1558 & n2767 ;
  assign n2770 = n2768 & ~n2769 ;
  buffer buf_n2771( .i (n2770), .o (n2771) );
  assign n2774 = ~n2742 & n2771 ;
  assign n2775 = n1324 & n2744 ;
  assign n2776 = n2747 & ~n2775 ;
  assign n2777 = ~n2774 & n2776 ;
  assign n2778 = n2754 | n2777 ;
  buffer buf_n2779( .i (n2778), .o (n2779) );
  inverter inv_n3924( .i (n2779), .o (n3924) );
  assign n2782 = G55 & n2724 ;
  buffer buf_n2763( .i (n2762), .o (n2763) );
  buffer buf_n2764( .i (n2763), .o (n2764) );
  buffer buf_n2765( .i (n2764), .o (n2765) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n2757( .i (n2756), .o (n2757) );
  buffer buf_n2758( .i (n2757), .o (n2758) );
  buffer buf_n2759( .i (n2758), .o (n2759) );
  buffer buf_n2760( .i (n2759), .o (n2760) );
  assign n2783 = n1506 | n2760 ;
  assign n2784 = ~n2765 & n2783 ;
  buffer buf_n2785( .i (n2784), .o (n2785) );
  assign n2786 = ~n2742 & n2785 ;
  assign n2787 = n1276 & n2744 ;
  assign n2788 = n2747 & ~n2787 ;
  assign n2789 = ~n2786 & n2788 ;
  assign n2790 = n2782 | n2789 ;
  buffer buf_n2791( .i (n2790), .o (n2791) );
  inverter inv_n3925( .i (n2791), .o (n3925) );
  buffer buf_n2185( .i (n2184), .o (n2185) );
  assign n2794 = n2185 & n2261 ;
  assign n2795 = n2185 | n2261 ;
  assign n2796 = ~n2794 & n2795 ;
  buffer buf_n2797( .i (n2796), .o (n2797) );
  buffer buf_n2798( .i (n2797), .o (n2798) );
  buffer buf_n2799( .i (n2798), .o (n2799) );
  buffer buf_n2800( .i (n2799), .o (n2800) );
  buffer buf_n2801( .i (n2800), .o (n2801) );
  buffer buf_n2802( .i (n2801), .o (n2802) );
  buffer buf_n2803( .i (n2802), .o (n2803) );
  buffer buf_n2804( .i (n2803), .o (n2804) );
  buffer buf_n2805( .i (n2804), .o (n2805) );
  buffer buf_n2806( .i (n2805), .o (n2806) );
  buffer buf_n2208( .i (n2207), .o (n2208) );
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n2211( .i (n2210), .o (n2211) );
  buffer buf_n2212( .i (n2211), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  buffer buf_n2214( .i (n2213), .o (n2214) );
  buffer buf_n2215( .i (n2214), .o (n2215) );
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n2221( .i (n2220), .o (n2221) );
  buffer buf_n2280( .i (n2279), .o (n2280) );
  assign n2807 = n2221 & n2280 ;
  assign n2808 = n2221 | n2280 ;
  assign n2809 = ~n2807 & n2808 ;
  buffer buf_n2810( .i (n2809), .o (n2810) );
  assign n2811 = ~n2806 & n2810 ;
  assign n2812 = n2806 & ~n2810 ;
  assign n2813 = n2811 | n2812 ;
  buffer buf_n2814( .i (n2813), .o (n2814) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  assign n2815 = n381 & n490 ;
  assign n2816 = G133 & ~n381 ;
  assign n2817 = n2815 | n2816 ;
  buffer buf_n2818( .i (n2817), .o (n2818) );
  buffer buf_n2020( .i (n2019), .o (n2020) );
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2028( .i (n2027), .o (n2028) );
  buffer buf_n2029( .i (n2028), .o (n2029) );
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n2031( .i (n2030), .o (n2031) );
  buffer buf_n2032( .i (n2031), .o (n2032) );
  buffer buf_n2033( .i (n2032), .o (n2033) );
  buffer buf_n2034( .i (n2033), .o (n2034) );
  buffer buf_n2035( .i (n2034), .o (n2035) );
  buffer buf_n2120( .i (n2119), .o (n2120) );
  buffer buf_n2121( .i (n2120), .o (n2121) );
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  buffer buf_n2129( .i (n2128), .o (n2129) );
  buffer buf_n2130( .i (n2129), .o (n2130) );
  buffer buf_n2131( .i (n2130), .o (n2131) );
  buffer buf_n2132( .i (n2131), .o (n2132) );
  buffer buf_n2133( .i (n2132), .o (n2133) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  assign n2819 = n2035 | n2135 ;
  assign n2820 = n2035 & n2135 ;
  assign n2821 = n2819 & ~n2820 ;
  buffer buf_n2822( .i (n2821), .o (n2822) );
  assign n2823 = n2818 | n2822 ;
  assign n2824 = n2818 & n2822 ;
  assign n2825 = n2823 & ~n2824 ;
  buffer buf_n2826( .i (n2825), .o (n2826) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n1969( .i (n1968), .o (n1969) );
  buffer buf_n1970( .i (n1969), .o (n1970) );
  buffer buf_n1971( .i (n1970), .o (n1971) );
  buffer buf_n1972( .i (n1971), .o (n1972) );
  buffer buf_n1973( .i (n1972), .o (n1973) );
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  buffer buf_n2307( .i (n2306), .o (n2307) );
  buffer buf_n2308( .i (n2307), .o (n2308) );
  buffer buf_n2309( .i (n2308), .o (n2309) );
  buffer buf_n2310( .i (n2309), .o (n2310) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  assign n2827 = n1982 & n2317 ;
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n2289( .i (n2288), .o (n2289) );
  buffer buf_n2290( .i (n2289), .o (n2290) );
  buffer buf_n2291( .i (n2290), .o (n2291) );
  buffer buf_n2292( .i (n2291), .o (n2292) );
  buffer buf_n2293( .i (n2292), .o (n2293) );
  buffer buf_n2294( .i (n2293), .o (n2294) );
  buffer buf_n2295( .i (n2294), .o (n2295) );
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n2297( .i (n2296), .o (n2297) );
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  assign n2828 = n422 | n2300 ;
  assign n2829 = ~n2827 & n2828 ;
  buffer buf_n2830( .i (n2829), .o (n2830) );
  assign n2831 = ~n2074 & n2830 ;
  assign n2832 = n2074 & ~n2830 ;
  assign n2833 = n2831 | n2832 ;
  buffer buf_n2834( .i (n2833), .o (n2834) );
  assign n2835 = n2826 & ~n2834 ;
  assign n2836 = ~n2826 & n2834 ;
  assign n2837 = n2835 | n2836 ;
  buffer buf_n2838( .i (n2837), .o (n2838) );
  assign n2839 = ~n2814 & n2838 ;
  assign n2840 = n2814 & ~n2838 ;
  assign n2841 = n2839 | n2840 ;
  buffer buf_n2842( .i (n2841), .o (n2842) );
  inverter inv_n3926( .i (n2842), .o (n3926) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n1522( .i (n1521), .o (n1522) );
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  buffer buf_n1534( .i (n1533), .o (n1534) );
  buffer buf_n1535( .i (n1534), .o (n1535) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  assign n2843 = n1535 & n1583 ;
  assign n2844 = n1535 | n1583 ;
  assign n2845 = ~n2843 & n2844 ;
  buffer buf_n2846( .i (n2845), .o (n2846) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  buffer buf_n1455( .i (n1454), .o (n1455) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  assign n2847 = ~n1393 & n1462 ;
  assign n2848 = n1393 & ~n1462 ;
  assign n2849 = n2847 | n2848 ;
  buffer buf_n2850( .i (n2849), .o (n2850) );
  assign n2851 = n2846 | n2850 ;
  assign n2852 = n2846 & n2850 ;
  assign n2853 = n2851 & ~n2852 ;
  buffer buf_n2854( .i (n2853), .o (n2854) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  buffer buf_n1813( .i (n1812), .o (n1813) );
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  buffer buf_n1821( .i (n1820), .o (n1821) );
  buffer buf_n1822( .i (n1821), .o (n1822) );
  buffer buf_n1823( .i (n1822), .o (n1823) );
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1825( .i (n1824), .o (n1825) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  assign n2855 = n1756 & n1832 ;
  assign n2856 = n1756 | n1832 ;
  assign n2857 = ~n2855 & n2856 ;
  buffer buf_n2858( .i (n2857), .o (n2858) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  buffer buf_n1872( .i (n1871), .o (n1872) );
  buffer buf_n1873( .i (n1872), .o (n1873) );
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  buffer buf_n1879( .i (n1878), .o (n1879) );
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  assign n2859 = n285 & n405 ;
  assign n2860 = G112 & ~n405 ;
  assign n2861 = n2859 | n2860 ;
  buffer buf_n2862( .i (n2861), .o (n2862) );
  assign n2863 = n1887 & ~n2862 ;
  assign n2864 = ~n1887 & n2862 ;
  assign n2865 = n2863 | n2864 ;
  buffer buf_n2866( .i (n2865), .o (n2866) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  buffer buf_n1658( .i (n1657), .o (n1658) );
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  assign n2867 = ~n1349 & n1667 ;
  assign n2868 = n1349 & ~n1667 ;
  assign n2869 = n2867 | n2868 ;
  buffer buf_n2870( .i (n2869), .o (n2870) );
  assign n2871 = ~n2866 & n2870 ;
  assign n2872 = n2866 & ~n2870 ;
  assign n2873 = n2871 | n2872 ;
  buffer buf_n2874( .i (n2873), .o (n2874) );
  assign n2875 = ~n2858 & n2874 ;
  assign n2876 = n2858 & ~n2874 ;
  assign n2877 = n2875 | n2876 ;
  buffer buf_n2878( .i (n2877), .o (n2878) );
  assign n2879 = ~n2854 & n2878 ;
  assign n2880 = n2854 & ~n2878 ;
  assign n2881 = n2879 | n2880 ;
  buffer buf_n2882( .i (n2881), .o (n2882) );
  inverter inv_n3927( .i (n2882), .o (n3927) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  assign n2883 = n2455 | n2687 ;
  buffer buf_n2884( .i (n2883), .o (n2884) );
  buffer buf_n2885( .i (n2884), .o (n2885) );
  buffer buf_n2886( .i (n2885), .o (n2886) );
  assign n2888 = n1962 & n2886 ;
  assign n2889 = n2499 | n2888 ;
  buffer buf_n2890( .i (n2889), .o (n2890) );
  assign n2891 = n1728 | n2890 ;
  assign n2892 = n1728 & n2890 ;
  assign n2893 = n2891 & ~n2892 ;
  buffer buf_n2894( .i (n2893), .o (n2894) );
  buffer buf_n2895( .i (n2894), .o (n2895) );
  buffer buf_n2896( .i (n2895), .o (n2896) );
  buffer buf_n2897( .i (n2896), .o (n2897) );
  buffer buf_n2898( .i (n2897), .o (n2898) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  buffer buf_n1930( .i (n1929), .o (n1930) );
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n1934( .i (n1933), .o (n1934) );
  buffer buf_n1935( .i (n1934), .o (n1935) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n2887( .i (n2886), .o (n2887) );
  assign n2899 = n1945 | n2887 ;
  assign n2900 = n1945 & n2887 ;
  assign n2901 = n2899 & ~n2900 ;
  buffer buf_n2902( .i (n2901), .o (n2902) );
  buffer buf_n2903( .i (n2902), .o (n2903) );
  buffer buf_n2904( .i (n2903), .o (n2904) );
  buffer buf_n2905( .i (n2904), .o (n2905) );
  buffer buf_n2906( .i (n2905), .o (n2906) );
  buffer buf_n2907( .i (n2906), .o (n2907) );
  buffer buf_n2712( .i (n2711), .o (n2712) );
  buffer buf_n2713( .i (n2712), .o (n2713) );
  buffer buf_n2714( .i (n2713), .o (n2714) );
  buffer buf_n2772( .i (n2771), .o (n2772) );
  buffer buf_n2773( .i (n2772), .o (n2773) );
  buffer buf_n2741( .i (n2740), .o (n2741) );
  assign n2908 = ~n2556 & n2785 ;
  assign n2909 = n2741 & n2908 ;
  assign n2910 = n2773 & n2909 ;
  assign n2911 = n2714 & n2910 ;
  assign n2912 = ~n2907 & n2911 ;
  assign n2913 = n2898 & n2912 ;
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n2474( .i (n2473), .o (n2474) );
  buffer buf_n2475( .i (n2474), .o (n2475) );
  buffer buf_n2476( .i (n2475), .o (n2476) );
  buffer buf_n2477( .i (n2476), .o (n2477) );
  buffer buf_n2478( .i (n2477), .o (n2478) );
  buffer buf_n2479( .i (n2478), .o (n2479) );
  buffer buf_n2480( .i (n2479), .o (n2480) );
  buffer buf_n2481( .i (n2480), .o (n2481) );
  buffer buf_n2482( .i (n2481), .o (n2482) );
  buffer buf_n2483( .i (n2482), .o (n2483) );
  buffer buf_n2484( .i (n2483), .o (n2484) );
  buffer buf_n2485( .i (n2484), .o (n2485) );
  assign n2914 = n1960 & n2884 ;
  assign n2915 = n2485 | n2914 ;
  buffer buf_n2916( .i (n2915), .o (n2916) );
  assign n2917 = ~n1802 & n2916 ;
  assign n2918 = n1802 & ~n2916 ;
  assign n2919 = n2917 | n2918 ;
  buffer buf_n2920( .i (n2919), .o (n2920) );
  buffer buf_n2921( .i (n2920), .o (n2921) );
  buffer buf_n2922( .i (n2921), .o (n2922) );
  buffer buf_n2923( .i (n2922), .o (n2923) );
  buffer buf_n2924( .i (n2923), .o (n2924) );
  buffer buf_n2925( .i (n2924), .o (n2925) );
  buffer buf_n2926( .i (n2925), .o (n2926) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  buffer buf_n1846( .i (n1845), .o (n1846) );
  buffer buf_n1847( .i (n1846), .o (n1847) );
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n1915( .i (n1914), .o (n1915) );
  buffer buf_n1916( .i (n1915), .o (n1916) );
  buffer buf_n1917( .i (n1916), .o (n1917) );
  buffer buf_n1918( .i (n1917), .o (n1918) );
  buffer buf_n1919( .i (n1918), .o (n1919) );
  buffer buf_n1920( .i (n1919), .o (n1920) );
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  assign n2927 = n1925 & n2884 ;
  buffer buf_n1890( .i (n1889), .o (n1890) );
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  assign n2928 = n1906 | n2884 ;
  assign n2929 = ~n2927 & n2928 ;
  buffer buf_n2930( .i (n2929), .o (n2930) );
  assign n2931 = n1861 | n2930 ;
  assign n2932 = n1861 & n2930 ;
  assign n2933 = n2931 & ~n2932 ;
  buffer buf_n2934( .i (n2933), .o (n2934) );
  buffer buf_n2935( .i (n2934), .o (n2935) );
  buffer buf_n2936( .i (n2935), .o (n2936) );
  buffer buf_n2937( .i (n2936), .o (n2937) );
  buffer buf_n2938( .i (n2937), .o (n2938) );
  buffer buf_n2939( .i (n2938), .o (n2939) );
  buffer buf_n2940( .i (n2939), .o (n2940) );
  assign n2941 = n2926 & ~n2940 ;
  assign n2942 = n2913 & n2941 ;
  buffer buf_n2200( .i (n2199), .o (n2200) );
  buffer buf_n2201( .i (n2200), .o (n2201) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  buffer buf_n2203( .i (n2202), .o (n2203) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  buffer buf_n2235( .i (n2234), .o (n2235) );
  buffer buf_n2236( .i (n2235), .o (n2236) );
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n2321( .i (n2320), .o (n2321) );
  buffer buf_n2322( .i (n2321), .o (n2322) );
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2325( .i (n2324), .o (n2325) );
  buffer buf_n2326( .i (n2325), .o (n2326) );
  buffer buf_n2329( .i (n2328), .o (n2329) );
  buffer buf_n2330( .i (n2329), .o (n2330) );
  buffer buf_n2331( .i (n2330), .o (n2331) );
  buffer buf_n2332( .i (n2331), .o (n2332) );
  buffer buf_n2333( .i (n2332), .o (n2333) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  assign n2943 = n2334 & n2600 ;
  assign n2944 = n2326 | n2943 ;
  buffer buf_n2945( .i (n2944), .o (n2945) );
  buffer buf_n2946( .i (n2945), .o (n2946) );
  assign n2950 = n2239 & n2946 ;
  buffer buf_n2224( .i (n2223), .o (n2224) );
  buffer buf_n2225( .i (n2224), .o (n2225) );
  buffer buf_n2226( .i (n2225), .o (n2226) );
  buffer buf_n2227( .i (n2226), .o (n2227) );
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  assign n2951 = n2230 | n2946 ;
  assign n2952 = ~n2950 & n2951 ;
  buffer buf_n2953( .i (n2952), .o (n2953) );
  assign n2954 = n2203 & n2953 ;
  assign n2955 = n2203 | n2953 ;
  assign n2956 = ~n2954 & n2955 ;
  buffer buf_n2957( .i (n2956), .o (n2957) );
  buffer buf_n2958( .i (n2957), .o (n2958) );
  buffer buf_n2959( .i (n2958), .o (n2959) );
  buffer buf_n2960( .i (n2959), .o (n2960) );
  buffer buf_n2961( .i (n2960), .o (n2961) );
  buffer buf_n2962( .i (n2961), .o (n2962) );
  buffer buf_n2963( .i (n2962), .o (n2963) );
  buffer buf_n2964( .i (n2963), .o (n2964) );
  buffer buf_n2965( .i (n2964), .o (n2965) );
  buffer buf_n2189( .i (n2188), .o (n2189) );
  buffer buf_n2190( .i (n2189), .o (n2190) );
  buffer buf_n2191( .i (n2190), .o (n2191) );
  buffer buf_n2192( .i (n2191), .o (n2192) );
  buffer buf_n2195( .i (n2194), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  buffer buf_n2197( .i (n2196), .o (n2197) );
  assign n2966 = n2197 & n2230 ;
  assign n2967 = n2192 | n2966 ;
  buffer buf_n2947( .i (n2946), .o (n2947) );
  assign n2968 = n2251 & n2947 ;
  assign n2969 = n2967 | n2968 ;
  buffer buf_n2970( .i (n2969), .o (n2970) );
  assign n2971 = n2279 | n2970 ;
  assign n2972 = n2279 & n2970 ;
  assign n2973 = n2971 & ~n2972 ;
  buffer buf_n2974( .i (n2973), .o (n2974) );
  buffer buf_n2975( .i (n2974), .o (n2975) );
  buffer buf_n2976( .i (n2975), .o (n2976) );
  buffer buf_n2977( .i (n2976), .o (n2977) );
  buffer buf_n2978( .i (n2977), .o (n2978) );
  buffer buf_n2979( .i (n2978), .o (n2979) );
  buffer buf_n2980( .i (n2979), .o (n2980) );
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  buffer buf_n2948( .i (n2947), .o (n2948) );
  buffer buf_n2949( .i (n2948), .o (n2949) );
  assign n2981 = n2249 & n2949 ;
  assign n2982 = n2249 | n2949 ;
  assign n2983 = ~n2981 & n2982 ;
  buffer buf_n2984( .i (n2983), .o (n2984) );
  buffer buf_n2985( .i (n2984), .o (n2985) );
  buffer buf_n2986( .i (n2985), .o (n2986) );
  buffer buf_n2987( .i (n2986), .o (n2987) );
  buffer buf_n2988( .i (n2987), .o (n2988) );
  buffer buf_n2989( .i (n2988), .o (n2989) );
  buffer buf_n2990( .i (n2989), .o (n2990) );
  buffer buf_n2612( .i (n2611), .o (n2612) );
  buffer buf_n2613( .i (n2612), .o (n2613) );
  buffer buf_n2614( .i (n2613), .o (n2614) );
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  buffer buf_n2636( .i (n2635), .o (n2636) );
  buffer buf_n2637( .i (n2636), .o (n2637) );
  buffer buf_n2638( .i (n2637), .o (n2638) );
  buffer buf_n2639( .i (n2638), .o (n2639) );
  buffer buf_n2640( .i (n2639), .o (n2640) );
  buffer buf_n2641( .i (n2640), .o (n2641) );
  buffer buf_n2659( .i (n2658), .o (n2659) );
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2660), .o (n2661) );
  buffer buf_n2534( .i (n2533), .o (n2534) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  assign n2991 = n2521 & n2567 ;
  assign n2992 = ~n2535 & n2991 ;
  assign n2993 = n2661 & n2992 ;
  assign n2994 = n2641 & n2993 ;
  assign n2995 = n2616 & n2994 ;
  assign n2996 = ~n2990 & n2995 ;
  assign n2997 = ~n2980 & n2996 ;
  assign n2998 = ~n2965 & n2997 ;
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n745( .i (G158), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  assign n2999 = n748 | n2563 ;
  buffer buf_n749( .i (G159), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  assign n3000 = n747 & ~n2527 ;
  assign n3001 = n752 & ~n3000 ;
  assign n3002 = n2999 & n3001 ;
  buffer buf_n862( .i (G81), .o (n862) );
  assign n3003 = n745 | n749 ;
  buffer buf_n3004( .i (n3003), .o (n3004) );
  buffer buf_n3005( .i (n3004), .o (n3005) );
  assign n3006 = n862 & ~n3005 ;
  buffer buf_n861( .i (G80), .o (n861) );
  assign n3007 = n745 & ~n749 ;
  buffer buf_n3008( .i (n3007), .o (n3008) );
  buffer buf_n3009( .i (n3008), .o (n3009) );
  assign n3010 = n861 & n3009 ;
  assign n3011 = n3006 | n3010 ;
  assign n3012 = n3002 | n3011 ;
  assign n3013 = n846 & n3012 ;
  buffer buf_n754( .i (G160), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  assign n3014 = n757 | n2563 ;
  buffer buf_n758( .i (G161), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  assign n3015 = n756 & ~n2527 ;
  assign n3016 = n761 & ~n3015 ;
  assign n3017 = n3014 & n3016 ;
  assign n3018 = n754 | n758 ;
  buffer buf_n3019( .i (n3018), .o (n3019) );
  buffer buf_n3020( .i (n3019), .o (n3020) );
  assign n3021 = n862 & ~n3020 ;
  assign n3022 = n754 & ~n758 ;
  buffer buf_n3023( .i (n3022), .o (n3023) );
  buffer buf_n3024( .i (n3023), .o (n3024) );
  assign n3025 = n861 & n3024 ;
  assign n3026 = n3021 | n3025 ;
  assign n3027 = n3017 | n3026 ;
  assign n3028 = n846 & n3027 ;
  buffer buf_n2721( .i (n2720), .o (n2721) );
  buffer buf_n2722( .i (n2721), .o (n2722) );
  assign n3029 = n791 | n2722 ;
  buffer buf_n2624( .i (n2623), .o (n2624) );
  buffer buf_n2625( .i (n2624), .o (n2625) );
  assign n3030 = n790 & ~n2625 ;
  assign n3031 = n787 & ~n3030 ;
  assign n3032 = n3029 & n3031 ;
  buffer buf_n753( .i (G16), .o (n753) );
  assign n3033 = n753 & n2581 ;
  buffer buf_n568( .i (G14), .o (n568) );
  assign n3034 = n568 & ~n2585 ;
  assign n3035 = n3033 | n3034 ;
  assign n3036 = n3032 | n3035 ;
  buffer buf_n2752( .i (n2751), .o (n2752) );
  buffer buf_n2753( .i (n2752), .o (n2753) );
  assign n3037 = n791 | n2753 ;
  buffer buf_n2648( .i (n2647), .o (n2648) );
  buffer buf_n2649( .i (n2648), .o (n2649) );
  buffer buf_n2650( .i (n2649), .o (n2650) );
  buffer buf_n2651( .i (n2650), .o (n2651) );
  assign n3038 = n790 & ~n2651 ;
  assign n3039 = n787 & ~n3038 ;
  assign n3040 = n3037 & n3039 ;
  buffer buf_n842( .i (G6), .o (n842) );
  assign n3041 = n842 & ~n2585 ;
  buffer buf_n829( .i (G27), .o (n829) );
  assign n3042 = n829 & n2581 ;
  assign n3043 = n3041 | n3042 ;
  assign n3044 = n3040 | n3043 ;
  buffer buf_n2780( .i (n2779), .o (n2780) );
  buffer buf_n2781( .i (n2780), .o (n2781) );
  assign n3045 = n791 | n2781 ;
  buffer buf_n2669( .i (n2668), .o (n2669) );
  buffer buf_n2670( .i (n2669), .o (n2670) );
  buffer buf_n3046( .i (n789), .o (n3046) );
  assign n3047 = ~n2670 & n3046 ;
  assign n3048 = n787 & ~n3047 ;
  assign n3049 = n3045 & n3048 ;
  buffer buf_n828( .i (G26), .o (n828) );
  assign n3050 = n828 & n2581 ;
  buffer buf_n837( .i (G5), .o (n837) );
  assign n3051 = n837 & ~n2585 ;
  assign n3052 = n3050 | n3051 ;
  assign n3053 = n3049 | n3052 ;
  buffer buf_n2792( .i (n2791), .o (n2792) );
  buffer buf_n2793( .i (n2792), .o (n2793) );
  buffer buf_n3054( .i (n3046), .o (n3054) );
  assign n3055 = n2793 | n3054 ;
  buffer buf_n2542( .i (n2541), .o (n2542) );
  buffer buf_n2543( .i (n2542), .o (n2543) );
  assign n3056 = ~n2543 & n3046 ;
  buffer buf_n3057( .i (n786), .o (n3057) );
  assign n3058 = ~n3056 & n3057 ;
  assign n3059 = n3055 & n3058 ;
  buffer buf_n826( .i (G24), .o (n826) );
  buffer buf_n3060( .i (n2580), .o (n3060) );
  assign n3061 = n826 & n3060 ;
  buffer buf_n827( .i (G25), .o (n827) );
  buffer buf_n3062( .i (n2584), .o (n3062) );
  assign n3063 = n827 & ~n3062 ;
  assign n3064 = n3061 | n3063 ;
  assign n3065 = n3059 | n3064 ;
  assign n3066 = n795 | n2722 ;
  assign n3067 = n794 & ~n2625 ;
  assign n3068 = n799 & ~n3067 ;
  assign n3069 = n3066 & n3068 ;
  assign n3070 = n568 & ~n2681 ;
  assign n3071 = n753 & n2677 ;
  assign n3072 = n3070 | n3071 ;
  assign n3073 = n3069 | n3072 ;
  assign n3074 = n795 | n2753 ;
  assign n3075 = n794 & ~n2651 ;
  assign n3076 = n799 & ~n3075 ;
  assign n3077 = n3074 & n3076 ;
  assign n3078 = n829 & n2677 ;
  assign n3079 = n842 & ~n2681 ;
  assign n3080 = n3078 | n3079 ;
  assign n3081 = n3077 | n3080 ;
  assign n3082 = n795 | n2781 ;
  buffer buf_n3083( .i (n793), .o (n3083) );
  assign n3084 = ~n2670 & n3083 ;
  assign n3085 = n799 & ~n3084 ;
  assign n3086 = n3082 & n3085 ;
  assign n3087 = n837 & ~n2681 ;
  assign n3088 = n828 & n2677 ;
  assign n3089 = n3087 | n3088 ;
  assign n3090 = n3086 | n3089 ;
  buffer buf_n3091( .i (n3083), .o (n3091) );
  assign n3092 = n2793 | n3091 ;
  assign n3093 = ~n2543 & n3083 ;
  buffer buf_n3094( .i (n798), .o (n3094) );
  assign n3095 = ~n3093 & n3094 ;
  assign n3096 = n3092 & n3095 ;
  buffer buf_n3097( .i (n2676), .o (n3097) );
  assign n3098 = n826 & n3097 ;
  buffer buf_n3099( .i (n2680), .o (n3099) );
  assign n3100 = n827 & ~n3099 ;
  assign n3101 = n3098 | n3100 ;
  assign n3102 = n3096 | n3101 ;
  assign n3103 = n748 | n2721 ;
  assign n3104 = n747 & ~n2624 ;
  assign n3105 = n752 & ~n3104 ;
  assign n3106 = n3103 & n3105 ;
  buffer buf_n857( .i (G76), .o (n857) );
  assign n3107 = n857 & ~n3005 ;
  buffer buf_n867( .i (G86), .o (n867) );
  assign n3108 = n867 & n3009 ;
  assign n3109 = n3107 | n3108 ;
  assign n3110 = n3106 | n3109 ;
  assign n3111 = n846 & n3110 ;
  assign n3112 = n748 | n2792 ;
  assign n3113 = n747 & ~n2542 ;
  assign n3114 = n752 & ~n3113 ;
  assign n3115 = n3112 & n3114 ;
  buffer buf_n853( .i (G72), .o (n853) );
  assign n3116 = n853 & ~n3005 ;
  buffer buf_n863( .i (G82), .o (n863) );
  assign n3117 = n863 & n3009 ;
  assign n3118 = n3116 | n3117 ;
  assign n3119 = n3115 | n3118 ;
  assign n3120 = n846 & n3119 ;
  assign n3121 = n748 | n2780 ;
  buffer buf_n3122( .i (n746), .o (n3122) );
  assign n3123 = ~n2669 & n3122 ;
  assign n3124 = n752 & ~n3123 ;
  assign n3125 = n3121 & n3124 ;
  buffer buf_n851( .i (G70), .o (n851) );
  assign n3126 = n851 & ~n3005 ;
  buffer buf_n852( .i (G71), .o (n852) );
  assign n3127 = n852 & n3009 ;
  assign n3128 = n3126 | n3127 ;
  assign n3129 = n3125 | n3128 ;
  buffer buf_n3130( .i (n845), .o (n3130) );
  assign n3131 = n3129 & n3130 ;
  buffer buf_n3132( .i (n3122), .o (n3132) );
  assign n3133 = n2752 | n3132 ;
  assign n3134 = ~n2650 & n3122 ;
  buffer buf_n3135( .i (n751), .o (n3135) );
  assign n3136 = ~n3134 & n3135 ;
  assign n3137 = n3133 & n3136 ;
  buffer buf_n849( .i (G68), .o (n849) );
  buffer buf_n3138( .i (n3004), .o (n3138) );
  assign n3139 = n849 & ~n3138 ;
  buffer buf_n850( .i (G69), .o (n850) );
  buffer buf_n3140( .i (n3008), .o (n3140) );
  assign n3141 = n850 & n3140 ;
  assign n3142 = n3139 | n3141 ;
  assign n3143 = n3137 | n3142 ;
  assign n3144 = n3130 & n3143 ;
  assign n3145 = n757 | n2721 ;
  assign n3146 = n756 & ~n2624 ;
  assign n3147 = n761 & ~n3146 ;
  assign n3148 = n3145 & n3147 ;
  assign n3149 = n857 & ~n3020 ;
  assign n3150 = n867 & n3024 ;
  assign n3151 = n3149 | n3150 ;
  assign n3152 = n3148 | n3151 ;
  assign n3153 = n3130 & n3152 ;
  assign n3154 = n757 | n2792 ;
  assign n3155 = n756 & ~n2542 ;
  assign n3156 = n761 & ~n3155 ;
  assign n3157 = n3154 & n3156 ;
  assign n3158 = n853 & ~n3020 ;
  assign n3159 = n863 & n3024 ;
  assign n3160 = n3158 | n3159 ;
  assign n3161 = n3157 | n3160 ;
  assign n3162 = n3130 & n3161 ;
  assign n3163 = n757 | n2780 ;
  buffer buf_n3164( .i (n755), .o (n3164) );
  assign n3165 = ~n2669 & n3164 ;
  assign n3166 = n761 & ~n3165 ;
  assign n3167 = n3163 & n3166 ;
  assign n3168 = n851 & ~n3020 ;
  assign n3169 = n852 & n3024 ;
  assign n3170 = n3168 | n3169 ;
  assign n3171 = n3167 | n3170 ;
  buffer buf_n3172( .i (n845), .o (n3172) );
  assign n3173 = n3171 & n3172 ;
  buffer buf_n3174( .i (n3164), .o (n3174) );
  assign n3175 = n2752 | n3174 ;
  assign n3176 = ~n2650 & n3164 ;
  buffer buf_n3177( .i (n760), .o (n3177) );
  assign n3178 = ~n3176 & n3177 ;
  assign n3179 = n3175 & n3178 ;
  buffer buf_n3180( .i (n3019), .o (n3180) );
  assign n3181 = n849 & ~n3180 ;
  buffer buf_n3182( .i (n3023), .o (n3182) );
  assign n3183 = n850 & n3182 ;
  assign n3184 = n3181 | n3183 ;
  assign n3185 = n3179 | n3184 ;
  assign n3186 = n3172 & n3185 ;
  buffer buf_n782( .i (G171), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n780( .i (G170), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n2568( .i (n2567), .o (n2568) );
  buffer buf_n2569( .i (n2568), .o (n2569) );
  buffer buf_n2570( .i (n2569), .o (n2570) );
  buffer buf_n2571( .i (n2570), .o (n2571) );
  buffer buf_n2572( .i (n2571), .o (n2572) );
  assign n3187 = n781 & n2572 ;
  buffer buf_n843( .i (G61), .o (n843) );
  buffer buf_n2270( .i (n2269), .o (n2270) );
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2273( .i (n2272), .o (n2273) );
  buffer buf_n2274( .i (n2273), .o (n2274) );
  assign n3188 = ~n843 & n2274 ;
  assign n3189 = n843 & ~n2274 ;
  assign n3190 = n3188 | n3189 ;
  buffer buf_n3191( .i (n3190), .o (n3191) );
  assign n3194 = n781 | n3191 ;
  assign n3195 = ~n3187 & n3194 ;
  assign n3196 = n783 & ~n3195 ;
  assign n3197 = G178 & G62 ;
  buffer buf_n838( .i (G54), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  assign n3198 = n780 & ~n841 ;
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  assign n3199 = n780 | n1126 ;
  assign n3200 = ~n3198 & n3199 ;
  assign n3201 = n782 | n3200 ;
  assign n3202 = ~n3197 & n3201 ;
  assign n3203 = ~n3196 & n3202 ;
  buffer buf_n2573( .i (n2572), .o (n2573) );
  buffer buf_n2574( .i (n2573), .o (n2574) );
  buffer buf_n3192( .i (n3191), .o (n3192) );
  buffer buf_n3193( .i (n3192), .o (n3193) );
  assign n3204 = n2574 & n3193 ;
  assign n3205 = n2574 | n3193 ;
  assign n3206 = n3204 | ~n3205 ;
  assign n3207 = n838 & n2724 ;
  assign n3208 = n2567 & ~n2742 ;
  assign n3209 = ~n1121 & n2744 ;
  assign n3210 = n2747 & ~n3209 ;
  assign n3211 = ~n3208 & n3210 ;
  assign n3212 = n3207 | n3211 ;
  buffer buf_n3213( .i (n3212), .o (n3213) );
  inverter inv_n3928( .i (n3213), .o (n3928) );
  buffer buf_n3215( .i (n2723), .o (n3215) );
  assign n3216 = G52 & n3215 ;
  buffer buf_n3217( .i (n2663), .o (n3217) );
  buffer buf_n3218( .i (n3217), .o (n3218) );
  assign n3219 = n2974 | n3218 ;
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  assign n3220 = ~n1140 & n3217 ;
  buffer buf_n3221( .i (n2746), .o (n3221) );
  assign n3222 = ~n3220 & n3221 ;
  assign n3223 = n3219 & n3222 ;
  assign n3224 = n3216 | n3223 ;
  buffer buf_n3225( .i (n3224), .o (n3225) );
  inverter inv_n3929( .i (n3225), .o (n3929) );
  assign n3228 = G47 & n2723 ;
  assign n3229 = n2957 | n3217 ;
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  assign n3230 = n1065 & n2663 ;
  assign n3231 = n2746 & ~n3230 ;
  assign n3232 = n3229 & n3231 ;
  assign n3233 = n3228 | n3232 ;
  buffer buf_n3234( .i (n3233), .o (n3234) );
  inverter inv_n3930( .i (n3234), .o (n3930) );
  assign n3238 = G43 & n2723 ;
  assign n3239 = n2984 | n3217 ;
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n3240( .i (n801), .o (n3240) );
  assign n3241 = n1085 & n3240 ;
  assign n3242 = n2746 & ~n3241 ;
  assign n3243 = n3239 & n3242 ;
  assign n3244 = n3238 | n3243 ;
  buffer buf_n3245( .i (n3244), .o (n3245) );
  inverter inv_n3931( .i (n3245), .o (n3931) );
  assign n3249 = n739 & n997 ;
  assign n3250 = n1005 & n3249 ;
  assign n3251 = n999 & n3250 ;
  assign n3252 = ~n2385 & n3251 ;
  assign n3253 = ~n2424 & n3252 ;
  assign n3254 = ~n2842 & n3253 ;
  assign n3255 = ~n2882 & n3254 ;
  buffer buf_n2511( .i (n2510), .o (n2511) );
  assign n3256 = G46 & n2511 ;
  buffer buf_n805( .i (n804), .o (n805) );
  assign n3257 = ~n805 & n2894 ;
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  assign n3258 = n1296 & n3218 ;
  assign n3259 = n811 & ~n3258 ;
  assign n3260 = ~n3257 & n3259 ;
  assign n3261 = n3256 | n3260 ;
  buffer buf_n3262( .i (n3261), .o (n3262) );
  inverter inv_n3932( .i (n3262), .o (n3932) );
  buffer buf_n3264( .i (n2508), .o (n3264) );
  assign n3265 = G45 & n3264 ;
  buffer buf_n3266( .i (n3240), .o (n3266) );
  assign n3267 = n2920 & ~n3266 ;
  assign n3268 = n1225 & n3240 ;
  buffer buf_n3269( .i (n808), .o (n3269) );
  assign n3270 = ~n3268 & n3269 ;
  assign n3271 = ~n3267 & n3270 ;
  assign n3272 = n3265 | n3271 ;
  buffer buf_n3273( .i (n3272), .o (n3273) );
  inverter inv_n3933( .i (n3273), .o (n3933) );
  assign n3277 = G20 & n3264 ;
  assign n3278 = n2934 | n3266 ;
  assign n3279 = n1238 & n3240 ;
  assign n3280 = n3269 & ~n3279 ;
  assign n3281 = n3278 & n3280 ;
  assign n3282 = n3277 | n3281 ;
  buffer buf_n3283( .i (n3282), .o (n3283) );
  inverter inv_n3934( .i (n3283), .o (n3934) );
  assign n3287 = G44 & n3264 ;
  assign n3288 = n2902 | n3266 ;
  buffer buf_n3289( .i (n800), .o (n3289) );
  buffer buf_n3290( .i (n3289), .o (n3290) );
  assign n3291 = n1211 & n3290 ;
  assign n3292 = n3269 & ~n3291 ;
  assign n3293 = n3288 & n3292 ;
  assign n3294 = n3287 | n3293 ;
  buffer buf_n3295( .i (n3294), .o (n3295) );
  inverter inv_n3935( .i (n3295), .o (n3935) );
  buffer buf_n3263( .i (n3262), .o (n3263) );
  assign n3299 = n3091 | n3263 ;
  buffer buf_n3214( .i (n3213), .o (n3214) );
  assign n3300 = n3083 & ~n3214 ;
  assign n3301 = n3094 & ~n3300 ;
  assign n3302 = n3299 & n3301 ;
  buffer buf_n835( .i (G41), .o (n835) );
  assign n3303 = n835 & ~n3099 ;
  buffer buf_n836( .i (G42), .o (n836) );
  assign n3304 = n836 & n3097 ;
  assign n3305 = n3303 | n3304 ;
  assign n3306 = n3302 | n3305 ;
  assign n3307 = n3054 | n3263 ;
  assign n3308 = n3046 & ~n3214 ;
  assign n3309 = n3057 & ~n3308 ;
  assign n3310 = n3307 & n3309 ;
  assign n3311 = n835 & ~n3062 ;
  assign n3312 = n836 & n3060 ;
  assign n3313 = n3311 | n3312 ;
  assign n3314 = n3310 | n3313 ;
  buffer buf_n3226( .i (n3225), .o (n3226) );
  buffer buf_n3227( .i (n3226), .o (n3227) );
  assign n3315 = n3054 & ~n3227 ;
  buffer buf_n3274( .i (n3273), .o (n3274) );
  buffer buf_n3275( .i (n3274), .o (n3275) );
  buffer buf_n3316( .i (n789), .o (n3316) );
  assign n3317 = n3275 | n3316 ;
  assign n3318 = n3057 & n3317 ;
  assign n3319 = ~n3315 & n3318 ;
  buffer buf_n779( .i (G17), .o (n779) );
  assign n3320 = n779 & n3060 ;
  buffer buf_n813( .i (G18), .o (n813) );
  assign n3321 = n813 & ~n3062 ;
  assign n3322 = n3320 | n3321 ;
  assign n3323 = n3319 | n3322 ;
  buffer buf_n3235( .i (n3234), .o (n3235) );
  buffer buf_n3236( .i (n3235), .o (n3236) );
  buffer buf_n3237( .i (n3236), .o (n3237) );
  assign n3324 = n3054 & ~n3237 ;
  buffer buf_n3284( .i (n3283), .o (n3284) );
  buffer buf_n3285( .i (n3284), .o (n3285) );
  assign n3325 = n3285 | n3316 ;
  assign n3326 = n3057 & n3325 ;
  assign n3327 = ~n3324 & n3326 ;
  buffer buf_n832( .i (G39), .o (n832) );
  assign n3328 = n832 & n3060 ;
  buffer buf_n834( .i (G40), .o (n834) );
  assign n3329 = n834 & ~n3062 ;
  assign n3330 = n3328 | n3329 ;
  assign n3331 = n3327 | n3330 ;
  buffer buf_n3246( .i (n3245), .o (n3246) );
  buffer buf_n3247( .i (n3246), .o (n3247) );
  buffer buf_n3248( .i (n3247), .o (n3248) );
  buffer buf_n3332( .i (n3316), .o (n3332) );
  assign n3333 = ~n3248 & n3332 ;
  buffer buf_n3296( .i (n3295), .o (n3296) );
  buffer buf_n3297( .i (n3296), .o (n3297) );
  assign n3334 = n3297 | n3316 ;
  buffer buf_n3335( .i (n786), .o (n3335) );
  assign n3336 = n3334 & n3335 ;
  assign n3337 = ~n3333 & n3336 ;
  buffer buf_n831( .i (G36), .o (n831) );
  buffer buf_n3338( .i (n2580), .o (n3338) );
  assign n3339 = n831 & n3338 ;
  buffer buf_n716( .i (G15), .o (n716) );
  buffer buf_n3340( .i (n2584), .o (n3340) );
  assign n3341 = n716 & ~n3340 ;
  assign n3342 = n3339 | n3341 ;
  assign n3343 = n3337 | n3342 ;
  buffer buf_n3276( .i (n3275), .o (n3276) );
  assign n3344 = n3091 | n3276 ;
  buffer buf_n3345( .i (n793), .o (n3345) );
  assign n3346 = ~n3226 & n3345 ;
  assign n3347 = n3094 & ~n3346 ;
  assign n3348 = n3344 & n3347 ;
  assign n3349 = n779 & n3097 ;
  assign n3350 = n813 & ~n3099 ;
  assign n3351 = n3349 | n3350 ;
  assign n3352 = n3348 | n3351 ;
  buffer buf_n3286( .i (n3285), .o (n3286) );
  assign n3353 = n3091 | n3286 ;
  assign n3354 = ~n3236 & n3345 ;
  assign n3355 = n3094 & ~n3354 ;
  assign n3356 = n3353 & n3355 ;
  assign n3357 = n832 & n3097 ;
  assign n3358 = n834 & ~n3099 ;
  assign n3359 = n3357 | n3358 ;
  assign n3360 = n3356 | n3359 ;
  buffer buf_n3298( .i (n3297), .o (n3298) );
  buffer buf_n3361( .i (n3345), .o (n3361) );
  assign n3362 = n3298 | n3361 ;
  assign n3363 = ~n3247 & n3345 ;
  buffer buf_n3364( .i (n798), .o (n3364) );
  assign n3365 = ~n3363 & n3364 ;
  assign n3366 = n3362 & n3365 ;
  buffer buf_n3367( .i (n2676), .o (n3367) );
  assign n3368 = n831 & n3367 ;
  buffer buf_n3369( .i (n2680), .o (n3369) );
  assign n3370 = n716 & ~n3369 ;
  assign n3371 = n3368 | n3370 ;
  assign n3372 = n3366 | n3371 ;
  assign n3373 = n3132 & ~n3247 ;
  assign n3374 = n3122 | n3296 ;
  assign n3375 = n3135 & n3374 ;
  assign n3376 = ~n3373 & n3375 ;
  buffer buf_n858( .i (G77), .o (n858) );
  assign n3377 = n858 & ~n3138 ;
  buffer buf_n868( .i (G87), .o (n868) );
  assign n3378 = n868 & n3140 ;
  assign n3379 = n3377 | n3378 ;
  assign n3380 = n3376 | n3379 ;
  assign n3381 = n3172 & n3380 ;
  assign n3382 = n3132 & ~n3236 ;
  buffer buf_n3383( .i (n746), .o (n3383) );
  assign n3384 = n3284 | n3383 ;
  assign n3385 = n3135 & n3384 ;
  assign n3386 = ~n3382 & n3385 ;
  buffer buf_n856( .i (G75), .o (n856) );
  assign n3387 = n856 & ~n3138 ;
  buffer buf_n866( .i (G85), .o (n866) );
  assign n3388 = n866 & n3140 ;
  assign n3389 = n3387 | n3388 ;
  assign n3390 = n3386 | n3389 ;
  assign n3391 = n3172 & n3390 ;
  assign n3392 = n3132 & ~n3226 ;
  assign n3393 = n3274 | n3383 ;
  assign n3394 = n3135 & n3393 ;
  assign n3395 = ~n3392 & n3394 ;
  buffer buf_n865( .i (G84), .o (n865) );
  assign n3396 = n865 & n3140 ;
  buffer buf_n855( .i (G74), .o (n855) );
  assign n3397 = n855 & ~n3138 ;
  assign n3398 = n3396 | n3397 ;
  assign n3399 = n3395 | n3398 ;
  buffer buf_n3400( .i (n845), .o (n3400) );
  assign n3401 = n3399 & n3400 ;
  buffer buf_n3402( .i (n3383), .o (n3402) );
  assign n3403 = n3262 | n3402 ;
  assign n3404 = ~n3213 & n3383 ;
  buffer buf_n3405( .i (n751), .o (n3405) );
  assign n3406 = ~n3404 & n3405 ;
  assign n3407 = n3403 & n3406 ;
  buffer buf_n854( .i (G73), .o (n854) );
  buffer buf_n3408( .i (n3004), .o (n3408) );
  assign n3409 = n854 & ~n3408 ;
  buffer buf_n864( .i (G83), .o (n864) );
  buffer buf_n3410( .i (n3008), .o (n3410) );
  assign n3411 = n864 & n3410 ;
  assign n3412 = n3409 | n3411 ;
  assign n3413 = n3407 | n3412 ;
  assign n3414 = n3400 & n3413 ;
  assign n3415 = n3174 | n3297 ;
  assign n3416 = n3164 & ~n3246 ;
  assign n3417 = n3177 & ~n3416 ;
  assign n3418 = n3415 & n3417 ;
  assign n3419 = n858 & ~n3180 ;
  assign n3420 = n868 & n3182 ;
  assign n3421 = n3419 | n3420 ;
  assign n3422 = n3418 | n3421 ;
  assign n3423 = n3400 & n3422 ;
  assign n3424 = n3174 | n3285 ;
  buffer buf_n3425( .i (n755), .o (n3425) );
  assign n3426 = ~n3235 & n3425 ;
  assign n3427 = n3177 & ~n3426 ;
  assign n3428 = n3424 & n3427 ;
  assign n3429 = n866 & n3182 ;
  assign n3430 = n856 & ~n3180 ;
  assign n3431 = n3429 | n3430 ;
  assign n3432 = n3428 | n3431 ;
  assign n3433 = n3400 & n3432 ;
  assign n3434 = n3174 & ~n3226 ;
  assign n3435 = n3274 | n3425 ;
  assign n3436 = n3177 & n3435 ;
  assign n3437 = ~n3434 & n3436 ;
  assign n3438 = n855 & ~n3180 ;
  assign n3439 = n865 & n3182 ;
  assign n3440 = n3438 | n3439 ;
  assign n3441 = n3437 | n3440 ;
  buffer buf_n3442( .i (n844), .o (n3442) );
  buffer buf_n3443( .i (n3442), .o (n3443) );
  assign n3444 = n3441 & n3443 ;
  buffer buf_n3445( .i (n3425), .o (n3445) );
  assign n3446 = n3262 | n3445 ;
  assign n3447 = ~n3213 & n3425 ;
  buffer buf_n3448( .i (n760), .o (n3448) );
  assign n3449 = ~n3447 & n3448 ;
  assign n3450 = n3446 & n3449 ;
  buffer buf_n3451( .i (n3019), .o (n3451) );
  assign n3452 = n854 & ~n3451 ;
  buffer buf_n3453( .i (n3023), .o (n3453) );
  assign n3454 = n864 & n3453 ;
  assign n3455 = n3452 | n3454 ;
  assign n3456 = n3450 | n3455 ;
  assign n3457 = n3443 & n3456 ;
  assign n3458 = ~n665 & n2182 ;
  buffer buf_n3459( .i (n3458), .o (n3459) );
  buffer buf_n3460( .i (n3459), .o (n3460) );
  assign n3461 = n2226 & ~n3460 ;
  assign n3462 = n666 & ~n2233 ;
  assign n3463 = n3459 | n3462 ;
  assign n3464 = n2184 & ~n2241 ;
  assign n3465 = n3463 & ~n3464 ;
  assign n3466 = n3461 | n3465 ;
  buffer buf_n3467( .i (n3466), .o (n3467) );
  assign n3468 = n2797 & n3467 ;
  assign n3469 = n2797 | n3467 ;
  assign n3470 = ~n3468 & n3469 ;
  assign n3471 = n2947 & ~n3470 ;
  assign n3472 = ~n2187 & n2226 ;
  assign n3473 = n2194 & ~n3472 ;
  buffer buf_n3474( .i (n3473), .o (n3474) );
  assign n3475 = ~n2235 & n2261 ;
  buffer buf_n3476( .i (n2260), .o (n3476) );
  assign n3477 = n2235 & ~n3476 ;
  assign n3478 = n3475 | n3477 ;
  buffer buf_n3479( .i (n3478), .o (n3479) );
  assign n3480 = n3474 & n3479 ;
  assign n3481 = n3474 | n3479 ;
  assign n3482 = ~n3480 & n3481 ;
  assign n3483 = n2947 | n3482 ;
  assign n3484 = ~n3471 & n3483 ;
  buffer buf_n3485( .i (n3484), .o (n3485) );
  buffer buf_n3486( .i (n3485), .o (n3486) );
  buffer buf_n1987( .i (n1986), .o (n1987) );
  buffer buf_n1988( .i (n1987), .o (n1988) );
  buffer buf_n1989( .i (n1988), .o (n1989) );
  buffer buf_n1990( .i (n1989), .o (n1990) );
  buffer buf_n1991( .i (n1990), .o (n1991) );
  buffer buf_n1992( .i (n1991), .o (n1992) );
  assign n3487 = n1992 & ~n2628 ;
  buffer buf_n1998( .i (n1997), .o (n1998) );
  buffer buf_n1999( .i (n1998), .o (n1999) );
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n2001( .i (n2000), .o (n2001) );
  buffer buf_n2002( .i (n2001), .o (n2002) );
  assign n3488 = ~n2002 & n2628 ;
  assign n3489 = n3487 | n3488 ;
  buffer buf_n3490( .i (n3489), .o (n3490) );
  buffer buf_n762( .i (G162), .o (n762) );
  assign n3491 = n762 & n2060 ;
  assign n3492 = n2041 & n3491 ;
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  buffer buf_n2098( .i (n2097), .o (n2098) );
  assign n3493 = n762 | n2040 ;
  assign n3494 = n2098 & n3493 ;
  assign n3495 = ~n3492 & n3494 ;
  buffer buf_n3496( .i (n3495), .o (n3496) );
  assign n3497 = ~n2004 & n2336 ;
  assign n3498 = n2004 & ~n2336 ;
  assign n3499 = n3497 | n3498 ;
  buffer buf_n3500( .i (n3499), .o (n3500) );
  assign n3501 = n3496 & n3500 ;
  assign n3502 = n3496 | n3500 ;
  assign n3503 = ~n3501 & n3502 ;
  buffer buf_n3504( .i (n3503), .o (n3504) );
  assign n3505 = ~n2152 & n3504 ;
  assign n3506 = n2152 & ~n3504 ;
  assign n3507 = n3505 | n3506 ;
  buffer buf_n3508( .i (n3507), .o (n3508) );
  assign n3509 = n3490 & ~n3508 ;
  assign n3510 = ~n3490 & n3508 ;
  assign n3511 = n3509 | n3510 ;
  buffer buf_n3512( .i (n3511), .o (n3512) );
  buffer buf_n3513( .i (n3512), .o (n3513) );
  assign n3514 = n3486 | n3513 ;
  assign n3515 = n3485 & n3512 ;
  assign n3516 = n3290 | n3515 ;
  assign n3517 = n3514 & ~n3516 ;
  assign n3518 = ~n689 & n994 ;
  buffer buf_n3519( .i (n180), .o (n3519) );
  assign n3520 = n689 & ~n3519 ;
  assign n3521 = n3518 | n3520 ;
  buffer buf_n3522( .i (n3521), .o (n3522) );
  assign n3523 = ~n1152 & n3522 ;
  assign n3524 = n1152 & ~n3522 ;
  assign n3525 = n3523 | n3524 ;
  buffer buf_n3526( .i (n3525), .o (n3526) );
  assign n3527 = n182 | n348 ;
  assign n3528 = ~n186 & n348 ;
  assign n3529 = n3527 & ~n3528 ;
  assign n3530 = n677 & ~n3529 ;
  assign n3531 = n190 & n348 ;
  buffer buf_n3532( .i (n347), .o (n3532) );
  assign n3533 = n995 & ~n3532 ;
  assign n3534 = n3531 | n3533 ;
  assign n3535 = ~n677 & n3534 ;
  assign n3536 = n3530 | n3535 ;
  buffer buf_n3537( .i (n3536), .o (n3537) );
  assign n3538 = n3526 | n3537 ;
  assign n3539 = n3526 & n3537 ;
  assign n3540 = n3538 & ~n3539 ;
  buffer buf_n3541( .i (n3540), .o (n3541) );
  assign n3542 = n182 | n456 ;
  assign n3543 = ~n186 & n456 ;
  assign n3544 = n3542 & ~n3543 ;
  assign n3545 = n727 & ~n3544 ;
  assign n3546 = n190 & n456 ;
  buffer buf_n3547( .i (n455), .o (n3547) );
  assign n3548 = n995 & ~n3547 ;
  assign n3549 = n3546 | n3548 ;
  assign n3550 = ~n727 & n3549 ;
  assign n3551 = n3545 | n3550 ;
  buffer buf_n3552( .i (n3551), .o (n3552) );
  assign n3553 = n182 | n432 ;
  assign n3554 = ~n186 & n432 ;
  assign n3555 = n3553 & ~n3554 ;
  assign n3556 = n707 & ~n3555 ;
  assign n3557 = n190 & n432 ;
  buffer buf_n3558( .i (n431), .o (n3558) );
  assign n3559 = n995 & ~n3558 ;
  assign n3560 = n3557 | n3559 ;
  assign n3561 = ~n707 & n3560 ;
  assign n3562 = n3556 | n3561 ;
  buffer buf_n3563( .i (n3562), .o (n3563) );
  assign n3564 = n3552 | n3563 ;
  assign n3565 = n3552 & n3563 ;
  assign n3566 = n3564 & ~n3565 ;
  buffer buf_n3567( .i (n3566), .o (n3567) );
  assign n3568 = n3541 | n3567 ;
  assign n3569 = n3541 & n3567 ;
  assign n3570 = n3568 & ~n3569 ;
  buffer buf_n3571( .i (n3570), .o (n3571) );
  buffer buf_n3572( .i (n3571), .o (n3572) );
  assign n3573 = n1057 | n1077 ;
  assign n3574 = ~n1087 & n3573 ;
  buffer buf_n3575( .i (n3574), .o (n3575) );
  assign n3576 = ~n1112 & n1131 ;
  assign n3577 = n1142 | n3576 ;
  buffer buf_n3578( .i (n3577), .o (n3578) );
  assign n3579 = n3575 | n3578 ;
  assign n3580 = n3575 & n3578 ;
  assign n3581 = n3579 & ~n3580 ;
  buffer buf_n3582( .i (n3581), .o (n3582) );
  buffer buf_n3583( .i (n3582), .o (n3583) );
  assign n3584 = n3572 | n3583 ;
  assign n3585 = n3571 & n3582 ;
  assign n3586 = n3289 & ~n3585 ;
  assign n3587 = n3584 & n3586 ;
  assign n3588 = n3269 & ~n3587 ;
  assign n3589 = ~n3517 & n3588 ;
  buffer buf_n3590( .i (n3589), .o (n3590) );
  buffer buf_n3591( .i (n3590), .o (n3591) );
  buffer buf_n3592( .i (n3591), .o (n3592) );
  buffer buf_n3593( .i (n3592), .o (n3593) );
  buffer buf_n3594( .i (n3593), .o (n3594) );
  buffer buf_n3595( .i (n3594), .o (n3595) );
  buffer buf_n3596( .i (n3595), .o (n3596) );
  buffer buf_n2512( .i (n2511), .o (n2512) );
  buffer buf_n2513( .i (n2512), .o (n2513) );
  buffer buf_n2514( .i (n2513), .o (n2514) );
  buffer buf_n2515( .i (n2514), .o (n2515) );
  buffer buf_n2516( .i (n2515), .o (n2516) );
  assign n3597 = ~G51 & n2516 ;
  assign n3598 = ~n3596 & ~n3597 ;
  assign n3599 = n1425 & n1482 ;
  assign n3600 = n1422 | n1493 ;
  assign n3601 = ~n1508 & n3600 ;
  buffer buf_n3602( .i (n3601), .o (n3602) );
  buffer buf_n2427( .i (n2426), .o (n2427) );
  buffer buf_n2428( .i (n2427), .o (n2428) );
  buffer buf_n2429( .i (n2428), .o (n2429) );
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  assign n3603 = n1401 | n1480 ;
  assign n3604 = ~n2431 & n3603 ;
  assign n3605 = n3602 | n3604 ;
  assign n3606 = ~n3599 & n3605 ;
  buffer buf_n3607( .i (n3606), .o (n3607) );
  assign n3608 = n2441 & ~n3607 ;
  assign n3609 = ~n2441 & n3607 ;
  assign n3610 = n3608 | n3609 ;
  buffer buf_n3611( .i (n3610), .o (n3611) );
  buffer buf_n3612( .i (n3611), .o (n3612) );
  assign n3613 = n2705 | n3612 ;
  buffer buf_n741( .i (G157), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  assign n3614 = n2704 & n3611 ;
  assign n3615 = n744 | n3614 ;
  assign n3616 = n3613 & ~n3615 ;
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  assign n3617 = n1417 & n1472 ;
  assign n3618 = n1417 | n1482 ;
  assign n3619 = ~n3617 & n3618 ;
  buffer buf_n3620( .i (n3619), .o (n3620) );
  assign n3621 = n2728 & ~n3620 ;
  assign n3622 = ~n2728 & n3620 ;
  assign n3623 = n3621 | n3622 ;
  buffer buf_n3624( .i (n3623), .o (n3624) );
  buffer buf_n3625( .i (n3624), .o (n3625) );
  assign n3626 = n1364 | n3602 ;
  assign n3627 = n1364 & n3602 ;
  assign n3628 = n3626 & ~n3627 ;
  buffer buf_n3629( .i (n3628), .o (n3629) );
  assign n3630 = n1625 | n2698 ;
  buffer buf_n3631( .i (n3630), .o (n3631) );
  assign n3632 = n3629 & ~n3631 ;
  assign n3633 = ~n3629 & n3631 ;
  assign n3634 = n3632 | n3633 ;
  buffer buf_n3635( .i (n3634), .o (n3635) );
  buffer buf_n3636( .i (n3635), .o (n3636) );
  assign n3637 = n3625 & n3636 ;
  assign n3638 = n3624 | n3635 ;
  assign n3639 = n744 & n3638 ;
  assign n3640 = ~n3637 & n3639 ;
  assign n3641 = n3616 | n3640 ;
  buffer buf_n3642( .i (n3641), .o (n3642) );
  buffer buf_n3643( .i (n3642), .o (n3643) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  assign n3644 = n1947 | n2471 ;
  buffer buf_n3645( .i (n3644), .o (n3645) );
  buffer buf_n3646( .i (n3645), .o (n3646) );
  buffer buf_n3647( .i (n3646), .o (n3647) );
  buffer buf_n3648( .i (n3647), .o (n3648) );
  assign n3649 = ~n1765 & n3648 ;
  assign n3650 = n1784 & ~n3649 ;
  buffer buf_n3651( .i (n3650), .o (n3651) );
  assign n3652 = n1710 | n1845 ;
  assign n3653 = n1710 & n1845 ;
  assign n3654 = n3652 & ~n3653 ;
  buffer buf_n3655( .i (n3654), .o (n3655) );
  buffer buf_n3656( .i (n3655), .o (n3656) );
  buffer buf_n3657( .i (n3656), .o (n3657) );
  buffer buf_n2465( .i (n2464), .o (n2465) );
  buffer buf_n2466( .i (n2465), .o (n2466) );
  buffer buf_n2467( .i (n2466), .o (n2467) );
  buffer buf_n2468( .i (n2467), .o (n2468) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  assign n3658 = n1895 | n3645 ;
  assign n3659 = ~n2469 & n3658 ;
  buffer buf_n3660( .i (n3659), .o (n3660) );
  assign n3661 = n3657 & n3660 ;
  assign n3662 = n3657 | n3660 ;
  assign n3663 = ~n3661 & n3662 ;
  buffer buf_n3664( .i (n3663), .o (n3664) );
  assign n3665 = n3651 & n3664 ;
  assign n3666 = n3651 | n3664 ;
  assign n3667 = ~n3665 & n3666 ;
  buffer buf_n3668( .i (n3667), .o (n3668) );
  assign n3669 = n2455 & n3668 ;
  assign n3670 = n1763 | n2474 ;
  assign n3671 = ~n2487 & n3670 ;
  buffer buf_n3672( .i (n3671), .o (n3672) );
  buffer buf_n3673( .i (n3672), .o (n3673) );
  assign n3674 = ~n1786 & n1912 ;
  assign n3675 = n1786 & ~n1912 ;
  assign n3676 = n3674 | n3675 ;
  buffer buf_n3677( .i (n3676), .o (n3677) );
  assign n3678 = n3655 & ~n3677 ;
  assign n3679 = ~n3655 & n3677 ;
  assign n3680 = n3678 | n3679 ;
  buffer buf_n3681( .i (n3680), .o (n3681) );
  buffer buf_n3682( .i (n3681), .o (n3682) );
  assign n3683 = n3673 | n3682 ;
  assign n3684 = n3672 & n3681 ;
  assign n3685 = n2451 | n3684 ;
  assign n3686 = n3683 & ~n3685 ;
  buffer buf_n3687( .i (n3686), .o (n3687) );
  buffer buf_n3688( .i (n3687), .o (n3688) );
  assign n3689 = n741 | n3688 ;
  assign n3690 = n3669 | n3689 ;
  assign n3691 = n1636 | n2454 ;
  assign n3692 = n3668 & n3691 ;
  assign n3693 = ~n1636 & n3687 ;
  assign n3694 = n741 & ~n3693 ;
  assign n3695 = ~n3692 & n3694 ;
  assign n3696 = n3690 & ~n3695 ;
  buffer buf_n3697( .i (n3696), .o (n3697) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  assign n3698 = n1553 | n1607 ;
  assign n3699 = ~n1622 & n3698 ;
  buffer buf_n3700( .i (n3699), .o (n3700) );
  assign n3701 = n3697 & ~n3700 ;
  assign n3702 = ~n3697 & n3700 ;
  assign n3703 = n3701 | n3702 ;
  buffer buf_n3704( .i (n3703), .o (n3704) );
  buffer buf_n3705( .i (n3704), .o (n3705) );
  assign n3706 = ~n3643 & n3705 ;
  assign n3707 = n3642 & ~n3704 ;
  assign n3708 = n3266 | n3707 ;
  assign n3709 = n3706 | n3708 ;
  assign n3710 = n183 | n907 ;
  assign n3711 = ~n187 & n907 ;
  assign n3712 = n3710 & ~n3711 ;
  assign n3713 = n634 & ~n3712 ;
  assign n3714 = n191 & n907 ;
  buffer buf_n3715( .i (n906), .o (n3715) );
  assign n3716 = n996 & ~n3715 ;
  assign n3717 = n3714 | n3716 ;
  assign n3718 = ~n634 & n3717 ;
  assign n3719 = n3713 | n3718 ;
  buffer buf_n3720( .i (n3719), .o (n3720) );
  assign n3721 = n183 | n935 ;
  assign n3722 = ~n187 & n935 ;
  assign n3723 = n3721 & ~n3722 ;
  assign n3724 = n657 & ~n3723 ;
  assign n3725 = n191 & n935 ;
  buffer buf_n3726( .i (n934), .o (n3726) );
  assign n3727 = n996 & ~n3726 ;
  assign n3728 = n3725 | n3727 ;
  assign n3729 = ~n657 & n3728 ;
  assign n3730 = n3724 | n3729 ;
  buffer buf_n3731( .i (n3730), .o (n3731) );
  assign n3732 = n3720 & ~n3731 ;
  assign n3733 = ~n3720 & n3731 ;
  assign n3734 = n3732 | n3733 ;
  buffer buf_n3735( .i (n3734), .o (n3735) );
  buffer buf_n3736( .i (n3519), .o (n3736) );
  buffer buf_n3737( .i (n3736), .o (n3737) );
  assign n3738 = n962 | n3737 ;
  buffer buf_n3739( .i (n184), .o (n3739) );
  buffer buf_n3740( .i (n3739), .o (n3740) );
  buffer buf_n3741( .i (n3740), .o (n3741) );
  assign n3742 = n962 & ~n3741 ;
  assign n3743 = n3738 & ~n3742 ;
  assign n3744 = n583 & ~n3743 ;
  buffer buf_n3745( .i (n189), .o (n3745) );
  buffer buf_n3746( .i (n3745), .o (n3746) );
  assign n3747 = n962 & n3746 ;
  buffer buf_n3748( .i (n961), .o (n3748) );
  buffer buf_n3749( .i (n993), .o (n3749) );
  buffer buf_n3750( .i (n3749), .o (n3750) );
  buffer buf_n3751( .i (n3750), .o (n3751) );
  assign n3752 = ~n3748 & n3751 ;
  assign n3753 = n3747 | n3752 ;
  assign n3754 = ~n583 & n3753 ;
  assign n3755 = n3744 | n3754 ;
  buffer buf_n3756( .i (n3755), .o (n3756) );
  assign n3757 = n1287 & n3756 ;
  assign n3758 = n1287 | n3756 ;
  assign n3759 = ~n3757 & n3758 ;
  buffer buf_n3760( .i (n3759), .o (n3760) );
  assign n3761 = ~n3735 & n3760 ;
  assign n3762 = n3735 & ~n3760 ;
  assign n3763 = n3761 | n3762 ;
  buffer buf_n3764( .i (n3763), .o (n3764) );
  buffer buf_n3765( .i (n3764), .o (n3765) );
  assign n3766 = n246 | n3737 ;
  assign n3767 = n246 & ~n3741 ;
  assign n3768 = n3766 & ~n3767 ;
  assign n3769 = n559 & ~n3768 ;
  assign n3770 = n246 & n3746 ;
  buffer buf_n3771( .i (n245), .o (n3771) );
  assign n3772 = n3751 & ~n3771 ;
  assign n3773 = n3770 | n3772 ;
  assign n3774 = ~n559 & n3773 ;
  assign n3775 = n3769 | n3774 ;
  buffer buf_n3776( .i (n3775), .o (n3776) );
  assign n3777 = n222 | n3737 ;
  assign n3778 = n222 & ~n3741 ;
  assign n3779 = n3777 & ~n3778 ;
  assign n3780 = n539 & ~n3779 ;
  assign n3781 = n222 & n3746 ;
  buffer buf_n3782( .i (n221), .o (n3782) );
  assign n3783 = n3751 & ~n3782 ;
  assign n3784 = n3781 | n3783 ;
  assign n3785 = ~n539 & n3784 ;
  assign n3786 = n3780 | n3785 ;
  buffer buf_n3787( .i (n3786), .o (n3787) );
  assign n3788 = n3776 & n3787 ;
  assign n3789 = n3776 | n3787 ;
  assign n3790 = ~n3788 & n3789 ;
  buffer buf_n3791( .i (n3790), .o (n3791) );
  assign n3792 = n984 | n3737 ;
  assign n3793 = n984 & ~n3741 ;
  assign n3794 = n3792 & ~n3793 ;
  assign n3795 = n600 & ~n3794 ;
  assign n3796 = n984 & n3746 ;
  buffer buf_n3797( .i (n983), .o (n3797) );
  assign n3798 = n3751 & ~n3797 ;
  assign n3799 = n3796 | n3798 ;
  assign n3800 = ~n600 & n3799 ;
  assign n3801 = n3795 | n3800 ;
  buffer buf_n3802( .i (n3801), .o (n3802) );
  assign n3803 = n180 | n267 ;
  assign n3804 = ~n184 & n267 ;
  assign n3805 = n3803 & ~n3804 ;
  assign n3806 = n499 & ~n3805 ;
  assign n3807 = n188 & n267 ;
  buffer buf_n3808( .i (n266), .o (n3808) );
  assign n3809 = n993 & ~n3808 ;
  assign n3810 = n3807 | n3809 ;
  assign n3811 = ~n499 & n3810 ;
  assign n3812 = n3806 | n3811 ;
  buffer buf_n3813( .i (n3812), .o (n3813) );
  assign n3814 = n180 | n199 ;
  assign n3815 = ~n184 & n199 ;
  assign n3816 = n3814 & ~n3815 ;
  assign n3817 = n517 & ~n3816 ;
  assign n3818 = n188 & n199 ;
  buffer buf_n3819( .i (n198), .o (n3819) );
  assign n3820 = n993 & ~n3819 ;
  assign n3821 = n3818 | n3820 ;
  assign n3822 = ~n517 & n3821 ;
  assign n3823 = n3817 | n3822 ;
  buffer buf_n3824( .i (n3823), .o (n3824) );
  assign n3825 = n3813 & n3824 ;
  assign n3826 = n3813 | n3824 ;
  assign n3827 = ~n3825 & n3826 ;
  buffer buf_n3828( .i (n3827), .o (n3828) );
  assign n3829 = n3802 & ~n3828 ;
  assign n3830 = ~n3802 & n3828 ;
  assign n3831 = n3829 | n3830 ;
  buffer buf_n3832( .i (n3831), .o (n3832) );
  assign n3833 = ~n3791 & n3832 ;
  assign n3834 = n3791 & ~n3832 ;
  assign n3835 = n3833 | n3834 ;
  buffer buf_n3836( .i (n3835), .o (n3836) );
  buffer buf_n3837( .i (n3836), .o (n3837) );
  assign n3838 = ~n3765 & n3837 ;
  assign n3839 = n3764 & ~n3836 ;
  assign n3840 = n3290 & ~n3839 ;
  assign n3841 = ~n3838 & n3840 ;
  assign n3842 = n3221 & ~n3841 ;
  assign n3843 = n3709 & n3842 ;
  buffer buf_n3844( .i (n3843), .o (n3844) );
  buffer buf_n3845( .i (n3844), .o (n3845) );
  buffer buf_n3846( .i (n3845), .o (n3846) );
  buffer buf_n3847( .i (n3846), .o (n3847) );
  buffer buf_n3848( .i (n3847), .o (n3848) );
  buffer buf_n3849( .i (n3848), .o (n3849) );
  assign n3850 = ~G49 & n2516 ;
  assign n3851 = ~n3849 & ~n3850 ;
  buffer buf_n812( .i (n811), .o (n812) );
  assign n3852 = G38 & ~n812 ;
  assign n3853 = n3844 | n3852 ;
  buffer buf_n3854( .i (n3853), .o (n3854) );
  buffer buf_n3855( .i (n3854), .o (n3855) );
  assign n3856 = n3332 | n3855 ;
  assign n3857 = G37 & ~n811 ;
  assign n3858 = n3590 | n3857 ;
  buffer buf_n3859( .i (n3858), .o (n3859) );
  buffer buf_n3860( .i (n3859), .o (n3860) );
  buffer buf_n3861( .i (n789), .o (n3861) );
  assign n3862 = ~n3860 & n3861 ;
  assign n3863 = n3335 & ~n3862 ;
  assign n3864 = n3856 & n3863 ;
  buffer buf_n825( .i (G23), .o (n825) );
  assign n3865 = n825 & ~n3340 ;
  buffer buf_n833( .i (G4), .o (n833) );
  assign n3866 = n833 & n3338 ;
  assign n3867 = n3865 | n3866 ;
  assign n3868 = n3864 | n3867 ;
  assign n3869 = n3361 | n3855 ;
  buffer buf_n3870( .i (n793), .o (n3870) );
  assign n3871 = ~n3860 & n3870 ;
  assign n3872 = n3364 & ~n3871 ;
  assign n3873 = n3869 & n3872 ;
  assign n3874 = n825 & ~n3369 ;
  assign n3875 = n833 & n3367 ;
  assign n3876 = n3874 | n3875 ;
  assign n3877 = n3873 | n3876 ;
  assign n3878 = n3402 | n3854 ;
  buffer buf_n3879( .i (n746), .o (n3879) );
  assign n3880 = ~n3859 & n3879 ;
  assign n3881 = n3405 & ~n3880 ;
  assign n3882 = n3878 & n3881 ;
  buffer buf_n860( .i (G79), .o (n860) );
  assign n3883 = n860 & ~n3408 ;
  buffer buf_n859( .i (G78), .o (n859) );
  assign n3884 = n859 & n3410 ;
  assign n3885 = n3883 | n3884 ;
  assign n3886 = n3882 | n3885 ;
  assign n3887 = ~n3443 | ~n3886 ;
  assign n3888 = n3445 | n3854 ;
  buffer buf_n3889( .i (n755), .o (n3889) );
  assign n3890 = ~n3859 & n3889 ;
  assign n3891 = n3448 & ~n3890 ;
  assign n3892 = n3888 & n3891 ;
  assign n3893 = n860 & ~n3451 ;
  assign n3894 = n859 & n3453 ;
  assign n3895 = n3893 | n3894 ;
  assign n3896 = n3892 | n3895 ;
  assign n3897 = ~n3443 | ~n3896 ;
  assign G5193 = n3898 ;
  assign G5194 = n3899 ;
  assign G5195 = n3900 ;
  assign G5196 = n736 ;
  assign G5197 = n3901 ;
  assign G5198 = n3902 ;
  assign G5199 = n999 ;
  assign G5200 = n3903 ;
  assign G5201 = n736 ;
  assign G5202 = n736 ;
  assign G5203 = n3904 ;
  assign G5204 = n3905 ;
  assign G5205 = n1000 ;
  assign G5206 = n3906 ;
  assign G5207 = n3907 ;
  assign G5208 = n3908 ;
  assign G5209 = n3909 ;
  assign G5210 = n1001 ;
  assign G5211 = n1002 ;
  assign G5212 = n1003 ;
  assign G5213 = n3910 ;
  assign G5214 = n844 ;
  assign G5215 = n847 ;
  assign G5216 = n179 ;
  assign G5217 = n737 ;
  assign G5218 = n299 ;
  assign G5219 = n737 ;
  assign G5220 = n1011 ;
  assign G5221 = n3913 ;
  assign G5222 = n3911 ;
  assign G5223 = n3911 ;
  assign G5224 = n3911 ;
  assign G5225 = n3911 ;
  assign G5226 = n3912 ;
  assign G5227 = n3912 ;
  assign G5228 = n1015 ;
  assign G5229 = n1020 ;
  assign G5230 = n1020 ;
  assign G5231 = n1021 ;
  assign G5232 = n1026 ;
  assign G5233 = n1032 ;
  assign G5234 = n1038 ;
  assign G5235 = n1045 ;
  assign G5236 = n1198 ;
  assign G5237 = n1328 ;
  assign G5238 = n1966 ;
  assign G5239 = n2353 ;
  assign G5240 = n2353 ;
  assign G5241 = n1966 ;
  assign G5242 = n3914 ;
  assign G5243 = n3915 ;
  assign G5244 = n2503 ;
  assign G5245 = n2505 ;
  assign G5246 = n2503 ;
  assign G5247 = n2505 ;
  assign G5248 = n3916 ;
  assign G5249 = n3917 ;
  assign G5250 = n3918 ;
  assign G5251 = n2567 ;
  assign G5252 = n2588 ;
  assign G5253 = n3919 ;
  assign G5254 = n3920 ;
  assign G5255 = n3921 ;
  assign G5256 = n2684 ;
  assign G5257 = n3922 ;
  assign G5258 = n3923 ;
  assign G5259 = n3924 ;
  assign G5260 = n3925 ;
  assign G5261 = n3926 ;
  assign G5262 = n3927 ;
  assign G5263 = n2942 ;
  assign G5264 = n2998 ;
  assign G5265 = n3013 ;
  assign G5266 = n3028 ;
  assign G5267 = n3036 ;
  assign G5268 = n3044 ;
  assign G5269 = n3053 ;
  assign G5270 = n3065 ;
  assign G5271 = n3073 ;
  assign G5272 = n3081 ;
  assign G5273 = n3090 ;
  assign G5274 = n3102 ;
  assign G5275 = n3111 ;
  assign G5276 = n3120 ;
  assign G5277 = n3131 ;
  assign G5278 = n3144 ;
  assign G5279 = n3153 ;
  assign G5280 = n3162 ;
  assign G5281 = n3173 ;
  assign G5282 = n3186 ;
  assign G5283 = n3203 ;
  assign G5284 = n3206 ;
  assign G5285 = n3928 ;
  assign G5286 = n3929 ;
  assign G5287 = n3930 ;
  assign G5288 = n3931 ;
  assign G5289 = n3255 ;
  assign G5290 = n3932 ;
  assign G5291 = n3933 ;
  assign G5292 = n3934 ;
  assign G5293 = n3935 ;
  assign G5294 = n3306 ;
  assign G5295 = n3314 ;
  assign G5296 = n3323 ;
  assign G5297 = n3331 ;
  assign G5298 = n3343 ;
  assign G5299 = n3352 ;
  assign G5300 = n3360 ;
  assign G5301 = n3372 ;
  assign G5302 = n3381 ;
  assign G5303 = n3391 ;
  assign G5304 = n3401 ;
  assign G5305 = n3414 ;
  assign G5306 = n3423 ;
  assign G5307 = n3433 ;
  assign G5308 = n3444 ;
  assign G5309 = n3457 ;
  assign G5310 = n3598 ;
  assign G5311 = n3851 ;
  assign G5312 = n3868 ;
  assign G5313 = n3877 ;
  assign G5314 = n3887 ;
  assign G5315 = n3897 ;
endmodule
