module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( b_4_ , a_1_ , a_2_ , b_1_ , b_7_ , a_6_ , a_4_ , b_2_ , a_7_ , a_5_ , b_5_ , b_3_ , b_6_ , b_0_ , a_3_ , a_0_ , s_1_ , s_8_ , s_3_ , s_5_ , s_9_ , s_2_ , s_11_ , s_15_ , s_4_ , s_10_ , s_14_ , s_7_ , s_13_ , s_12_ , s_6_ , s_0_ );
  input b_4_ , a_1_ , a_2_ , b_1_ , b_7_ , a_6_ , a_4_ , b_2_ , a_7_ , a_5_ , b_5_ , b_3_ , b_6_ , b_0_ , a_3_ , a_0_ ;
  output s_1_ , s_8_ , s_3_ , s_5_ , s_9_ , s_2_ , s_11_ , s_15_ , s_4_ , s_10_ , s_14_ , s_7_ , s_13_ , s_12_ , s_6_ , s_0_ ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 ;
  assign n17 = a_1_ & b_0_ ;
  buffer buf_n18( .i (n17), .o (n18) );
  assign n19 = b_1_ & a_0_ ;
  buffer buf_n20( .i (n19), .o (n20) );
  assign n21 = n18 & n20 ;
  buffer buf_n22( .i (n21), .o (n22) );
  assign n23 = n18 | n20 ;
  buffer buf_n24( .i (n23), .o (n24) );
  assign n25 = ~n22 & n24 ;
  assign n26 = a_1_ & b_6_ ;
  buffer buf_n27( .i (n26), .o (n27) );
  assign n28 = b_4_ & a_2_ ;
  buffer buf_n29( .i (n28), .o (n29) );
  assign n30 = b_3_ & a_3_ ;
  buffer buf_n31( .i (n30), .o (n31) );
  assign n32 = n29 & n31 ;
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  assign n38 = a_1_ & b_5_ ;
  buffer buf_n39( .i (n38), .o (n39) );
  assign n40 = n29 | n31 ;
  buffer buf_n41( .i (n40), .o (n41) );
  assign n42 = ~n33 & n41 ;
  buffer buf_n43( .i (n42), .o (n43) );
  assign n44 = n39 & n43 ;
  buffer buf_n45( .i (n44), .o (n45) );
  assign n46 = n37 | n45 ;
  buffer buf_n47( .i (n46), .o (n47) );
  assign n48 = n27 & n47 ;
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  assign n54 = b_7_ & a_0_ ;
  buffer buf_n55( .i (n54), .o (n55) );
  assign n56 = n27 | n47 ;
  buffer buf_n57( .i (n56), .o (n57) );
  assign n58 = ~n49 & n57 ;
  buffer buf_n59( .i (n58), .o (n59) );
  assign n60 = n55 & n59 ;
  buffer buf_n61( .i (n60), .o (n61) );
  assign n62 = n53 | n61 ;
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  assign n72 = a_1_ & b_7_ ;
  buffer buf_n73( .i (n72), .o (n73) );
  assign n74 = a_2_ & b_6_ ;
  buffer buf_n75( .i (n74), .o (n75) );
  assign n76 = b_4_ & a_3_ ;
  buffer buf_n77( .i (n76), .o (n77) );
  assign n78 = a_4_ & b_3_ ;
  buffer buf_n79( .i (n78), .o (n79) );
  assign n80 = n77 & n79 ;
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  assign n86 = n77 | n79 ;
  buffer buf_n87( .i (n86), .o (n87) );
  assign n88 = ~n81 & n87 ;
  buffer buf_n89( .i (n88), .o (n89) );
  assign n90 = a_2_ & b_5_ ;
  buffer buf_n91( .i (n90), .o (n91) );
  assign n92 = n89 & n91 ;
  buffer buf_n93( .i (n92), .o (n93) );
  assign n94 = n85 | n93 ;
  buffer buf_n95( .i (n94), .o (n95) );
  assign n96 = n75 & n95 ;
  buffer buf_n97( .i (n96), .o (n97) );
  assign n102 = n75 | n95 ;
  buffer buf_n103( .i (n102), .o (n103) );
  assign n104 = ~n97 & n103 ;
  buffer buf_n105( .i (n104), .o (n105) );
  assign n106 = n73 & n105 ;
  buffer buf_n107( .i (n106), .o (n107) );
  assign n108 = n73 | n105 ;
  buffer buf_n109( .i (n108), .o (n109) );
  assign n110 = ~n107 & n109 ;
  buffer buf_n111( .i (n110), .o (n111) );
  assign n112 = b_5_ & a_3_ ;
  buffer buf_n113( .i (n112), .o (n113) );
  assign n114 = b_4_ & a_4_ ;
  buffer buf_n115( .i (n114), .o (n115) );
  assign n116 = a_5_ & b_3_ ;
  buffer buf_n117( .i (n116), .o (n117) );
  assign n118 = n115 & n117 ;
  buffer buf_n119( .i (n118), .o (n119) );
  assign n124 = n115 | n117 ;
  buffer buf_n125( .i (n124), .o (n125) );
  assign n126 = ~n119 & n125 ;
  buffer buf_n127( .i (n126), .o (n127) );
  assign n128 = n113 & n127 ;
  buffer buf_n129( .i (n128), .o (n129) );
  assign n130 = n113 | n127 ;
  buffer buf_n131( .i (n130), .o (n131) );
  assign n132 = ~n129 & n131 ;
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  assign n139 = b_1_ & a_6_ ;
  buffer buf_n140( .i (n139), .o (n140) );
  assign n145 = a_7_ & b_0_ ;
  buffer buf_n146( .i (n145), .o (n146) );
  assign n147 = n140 & n146 ;
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  assign n153 = b_2_ & a_5_ ;
  buffer buf_n154( .i (n153), .o (n154) );
  assign n155 = n140 | n146 ;
  buffer buf_n156( .i (n155), .o (n156) );
  assign n157 = ~n148 & n156 ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n159 = n154 & n158 ;
  buffer buf_n160( .i (n159), .o (n160) );
  assign n161 = n152 | n160 ;
  buffer buf_n162( .i (n161), .o (n162) );
  assign n163 = b_1_ & a_7_ ;
  assign n164 = a_6_ & b_2_ ;
  assign n165 = n163 | n164 ;
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  assign n166 = b_2_ & a_7_ ;
  buffer buf_n167( .i (n166), .o (n167) );
  assign n168 = n144 & n167 ;
  buffer buf_n169( .i (n168), .o (n169) );
  assign n173 = n165 & ~n169 ;
  buffer buf_n174( .i (n173), .o (n174) );
  assign n175 = n162 & n174 ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n181 = n162 | n174 ;
  buffer buf_n182( .i (n181), .o (n182) );
  assign n183 = ~n176 & n182 ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n185 = n138 & n184 ;
  buffer buf_n186( .i (n185), .o (n186) );
  assign n187 = n138 | n184 ;
  buffer buf_n188( .i (n187), .o (n188) );
  assign n189 = ~n186 & n188 ;
  buffer buf_n190( .i (n189), .o (n190) );
  assign n191 = n154 | n158 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = ~n160 & n192 ;
  buffer buf_n194( .i (n193), .o (n194) );
  assign n195 = a_5_ & b_0_ ;
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  assign n198 = n140 & n197 ;
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  assign n204 = a_4_ & b_2_ ;
  buffer buf_n205( .i (n204), .o (n205) );
  assign n206 = b_1_ & a_5_ ;
  assign n207 = a_6_ & b_0_ ;
  assign n208 = n206 | n207 ;
  assign n209 = ~n199 & n208 ;
  buffer buf_n210( .i (n209), .o (n210) );
  assign n211 = n205 & n210 ;
  buffer buf_n212( .i (n211), .o (n212) );
  assign n213 = n203 | n212 ;
  buffer buf_n214( .i (n213), .o (n214) );
  assign n215 = n194 & n214 ;
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  assign n221 = n89 | n91 ;
  buffer buf_n222( .i (n221), .o (n222) );
  assign n223 = ~n93 & n222 ;
  buffer buf_n224( .i (n223), .o (n224) );
  assign n225 = n194 | n214 ;
  buffer buf_n226( .i (n225), .o (n226) );
  assign n227 = ~n216 & n226 ;
  buffer buf_n228( .i (n227), .o (n228) );
  assign n229 = n224 & n228 ;
  buffer buf_n230( .i (n229), .o (n230) );
  assign n231 = n220 | n230 ;
  buffer buf_n232( .i (n231), .o (n232) );
  assign n233 = n190 & n232 ;
  buffer buf_n234( .i (n233), .o (n234) );
  assign n239 = n190 | n232 ;
  buffer buf_n240( .i (n239), .o (n240) );
  assign n241 = ~n234 & n240 ;
  buffer buf_n242( .i (n241), .o (n242) );
  assign n243 = n111 & n242 ;
  buffer buf_n244( .i (n243), .o (n244) );
  assign n245 = n111 | n242 ;
  buffer buf_n246( .i (n245), .o (n246) );
  assign n247 = ~n244 & n246 ;
  buffer buf_n248( .i (n247), .o (n248) );
  assign n249 = n224 | n228 ;
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = ~n230 & n250 ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n253 = n205 | n210 ;
  buffer buf_n254( .i (n253), .o (n254) );
  assign n255 = ~n212 & n254 ;
  buffer buf_n256( .i (n255), .o (n256) );
  assign n257 = b_1_ & a_4_ ;
  buffer buf_n258( .i (n257), .o (n258) );
  assign n259 = n196 & n258 ;
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  assign n265 = b_2_ & a_3_ ;
  buffer buf_n266( .i (n265), .o (n266) );
  assign n267 = n196 | n258 ;
  buffer buf_n268( .i (n267), .o (n268) );
  assign n269 = ~n260 & n268 ;
  buffer buf_n270( .i (n269), .o (n270) );
  assign n271 = n266 & n270 ;
  buffer buf_n272( .i (n271), .o (n272) );
  assign n273 = n264 | n272 ;
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  assign n276 = n256 & n275 ;
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  assign n282 = n39 | n43 ;
  buffer buf_n283( .i (n282), .o (n283) );
  assign n284 = ~n45 & n283 ;
  buffer buf_n285( .i (n284), .o (n285) );
  assign n286 = n256 | n275 ;
  buffer buf_n287( .i (n286), .o (n287) );
  assign n288 = ~n277 & n287 ;
  buffer buf_n289( .i (n288), .o (n289) );
  assign n290 = n285 & n289 ;
  buffer buf_n291( .i (n290), .o (n291) );
  assign n292 = n281 | n291 ;
  buffer buf_n293( .i (n292), .o (n293) );
  assign n294 = n252 & n293 ;
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  assign n300 = n55 | n59 ;
  buffer buf_n301( .i (n300), .o (n301) );
  assign n302 = ~n61 & n301 ;
  buffer buf_n303( .i (n302), .o (n303) );
  assign n304 = n252 | n293 ;
  buffer buf_n305( .i (n304), .o (n305) );
  assign n306 = ~n295 & n305 ;
  buffer buf_n307( .i (n306), .o (n307) );
  assign n308 = n303 & n307 ;
  buffer buf_n309( .i (n308), .o (n309) );
  assign n310 = n299 | n309 ;
  buffer buf_n311( .i (n310), .o (n311) );
  assign n312 = n248 & n311 ;
  buffer buf_n313( .i (n312), .o (n313) );
  assign n318 = n248 | n311 ;
  buffer buf_n319( .i (n318), .o (n319) );
  assign n320 = ~n313 & n319 ;
  buffer buf_n321( .i (n320), .o (n321) );
  assign n322 = n71 & n321 ;
  buffer buf_n323( .i (n322), .o (n323) );
  assign n324 = n71 | n321 ;
  buffer buf_n325( .i (n324), .o (n325) );
  assign n326 = ~n323 & n325 ;
  buffer buf_n327( .i (n326), .o (n327) );
  assign n328 = n303 | n307 ;
  buffer buf_n329( .i (n328), .o (n329) );
  assign n330 = ~n309 & n329 ;
  buffer buf_n331( .i (n330), .o (n331) );
  assign n332 = n285 | n289 ;
  buffer buf_n333( .i (n332), .o (n333) );
  assign n334 = ~n291 & n333 ;
  buffer buf_n335( .i (n334), .o (n335) );
  assign n336 = n266 | n270 ;
  buffer buf_n337( .i (n336), .o (n337) );
  assign n338 = ~n272 & n337 ;
  buffer buf_n339( .i (n338), .o (n339) );
  assign n340 = a_4_ & b_0_ ;
  buffer buf_n341( .i (n340), .o (n341) );
  assign n342 = b_1_ & a_3_ ;
  buffer buf_n343( .i (n342), .o (n343) );
  assign n344 = n341 & n343 ;
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  assign n350 = a_2_ & b_2_ ;
  buffer buf_n351( .i (n350), .o (n351) );
  assign n352 = n341 | n343 ;
  buffer buf_n353( .i (n352), .o (n353) );
  assign n354 = ~n345 & n353 ;
  buffer buf_n355( .i (n354), .o (n355) );
  assign n356 = n351 & n355 ;
  buffer buf_n357( .i (n356), .o (n357) );
  assign n358 = n349 | n357 ;
  buffer buf_n359( .i (n358), .o (n359) );
  assign n360 = n339 & n359 ;
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  assign n366 = b_5_ & a_0_ ;
  buffer buf_n367( .i (n366), .o (n367) );
  assign n368 = b_4_ & a_1_ ;
  buffer buf_n369( .i (n368), .o (n369) );
  assign n370 = a_2_ & b_3_ ;
  buffer buf_n371( .i (n370), .o (n371) );
  assign n372 = n369 | n371 ;
  buffer buf_n373( .i (n372), .o (n373) );
  assign n374 = n369 & n371 ;
  buffer buf_n375( .i (n374), .o (n375) );
  assign n380 = n373 & ~n375 ;
  buffer buf_n381( .i (n380), .o (n381) );
  assign n382 = n367 & n381 ;
  buffer buf_n383( .i (n382), .o (n383) );
  assign n384 = n367 | n381 ;
  buffer buf_n385( .i (n384), .o (n385) );
  assign n386 = ~n383 & n385 ;
  buffer buf_n387( .i (n386), .o (n387) );
  assign n388 = n339 | n359 ;
  buffer buf_n389( .i (n388), .o (n389) );
  assign n390 = ~n361 & n389 ;
  buffer buf_n391( .i (n390), .o (n391) );
  assign n392 = n387 & n391 ;
  buffer buf_n393( .i (n392), .o (n393) );
  assign n394 = n365 | n393 ;
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  assign n397 = n335 & n396 ;
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  assign n403 = b_6_ & a_0_ ;
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  assign n405 = n379 | n383 ;
  buffer buf_n406( .i (n405), .o (n406) );
  assign n407 = n404 & n406 ;
  buffer buf_n408( .i (n407), .o (n408) );
  assign n424 = n404 | n406 ;
  buffer buf_n425( .i (n424), .o (n425) );
  assign n426 = ~n408 & n425 ;
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  assign n433 = n335 | n396 ;
  buffer buf_n434( .i (n433), .o (n434) );
  assign n435 = ~n398 & n434 ;
  buffer buf_n436( .i (n435), .o (n436) );
  assign n437 = n432 & n436 ;
  buffer buf_n438( .i (n437), .o (n438) );
  assign n439 = n402 | n438 ;
  buffer buf_n440( .i (n439), .o (n440) );
  assign n441 = n331 & n440 ;
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  assign n447 = n331 | n440 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = ~n442 & n448 ;
  buffer buf_n450( .i (n449), .o (n450) );
  assign n451 = n423 & n450 ;
  buffer buf_n452( .i (n451), .o (n452) );
  assign n453 = n446 | n452 ;
  buffer buf_n454( .i (n453), .o (n454) );
  assign n455 = n327 | n454 ;
  buffer buf_n456( .i (n455), .o (n456) );
  assign n457 = n327 & n454 ;
  buffer buf_n458( .i (n457), .o (n458) );
  assign n467 = n456 & ~n458 ;
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  assign n473 = n423 | n450 ;
  buffer buf_n474( .i (n473), .o (n474) );
  assign n475 = ~n452 & n474 ;
  buffer buf_n476( .i (n475), .o (n476) );
  assign n477 = n432 | n436 ;
  buffer buf_n478( .i (n477), .o (n478) );
  assign n479 = ~n438 & n478 ;
  buffer buf_n480( .i (n479), .o (n480) );
  assign n481 = n387 | n391 ;
  buffer buf_n482( .i (n481), .o (n482) );
  assign n483 = ~n393 & n482 ;
  buffer buf_n484( .i (n483), .o (n484) );
  assign n485 = n351 | n355 ;
  buffer buf_n486( .i (n485), .o (n486) );
  assign n487 = ~n357 & n486 ;
  buffer buf_n488( .i (n487), .o (n488) );
  assign n489 = a_2_ & b_1_ ;
  buffer buf_n490( .i (n489), .o (n490) );
  assign n491 = b_0_ & a_3_ ;
  buffer buf_n492( .i (n491), .o (n492) );
  assign n493 = n490 & n492 ;
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  assign n499 = a_1_ & b_2_ ;
  buffer buf_n500( .i (n499), .o (n500) );
  assign n501 = n490 | n492 ;
  buffer buf_n502( .i (n501), .o (n502) );
  assign n503 = ~n494 & n502 ;
  buffer buf_n504( .i (n503), .o (n504) );
  assign n505 = n500 & n504 ;
  buffer buf_n506( .i (n505), .o (n506) );
  assign n507 = n498 | n506 ;
  buffer buf_n508( .i (n507), .o (n508) );
  assign n509 = n488 & n508 ;
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  assign n515 = a_1_ & b_3_ ;
  assign n516 = b_4_ & a_0_ ;
  assign n517 = n515 | n516 ;
  assign n518 = b_3_ & a_0_ ;
  buffer buf_n519( .i (n518), .o (n519) );
  assign n528 = n369 & n519 ;
  buffer buf_n529( .i (n528), .o (n529) );
  assign n544 = n517 & ~n529 ;
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  assign n550 = n488 | n508 ;
  buffer buf_n551( .i (n550), .o (n551) );
  assign n552 = ~n510 & n551 ;
  buffer buf_n553( .i (n552), .o (n553) );
  assign n554 = n549 & n553 ;
  buffer buf_n555( .i (n554), .o (n555) );
  assign n556 = n514 | n555 ;
  buffer buf_n557( .i (n556), .o (n557) );
  assign n558 = n484 & n557 ;
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  assign n564 = n484 | n557 ;
  buffer buf_n565( .i (n564), .o (n565) );
  assign n566 = ~n559 & n565 ;
  buffer buf_n567( .i (n566), .o (n567) );
  assign n568 = n543 & n567 ;
  buffer buf_n569( .i (n568), .o (n569) );
  assign n570 = n563 | n569 ;
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  assign n573 = n480 & n572 ;
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  assign n581 = n476 & n580 ;
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  assign n587 = n476 | n580 ;
  buffer buf_n588( .i (n587), .o (n588) );
  assign n589 = ~n582 & n588 ;
  buffer buf_n590( .i (n589), .o (n590) );
  assign n591 = n480 | n572 ;
  buffer buf_n592( .i (n591), .o (n592) );
  assign n593 = ~n574 & n592 ;
  buffer buf_n594( .i (n593), .o (n594) );
  assign n595 = n543 | n567 ;
  buffer buf_n596( .i (n595), .o (n596) );
  assign n597 = ~n569 & n596 ;
  buffer buf_n598( .i (n597), .o (n598) );
  assign n599 = n549 | n553 ;
  buffer buf_n600( .i (n599), .o (n600) );
  assign n601 = ~n555 & n600 ;
  buffer buf_n602( .i (n601), .o (n602) );
  assign n603 = a_1_ & b_1_ ;
  buffer buf_n604( .i (n603), .o (n604) );
  assign n605 = a_2_ & b_0_ ;
  buffer buf_n606( .i (n605), .o (n606) );
  assign n607 = n604 & n606 ;
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  assign n613 = b_2_ & a_0_ ;
  buffer buf_n614( .i (n613), .o (n614) );
  assign n615 = n604 | n606 ;
  buffer buf_n616( .i (n615), .o (n616) );
  assign n617 = ~n608 & n616 ;
  buffer buf_n618( .i (n617), .o (n618) );
  assign n619 = n614 & n618 ;
  buffer buf_n620( .i (n619), .o (n620) );
  assign n621 = n612 | n620 ;
  buffer buf_n622( .i (n621), .o (n622) );
  assign n623 = n500 | n504 ;
  buffer buf_n624( .i (n623), .o (n624) );
  assign n625 = ~n506 & n624 ;
  buffer buf_n626( .i (n625), .o (n626) );
  assign n627 = n622 & n626 ;
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  assign n633 = n622 | n626 ;
  buffer buf_n634( .i (n633), .o (n634) );
  assign n635 = ~n628 & n634 ;
  buffer buf_n636( .i (n635), .o (n636) );
  assign n637 = n527 & n636 ;
  buffer buf_n638( .i (n637), .o (n638) );
  assign n639 = n632 | n638 ;
  buffer buf_n640( .i (n639), .o (n640) );
  assign n641 = n602 & n640 ;
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  assign n649 = n598 & n648 ;
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  assign n654 = n594 & n653 ;
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  assign n660 = n594 | n653 ;
  buffer buf_n661( .i (n660), .o (n661) );
  assign n662 = ~n655 & n661 ;
  buffer buf_n663( .i (n662), .o (n663) );
  assign n664 = n598 | n648 ;
  buffer buf_n665( .i (n664), .o (n665) );
  assign n666 = ~n650 & n665 ;
  buffer buf_n667( .i (n666), .o (n667) );
  assign n668 = n602 | n640 ;
  buffer buf_n669( .i (n668), .o (n669) );
  assign n670 = ~n642 & n669 ;
  buffer buf_n671( .i (n670), .o (n671) );
  assign n672 = n614 | n618 ;
  buffer buf_n673( .i (n672), .o (n673) );
  assign n674 = ~n620 & n673 ;
  buffer buf_n675( .i (n674), .o (n675) );
  assign n676 = n22 & n675 ;
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  assign n684 = n527 | n636 ;
  buffer buf_n685( .i (n684), .o (n685) );
  assign n686 = ~n638 & n685 ;
  buffer buf_n687( .i (n686), .o (n687) );
  assign n688 = n683 & n687 ;
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  assign n692 = n671 & n691 ;
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  assign n700 = n667 & n699 ;
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  assign n705 = n663 & n704 ;
  buffer buf_n706( .i (n705), .o (n706) );
  assign n707 = n659 | n706 ;
  buffer buf_n708( .i (n707), .o (n708) );
  assign n709 = n590 & n708 ;
  buffer buf_n710( .i (n709), .o (n710) );
  assign n711 = n586 | n710 ;
  buffer buf_n712( .i (n711), .o (n712) );
  assign n713 = n472 & n712 ;
  buffer buf_n714( .i (n713), .o (n714) );
  assign n715 = n472 | n712 ;
  buffer buf_n716( .i (n715), .o (n716) );
  assign n717 = ~n714 & n716 ;
  assign n718 = n683 | n687 ;
  buffer buf_n719( .i (n718), .o (n719) );
  assign n720 = ~n689 & n719 ;
  assign n721 = n667 | n699 ;
  buffer buf_n722( .i (n721), .o (n722) );
  assign n723 = ~n701 & n722 ;
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  assign n724 = n466 | n714 ;
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  assign n726 = n317 | n323 ;
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  assign n728 = n101 | n107 ;
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  assign n738 = a_2_ & b_7_ ;
  buffer buf_n739( .i (n738), .o (n739) );
  assign n740 = b_6_ & a_3_ ;
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  assign n742 = n123 | n129 ;
  buffer buf_n743( .i (n742), .o (n743) );
  assign n744 = n741 & n743 ;
  buffer buf_n745( .i (n744), .o (n745) );
  assign n750 = n741 | n743 ;
  buffer buf_n751( .i (n750), .o (n751) );
  assign n752 = ~n745 & n751 ;
  buffer buf_n753( .i (n752), .o (n753) );
  assign n754 = n739 & n753 ;
  buffer buf_n755( .i (n754), .o (n755) );
  assign n756 = n739 | n753 ;
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = ~n755 & n757 ;
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  assign n765 = a_4_ & b_5_ ;
  buffer buf_n766( .i (n765), .o (n766) );
  assign n767 = b_4_ & a_5_ ;
  assign n768 = a_6_ & b_3_ ;
  buffer buf_n769( .i (n768), .o (n769) );
  assign n770 = n767 | n769 ;
  buffer buf_n771( .i (n770), .o (n771) );
  assign n772 = b_4_ & a_6_ ;
  buffer buf_n773( .i (n772), .o (n773) );
  assign n774 = n117 & n773 ;
  buffer buf_n775( .i (n774), .o (n775) );
  assign n780 = n771 & ~n775 ;
  buffer buf_n781( .i (n780), .o (n781) );
  assign n782 = n766 & n781 ;
  buffer buf_n783( .i (n782), .o (n783) );
  assign n784 = n766 | n781 ;
  buffer buf_n785( .i (n784), .o (n785) );
  assign n786 = ~n783 & n785 ;
  buffer buf_n787( .i (n786), .o (n787) );
  assign n788 = ~n144 & n167 ;
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  assign n791 = n787 & n790 ;
  buffer buf_n792( .i (n791), .o (n792) );
  assign n793 = n787 | n790 ;
  buffer buf_n794( .i (n793), .o (n794) );
  assign n795 = ~n792 & n794 ;
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  assign n802 = n180 | n186 ;
  buffer buf_n803( .i (n802), .o (n803) );
  assign n804 = n801 & n803 ;
  buffer buf_n805( .i (n804), .o (n805) );
  assign n810 = n801 | n803 ;
  buffer buf_n811( .i (n810), .o (n811) );
  assign n812 = ~n805 & n811 ;
  buffer buf_n813( .i (n812), .o (n813) );
  assign n814 = n764 & n813 ;
  buffer buf_n815( .i (n814), .o (n815) );
  assign n816 = n764 | n813 ;
  buffer buf_n817( .i (n816), .o (n817) );
  assign n818 = ~n815 & n817 ;
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  assign n820 = n238 | n244 ;
  buffer buf_n821( .i (n820), .o (n821) );
  assign n822 = n819 & n821 ;
  buffer buf_n823( .i (n822), .o (n823) );
  assign n828 = n819 | n821 ;
  buffer buf_n829( .i (n828), .o (n829) );
  assign n830 = ~n823 & n829 ;
  buffer buf_n831( .i (n830), .o (n831) );
  assign n832 = n737 & n831 ;
  buffer buf_n833( .i (n832), .o (n833) );
  assign n834 = n737 | n831 ;
  buffer buf_n835( .i (n834), .o (n835) );
  assign n836 = ~n833 & n835 ;
  buffer buf_n837( .i (n836), .o (n837) );
  assign n838 = n727 & n837 ;
  buffer buf_n839( .i (n838), .o (n839) );
  assign n850 = n727 | n837 ;
  buffer buf_n851( .i (n850), .o (n851) );
  assign n863 = ~n839 & n851 ;
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  assign n873 = n725 | n872 ;
  assign n874 = n725 & n872 ;
  assign n875 = n873 & ~n874 ;
  assign n876 = n22 | n675 ;
  buffer buf_n877( .i (n876), .o (n877) );
  assign n878 = ~n677 & n877 ;
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  assign n879 = n779 | n783 ;
  buffer buf_n880( .i (n879), .o (n880) );
  assign n881 = a_4_ & b_6_ ;
  buffer buf_n882( .i (n881), .o (n882) );
  assign n883 = n880 & n882 ;
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  assign n889 = b_7_ & a_3_ ;
  buffer buf_n890( .i (n889), .o (n890) );
  assign n891 = n880 | n882 ;
  buffer buf_n892( .i (n891), .o (n892) );
  assign n893 = ~n884 & n892 ;
  buffer buf_n894( .i (n893), .o (n894) );
  assign n895 = n890 & n894 ;
  buffer buf_n896( .i (n895), .o (n896) );
  assign n897 = n888 | n896 ;
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  assign n907 = a_7_ & b_5_ ;
  buffer buf_n908( .i (n907), .o (n908) );
  assign n919 = n773 & n908 ;
  buffer buf_n920( .i (n919), .o (n920) );
  assign n921 = b_4_ & a_7_ ;
  buffer buf_n922( .i (n921), .o (n922) );
  assign n923 = a_6_ & b_5_ ;
  assign n924 = n922 | n923 ;
  buffer buf_n925( .i (n924), .o (n925) );
  assign n926 = ~n920 & n925 ;
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  assign n940 = b_7_ & a_4_ ;
  buffer buf_n941( .i (n940), .o (n941) );
  assign n942 = n769 & n922 ;
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  assign n948 = a_5_ & b_5_ ;
  buffer buf_n949( .i (n948), .o (n949) );
  assign n950 = a_7_ & b_3_ ;
  assign n951 = n773 | n950 ;
  buffer buf_n952( .i (n951), .o (n952) );
  assign n953 = ~n943 & n952 ;
  buffer buf_n954( .i (n953), .o (n954) );
  assign n955 = n949 & n954 ;
  buffer buf_n956( .i (n955), .o (n956) );
  assign n957 = n947 | n956 ;
  buffer buf_n958( .i (n957), .o (n958) );
  assign n959 = a_5_ & b_6_ ;
  buffer buf_n960( .i (n959), .o (n960) );
  assign n961 = n958 & n960 ;
  buffer buf_n962( .i (n961), .o (n962) );
  assign n967 = n958 | n960 ;
  buffer buf_n968( .i (n967), .o (n968) );
  assign n969 = ~n962 & n968 ;
  buffer buf_n970( .i (n969), .o (n970) );
  assign n971 = n941 & n970 ;
  buffer buf_n972( .i (n971), .o (n972) );
  assign n973 = n941 | n970 ;
  buffer buf_n974( .i (n973), .o (n974) );
  assign n975 = ~n972 & n974 ;
  buffer buf_n976( .i (n975), .o (n976) );
  assign n977 = n939 & n976 ;
  buffer buf_n978( .i (n977), .o (n978) );
  assign n979 = n939 | n976 ;
  buffer buf_n980( .i (n979), .o (n980) );
  assign n981 = ~n978 & n980 ;
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  assign n983 = n172 | n792 ;
  buffer buf_n984( .i (n983), .o (n984) );
  assign n985 = n949 | n954 ;
  buffer buf_n986( .i (n985), .o (n986) );
  assign n987 = ~n956 & n986 ;
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  assign n993 = n984 & n992 ;
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  assign n999 = n984 | n992 ;
  buffer buf_n1000( .i (n999), .o (n1000) );
  assign n1001 = ~n994 & n1000 ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  assign n1003 = n890 | n894 ;
  buffer buf_n1004( .i (n1003), .o (n1004) );
  assign n1005 = ~n896 & n1004 ;
  buffer buf_n1006( .i (n1005), .o (n1006) );
  assign n1007 = n1002 & n1006 ;
  buffer buf_n1008( .i (n1007), .o (n1008) );
  assign n1009 = n998 | n1008 ;
  buffer buf_n1010( .i (n1009), .o (n1010) );
  assign n1011 = n982 & n1010 ;
  buffer buf_n1012( .i (n1011), .o (n1012) );
  assign n1017 = n982 | n1010 ;
  buffer buf_n1018( .i (n1017), .o (n1018) );
  assign n1019 = ~n1012 & n1018 ;
  buffer buf_n1020( .i (n1019), .o (n1020) );
  assign n1021 = n906 & n1020 ;
  buffer buf_n1022( .i (n1021), .o (n1022) );
  assign n1023 = n906 | n1020 ;
  buffer buf_n1024( .i (n1023), .o (n1024) );
  assign n1025 = ~n1022 & n1024 ;
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  assign n1032 = n809 | n815 ;
  buffer buf_n1033( .i (n1032), .o (n1033) );
  assign n1034 = n1002 | n1006 ;
  buffer buf_n1035( .i (n1034), .o (n1035) );
  assign n1036 = ~n1008 & n1035 ;
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  assign n1043 = n1033 & n1042 ;
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  assign n1049 = n749 | n755 ;
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  assign n1064 = n1033 | n1042 ;
  buffer buf_n1065( .i (n1064), .o (n1065) );
  assign n1066 = ~n1044 & n1065 ;
  buffer buf_n1067( .i (n1066), .o (n1067) );
  assign n1068 = n1063 & n1067 ;
  buffer buf_n1069( .i (n1068), .o (n1069) );
  assign n1070 = n1048 | n1069 ;
  buffer buf_n1071( .i (n1070), .o (n1071) );
  assign n1072 = n1031 & n1071 ;
  buffer buf_n1073( .i (n1072), .o (n1073) );
  assign n1093 = n1031 | n1071 ;
  buffer buf_n1094( .i (n1093), .o (n1094) );
  assign n1095 = ~n1073 & n1094 ;
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  assign n1112 = n827 | n833 ;
  buffer buf_n1113( .i (n1112), .o (n1113) );
  assign n1114 = n1063 | n1067 ;
  buffer buf_n1115( .i (n1114), .o (n1115) );
  assign n1116 = ~n1069 & n1115 ;
  buffer buf_n1117( .i (n1116), .o (n1117) );
  assign n1118 = n1113 & n1117 ;
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  assign n1135 = n725 | n849 ;
  assign n1136 = n862 & n1135 ;
  buffer buf_n1137( .i (n1136), .o (n1137) );
  assign n1138 = n1113 | n1117 ;
  buffer buf_n1139( .i (n1138), .o (n1139) );
  assign n1140 = ~n1119 & n1139 ;
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  assign n1153 = n1137 & n1152 ;
  buffer buf_n1154( .i (n1153), .o (n1154) );
  assign n1155 = n1134 | n1154 ;
  buffer buf_n1156( .i (n1155), .o (n1156) );
  assign n1157 = n1111 | n1156 ;
  buffer buf_n1158( .i (n1157), .o (n1158) );
  assign n1159 = n1111 & n1156 ;
  buffer buf_n1160( .i (n1159), .o (n1160) );
  assign n1161 = n1158 & ~n1160 ;
  assign n1162 = a_6_ & b_6_ ;
  buffer buf_n1163( .i (n1162), .o (n1163) );
  assign n1164 = b_7_ & a_7_ ;
  buffer buf_n1165( .i (n1164), .o (n1165) );
  assign n1166 = n1163 & n1165 ;
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  assign n1186 = ~n1163 & n1165 ;
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  assign n1204 = a_7_ & b_6_ ;
  assign n1205 = b_7_ & a_6_ ;
  assign n1206 = n1204 | n1205 ;
  assign n1207 = ~n1167 & n1206 ;
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  assign n1215 = b_7_ & a_5_ ;
  buffer buf_n1216( .i (n1215), .o (n1216) );
  assign n1217 = b_6_ & n920 ;
  buffer buf_n1218( .i (n1217), .o (n1218) );
  assign n1223 = n920 | n1163 ;
  buffer buf_n1224( .i (n1223), .o (n1224) );
  assign n1225 = ~n1218 & n1224 ;
  buffer buf_n1226( .i (n1225), .o (n1226) );
  assign n1227 = n1216 & n1226 ;
  buffer buf_n1228( .i (n1227), .o (n1228) );
  assign n1229 = n1216 | n1226 ;
  buffer buf_n1230( .i (n1229), .o (n1230) );
  assign n1231 = ~n1228 & n1230 ;
  buffer buf_n1232( .i (n1231), .o (n1232) );
  assign n1233 = n918 & n1232 ;
  buffer buf_n1234( .i (n1233), .o (n1234) );
  assign n1235 = n1214 & n1234 ;
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  assign n1241 = n1222 | n1228 ;
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n1247( .i (n1246), .o (n1247) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  assign n1249 = n1214 | n1234 ;
  buffer buf_n1250( .i (n1249), .o (n1250) );
  assign n1251 = ~n1236 & n1250 ;
  buffer buf_n1252( .i (n1251), .o (n1252) );
  assign n1253 = n1248 & n1252 ;
  buffer buf_n1254( .i (n1253), .o (n1254) );
  assign n1255 = n1240 | n1254 ;
  buffer buf_n1256( .i (n1255), .o (n1256) );
  assign n1257 = n1203 & n1256 ;
  buffer buf_n1258( .i (n1257), .o (n1258) );
  assign n1259 = n1185 | n1258 ;
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  assign n1303 = n1203 | n1256 ;
  buffer buf_n1304( .i (n1303), .o (n1304) );
  assign n1305 = ~n1258 & n1304 ;
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  assign n1347 = n1248 | n1252 ;
  buffer buf_n1348( .i (n1347), .o (n1348) );
  assign n1349 = ~n1254 & n1348 ;
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  assign n1357 = n918 | n1232 ;
  buffer buf_n1358( .i (n1357), .o (n1358) );
  assign n1359 = ~n1234 & n1358 ;
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  assign n1365 = n978 & n1364 ;
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  assign n1371 = n966 | n972 ;
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  assign n1379 = n978 | n1364 ;
  buffer buf_n1380( .i (n1379), .o (n1380) );
  assign n1381 = ~n1366 & n1380 ;
  buffer buf_n1382( .i (n1381), .o (n1382) );
  assign n1383 = n1378 & n1382 ;
  buffer buf_n1384( .i (n1383), .o (n1384) );
  assign n1385 = n1370 | n1384 ;
  buffer buf_n1386( .i (n1385), .o (n1386) );
  assign n1387 = n1356 & n1386 ;
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  assign n1423 = n1356 | n1386 ;
  buffer buf_n1424( .i (n1423), .o (n1424) );
  assign n1425 = ~n1388 & n1424 ;
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  buffer buf_n1455( .i (n1454), .o (n1455) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  assign n1457 = n1378 | n1382 ;
  buffer buf_n1458( .i (n1457), .o (n1458) );
  assign n1459 = ~n1384 & n1458 ;
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  assign n1463 = n1016 | n1022 ;
  buffer buf_n1464( .i (n1463), .o (n1464) );
  assign n1465 = n1462 & n1464 ;
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n1488( .i (n1487), .o (n1488) );
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  assign n1495 = n1462 | n1464 ;
  buffer buf_n1496( .i (n1495), .o (n1496) );
  assign n1497 = ~n1466 & n1496 ;
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n1522( .i (n1521), .o (n1522) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  assign n1523 = n1092 | n1160 ;
  buffer buf_n1524( .i (n1523), .o (n1524) );
  assign n1525 = n1522 & n1524 ;
  buffer buf_n1526( .i (n1525), .o (n1526) );
  assign n1527 = n1494 | n1526 ;
  buffer buf_n1528( .i (n1527), .o (n1528) );
  assign n1529 = n1456 & n1528 ;
  buffer buf_n1530( .i (n1529), .o (n1530) );
  assign n1531 = n1422 | n1530 ;
  buffer buf_n1532( .i (n1531), .o (n1532) );
  assign n1533 = n1346 & n1532 ;
  buffer buf_n1534( .i (n1533), .o (n1534) );
  assign n1535 = n1302 | n1534 ;
  assign n1536 = n671 | n691 ;
  buffer buf_n1537( .i (n1536), .o (n1537) );
  assign n1538 = ~n693 & n1537 ;
  assign n1539 = n1137 | n1152 ;
  buffer buf_n1540( .i (n1539), .o (n1540) );
  assign n1541 = ~n1154 & n1540 ;
  assign n1542 = n1346 | n1532 ;
  buffer buf_n1543( .i (n1542), .o (n1543) );
  assign n1544 = ~n1534 & n1543 ;
  assign n1545 = n590 | n708 ;
  buffer buf_n1546( .i (n1545), .o (n1546) );
  assign n1547 = ~n710 & n1546 ;
  assign n1548 = n1456 | n1528 ;
  buffer buf_n1549( .i (n1548), .o (n1549) );
  assign n1550 = ~n1530 & n1549 ;
  assign n1551 = n1522 | n1524 ;
  buffer buf_n1552( .i (n1551), .o (n1552) );
  assign n1553 = ~n1526 & n1552 ;
  assign n1554 = n663 | n704 ;
  buffer buf_n1555( .i (n1554), .o (n1555) );
  assign n1556 = ~n706 & n1555 ;
  assign n1557 = b_0_ & a_0_ ;
  assign s_1_ = n25 ;
  assign s_8_ = n717 ;
  assign s_3_ = n720 ;
  assign s_5_ = n723 ;
  assign s_9_ = n875 ;
  assign s_2_ = n878 ;
  assign s_11_ = n1161 ;
  assign s_15_ = n1535 ;
  assign s_4_ = n1538 ;
  assign s_10_ = n1541 ;
  assign s_14_ = n1544 ;
  assign s_7_ = n1547 ;
  assign s_13_ = n1550 ;
  assign s_12_ = n1553 ;
  assign s_6_ = n1556 ;
  assign s_0_ = n1557 ;
endmodule
