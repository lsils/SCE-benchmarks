module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( in_6_ , in_15_ , in_13_ , in_14_ , in_2_ , in_10_ , in_24_ , in_8_ , in_22_ , in_20_ , in_7_ , in_25_ , in_5_ , in_4_ , in_23_ , in_27_ , in_1_ , in_0_ , in_16_ , in_30_ , in_26_ , in_12_ , in_11_ , in_17_ , in_19_ , in_18_ , in_21_ , in_31_ , in_29_ , in_28_ , in_9_ , in_3_ , out_2_ , out_1_ , out_3_ , out_0_ , out_5_ , out_4_ );
  input in_6_ , in_15_ , in_13_ , in_14_ , in_2_ , in_10_ , in_24_ , in_8_ , in_22_ , in_20_ , in_7_ , in_25_ , in_5_ , in_4_ , in_23_ , in_27_ , in_1_ , in_0_ , in_16_ , in_30_ , in_26_ , in_12_ , in_11_ , in_17_ , in_19_ , in_18_ , in_21_ , in_31_ , in_29_ , in_28_ , in_9_ , in_3_ ;
  output out_2_ , out_1_ , out_3_ , out_0_ , out_5_ , out_4_ ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 ;
  assign n33 = in_29_ | in_28_ ;
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  assign n42 = in_20_ | in_21_ ;
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  assign n46 = in_16_ | in_17_ ;
  buffer buf_n47( .i (n46), .o (n47) );
  assign n48 = in_19_ & in_18_ ;
  buffer buf_n49( .i (n48), .o (n49) );
  assign n50 = ( n43 & n47 ) | ( n43 & n49 ) | ( n47 & n49 ) ;
  buffer buf_n51( .i (n50), .o (n51) );
  assign n57 = ( ~n43 & n47 ) | ( ~n43 & n49 ) | ( n47 & n49 ) ;
  buffer buf_n58( .i (n57), .o (n58) );
  assign n59 = ( n45 & ~n51 ) | ( n45 & n58 ) | ( ~n51 & n58 ) ;
  buffer buf_n60( .i (n59), .o (n60) );
  assign n61 = in_27_ & in_26_ ;
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  assign n65 = in_22_ & in_23_ ;
  buffer buf_n66( .i (n65), .o (n66) );
  assign n67 = in_24_ | in_25_ ;
  buffer buf_n68( .i (n67), .o (n68) );
  assign n69 = ( n62 & n66 ) | ( n62 & n68 ) | ( n66 & n68 ) ;
  buffer buf_n70( .i (n69), .o (n70) );
  assign n76 = ( ~n62 & n66 ) | ( ~n62 & n68 ) | ( n66 & n68 ) ;
  buffer buf_n77( .i (n76), .o (n77) );
  assign n78 = ( n64 & ~n70 ) | ( n64 & n77 ) | ( ~n70 & n77 ) ;
  buffer buf_n79( .i (n78), .o (n79) );
  assign n80 = ( n38 & n60 ) | ( n38 & n79 ) | ( n60 & n79 ) ;
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  assign n85 = ( n56 & n75 ) | ( n56 & n82 ) | ( n75 & n82 ) ;
  buffer buf_n86( .i (n85), .o (n86) );
  assign n91 = ( n56 & n75 ) | ( n56 & ~n82 ) | ( n75 & ~n82 ) ;
  buffer buf_n92( .i (n91), .o (n92) );
  assign n93 = ( n84 & ~n86 ) | ( n84 & n92 ) | ( ~n86 & n92 ) ;
  buffer buf_n94( .i (n93), .o (n94) );
  assign n95 = in_30_ & in_31_ ;
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  assign n106 = ( ~n38 & n60 ) | ( ~n38 & n79 ) | ( n60 & n79 ) ;
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n81), .o (n109) );
  assign n110 = ( n41 & n108 ) | ( n41 & ~n109 ) | ( n108 & ~n109 ) ;
  buffer buf_n111( .i (n110), .o (n111) );
  assign n112 = n105 & n111 ;
  buffer buf_n113( .i (n112), .o (n113) );
  assign n114 = n94 & n113 ;
  buffer buf_n115( .i (n114), .o (n115) );
  assign n116 = n94 | n113 ;
  buffer buf_n117( .i (n116), .o (n117) );
  assign n118 = ~n115 & n117 ;
  buffer buf_n119( .i (n118), .o (n119) );
  assign n121 = in_13_ | in_12_ ;
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  assign n130 = in_5_ | in_4_ ;
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  assign n134 = in_1_ | in_0_ ;
  buffer buf_n135( .i (n134), .o (n135) );
  assign n136 = in_2_ & in_3_ ;
  buffer buf_n137( .i (n136), .o (n137) );
  assign n138 = ( n131 & n135 ) | ( n131 & n137 ) | ( n135 & n137 ) ;
  buffer buf_n139( .i (n138), .o (n139) );
  assign n145 = ( ~n131 & n135 ) | ( ~n131 & n137 ) | ( n135 & n137 ) ;
  buffer buf_n146( .i (n145), .o (n146) );
  assign n147 = ( n133 & ~n139 ) | ( n133 & n146 ) | ( ~n139 & n146 ) ;
  buffer buf_n148( .i (n147), .o (n148) );
  assign n149 = in_10_ & in_11_ ;
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  assign n153 = in_6_ & in_7_ ;
  buffer buf_n154( .i (n153), .o (n154) );
  assign n155 = in_8_ | in_9_ ;
  buffer buf_n156( .i (n155), .o (n156) );
  assign n157 = ( n150 & n154 ) | ( n150 & n156 ) | ( n154 & n156 ) ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n164 = ( ~n150 & n154 ) | ( ~n150 & n156 ) | ( n154 & n156 ) ;
  buffer buf_n165( .i (n164), .o (n165) );
  assign n166 = ( n152 & ~n158 ) | ( n152 & n165 ) | ( ~n158 & n165 ) ;
  buffer buf_n167( .i (n166), .o (n167) );
  assign n168 = ( n126 & n148 ) | ( n126 & n167 ) | ( n148 & n167 ) ;
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  assign n173 = ( n144 & n163 ) | ( n144 & n170 ) | ( n163 & n170 ) ;
  buffer buf_n174( .i (n173), .o (n174) );
  assign n179 = ( n144 & n163 ) | ( n144 & ~n170 ) | ( n163 & ~n170 ) ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = ( n172 & ~n174 ) | ( n172 & n180 ) | ( ~n174 & n180 ) ;
  buffer buf_n182( .i (n181), .o (n182) );
  assign n183 = in_15_ & in_14_ ;
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  assign n194 = ( ~n126 & n148 ) | ( ~n126 & n167 ) | ( n148 & n167 ) ;
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n169), .o (n197) );
  assign n198 = ( n129 & n196 ) | ( n129 & ~n197 ) | ( n196 & ~n197 ) ;
  buffer buf_n199( .i (n198), .o (n199) );
  assign n200 = n193 & n199 ;
  buffer buf_n201( .i (n200), .o (n201) );
  assign n202 = n182 & n201 ;
  buffer buf_n203( .i (n202), .o (n203) );
  assign n204 = n182 | n201 ;
  buffer buf_n205( .i (n204), .o (n205) );
  assign n206 = ~n203 & n205 ;
  buffer buf_n207( .i (n206), .o (n207) );
  assign n209 = n119 & n207 ;
  assign n210 = n119 | n207 ;
  assign n211 = ~n209 & n210 ;
  buffer buf_n212( .i (n211), .o (n212) );
  assign n213 = n105 | n111 ;
  buffer buf_n214( .i (n213), .o (n214) );
  assign n215 = ~n113 & n214 ;
  buffer buf_n216( .i (n215), .o (n216) );
  assign n217 = n193 | n199 ;
  buffer buf_n218( .i (n217), .o (n218) );
  assign n219 = ~n201 & n218 ;
  buffer buf_n220( .i (n219), .o (n220) );
  assign n221 = n216 & n220 ;
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  assign n226 = n212 & n225 ;
  assign n227 = n212 | n225 ;
  assign n228 = ~n226 & n227 ;
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  assign n232 = n216 | n220 ;
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  assign n235 = ~n223 & n234 ;
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  assign n242 = n90 & n115 ;
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  assign n249 = n90 | n115 ;
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  assign n252 = ~n244 & n251 ;
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  assign n254 = n178 & n203 ;
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  assign n261 = n178 | n203 ;
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  assign n264 = ~n256 & n263 ;
  buffer buf_n265( .i (n264), .o (n265) );
  assign n266 = n253 & n265 ;
  assign n267 = n253 | n265 ;
  assign n268 = ~n266 & n267 ;
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n208( .i (n207), .o (n208) );
  assign n270 = ( n120 & n208 ) | ( n120 & n223 ) | ( n208 & n223 ) ;
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  assign n275 = n269 & n274 ;
  assign n276 = n269 | n274 ;
  assign n277 = ~n275 & n276 ;
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  assign n278 = ( n253 & n265 ) | ( n253 & n271 ) | ( n265 & n271 ) ;
  buffer buf_n279( .i (n278), .o (n279) );
  assign n280 = ( n248 & n260 ) | ( n248 & n279 ) | ( n260 & n279 ) ;
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  assign n283 = n245 | n257 ;
  assign n284 = n245 & n257 ;
  assign n285 = n283 & ~n284 ;
  buffer buf_n286( .i (n285), .o (n286) );
  assign n287 = n279 & n286 ;
  assign n288 = n279 | n286 ;
  assign n289 = ~n287 & n288 ;
  buffer buf_n290( .i (n289), .o (n290) );
  assign out_2_ = n231 ;
  assign out_1_ = n241 ;
  assign out_3_ = n277 ;
  assign out_0_ = 1'b0 ;
  assign out_5_ = n282 ;
  assign out_4_ = n290 ;
endmodule
