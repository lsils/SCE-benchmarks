module top( G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 );
  input G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 ;
  output G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 ;
  wire n1250 , n1251 , n1252 , n1280 , n1281 , n1309 , n1337 , n1366 , n1393 , n1420 , n1421 , n1422 , n1424 , n1425 , n1426 , n1428 , n1454 , n1455 , n1456 , n1481 , n1485 , n1486 , n1487 , n1488 , n1490 , n1491 , n1492 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1547 , n1548 , n1549 , n1550 , n1552 , n1553 , n1554 , n1579 , n1581 , n1582 , n1583 , n1585 , n1589 , n1590 , n1591 , n1592 , n1615 , n1618 , n1619 , n1620 , n1623 , n1624 , n1625 , n1626 , n1648 , n1650 , n1651 , n1652 , n1655 , n1657 , n1658 , n1659 , n1681 , n1684 , n1685 , n1686 , n1690 , n1691 , n1692 , n1693 , n1700 , n1719 , n1725 , n1727 , n1748 , n1757 , n1778 , n1780 , n1782 , n1783 , n1787 , n1788 , n1789 , n1790 , n1811 , n1812 , n1815 , n1816 , n1817 , n1819 , n1842 , n1844 , n1845 , n1846 , n1851 , n1852 , n1853 , n1854 , n1875 , n1879 , n1880 , n1881 , n1885 , n1886 , n1887 , n1888 , n1909 , n1911 , n1913 , n1914 , n1919 , n1920 , n1921 , n1922 , n1930 , n1931 , n1932 , n1949 , n1950 , n1951 , n1968 , n1969 , n1987 , n1989 , n1990 , n1991 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2018 , n2019 , n2020 , n2021 , n2040 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2056 , n2057 , n2058 , n2064 , n2073 , n2074 , n2075 , n2077 , n2086 , n2087 , n2088 , n2090 , n2091 , n2093 , n2102 , n2103 , n2104 , n2106 , n2112 , n2113 , n2114 , n2120 , n2121 , n2128 , n2129 , n2130 , n2135 , n2139 , n2141 , n2150 , n2151 , n2152 , n2154 , n2164 , n2165 , n2166 , n2168 , n2170 , n2178 , n2179 , n2180 , n2184 , n2187 , n2188 , n2189 , n2191 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2207 , n2208 , n2210 , n2211 , n2212 , n2215 , n2222 , n2223 , n2225 , n2226 , n2227 , n2228 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2246 , n2247 , n2249 , n2250 , n2251 , n2253 , n2254 , n2258 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2280 , n2281 , n2290 , n2291 , n2292 , n2294 , n2295 , n2297 , n2306 , n2307 , n2308 , n2310 , n2311 , n2312 , n2320 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2340 , n2341 , n2342 , n2347 , n2348 , n2349 , n2350 , n2351 , n2361 , n2364 , n2365 , n2366 , n2370 , n2371 , n2372 , n2373 , n2375 , n2376 , n2394 , n2395 , n2396 , n2398 , n2399 , n2400 , n2401 , n2418 , n2421 , n2439 , n2443 , n2445 , n2448 , n2450 , n2461 , n2463 , n2473 , n2482 , n2483 , n2484 , n2485 , n2491 , n2492 , n2493 , n2495 , n2498 , n2499 , n2500 , n2502 , n2504 , n2505 , n2506 , n2507 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2522 , n2524 , n2525 , n2534 , n2535 , n2536 , n2537 , n2539 , n2542 , n2543 , n2547 , n2551 , n2552 , n2553 , n2554 , n2555 , n2558 , n2564 , n2566 , n2572 , n2577 , n2579 , n2587 , n2588 , n2590 , n2592 , n2593 , n2595 , n2599 , n2602 , n2606 , n2608 , n2609 , n2610 , n2620 , n2621 , n2622 , n2623 , n2624 , n2634 , n2635 , n2643 ;
  buffer buf_n265( .i (G115), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n354( .i (G124), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n551( .i (G137), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n753( .i (G32), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n207( .i (G106), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n1006( .i (G64), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1070( .i (G76), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n912( .i (G53), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n1209( .i (G96), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n820( .i (G43), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n1147( .i (G86), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n626( .i (G141), .o (n626) );
  buffer buf_n642( .i (G142), .o (n642) );
  assign n1250 = n626 | n642 ;
  buffer buf_n595( .i (G139), .o (n595) );
  buffer buf_n612( .i (G140), .o (n612) );
  assign n1251 = n595 | n612 ;
  assign n1252 = n1250 | n1251 ;
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n248( .i (G11), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n329( .i (G121), .o (n329) );
  buffer buf_n696( .i (G2), .o (n696) );
  assign n1280 = n329 | n696 ;
  assign n1281 = n249 | n1280 ;
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1064( .i (G74), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  assign n1309 = n266 & ~n1065 ;
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1051( .i (G7), .o (n1051) );
  assign n1337 = n329 | n1051 ;
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n310( .i (G119), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  assign n1366 = n312 | n1338 ;
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n678( .i (G147), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  assign n1393 = n680 | n1338 ;
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  assign n1420 = n912 & ~n1209 ;
  assign n1421 = n820 | n1147 ;
  assign n1422 = n1420 & ~n1421 ;
  buffer buf_n1423( .i (n1422), .o (n1423) );
  assign n1424 = ~n207 & n753 ;
  assign n1425 = n1006 | n1070 ;
  assign n1426 = n1424 & ~n1425 ;
  buffer buf_n1427( .i (n1426), .o (n1427) );
  assign n1428 = n1423 | n1427 ;
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n681( .i (n680), .o (n681) );
  assign n1454 = n681 & ~n1427 ;
  buffer buf_n313( .i (n312), .o (n313) );
  assign n1455 = n313 & ~n1423 ;
  assign n1456 = n1454 | n1455 ;
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n245( .i (G109), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  assign n1481 = G145 | G146 ;
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  assign n1485 = n247 & ~n1483 ;
  buffer buf_n1108( .i (G79), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  assign n1486 = n1110 & ~n1483 ;
  assign n1487 = n1485 | n1486 ;
  buffer buf_n1185( .i (G89), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  assign n1488 = n1187 & ~n1483 ;
  buffer buf_n1247( .i (G99), .o (n1247) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1489( .i (n1482), .o (n1489) );
  assign n1490 = n1249 & ~n1489 ;
  assign n1491 = n1488 | n1490 ;
  assign n1492 = n1487 | n1491 ;
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n241( .i (G108), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  assign n1517 = n244 | n1484 ;
  buffer buf_n1243( .i (G98), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  assign n1518 = n1246 & ~n1484 ;
  assign n1519 = n1517 & ~n1518 ;
  buffer buf_n1181( .i (G88), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  assign n1520 = n1184 & ~n1484 ;
  buffer buf_n1104( .i (G78), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  assign n1521 = n1107 & ~n1484 ;
  assign n1522 = n1520 | n1521 ;
  assign n1523 = n1519 & ~n1522 ;
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  buffer buf_n1534( .i (n1533), .o (n1534) );
  buffer buf_n1535( .i (n1534), .o (n1535) );
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1128( .i (G80), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n1547 = n1130 | n1489 ;
  buffer buf_n1190( .i (G90), .o (n1190) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  assign n1548 = n1192 & ~n1489 ;
  assign n1549 = n1547 & ~n1548 ;
  buffer buf_n188( .i (G100), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  assign n1550 = n190 & ~n1489 ;
  buffer buf_n250( .i (G110), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n1551( .i (n1482), .o (n1551) );
  assign n1552 = n252 & ~n1551 ;
  assign n1553 = n1550 | n1552 ;
  assign n1554 = n1549 & ~n1553 ;
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n1556( .i (n1555), .o (n1556) );
  buffer buf_n1557( .i (n1556), .o (n1557) );
  buffer buf_n1558( .i (n1557), .o (n1558) );
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n296( .i (G117), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n792( .i (G36), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  assign n1579 = n298 & ~n794 ;
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n325( .i (G120), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n1045( .i (G68), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  assign n1581 = n298 & ~n1047 ;
  assign n1582 = n328 | n1581 ;
  assign n1583 = n1580 & ~n1582 ;
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n864( .i (G46), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  assign n1585 = n298 | n327 ;
  buffer buf_n1586( .i (n1585), .o (n1586) );
  assign n1589 = n868 & ~n1586 ;
  buffer buf_n962( .i (G57), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  assign n1590 = n966 & ~n1586 ;
  assign n1591 = n1589 | n1590 ;
  assign n1592 = n1584 & ~n1591 ;
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n795( .i (G37), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  assign n1615 = n298 & ~n797 ;
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1048( .i (G69), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1617( .i (n297), .o (n1617) );
  assign n1618 = ~n1050 & n1617 ;
  assign n1619 = n328 | n1618 ;
  assign n1620 = n1616 & ~n1619 ;
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n869( .i (G47), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  assign n1623 = n874 & ~n1587 ;
  buffer buf_n967( .i (G58), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  assign n1624 = n972 & ~n1587 ;
  assign n1625 = n1623 | n1624 ;
  assign n1626 = n1622 & ~n1625 ;
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n1633( .i (n1632), .o (n1633) );
  buffer buf_n1634( .i (n1633), .o (n1634) );
  buffer buf_n1635( .i (n1634), .o (n1635) );
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n1637( .i (n1636), .o (n1637) );
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n798( .i (G38), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  assign n1648 = ~n800 & n1617 ;
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1052( .i (G70), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  assign n1650 = ~n1054 & n1617 ;
  assign n1651 = n328 | n1650 ;
  assign n1652 = n1649 & ~n1651 ;
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n875( .i (G48), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  assign n1655 = n880 & ~n1587 ;
  buffer buf_n973( .i (G59), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n1656( .i (n1586), .o (n1656) );
  assign n1657 = n978 & ~n1656 ;
  assign n1658 = n1655 | n1657 ;
  assign n1659 = n1654 & ~n1658 ;
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n330( .i (G122), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n750( .i (G31), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  assign n1681 = ~n752 & n1617 ;
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1003( .i (G63), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1683( .i (n297), .o (n1683) );
  assign n1684 = ~n1005 & n1683 ;
  assign n1685 = n328 | n1684 ;
  assign n1686 = n1682 & ~n1685 ;
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n813( .i (G42), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  assign n1690 = n819 & ~n1588 ;
  buffer buf_n905( .i (G52), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  assign n1691 = n911 & ~n1588 ;
  assign n1692 = n1690 | n1691 ;
  assign n1693 = n1689 & ~n1692 ;
  buffer buf_n1694( .i (n1693), .o (n1694) );
  assign n1700 = n340 | n1694 ;
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n719( .i (G28), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n295( .i (G116), .o (n295) );
  assign n1719 = n295 | n329 ;
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  assign n1725 = n1457 | n1724 ;
  buffer buf_n1726( .i (n1725), .o (n1726) );
  assign n1727 = n727 | n1726 ;
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  assign n1748 = G1 & ~G3 ;
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  assign n1757 = n1726 | n1756 ;
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n801( .i (G39), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  assign n1778 = n803 | n1683 ;
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1055( .i (G71), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  assign n1780 = ~n1057 & n1683 ;
  buffer buf_n1781( .i (n327), .o (n1781) );
  assign n1782 = n1780 | n1781 ;
  assign n1783 = n1779 & ~n1782 ;
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n881( .i (G49), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  assign n1787 = n887 & ~n1588 ;
  buffer buf_n982( .i (G60), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  assign n1788 = n988 & ~n1588 ;
  assign n1789 = n1787 | n1788 ;
  assign n1790 = n1786 | n1789 ;
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n956( .i (G56), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  assign n1811 = n961 & ~n1656 ;
  buffer buf_n789( .i (G35), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  assign n1812 = n791 | n1683 ;
  buffer buf_n1813( .i (n1812), .o (n1813) );
  buffer buf_n1042( .i (G67), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1814( .i (n297), .o (n1814) );
  assign n1815 = ~n1044 & n1814 ;
  assign n1816 = n1781 | n1815 ;
  assign n1817 = n1813 & ~n1816 ;
  buffer buf_n1818( .i (n1817), .o (n1818) );
  assign n1819 = n1811 & ~n1818 ;
  buffer buf_n1820( .i (n1819), .o (n1820) );
  buffer buf_n1821( .i (n1820), .o (n1821) );
  buffer buf_n1822( .i (n1821), .o (n1822) );
  buffer buf_n1823( .i (n1822), .o (n1823) );
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1825( .i (n1824), .o (n1825) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n786( .i (G34), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  assign n1842 = ~n788 & n1814 ;
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1039( .i (G66), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  assign n1844 = ~n1041 & n1814 ;
  assign n1845 = n1781 | n1844 ;
  assign n1846 = n1843 & ~n1845 ;
  buffer buf_n1847( .i (n1846), .o (n1847) );
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n857( .i (G45), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n1850( .i (n1656), .o (n1850) );
  assign n1851 = n863 & ~n1850 ;
  buffer buf_n949( .i (G55), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  assign n1852 = n955 & ~n1850 ;
  assign n1853 = n1851 | n1852 ;
  assign n1854 = n1849 & ~n1853 ;
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  buffer buf_n1872( .i (n1871), .o (n1872) );
  buffer buf_n1873( .i (n1872), .o (n1873) );
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n783( .i (G33), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  assign n1875 = ~n785 & n1814 ;
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1036( .i (G65), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1877( .i (n296), .o (n1877) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  assign n1879 = ~n1038 & n1878 ;
  assign n1880 = n1781 | n1879 ;
  assign n1881 = n1876 & ~n1880 ;
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n850( .i (G44), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  assign n1885 = n856 & ~n1850 ;
  buffer buf_n942( .i (G54), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  assign n1886 = n948 & ~n1850 ;
  assign n1887 = n1885 | n1886 ;
  assign n1888 = n1884 & ~n1887 ;
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1907( .i (n1906), .o (n1907) );
  buffer buf_n1908( .i (n1907), .o (n1908) );
  buffer buf_n342( .i (G123), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n807( .i (G40), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  assign n1909 = ~n809 & n1878 ;
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1058( .i (G72), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1911 = ~n1060 & n1878 ;
  buffer buf_n1912( .i (n327), .o (n1912) );
  assign n1913 = n1911 | n1912 ;
  assign n1914 = n1910 & ~n1913 ;
  buffer buf_n1915( .i (n1914), .o (n1915) );
  buffer buf_n1916( .i (n1915), .o (n1916) );
  buffer buf_n1917( .i (n1916), .o (n1917) );
  buffer buf_n891( .i (G50), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n1918( .i (n1656), .o (n1918) );
  assign n1919 = n897 & ~n1918 ;
  buffer buf_n989( .i (G61), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  assign n1920 = n995 & ~n1918 ;
  assign n1921 = n1919 | n1920 ;
  assign n1922 = n1917 & ~n1921 ;
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  assign n1930 = n353 | n1924 ;
  assign n1931 = n353 & ~n1662 ;
  assign n1932 = n1930 & ~n1931 ;
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n1934( .i (n1933), .o (n1934) );
  buffer buf_n1935( .i (n1934), .o (n1935) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  assign n1949 = n353 | n1792 ;
  assign n1950 = ~n353 & n1629 ;
  assign n1951 = n1949 & ~n1950 ;
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  buffer buf_n1954( .i (n1953), .o (n1954) );
  buffer buf_n1955( .i (n1954), .o (n1955) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  buffer buf_n1960( .i (n1959), .o (n1960) );
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n1967( .i (n1966), .o (n1967) );
  buffer buf_n299( .i (G118), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  assign n1968 = n309 & ~n340 ;
  assign n1969 = n1924 | n1968 ;
  buffer buf_n1970( .i (n1969), .o (n1970) );
  buffer buf_n1971( .i (n1970), .o (n1971) );
  buffer buf_n1972( .i (n1971), .o (n1972) );
  buffer buf_n1973( .i (n1972), .o (n1973) );
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  buffer buf_n1983( .i (n1982), .o (n1983) );
  buffer buf_n1984( .i (n1983), .o (n1984) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n1986( .i (n1985), .o (n1986) );
  assign n1987 = n352 & ~n1694 ;
  buffer buf_n1988( .i (n1987), .o (n1988) );
  assign n1989 = n309 | n352 ;
  assign n1990 = n1924 & ~n1989 ;
  assign n1991 = n1988 | n1990 ;
  buffer buf_n1992( .i (n1991), .o (n1992) );
  buffer buf_n1993( .i (n1992), .o (n1993) );
  buffer buf_n1994( .i (n1993), .o (n1994) );
  buffer buf_n1995( .i (n1994), .o (n1995) );
  buffer buf_n1996( .i (n1995), .o (n1996) );
  buffer buf_n1997( .i (n1996), .o (n1997) );
  buffer buf_n1998( .i (n1997), .o (n1998) );
  buffer buf_n1999( .i (n1998), .o (n1999) );
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n2001( .i (n2000), .o (n2001) );
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n2003), .o (n2004) );
  buffer buf_n2005( .i (n2004), .o (n2005) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n2007( .i (n2006), .o (n2007) );
  buffer buf_n667( .i (G144), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n658( .i (G143), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n1100( .i (G77), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n2008( .i (n1551), .o (n2008) );
  assign n2009 = n1103 & ~n2008 ;
  buffer buf_n1239( .i (G97), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  assign n2010 = n1242 & ~n2008 ;
  assign n2011 = n2009 & ~n2010 ;
  buffer buf_n237( .i (G107), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  assign n2012 = n240 & ~n2008 ;
  buffer buf_n1177( .i (G87), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  assign n2013 = n1180 & ~n2008 ;
  assign n2014 = n2012 | n2013 ;
  assign n2015 = n2011 & ~n2014 ;
  buffer buf_n2016( .i (n2015), .o (n2016) );
  buffer buf_n2017( .i (n2016), .o (n2017) );
  assign n2018 = n666 | n2017 ;
  assign n2019 = n666 & ~n2017 ;
  assign n2020 = n2018 & ~n2019 ;
  assign n2021 = n677 | n2020 ;
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2028( .i (n2027), .o (n2028) );
  buffer buf_n2029( .i (n2028), .o (n2029) );
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n2031( .i (n2030), .o (n2031) );
  buffer buf_n2032( .i (n2031), .o (n2032) );
  buffer buf_n2033( .i (n2032), .o (n2033) );
  buffer buf_n2034( .i (n2033), .o (n2034) );
  buffer buf_n2035( .i (n2034), .o (n2035) );
  buffer buf_n2036( .i (n2035), .o (n2036) );
  buffer buf_n2037( .i (n2036), .o (n2037) );
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n158( .i (G10), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n527( .i (G135), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n694( .i (G19), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n702( .i (G23), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  assign n2040 = ~n695 & n703 ;
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n1066( .i (G75), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n2047( .i (n1551), .o (n2047) );
  assign n2048 = n1069 & ~n2047 ;
  buffer buf_n1143( .i (G85), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  assign n2049 = n1146 & ~n2047 ;
  assign n2050 = n2048 & ~n2049 ;
  buffer buf_n1205( .i (G95), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  assign n2051 = n1208 & ~n2047 ;
  buffer buf_n203( .i (G105), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  assign n2052 = n206 & ~n2047 ;
  assign n2053 = n2051 | n2052 ;
  assign n2054 = n2050 & ~n2053 ;
  buffer buf_n2055( .i (n2054), .o (n2055) );
  assign n2056 = n709 & ~n2055 ;
  assign n2057 = n2046 & ~n2056 ;
  assign n2058 = n536 & ~n2057 ;
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  buffer buf_n384( .i (G125), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n314( .i (G12), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n447( .i (G13), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  assign n2064 = n316 & ~n449 ;
  buffer buf_n2065( .i (n2064), .o (n2065) );
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  assign n2073 = n324 & ~n1694 ;
  assign n2074 = n2072 & ~n2073 ;
  assign n2075 = n396 & ~n2074 ;
  buffer buf_n2076( .i (n2075), .o (n2076) );
  buffer buf_n450( .i (G130), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n682( .i (G15), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  assign n2077 = n316 & ~n684 ;
  buffer buf_n2078( .i (n2077), .o (n2078) );
  buffer buf_n2079( .i (n2078), .o (n2079) );
  buffer buf_n2080( .i (n2079), .o (n2080) );
  buffer buf_n2081( .i (n2080), .o (n2081) );
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  assign n2086 = ~n324 & n1628 ;
  assign n2087 = n2085 & ~n2086 ;
  assign n2088 = n462 & ~n2087 ;
  buffer buf_n2089( .i (n2088), .o (n2089) );
  assign n2090 = n2076 | n2089 ;
  assign n2091 = n2063 | n2090 ;
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n433( .i (G129), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n888( .i (G5), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  assign n2093 = n316 & ~n890 ;
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n2099( .i (n2098), .o (n2099) );
  buffer buf_n2100( .i (n2099), .o (n2100) );
  buffer buf_n2101( .i (n2100), .o (n2101) );
  assign n2102 = n324 & ~n1661 ;
  assign n2103 = n2101 & ~n2102 ;
  assign n2104 = n445 & ~n2103 ;
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n699( .i (G21), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  assign n2106 = ~n700 & n703 ;
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n2111( .i (n2110), .o (n2111) );
  assign n2112 = n708 & ~n1555 ;
  assign n2113 = n2111 & ~n2112 ;
  assign n2114 = n620 & ~n2113 ;
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  buffer buf_n2119( .i (n2118), .o (n2119) );
  assign n2120 = n2105 | n2119 ;
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n717( .i (G27), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  assign n2121 = n703 & ~n718 ;
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  assign n2128 = n709 & ~n1524 ;
  assign n2129 = n2127 & ~n2128 ;
  assign n2130 = n651 & ~n2129 ;
  buffer buf_n2131( .i (n2130), .o (n2131) );
  assign n2135 = n2059 | n2131 ;
  buffer buf_n2136( .i (n2135), .o (n2136) );
  buffer buf_n2137( .i (n2136), .o (n2137) );
  buffer buf_n2138( .i (n2137), .o (n2138) );
  assign n2139 = n2120 | n2138 ;
  buffer buf_n419( .i (G128), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n609( .i (G14), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n2140( .i (n315), .o (n2140) );
  assign n2141 = ~n611 & n2140 ;
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n2143( .i (n2142), .o (n2143) );
  buffer buf_n2144( .i (n2143), .o (n2144) );
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  assign n2150 = ~n324 & n1791 ;
  assign n2151 = n2149 & ~n2150 ;
  assign n2152 = n431 & ~n2151 ;
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n398( .i (G126), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n804( .i (G4), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  assign n2154 = ~n806 & n2140 ;
  buffer buf_n2155( .i (n2154), .o (n2155) );
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n2158( .i (n2157), .o (n2158) );
  buffer buf_n2159( .i (n2158), .o (n2159) );
  buffer buf_n2160( .i (n2159), .o (n2160) );
  buffer buf_n2161( .i (n2160), .o (n2161) );
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n2163( .i (n323), .o (n2163) );
  assign n2164 = ~n1923 & n2163 ;
  assign n2165 = n2162 & ~n2164 ;
  assign n2166 = n410 & ~n2165 ;
  buffer buf_n2167( .i (n2166), .o (n2167) );
  assign n2168 = n2153 | n2167 ;
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n715( .i (G26), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n2169( .i (n702), .o (n2169) );
  assign n2170 = ~n716 & n2169 ;
  buffer buf_n2171( .i (n2170), .o (n2171) );
  buffer buf_n2172( .i (n2171), .o (n2172) );
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n2175( .i (n2174), .o (n2175) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n710( .i (n709), .o (n710) );
  assign n2178 = n710 & ~n1495 ;
  assign n2179 = n2177 & ~n2178 ;
  assign n2180 = n636 & ~n2179 ;
  buffer buf_n2181( .i (n2180), .o (n2181) );
  assign n2184 = n2117 | n2181 ;
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  assign n2187 = n2168 | n2186 ;
  assign n2188 = n2139 | n2187 ;
  assign n2189 = n2092 | n2188 ;
  buffer buf_n2190( .i (n2189), .o (n2190) );
  buffer buf_n537( .i (G136), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n711( .i (G24), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  assign n2191 = ~n712 & n2169 ;
  buffer buf_n2192( .i (n2191), .o (n2192) );
  buffer buf_n2193( .i (n2192), .o (n2193) );
  buffer buf_n2194( .i (n2193), .o (n2194) );
  buffer buf_n2195( .i (n2194), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  buffer buf_n2197( .i (n2196), .o (n2197) );
  buffer buf_n1201( .i (G93), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n2198( .i (n1551), .o (n2198) );
  assign n2199 = n1204 & ~n2198 ;
  buffer buf_n199( .i (G103), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  assign n2200 = n202 & ~n2198 ;
  assign n2201 = n2199 & ~n2200 ;
  buffer buf_n261( .i (G113), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  assign n2202 = n264 & ~n2198 ;
  buffer buf_n1139( .i (G83), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  assign n2203 = n1142 & ~n2198 ;
  assign n2204 = n2202 | n2203 ;
  assign n2205 = n2201 & ~n2204 ;
  buffer buf_n2206( .i (n2205), .o (n2206) );
  assign n2207 = n709 & ~n2206 ;
  assign n2208 = n2197 & ~n2207 ;
  buffer buf_n2209( .i (n2208), .o (n2209) );
  assign n2210 = n547 | n2209 ;
  assign n2211 = n547 & ~n2209 ;
  assign n2212 = n2210 & ~n2211 ;
  buffer buf_n2213( .i (n2212), .o (n2213) );
  buffer buf_n2214( .i (n2213), .o (n2214) );
  buffer buf_n466( .i (G131), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n685( .i (G16), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  assign n2215 = ~n687 & n2140 ;
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n2221( .i (n2220), .o (n2221) );
  assign n2222 = n322 & ~n1593 ;
  assign n2223 = n2221 & ~n2222 ;
  buffer buf_n2224( .i (n2223), .o (n2224) );
  assign n2225 = n477 | n2224 ;
  assign n2226 = n477 & ~n2224 ;
  assign n2227 = n2225 & ~n2226 ;
  buffer buf_n581( .i (G138), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n697( .i (G20), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  assign n2228 = ~n698 & n2169 ;
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  buffer buf_n2231( .i (n2230), .o (n2231) );
  buffer buf_n2232( .i (n2231), .o (n2232) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  buffer buf_n1135( .i (G82), .o (n1135) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n2235( .i (n1482), .o (n2235) );
  buffer buf_n2236( .i (n2235), .o (n2236) );
  assign n2237 = n1138 & ~n2236 ;
  buffer buf_n195( .i (G102), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  assign n2238 = n198 & ~n2236 ;
  assign n2239 = n2237 & ~n2238 ;
  buffer buf_n257( .i (G112), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  assign n2240 = n260 & ~n2236 ;
  buffer buf_n1197( .i (G92), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  assign n2241 = n1200 & ~n2236 ;
  assign n2242 = n2240 | n2241 ;
  assign n2243 = n2239 & ~n2242 ;
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n708), .o (n2245) );
  assign n2246 = ~n2244 & n2245 ;
  assign n2247 = n2234 & ~n2246 ;
  buffer buf_n2248( .i (n2247), .o (n2248) );
  assign n2249 = n591 | n2248 ;
  assign n2250 = n591 & ~n2248 ;
  assign n2251 = n2249 & ~n2250 ;
  buffer buf_n2252( .i (n2251), .o (n2252) );
  assign n2253 = n2227 | n2252 ;
  assign n2254 = n2214 | n2253 ;
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n713( .i (G25), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  assign n2258 = ~n714 & n2169 ;
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n1131( .i (G81), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n2264( .i (n2235), .o (n2264) );
  assign n2265 = n1134 & ~n2264 ;
  buffer buf_n191( .i (G101), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  assign n2266 = n194 & ~n2264 ;
  assign n2267 = n2265 & ~n2266 ;
  buffer buf_n253( .i (G111), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  assign n2268 = n256 & ~n2264 ;
  buffer buf_n1193( .i (G91), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  assign n2269 = n1196 & ~n2264 ;
  assign n2270 = n2268 | n2269 ;
  assign n2271 = n2267 & ~n2270 ;
  assign n2272 = n708 & ~n2271 ;
  assign n2273 = n2263 & ~n2272 ;
  assign n2274 = n603 & ~n2273 ;
  buffer buf_n2275( .i (n2274), .o (n2275) );
  buffer buf_n2276( .i (n2275), .o (n2276) );
  buffer buf_n2277( .i (n2276), .o (n2277) );
  buffer buf_n2278( .i (n2277), .o (n2278) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  assign n2280 = n2089 | n2279 ;
  buffer buf_n514( .i (G134), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n691( .i (G18), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  assign n2281 = ~n693 & n2140 ;
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n2289( .i (n2288), .o (n2289) );
  assign n2290 = ~n1889 & n2163 ;
  assign n2291 = n2289 & ~n2290 ;
  assign n2292 = n526 & ~n2291 ;
  buffer buf_n2293( .i (n2292), .o (n2293) );
  assign n2294 = n2167 | n2293 ;
  assign n2295 = n2280 | n2294 ;
  buffer buf_n498( .i (G133), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n979( .i (G6), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n2296( .i (n315), .o (n2296) );
  assign n2297 = ~n981 & n2296 ;
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  assign n2306 = ~n1855 & n2163 ;
  assign n2307 = n2305 & ~n2306 ;
  assign n2308 = n510 & ~n2307 ;
  buffer buf_n2309( .i (n2308), .o (n2309) );
  assign n2310 = n710 & ~n2017 ;
  buffer buf_n1188( .i (G9), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n701( .i (G22), .o (n701) );
  assign n2311 = ~n701 & n702 ;
  assign n2312 = n1189 | n2311 ;
  buffer buf_n2313( .i (n2312), .o (n2313) );
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  assign n2320 = n2310 | n2319 ;
  buffer buf_n2321( .i (n2320), .o (n2321) );
  buffer buf_n2322( .i (n2321), .o (n2322) );
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  assign n2325 = n2309 | n2324 ;
  buffer buf_n2132( .i (n2131), .o (n2132) );
  buffer buf_n2133( .i (n2132), .o (n2133) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  assign n2326 = n2134 | n2309 ;
  assign n2327 = n2325 | n2326 ;
  assign n2328 = n2295 | n2327 ;
  buffer buf_n2182( .i (n2181), .o (n2182) );
  buffer buf_n2183( .i (n2182), .o (n2183) );
  assign n2329 = n2105 | n2183 ;
  assign n2330 = n2076 | n2153 ;
  assign n2331 = n2329 | n2330 ;
  assign n2332 = n2279 | n2293 ;
  buffer buf_n482( .i (G132), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n688( .i (G17), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  assign n2333 = ~n690 & n2296 ;
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n2335( .i (n2334), .o (n2335) );
  buffer buf_n2336( .i (n2335), .o (n2336) );
  buffer buf_n2337( .i (n2336), .o (n2337) );
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  assign n2340 = n322 & ~n1820 ;
  assign n2341 = n2339 & ~n2340 ;
  assign n2342 = n492 & ~n2341 ;
  buffer buf_n2343( .i (n2342), .o (n2343) );
  buffer buf_n2344( .i (n2343), .o (n2344) );
  buffer buf_n2345( .i (n2344), .o (n2345) );
  buffer buf_n2346( .i (n2345), .o (n2346) );
  assign n2347 = n2332 | n2346 ;
  assign n2348 = n2331 | n2347 ;
  assign n2349 = n2328 | n2348 ;
  assign n2350 = n2257 | n2349 ;
  assign n2351 = n2190 | n2350 ;
  buffer buf_n2352( .i (n2351), .o (n2352) );
  buffer buf_n2353( .i (n2352), .o (n2353) );
  buffer buf_n2354( .i (n2353), .o (n2354) );
  buffer buf_n2355( .i (n2354), .o (n2355) );
  buffer buf_n2356( .i (n2355), .o (n2356) );
  buffer buf_n2357( .i (n2356), .o (n2357) );
  buffer buf_n2358( .i (n2357), .o (n2358) );
  buffer buf_n2359( .i (n2358), .o (n2359) );
  buffer buf_n2360( .i (n2359), .o (n2360) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n810( .i (G41), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  assign n2361 = ~n812 & n1878 ;
  buffer buf_n2362( .i (n2361), .o (n2362) );
  buffer buf_n1061( .i (G73), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n2363( .i (n1877), .o (n2363) );
  assign n2364 = ~n1063 & n2363 ;
  assign n2365 = n1912 | n2364 ;
  assign n2366 = n2362 & ~n2365 ;
  buffer buf_n2367( .i (n2366), .o (n2367) );
  buffer buf_n2368( .i (n2367), .o (n2368) );
  buffer buf_n2369( .i (n2368), .o (n2369) );
  buffer buf_n898( .i (G51), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  assign n2370 = n904 & ~n1918 ;
  buffer buf_n996( .i (G62), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  assign n2371 = n1002 & ~n1918 ;
  assign n2372 = n2370 | n2371 ;
  assign n2373 = n2369 & ~n2372 ;
  buffer buf_n2374( .i (n2373), .o (n2374) );
  assign n2375 = n340 & ~n2374 ;
  assign n2376 = n341 | n2375 ;
  buffer buf_n2377( .i (n2376), .o (n2377) );
  buffer buf_n2378( .i (n2377), .o (n2378) );
  buffer buf_n2379( .i (n2378), .o (n2379) );
  buffer buf_n2380( .i (n2379), .o (n2380) );
  buffer buf_n2381( .i (n2380), .o (n2381) );
  buffer buf_n2382( .i (n2381), .o (n2382) );
  buffer buf_n2383( .i (n2382), .o (n2383) );
  buffer buf_n2384( .i (n2383), .o (n2384) );
  buffer buf_n2385( .i (n2384), .o (n2385) );
  buffer buf_n2386( .i (n2385), .o (n2386) );
  buffer buf_n2387( .i (n2386), .o (n2387) );
  buffer buf_n2388( .i (n2387), .o (n2388) );
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2391( .i (n2390), .o (n2391) );
  buffer buf_n2392( .i (n2391), .o (n2392) );
  buffer buf_n2393( .i (n2392), .o (n2393) );
  buffer buf_n728( .i (G29), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  assign n2394 = n1524 | n2016 ;
  assign n2395 = n1524 & ~n2016 ;
  assign n2396 = n2394 & ~n2395 ;
  buffer buf_n2397( .i (n2396), .o (n2397) );
  assign n2398 = n1497 | n2397 ;
  assign n2399 = ~n1497 & n2397 ;
  assign n2400 = n2398 & ~n2399 ;
  assign n2401 = n740 | n2400 ;
  buffer buf_n2402( .i (n2401), .o (n2402) );
  buffer buf_n2403( .i (n2402), .o (n2403) );
  buffer buf_n2404( .i (n2403), .o (n2404) );
  buffer buf_n2405( .i (n2404), .o (n2405) );
  buffer buf_n2406( .i (n2405), .o (n2406) );
  buffer buf_n2407( .i (n2406), .o (n2407) );
  buffer buf_n2408( .i (n2407), .o (n2408) );
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  buffer buf_n2411( .i (n2410), .o (n2411) );
  buffer buf_n2412( .i (n2411), .o (n2412) );
  buffer buf_n2413( .i (n2412), .o (n2413) );
  buffer buf_n2414( .i (n2413), .o (n2414) );
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n2416( .i (n2415), .o (n2416) );
  buffer buf_n2417( .i (n2416), .o (n2417) );
  assign n2418 = n352 & ~n2374 ;
  buffer buf_n2419( .i (n351), .o (n2419) );
  buffer buf_n2420( .i (n2419), .o (n2420) );
  assign n2421 = n2418 | n2420 ;
  buffer buf_n2422( .i (n2421), .o (n2422) );
  buffer buf_n2423( .i (n2422), .o (n2423) );
  buffer buf_n2424( .i (n2423), .o (n2424) );
  buffer buf_n2425( .i (n2424), .o (n2425) );
  buffer buf_n2426( .i (n2425), .o (n2426) );
  buffer buf_n2427( .i (n2426), .o (n2427) );
  buffer buf_n2428( .i (n2427), .o (n2428) );
  buffer buf_n2429( .i (n2428), .o (n2429) );
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  buffer buf_n2432( .i (n2431), .o (n2432) );
  buffer buf_n2433( .i (n2432), .o (n2433) );
  buffer buf_n2434( .i (n2433), .o (n2434) );
  buffer buf_n2435( .i (n2434), .o (n2435) );
  buffer buf_n2436( .i (n2435), .o (n2436) );
  buffer buf_n2437( .i (n2436), .o (n2437) );
  buffer buf_n2438( .i (n2437), .o (n2438) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n1111( .i (G8), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n412( .i (G127), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  assign n2439 = n418 | n1555 ;
  buffer buf_n2440( .i (n2439), .o (n2440) );
  buffer buf_n2441( .i (n2440), .o (n2441) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  buffer buf_n741( .i (G30), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  assign n2443 = n749 | n1495 ;
  buffer buf_n2444( .i (n2443), .o (n2444) );
  assign n2445 = n2442 | n2444 ;
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  assign n2448 = ~n1124 & n2447 ;
  buffer buf_n2449( .i (n2448), .o (n2449) );
  assign n2450 = ~n513 & n2449 ;
  buffer buf_n2451( .i (n2450), .o (n2451) );
  buffer buf_n2452( .i (n2451), .o (n2452) );
  buffer buf_n2453( .i (n2452), .o (n2453) );
  buffer buf_n2454( .i (n2453), .o (n2454) );
  buffer buf_n2455( .i (n2454), .o (n2455) );
  buffer buf_n2456( .i (n2455), .o (n2456) );
  buffer buf_n2457( .i (n2456), .o (n2457) );
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n2460( .i (n2459), .o (n2460) );
  assign n2461 = n1124 | n2447 ;
  buffer buf_n2462( .i (n2461), .o (n2462) );
  assign n2463 = n1860 | n2462 ;
  buffer buf_n2464( .i (n2463), .o (n2464) );
  buffer buf_n2465( .i (n2464), .o (n2465) );
  buffer buf_n2466( .i (n2465), .o (n2466) );
  buffer buf_n2467( .i (n2466), .o (n2467) );
  buffer buf_n2468( .i (n2467), .o (n2468) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  buffer buf_n2470( .i (n2469), .o (n2470) );
  buffer buf_n2471( .i (n2470), .o (n2471) );
  buffer buf_n2472( .i (n2471), .o (n2472) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  assign n2473 = ~n497 & n2449 ;
  buffer buf_n2474( .i (n2473), .o (n2474) );
  buffer buf_n2475( .i (n2474), .o (n2475) );
  buffer buf_n2476( .i (n2475), .o (n2476) );
  buffer buf_n2477( .i (n2476), .o (n2477) );
  buffer buf_n2478( .i (n2477), .o (n2478) );
  buffer buf_n2479( .i (n2478), .o (n2479) );
  buffer buf_n2480( .i (n2479), .o (n2480) );
  buffer buf_n2481( .i (n2480), .o (n2481) );
  buffer buf_n446( .i (n445), .o (n446) );
  assign n2482 = n446 & n2447 ;
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  assign n2483 = n625 & ~n2447 ;
  assign n2484 = n2482 & ~n2483 ;
  assign n2485 = n1666 & ~n2484 ;
  buffer buf_n2486( .i (n2485), .o (n2486) );
  buffer buf_n2487( .i (n2486), .o (n2487) );
  buffer buf_n2488( .i (n2487), .o (n2488) );
  buffer buf_n2489( .i (n2488), .o (n2489) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n2490( .i (n2446), .o (n2490) );
  assign n2491 = ~n432 & n2490 ;
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  assign n2492 = n608 & ~n2490 ;
  assign n2493 = n2491 | n2492 ;
  buffer buf_n2494( .i (n2493), .o (n2494) );
  assign n2495 = ~n1797 & n2494 ;
  buffer buf_n2496( .i (n2495), .o (n2496) );
  buffer buf_n2497( .i (n2496), .o (n2497) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  buffer buf_n411( .i (n410), .o (n411) );
  assign n2498 = ~n411 & n2490 ;
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  assign n2499 = n594 & ~n2490 ;
  assign n2500 = n2498 | n2499 ;
  buffer buf_n2501( .i (n2500), .o (n2501) );
  assign n2502 = n1929 | n2501 ;
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n2503( .i (n2446), .o (n2503) );
  assign n2504 = ~n397 & n2503 ;
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  assign n2505 = n550 & ~n2503 ;
  assign n2506 = n2504 | n2505 ;
  assign n2507 = ~n1699 & n2506 ;
  buffer buf_n2508( .i (n2507), .o (n2508) );
  assign n2509 = n2502 & n2508 ;
  assign n2510 = n1929 & n2501 ;
  assign n2511 = n1797 & n2494 ;
  assign n2512 = n2510 | n2511 ;
  assign n2513 = n2509 | n2512 ;
  assign n2514 = ~n2497 & n2513 ;
  assign n2515 = n2489 | n2514 ;
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  assign n2516 = n1127 & ~n1634 ;
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  assign n2517 = n465 & n2449 ;
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  assign n2518 = n641 & ~n2462 ;
  assign n2519 = n2517 & ~n2518 ;
  assign n2520 = n2516 & ~n2519 ;
  buffer buf_n2521( .i (n2520), .o (n2521) );
  assign n2522 = n2488 | n2521 ;
  buffer buf_n2523( .i (n2522), .o (n2523) );
  assign n2524 = n2515 & ~n2523 ;
  assign n2525 = n1119 & ~n1593 ;
  buffer buf_n2526( .i (n2525), .o (n2526) );
  buffer buf_n2527( .i (n2526), .o (n2527) );
  buffer buf_n2528( .i (n2527), .o (n2528) );
  buffer buf_n2529( .i (n2528), .o (n2529) );
  buffer buf_n2530( .i (n2529), .o (n2530) );
  buffer buf_n2531( .i (n2530), .o (n2531) );
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n2532), .o (n2533) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  assign n2534 = n481 & n2449 ;
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  assign n2535 = n657 & ~n2462 ;
  assign n2536 = n2534 & ~n2535 ;
  assign n2537 = n2533 & ~n2536 ;
  buffer buf_n2538( .i (n2537), .o (n2538) );
  assign n2539 = n2521 | n2538 ;
  buffer buf_n2540( .i (n2539), .o (n2540) );
  buffer buf_n2541( .i (n2540), .o (n2541) );
  assign n2542 = n2524 | n2541 ;
  assign n2543 = n1827 & ~n2462 ;
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  assign n2547 = n2538 | n2546 ;
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  assign n2551 = n2542 & ~n2550 ;
  assign n2552 = n2481 | n2551 ;
  assign n2553 = n2472 & n2552 ;
  assign n2554 = n2460 | n2553 ;
  assign n2555 = n2442 & ~n2444 ;
  buffer buf_n2556( .i (n2555), .o (n2556) );
  buffer buf_n2557( .i (n2556), .o (n2557) );
  assign n2558 = n544 | n2206 ;
  buffer buf_n2559( .i (n2558), .o (n2559) );
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  buffer buf_n2563( .i (n2562), .o (n2563) );
  assign n2564 = n2557 & ~n2563 ;
  buffer buf_n2565( .i (n2564), .o (n2565) );
  assign n2566 = n588 | n2244 ;
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n2568( .i (n2567), .o (n2568) );
  buffer buf_n2569( .i (n2568), .o (n2569) );
  buffer buf_n2570( .i (n2569), .o (n2570) );
  buffer buf_n2571( .i (n2570), .o (n2571) );
  assign n2572 = n2557 & ~n2571 ;
  buffer buf_n2573( .i (n2572), .o (n2573) );
  assign n2577 = n2565 & ~n2573 ;
  buffer buf_n2578( .i (n2577), .o (n2578) );
  assign n2579 = n534 | n2055 ;
  buffer buf_n2580( .i (n2579), .o (n2580) );
  buffer buf_n2581( .i (n2580), .o (n2581) );
  buffer buf_n2582( .i (n2581), .o (n2582) );
  assign n2587 = n524 & ~n1889 ;
  assign n2588 = n2582 & ~n2587 ;
  buffer buf_n2589( .i (n2588), .o (n2589) );
  assign n2590 = n2557 & ~n2589 ;
  buffer buf_n2591( .i (n2590), .o (n2591) );
  assign n2592 = n2573 | n2591 ;
  assign n2593 = n534 & ~n2055 ;
  buffer buf_n2594( .i (n2593), .o (n2594) );
  assign n2595 = n2559 & ~n2594 ;
  buffer buf_n2596( .i (n2595), .o (n2596) );
  buffer buf_n2597( .i (n2596), .o (n2597) );
  buffer buf_n2598( .i (n2597), .o (n2598) );
  assign n2599 = n2557 & ~n2598 ;
  buffer buf_n2600( .i (n2599), .o (n2600) );
  assign n2602 = n524 | n1889 ;
  buffer buf_n2603( .i (n2602), .o (n2603) );
  buffer buf_n2604( .i (n2603), .o (n2604) );
  buffer buf_n2605( .i (n2556), .o (n2605) );
  assign n2606 = ~n2604 & n2605 ;
  buffer buf_n2607( .i (n2606), .o (n2607) );
  assign n2608 = n2600 | n2607 ;
  assign n2609 = n2592 | n2608 ;
  assign n2610 = n2578 & ~n2609 ;
  buffer buf_n2611( .i (n2610), .o (n2611) );
  buffer buf_n2612( .i (n2611), .o (n2612) );
  buffer buf_n2613( .i (n2612), .o (n2613) );
  buffer buf_n2614( .i (n2613), .o (n2614) );
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  buffer buf_n2617( .i (n2616), .o (n2617) );
  buffer buf_n2618( .i (n2617), .o (n2618) );
  buffer buf_n2619( .i (n2618), .o (n2619) );
  assign n2620 = n2554 & n2619 ;
  buffer buf_n2574( .i (n2573), .o (n2574) );
  buffer buf_n2575( .i (n2574), .o (n2575) );
  buffer buf_n2576( .i (n2575), .o (n2576) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  buffer buf_n2583( .i (n2582), .o (n2583) );
  buffer buf_n2584( .i (n2583), .o (n2584) );
  buffer buf_n2585( .i (n2584), .o (n2585) );
  buffer buf_n2586( .i (n2585), .o (n2586) );
  assign n2621 = n2586 & ~n2607 ;
  assign n2622 = n2601 & ~n2621 ;
  assign n2623 = n2578 & ~n2622 ;
  assign n2624 = n2576 | n2623 ;
  buffer buf_n2625( .i (n2624), .o (n2625) );
  buffer buf_n2626( .i (n2625), .o (n2626) );
  buffer buf_n2627( .i (n2626), .o (n2627) );
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  buffer buf_n2631( .i (n2630), .o (n2631) );
  buffer buf_n2632( .i (n2631), .o (n2632) );
  buffer buf_n2633( .i (n2632), .o (n2633) );
  assign n2634 = n2620 | n2633 ;
  assign n2635 = n164 & ~n1457 ;
  buffer buf_n2636( .i (n2635), .o (n2636) );
  buffer buf_n2637( .i (n2636), .o (n2637) );
  buffer buf_n2638( .i (n2637), .o (n2638) );
  buffer buf_n2639( .i (n2638), .o (n2639) );
  buffer buf_n2640( .i (n2639), .o (n2640) );
  buffer buf_n2641( .i (n2640), .o (n2641) );
  buffer buf_n2642( .i (n2641), .o (n2642) );
  assign n2643 = n2402 & n2642 ;
  buffer buf_n2644( .i (n2643), .o (n2644) );
  buffer buf_n2645( .i (n2644), .o (n2645) );
  buffer buf_n2646( .i (n2645), .o (n2646) );
  buffer buf_n2647( .i (n2646), .o (n2647) );
  buffer buf_n2648( .i (n2647), .o (n2648) );
  buffer buf_n2649( .i (n2648), .o (n2649) );
  buffer buf_n2650( .i (n2649), .o (n2650) );
  buffer buf_n2651( .i (n2650), .o (n2651) );
  buffer buf_n2652( .i (n2651), .o (n2652) );
  buffer buf_n2653( .i (n2652), .o (n2653) );
  buffer buf_n2654( .i (n2653), .o (n2654) );
  buffer buf_n2655( .i (n2654), .o (n2655) );
  buffer buf_n2656( .i (n2655), .o (n2656) );
  buffer buf_n2657( .i (n2656), .o (n2657) );
  assign G2531 = n294 ;
  assign G2532 = n294 ;
  assign G2533 = n294 ;
  assign G2534 = n383 ;
  assign G2535 = n383 ;
  assign G2536 = n580 ;
  assign G2537 = n580 ;
  assign G2538 = n580 ;
  assign G2539 = n782 ;
  assign G2540 = n236 ;
  assign G2541 = n1035 ;
  assign G2542 = n1099 ;
  assign G2543 = n941 ;
  assign G2544 = n1238 ;
  assign G2545 = n849 ;
  assign G2546 = n1176 ;
  assign G2547 = n1279 ;
  assign G2548 = n1308 ;
  assign G2549 = n294 ;
  assign G2550 = n1336 ;
  assign G2551 = n1365 ;
  assign G2552 = n1392 ;
  assign G2553 = n1419 ;
  assign G2554 = n1453 ;
  assign G2555 = n1453 ;
  assign G2556 = n1480 ;
  assign G2557 = n1516 ;
  assign G2558 = n1546 ;
  assign G2559 = n1578 ;
  assign G2560 = n1614 ;
  assign G2561 = n1647 ;
  assign G2562 = n1680 ;
  assign G2563 = n1718 ;
  assign G2564 = n1747 ;
  assign G2565 = n1777 ;
  assign G2566 = n1810 ;
  assign G2567 = n1680 ;
  assign G2568 = n1647 ;
  assign G2569 = n1614 ;
  assign G2570 = n1841 ;
  assign G2571 = n1874 ;
  assign G2572 = n1908 ;
  assign G2573 = n1948 ;
  assign G2574 = n1948 ;
  assign G2575 = n1967 ;
  assign G2576 = n1967 ;
  assign G2577 = n1986 ;
  assign G2578 = n2007 ;
  assign G2579 = n2007 ;
  assign G2580 = n2039 ;
  assign G2581 = ~n187 ;
  assign G2582 = 1'b0 ;
  assign G2583 = 1'b0 ;
  assign G2584 = n2360 ;
  assign G2585 = n2360 ;
  assign G2586 = n2393 ;
  assign G2587 = ~n2417 ;
  assign G2588 = n2438 ;
  assign G2589 = n2438 ;
  assign G2590 = 1'b0 ;
  assign G2591 = ~n2634 ;
  assign G2592 = 1'b0 ;
  assign G2593 = ~n2657 ;
  assign G2594 = ~n2657 ;
endmodule
