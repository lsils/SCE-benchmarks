module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G6 , G7 , G8 , G9 , G3519 , G3520 , G3521 , G3522 , G3523 , G3524 , G3525 , G3526 , G3527 , G3528 , G3529 , G3530 , G3531 , G3532 , G3533 , G3534 , G3535 , G3536 , G3537 , G3538 , G3539 , G3540 );
  input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G6 , G7 , G8 , G9 ;
  output G3519 , G3520 , G3521 , G3522 , G3523 , G3524 , G3525 , G3526 , G3527 , G3528 , G3529 , G3530 , G3531 , G3532 , G3533 , G3534 , G3535 , G3536 , G3537 , G3538 , G3539 , G3540 ;
  wire n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 ;
  assign n51 = G8 | G9 ;
  buffer buf_n52( .i (n51), .o (n52) );
  assign n53 = G10 | G7 ;
  buffer buf_n54( .i (n53), .o (n54) );
  assign n57 = ~n52 & ~n54 ;
  assign n58 = G12 | G13 ;
  buffer buf_n59( .i (n58), .o (n59) );
  assign n60 = ~G11 | ~n59 ;
  assign n61 = G1 | G3 ;
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  assign n64 = G32 & ~G9 ;
  assign n65 = G31 & ~G8 ;
  assign n66 = n64 | n65 ;
  assign n67 = ~G13 & G36 ;
  assign n68 = ~G14 & G37 ;
  assign n69 = n67 | n68 ;
  assign n70 = n66 | n69 ;
  assign n71 = ~G11 & G34 ;
  assign n72 = ~G12 & G35 ;
  assign n73 = n71 | n72 ;
  assign n74 = ~G10 & G33 ;
  assign n75 = G30 & ~G7 ;
  assign n76 = n74 | n75 ;
  assign n77 = n73 | n76 ;
  assign n78 = n70 | n77 ;
  assign n79 = n63 & n78 ;
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  assign n82 = ~G1 & G2 ;
  buffer buf_n83( .i (n82), .o (n83) );
  assign n84 = ~G3 & n83 ;
  buffer buf_n85( .i (n84), .o (n85) );
  assign n86 = ~G7 & n52 ;
  buffer buf_n87( .i (n86), .o (n87) );
  assign n90 = n85 & n87 ;
  assign n91 = G2 | n62 ;
  buffer buf_n92( .i (n91), .o (n92) );
  assign n93 = G35 | G36 ;
  assign n94 = G34 & n93 ;
  assign n95 = ~n92 & n94 ;
  assign n96 = n90 | n95 ;
  assign n97 = ~n81 & ~n96 ;
  assign n98 = G36 | G37 ;
  assign n99 = G36 & G37 ;
  assign n100 = n98 & ~n99 ;
  buffer buf_n101( .i (n100), .o (n101) );
  assign n102 = G34 & ~G35 ;
  assign n103 = ~G34 & G35 ;
  assign n104 = n102 | n103 ;
  buffer buf_n105( .i (n104), .o (n105) );
  assign n106 = n101 | n105 ;
  assign n107 = n101 & n105 ;
  assign n108 = n106 & ~n107 ;
  buffer buf_n109( .i (n108), .o (n109) );
  assign n110 = G30 & ~G31 ;
  assign n111 = ~G30 & G31 ;
  assign n112 = n110 | n111 ;
  buffer buf_n113( .i (n112), .o (n113) );
  assign n114 = G32 | G33 ;
  assign n115 = G32 & G33 ;
  assign n116 = n114 & ~n115 ;
  buffer buf_n117( .i (n116), .o (n117) );
  assign n118 = n113 | n117 ;
  assign n119 = n113 & n117 ;
  assign n120 = n118 & ~n119 ;
  buffer buf_n121( .i (n120), .o (n121) );
  assign n122 = n109 | n121 ;
  assign n123 = n109 & n121 ;
  assign n124 = n122 & ~n123 ;
  assign n125 = G8 & G9 ;
  assign n126 = n52 & ~n125 ;
  buffer buf_n127( .i (n126), .o (n127) );
  assign n128 = G10 & G7 ;
  assign n129 = n54 & ~n128 ;
  buffer buf_n130( .i (n129), .o (n130) );
  assign n131 = ~n127 & n130 ;
  assign n132 = n127 & ~n130 ;
  assign n133 = n131 | n132 ;
  buffer buf_n134( .i (n133), .o (n134) );
  assign n135 = ~G11 & G13 ;
  assign n136 = G11 & ~G13 ;
  assign n137 = n135 | n136 ;
  buffer buf_n138( .i (n137), .o (n138) );
  assign n139 = G12 | G14 ;
  assign n140 = G12 & G14 ;
  assign n141 = n139 & ~n140 ;
  buffer buf_n142( .i (n141), .o (n142) );
  assign n143 = n138 & ~n142 ;
  assign n144 = ~n138 & n142 ;
  assign n145 = n143 | n144 ;
  buffer buf_n146( .i (n145), .o (n146) );
  assign n147 = n134 & n146 ;
  assign n148 = n134 | n146 ;
  assign n149 = ~n147 & n148 ;
  assign n150 = G3 & n83 ;
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  assign n155 = G7 | n153 ;
  assign n156 = ~G1 & G3 ;
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  assign n161 = G1 & G2 ;
  buffer buf_n162( .i (n161), .o (n162) );
  assign n163 = G1 & G3 ;
  assign n164 = G4 & n163 ;
  assign n165 = n162 | n164 ;
  buffer buf_n166( .i (n165), .o (n166) );
  assign n169 = n160 | n166 ;
  buffer buf_n170( .i (n169), .o (n170) );
  assign n171 = G7 & n170 ;
  assign n172 = n155 & ~n171 ;
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  assign n173 = G7 | n52 ;
  assign n174 = G3 & n173 ;
  buffer buf_n175( .i (n174), .o (n175) );
  assign n176 = G3 | G4 ;
  buffer buf_n177( .i (n176), .o (n177) );
  assign n178 = G21 & ~n177 ;
  assign n179 = ~G3 & G4 ;
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  assign n196 = ~G8 & n182 ;
  assign n197 = n178 | n196 ;
  assign n198 = n175 | n197 ;
  assign n199 = n168 & n198 ;
  buffer buf_n200( .i (n199), .o (n200) );
  assign n201 = n172 | n200 ;
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  assign n204 = G25 | G26 ;
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  assign n213 = G5 | G6 ;
  assign n214 = ~G1 & n213 ;
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  assign n219 = G4 & G5 ;
  buffer buf_n220( .i (n219), .o (n220) );
  assign n226 = n162 & ~n220 ;
  buffer buf_n227( .i (n226), .o (n227) );
  assign n230 = G38 & ~n227 ;
  buffer buf_n231( .i (n230), .o (n231) );
  assign n232 = n218 & n231 ;
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  assign n234 = G30 & ~n216 ;
  assign n235 = G4 | G49 ;
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  assign n239 = G28 & ~n238 ;
  assign n240 = G10 & ~G4 ;
  buffer buf_n241( .i (n240), .o (n241) );
  assign n242 = G29 & G4 ;
  assign n243 = n241 | n242 ;
  assign n244 = n239 | n243 ;
  assign n245 = n234 | n244 ;
  assign n246 = ~n229 & n245 ;
  buffer buf_n247( .i (n246), .o (n247) );
  assign n248 = n233 | n247 ;
  buffer buf_n249( .i (n248), .o (n249) );
  assign n250 = n212 & ~n249 ;
  assign n251 = n203 | n250 ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n253 = G23 | G24 ;
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  assign n258 = ~n249 & n257 ;
  assign n259 = n203 & n258 ;
  buffer buf_n260( .i (n259), .o (n260) );
  assign n262 = n252 & ~n260 ;
  buffer buf_n263( .i (n262), .o (n263) );
  assign n264 = G8 & n170 ;
  assign n265 = G8 | n153 ;
  assign n266 = ~n264 & n265 ;
  assign n267 = G3 & n127 ;
  assign n268 = ~G9 & n182 ;
  assign n269 = G22 & ~G3 ;
  buffer buf_n270( .i (n269), .o (n270) );
  assign n276 = ~G4 & n270 ;
  assign n277 = n268 | n276 ;
  assign n278 = n267 | n277 ;
  assign n279 = n168 & n278 ;
  buffer buf_n280( .i (n279), .o (n280) );
  assign n281 = n266 | n280 ;
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  assign n284 = G31 & ~n216 ;
  assign n285 = G29 & ~n238 ;
  assign n286 = G11 | G4 ;
  buffer buf_n287( .i (n286), .o (n287) );
  assign n288 = ~G30 & G4 ;
  assign n289 = n287 & ~n288 ;
  assign n290 = n285 | n289 ;
  assign n291 = n284 | n290 ;
  assign n292 = ~n229 & n291 ;
  buffer buf_n293( .i (n292), .o (n293) );
  assign n294 = n233 | n293 ;
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = n212 & ~n295 ;
  assign n297 = n283 | n296 ;
  buffer buf_n298( .i (n297), .o (n298) );
  assign n299 = n257 & ~n295 ;
  assign n300 = n283 & n299 ;
  buffer buf_n301( .i (n300), .o (n301) );
  assign n302 = n298 & ~n301 ;
  buffer buf_n303( .i (n302), .o (n303) );
  assign n304 = n263 & n303 ;
  buffer buf_n305( .i (n304), .o (n305) );
  assign n306 = G3 & n166 ;
  buffer buf_n307( .i (n306), .o (n307) );
  assign n309 = n170 & ~n307 ;
  assign n310 = G10 & ~n309 ;
  assign n311 = ~G10 & n152 ;
  assign n312 = G8 | n177 ;
  assign n313 = ~G11 & n182 ;
  assign n314 = n312 & ~n313 ;
  assign n315 = n167 & ~n314 ;
  assign n316 = n311 | n315 ;
  buffer buf_n317( .i (n316), .o (n317) );
  assign n318 = n310 | n317 ;
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  assign n321 = G33 & ~n215 ;
  assign n322 = G31 & ~n237 ;
  assign n323 = G13 | G4 ;
  assign n324 = ~G32 & G4 ;
  assign n325 = n323 & ~n324 ;
  assign n326 = n322 | n325 ;
  assign n327 = n321 | n326 ;
  assign n328 = ~n228 & n327 ;
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  assign n331 = n233 | n330 ;
  buffer buf_n332( .i (n331), .o (n332) );
  assign n333 = n212 & ~n332 ;
  assign n334 = n320 | n333 ;
  buffer buf_n335( .i (n334), .o (n335) );
  assign n336 = n257 & ~n332 ;
  assign n337 = n320 & n336 ;
  buffer buf_n338( .i (n337), .o (n338) );
  assign n339 = n335 & ~n338 ;
  buffer buf_n340( .i (n339), .o (n340) );
  assign n351 = n153 | n307 ;
  buffer buf_n352( .i (n351), .o (n352) );
  assign n353 = ~G9 & n352 ;
  assign n354 = G7 & ~n177 ;
  buffer buf_n355( .i (n181), .o (n355) );
  assign n356 = G10 & n355 ;
  assign n357 = n354 | n356 ;
  assign n358 = n167 & n357 ;
  buffer buf_n359( .i (n358), .o (n359) );
  assign n360 = G9 & ~n170 ;
  assign n361 = n359 | n360 ;
  buffer buf_n362( .i (n361), .o (n362) );
  assign n363 = n353 | n362 ;
  buffer buf_n364( .i (n363), .o (n364) );
  assign n365 = G32 & ~n216 ;
  assign n366 = G30 & ~n238 ;
  assign n367 = G12 | G4 ;
  buffer buf_n368( .i (n367), .o (n368) );
  assign n369 = ~G31 & G4 ;
  assign n370 = n368 & ~n369 ;
  assign n371 = n366 | n370 ;
  assign n372 = n365 | n371 ;
  assign n373 = ~n229 & n372 ;
  buffer buf_n374( .i (n373), .o (n374) );
  assign n375 = n233 | n374 ;
  buffer buf_n376( .i (n375), .o (n376) );
  assign n377 = n212 & ~n376 ;
  assign n378 = n364 | n377 ;
  buffer buf_n379( .i (n378), .o (n379) );
  assign n380 = n257 & ~n376 ;
  assign n381 = n364 & n380 ;
  buffer buf_n382( .i (n381), .o (n382) );
  assign n384 = n379 & ~n382 ;
  buffer buf_n385( .i (n384), .o (n385) );
  assign n386 = n340 & n385 ;
  buffer buf_n387( .i (n386), .o (n387) );
  assign n388 = n305 & n387 ;
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  assign n395 = G11 | n59 ;
  assign n396 = G3 & n395 ;
  assign n397 = G9 | n177 ;
  assign n398 = ~G12 & n355 ;
  assign n399 = n397 & ~n398 ;
  assign n400 = ~n396 & n399 ;
  assign n401 = n168 & ~n400 ;
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  assign n404 = ~G1 & G4 ;
  assign n405 = n151 | n404 ;
  assign n406 = n167 | n405 ;
  buffer buf_n407( .i (n406), .o (n407) );
  assign n408 = G11 & ~n407 ;
  buffer buf_n154( .i (n153), .o (n154) );
  assign n409 = ~G11 & n154 ;
  assign n410 = n408 | n409 ;
  assign n411 = n403 | n410 ;
  buffer buf_n412( .i (n411), .o (n412) );
  assign n413 = G32 & ~n237 ;
  assign n414 = G14 | G4 ;
  assign n415 = ~G33 & G4 ;
  assign n416 = n414 & ~n415 ;
  assign n417 = n413 | n416 ;
  assign n418 = G1 | G6 ;
  buffer buf_n419( .i (n418), .o (n419) );
  assign n420 = G38 | n419 ;
  assign n421 = ~G34 & n419 ;
  assign n422 = n420 & ~n421 ;
  buffer buf_n423( .i (n422), .o (n423) );
  assign n424 = n417 | n423 ;
  assign n425 = ~n228 & n424 ;
  buffer buf_n426( .i (n425), .o (n426) );
  assign n427 = n254 & ~n426 ;
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  assign n431 = n412 & n430 ;
  buffer buf_n432( .i (n431), .o (n432) );
  assign n434 = n209 & ~n426 ;
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  assign n438 = n412 | n437 ;
  buffer buf_n439( .i (n438), .o (n439) );
  assign n440 = ~n432 & n439 ;
  buffer buf_n441( .i (n440), .o (n441) );
  assign n442 = G12 | n154 ;
  assign n443 = G12 & n407 ;
  assign n444 = n442 & ~n443 ;
  assign n445 = G12 & G13 ;
  assign n446 = n59 & ~n445 ;
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = n307 & n448 ;
  assign n450 = ~G3 & n162 ;
  buffer buf_n451( .i (n450), .o (n451) );
  assign n452 = G13 & G4 ;
  assign n453 = n241 | n452 ;
  assign n454 = n451 & n453 ;
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  assign n457 = n449 | n456 ;
  buffer buf_n458( .i (n457), .o (n458) );
  assign n459 = n444 | n458 ;
  buffer buf_n460( .i (n459), .o (n460) );
  assign n461 = G5 | n419 ;
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  assign n466 = n231 & ~n465 ;
  buffer buf_n467( .i (n466), .o (n467) );
  assign n468 = G35 & n462 ;
  assign n469 = G33 & ~n237 ;
  assign n470 = G39 | G4 ;
  assign n471 = ~G34 & G4 ;
  assign n472 = n470 & ~n471 ;
  assign n473 = n469 | n472 ;
  assign n474 = n468 | n473 ;
  assign n475 = ~n228 & n474 ;
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  assign n478 = n467 | n477 ;
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n256), .o (n480) );
  assign n481 = ~n479 & n480 ;
  assign n482 = n460 & n481 ;
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n211), .o (n484) );
  assign n485 = ~n479 & n484 ;
  assign n486 = n460 | n485 ;
  buffer buf_n487( .i (n486), .o (n487) );
  assign n488 = ~n483 & n487 ;
  buffer buf_n489( .i (n488), .o (n489) );
  assign n490 = n441 & n489 ;
  buffer buf_n491( .i (n490), .o (n491) );
  assign n492 = ~G13 & n352 ;
  assign n493 = G13 & ~n407 ;
  assign n494 = G14 & G4 ;
  assign n495 = n287 & ~n494 ;
  assign n496 = n451 & ~n495 ;
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  assign n500 = n493 | n499 ;
  assign n501 = n492 | n500 ;
  buffer buf_n502( .i (n501), .o (n502) );
  assign n503 = G36 & n462 ;
  assign n504 = G35 & G4 ;
  assign n505 = ~G4 & G40 ;
  assign n506 = n504 | n505 ;
  buffer buf_n507( .i (n236), .o (n507) );
  assign n508 = G34 & ~n507 ;
  assign n509 = n506 | n508 ;
  assign n510 = n503 | n509 ;
  buffer buf_n511( .i (n227), .o (n511) );
  assign n512 = n510 & ~n511 ;
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  assign n515 = n467 | n514 ;
  buffer buf_n516( .i (n515), .o (n516) );
  assign n517 = n480 & ~n516 ;
  assign n518 = n502 & n517 ;
  buffer buf_n519( .i (n518), .o (n519) );
  assign n524 = n484 & ~n516 ;
  assign n525 = n502 | n524 ;
  buffer buf_n526( .i (n525), .o (n526) );
  assign n527 = ~n519 & n526 ;
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  assign n531 = n491 & n530 ;
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n308( .i (n307), .o (n308) );
  assign n533 = ~n308 & n407 ;
  assign n534 = G14 & ~n533 ;
  assign n535 = ~G14 & n151 ;
  assign n536 = G39 & G4 ;
  assign n537 = n368 & ~n536 ;
  assign n538 = n451 & ~n537 ;
  assign n539 = n535 | n538 ;
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  assign n543 = n534 | n542 ;
  buffer buf_n544( .i (n543), .o (n544) );
  assign n545 = G37 & n462 ;
  assign n546 = G36 & G4 ;
  assign n547 = ~G4 & G41 ;
  assign n548 = n546 | n547 ;
  assign n549 = G35 & ~n507 ;
  assign n550 = n548 | n549 ;
  assign n551 = n545 | n550 ;
  assign n552 = ~n511 & n551 ;
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  assign n555 = n467 | n554 ;
  buffer buf_n556( .i (n555), .o (n556) );
  assign n557 = n480 & ~n556 ;
  assign n558 = n544 & n557 ;
  buffer buf_n559( .i (n558), .o (n559) );
  assign n566 = n484 & ~n556 ;
  assign n567 = n544 | n566 ;
  buffer buf_n568( .i (n567), .o (n568) );
  assign n569 = ~n559 & n568 ;
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  assign n575 = n532 & n574 ;
  buffer buf_n576( .i (n575), .o (n576) );
  assign n577 = n391 & n576 ;
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  assign n578 = n532 & n565 ;
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  assign n579 = n491 & n523 ;
  buffer buf_n433( .i (n432), .o (n433) );
  assign n580 = n439 & n483 ;
  assign n581 = n433 | n580 ;
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  assign n585 = n579 | n584 ;
  buffer buf_n586( .i (n585), .o (n586) );
  assign n587 = n578 | n586 ;
  buffer buf_n588( .i (n587), .o (n588) );
  assign n589 = n392 & n588 ;
  buffer buf_n383( .i (n382), .o (n383) );
  assign n590 = n338 & n379 ;
  assign n591 = n383 | n590 ;
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  assign n594 = n305 & n593 ;
  buffer buf_n261( .i (n260), .o (n261) );
  assign n595 = n252 & n301 ;
  assign n596 = n261 | n595 ;
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  assign n600 = n594 | n599 ;
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  assign n607 = n589 | n604 ;
  assign n608 = G27 & G48 ;
  buffer buf_n609( .i (n608), .o (n609) );
  assign n652 = ~n92 & n609 ;
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  assign n670 = n502 & n658 ;
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  assign n674 = n528 | n673 ;
  assign n675 = n528 & n673 ;
  assign n676 = n674 & ~n675 ;
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  assign n679 = n544 & n658 ;
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  assign n683 = n570 | n682 ;
  assign n684 = n570 & n682 ;
  assign n685 = n683 & ~n684 ;
  buffer buf_n686( .i (n685), .o (n686) );
  assign n687 = G47 & n686 ;
  assign n688 = ~n678 & n687 ;
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  assign n695 = G5 & ~n92 ;
  buffer buf_n696( .i (n695), .o (n696) );
  assign n726 = n89 & ~n696 ;
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  assign n746 = n588 & ~n669 ;
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  assign n754 = ~G1 & n748 ;
  assign n755 = n745 | n754 ;
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  assign n756 = ~G2 & n195 ;
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = n686 & n757 ;
  assign n759 = ~G6 & n696 ;
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  assign n782 = ~G23 & G3 ;
  assign n783 = n83 & ~n782 ;
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  assign n796 = G25 & G3 ;
  buffer buf_n797( .i (n796), .o (n797) );
  assign n798 = G24 & G3 ;
  buffer buf_n799( .i (n798), .o (n799) );
  assign n800 = G26 & ~n799 ;
  buffer buf_n801( .i (n800), .o (n801) );
  assign n802 = n797 & n801 ;
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  assign n809 = G39 | G43 ;
  buffer buf_n810( .i (n809), .o (n810) );
  assign n811 = ~n807 & n810 ;
  assign n812 = ~G3 & G41 ;
  assign n813 = G4 & ~n812 ;
  assign n814 = ~n811 & n813 ;
  assign n815 = G24 | n205 ;
  assign n816 = G3 & n815 ;
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  assign n821 = G40 & n819 ;
  assign n822 = G26 | n799 ;
  buffer buf_n823( .i (n822), .o (n823) );
  assign n824 = n797 | n823 ;
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  assign n830 = G44 & n828 ;
  assign n831 = n821 | n830 ;
  assign n832 = ~n797 & n801 ;
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  assign n839 = G41 | G45 ;
  buffer buf_n840( .i (n839), .o (n840) );
  assign n841 = ~n836 & n840 ;
  assign n842 = n797 & ~n823 ;
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  assign n848 = G42 | G46 ;
  assign n849 = ~n846 & n848 ;
  assign n850 = n841 | n849 ;
  assign n851 = n831 | n850 ;
  assign n852 = n814 & ~n851 ;
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  assign n855 = G3 & n835 ;
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  assign n858 = G11 | n857 ;
  buffer buf_n859( .i (n858), .o (n859) );
  assign n860 = G13 | n805 ;
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  assign n865 = n859 & n864 ;
  assign n866 = G9 | n805 ;
  buffer buf_n867( .i (n866), .o (n867) );
  assign n868 = G7 | n836 ;
  assign n869 = n867 & n868 ;
  assign n870 = G10 | n846 ;
  assign n871 = ~G8 & n828 ;
  assign n872 = n870 & ~n871 ;
  assign n873 = n869 & n872 ;
  assign n874 = G22 & ~n845 ;
  assign n875 = G4 | n874 ;
  buffer buf_n876( .i (n875), .o (n876) );
  assign n877 = ~G12 & n819 ;
  buffer buf_n878( .i (n877), .o (n878) );
  assign n879 = n876 | n878 ;
  assign n880 = n873 & ~n879 ;
  buffer buf_n881( .i (n880), .o (n881) );
  assign n882 = n865 & n881 ;
  assign n883 = n854 | n882 ;
  assign n884 = ~n795 & n883 ;
  assign n885 = n768 & ~n884 ;
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  assign n888 = ~n758 & n887 ;
  buffer buf_n889( .i (n888), .o (n889) );
  assign n890 = G47 & ~n686 ;
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  assign n894 = ~G47 & n686 ;
  assign n895 = n771 | n894 ;
  assign n896 = n891 | n895 ;
  assign n897 = ~n889 & n896 ;
  buffer buf_n898( .i (n897), .o (n898) );
  inverter inv_n1894( .i (n898), .o (n1894) );
  assign n907 = n319 & n657 ;
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  assign n912 = n340 | n911 ;
  assign n913 = n340 & n911 ;
  assign n914 = n912 & ~n913 ;
  buffer buf_n915( .i (n914), .o (n915) );
  assign n924 = ~G2 & G4 ;
  buffer buf_n925( .i (n924), .o (n925) );
  assign n926 = n915 & n925 ;
  assign n927 = G20 & n827 ;
  assign n928 = ~G8 & n817 ;
  assign n929 = G19 & ~n834 ;
  assign n930 = n928 | n929 ;
  assign n931 = n927 | n930 ;
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  assign n935 = G7 | n857 ;
  assign n936 = G18 & ~n845 ;
  assign n937 = ~G21 & G9 ;
  assign n938 = n805 | n937 ;
  assign n939 = ~n936 & n938 ;
  buffer buf_n940( .i (n939), .o (n940) );
  assign n941 = ~n876 & n940 ;
  assign n942 = n935 & n941 ;
  assign n943 = ~n934 & n942 ;
  buffer buf_n829( .i (n828), .o (n829) );
  assign n944 = G40 & n829 ;
  assign n945 = n878 | n944 ;
  buffer buf_n837( .i (n836), .o (n837) );
  assign n946 = G41 & ~n837 ;
  assign n947 = G11 & ~G39 ;
  buffer buf_n948( .i (n947), .o (n948) );
  assign n949 = n807 | n948 ;
  assign n950 = ~n946 & n949 ;
  assign n951 = ~n945 & n950 ;
  assign n952 = G13 | n857 ;
  assign n953 = G14 & ~G42 ;
  buffer buf_n954( .i (n953), .o (n954) );
  assign n955 = n846 | n954 ;
  assign n956 = G4 & n955 ;
  buffer buf_n957( .i (n956), .o (n957) );
  assign n958 = n952 & n957 ;
  assign n959 = n951 & n958 ;
  assign n960 = n943 | n959 ;
  assign n961 = ~n794 & n960 ;
  assign n962 = n767 & ~n961 ;
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  assign n966 = ~n926 & n965 ;
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  assign n978 = n513 | n553 ;
  assign n979 = G24 | n426 ;
  assign n980 = n978 | n979 ;
  buffer buf_n981( .i (n980), .o (n981) );
  assign n982 = n479 | n981 ;
  buffer buf_n983( .i (n982), .o (n983) );
  assign n984 = n516 & n556 ;
  assign n985 = G24 & n426 ;
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  assign n988 = n479 & n987 ;
  assign n989 = n984 & n988 ;
  assign n990 = n983 & ~n989 ;
  assign n991 = n660 | n990 ;
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  assign n1000 = n576 & n668 ;
  assign n1001 = n999 & ~n1000 ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  assign n1003 = G47 & ~n1002 ;
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  assign n1007 = ~n747 & n921 ;
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  assign n1009 = ~n350 & n748 ;
  assign n1010 = n1008 | n1009 ;
  buffer buf_n1011( .i (n1010), .o (n1011) );
  assign n1012 = n1006 | n1011 ;
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  assign n1014 = n1006 & n1011 ;
  assign n1015 = n781 | n1014 ;
  assign n1016 = n1013 & ~n1015 ;
  assign n1017 = n977 | n1016 ;
  buffer buf_n1018( .i (n1017), .o (n1018) );
  assign n1026 = G47 & n1002 ;
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  assign n1029 = n364 & n658 ;
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  assign n1033 = n385 & ~n1032 ;
  assign n1034 = ~n385 & n1032 ;
  assign n1035 = n1033 | n1034 ;
  buffer buf_n1036( .i (n1035), .o (n1036) );
  assign n1046 = n915 & n1036 ;
  buffer buf_n1047( .i (n1046), .o (n1047) );
  assign n1054 = G27 & ~n92 ;
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  assign n1063 = n282 & n1059 ;
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  assign n1068 = n303 | n1067 ;
  assign n1069 = n303 & n1067 ;
  assign n1070 = n1068 & ~n1069 ;
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  assign n1075 = n1047 & n1073 ;
  buffer buf_n1076( .i (n1075), .o (n1076) );
  assign n1082 = n392 & n1076 ;
  assign n1083 = n392 | n1076 ;
  assign n1084 = ~n1082 & n1083 ;
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  assign n1088 = n1028 & ~n1087 ;
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  assign n1091 = n394 | n747 ;
  assign n1092 = ~n606 & n1091 ;
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  assign n1094 = n382 & ~n660 ;
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  assign n1100 = n338 & ~n660 ;
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  assign n1113 = n1036 & ~n1104 ;
  assign n1114 = n1099 | n1113 ;
  buffer buf_n1115( .i (n1114), .o (n1115) );
  assign n1116 = n1074 & n1115 ;
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  assign n1118 = n301 & ~n1062 ;
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  assign n1128 = n1117 | n1127 ;
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  assign n1132 = n1093 & n1131 ;
  assign n1133 = n1093 | n1131 ;
  assign n1134 = ~n1132 & n1133 ;
  buffer buf_n1135( .i (n1134), .o (n1135) );
  assign n1136 = n1090 & n1135 ;
  assign n1137 = n1090 | n1135 ;
  assign n1138 = ~n1136 & n1137 ;
  assign n1139 = G1 | G2 ;
  buffer buf_n1140( .i (n1139), .o (n1140) );
  assign n1145 = n62 & n1140 ;
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  assign n1175 = ~n1138 & n1174 ;
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  assign n1176 = G7 & ~G9 ;
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  assign n1177 = n56 | n127 ;
  assign n1178 = ~n1176 & n1177 ;
  assign n1179 = n1144 | n1178 ;
  assign n1180 = ~G14 & n85 ;
  assign n1181 = ~n447 & n1180 ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  assign n1183 = n1179 & ~n1182 ;
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  assign n1209 = n1175 | ~n1208 ;
  assign n1210 = ~n157 & n419 ;
  assign n1211 = ~n83 & n1210 ;
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n1245( .i (n659), .o (n1245) );
  assign n1246 = n559 & ~n1245 ;
  buffer buf_n1247( .i (n1246), .o (n1247) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  assign n1251 = n677 | n1250 ;
  buffer buf_n1252( .i (n1251), .o (n1252) );
  assign n1253 = n528 & n1247 ;
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  assign n1258 = n1252 & ~n1257 ;
  buffer buf_n1259( .i (n1258), .o (n1259) );
  assign n1260 = n893 | n1259 ;
  assign n1261 = n893 & n1259 ;
  assign n1262 = n1260 & ~n1261 ;
  buffer buf_n1263( .i (n1262), .o (n1263) );
  assign n1264 = n748 & n1263 ;
  assign n1265 = n716 | n1264 ;
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n1270( .i (n657), .o (n1270) );
  assign n1271 = n460 & n1270 ;
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  assign n1275 = n489 | n1274 ;
  assign n1276 = n489 & n1274 ;
  assign n1277 = n1275 & ~n1276 ;
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  assign n1283 = n519 & ~n1245 ;
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  assign n1290 = n1252 & ~n1289 ;
  buffer buf_n1291( .i (n1290), .o (n1291) );
  assign n1292 = n1282 | n1291 ;
  buffer buf_n1293( .i (n1292), .o (n1293) );
  assign n1294 = n1282 & n1291 ;
  buffer buf_n1295( .i (n1294), .o (n1295) );
  assign n1296 = n1293 & ~n1295 ;
  buffer buf_n1297( .i (n1296), .o (n1297) );
  assign n1298 = ~n694 & n1297 ;
  buffer buf_n1299( .i (n1298), .o (n1299) );
  assign n1300 = n694 & ~n1297 ;
  buffer buf_n1301( .i (n1300), .o (n1301) );
  assign n1303 = n1299 | n1301 ;
  buffer buf_n1304( .i (n1303), .o (n1304) );
  assign n1305 = n753 & ~n1304 ;
  assign n1306 = n1269 | n1305 ;
  assign n1307 = ~n1240 & n1306 ;
  buffer buf_n1302( .i (n1301), .o (n1302) );
  assign n1308 = n483 & ~n1245 ;
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  assign n1319 = n1293 & ~n1318 ;
  buffer buf_n1320( .i (n1319), .o (n1320) );
  assign n1321 = n412 & n1270 ;
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  assign n1325 = n441 | n1324 ;
  assign n1326 = n441 & n1324 ;
  assign n1327 = n1325 & ~n1326 ;
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  assign n1337 = n1320 & ~n1336 ;
  assign n1338 = ~n1320 & n1336 ;
  assign n1339 = n1337 | n1338 ;
  buffer buf_n1340( .i (n1339), .o (n1340) );
  assign n1341 = n1302 & ~n1340 ;
  assign n1342 = ~n1302 & n1340 ;
  assign n1343 = n1341 | n1342 ;
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  assign n1346 = ~n1307 & n1345 ;
  assign n1347 = n757 & n1328 ;
  buffer buf_n847( .i (n846), .o (n847) );
  assign n1348 = ~G19 & G7 ;
  buffer buf_n1349( .i (n1348), .o (n1349) );
  assign n1350 = n847 | n1349 ;
  assign n1351 = G21 & n828 ;
  assign n1352 = G20 & ~n836 ;
  assign n1353 = n1351 | n1352 ;
  assign n1354 = n1350 & ~n1353 ;
  buffer buf_n808( .i (n807), .o (n808) );
  assign n1355 = G10 & ~G22 ;
  assign n1356 = n808 | n1355 ;
  assign n1357 = n1354 & n1356 ;
  buffer buf_n1358( .i (n1357), .o (n1358) );
  assign n1359 = ~G9 & n818 ;
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  assign n1363 = G8 | n857 ;
  assign n1364 = ~n1362 & n1363 ;
  assign n1365 = ~G4 & n1364 ;
  assign n1366 = n1358 & n1365 ;
  assign n1367 = n810 & ~n847 ;
  assign n1368 = G12 & ~G40 ;
  buffer buf_n1369( .i (n1368), .o (n1369) );
  assign n1370 = n807 | n1369 ;
  assign n1371 = ~n1367 & n1370 ;
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  assign n1374 = G42 & ~n835 ;
  assign n1375 = G41 & n826 ;
  buffer buf_n1376( .i (n1375), .o (n1376) );
  assign n1377 = n1374 | n1376 ;
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n856), .o (n1381) );
  assign n1382 = G14 | n1381 ;
  buffer buf_n820( .i (n819), .o (n820) );
  assign n1383 = ~G13 & n820 ;
  assign n1384 = G4 & ~n1383 ;
  assign n1385 = n1382 & n1384 ;
  assign n1386 = ~n1380 & n1385 ;
  assign n1387 = n1373 & n1386 ;
  assign n1388 = n1366 | n1387 ;
  assign n1389 = ~n795 & n1388 ;
  assign n1390 = n768 & ~n1389 ;
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  assign n1393 = ~n1347 & n1392 ;
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  assign n1408 = n1346 | n1407 ;
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n747), .o (n1410) );
  assign n1411 = n1263 | n1410 ;
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  assign n1414 = ~n1266 & n1413 ;
  assign n1415 = n1233 & ~n1263 ;
  assign n1416 = n677 & n757 ;
  assign n1417 = G39 & n819 ;
  buffer buf_n1418( .i (n835), .o (n1418) );
  assign n1419 = G44 & ~n1418 ;
  assign n1420 = n1417 | n1419 ;
  buffer buf_n1421( .i (n845), .o (n1421) );
  assign n1422 = n840 & ~n1421 ;
  buffer buf_n1423( .i (n827), .o (n1423) );
  assign n1424 = G43 & n1423 ;
  assign n1425 = n1422 | n1424 ;
  assign n1426 = n1420 | n1425 ;
  assign n1427 = G40 & ~n856 ;
  assign n1428 = n806 | n954 ;
  assign n1429 = G4 & n1428 ;
  assign n1430 = ~n1427 & n1429 ;
  assign n1431 = ~n1426 & n1430 ;
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  assign n1434 = ~G7 & n1423 ;
  assign n1435 = G22 & ~n1418 ;
  assign n1436 = n1434 | n1435 ;
  buffer buf_n1437( .i (n804), .o (n1437) );
  assign n1438 = G12 | n1437 ;
  buffer buf_n1439( .i (n1438), .o (n1439) );
  assign n1440 = G9 | n1421 ;
  assign n1441 = n1439 & n1440 ;
  assign n1442 = ~n1436 & n1441 ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  assign n1445 = G10 | n1381 ;
  buffer buf_n1446( .i (n1445), .o (n1446) );
  assign n1447 = G8 | n1437 ;
  assign n1448 = ~G4 & n1447 ;
  buffer buf_n1449( .i (n1448), .o (n1449) );
  assign n1450 = ~G11 & n818 ;
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n844), .o (n1452) );
  assign n1453 = G21 & ~n1452 ;
  buffer buf_n1454( .i (n1453), .o (n1454) );
  assign n1455 = n1451 | n1454 ;
  assign n1456 = n1449 & ~n1455 ;
  buffer buf_n1457( .i (n1456), .o (n1457) );
  assign n1458 = n1446 & n1457 ;
  assign n1459 = n1444 & n1458 ;
  assign n1460 = n1433 | n1459 ;
  assign n1461 = ~n795 & n1460 ;
  assign n1462 = n768 & ~n1461 ;
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  assign n1465 = ~n1416 & n1464 ;
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  assign n1472 = n1415 | n1471 ;
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  assign n1475 = n1414 | n1474 ;
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n717( .i (n716), .o (n717) );
  assign n1477 = ~n717 & n1412 ;
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  assign n1480 = ~n1304 & n1479 ;
  buffer buf_n1481( .i (n1480), .o (n1481) );
  assign n1482 = n757 & n1278 ;
  buffer buf_n838( .i (n837), .o (n838) );
  assign n1483 = G21 & ~n838 ;
  assign n1484 = G8 | n847 ;
  assign n1485 = G11 & G7 ;
  buffer buf_n1486( .i (n806), .o (n1486) );
  assign n1487 = n1485 | n1486 ;
  assign n1488 = n1484 & n1487 ;
  assign n1489 = ~n1483 & n1488 ;
  assign n1490 = G9 | n1381 ;
  assign n1491 = G20 & ~n1452 ;
  assign n1492 = G4 | n1491 ;
  buffer buf_n1493( .i (n1492), .o (n1493) );
  assign n1496 = ~G10 & n818 ;
  buffer buf_n1497( .i (n1496), .o (n1497) );
  assign n1498 = G22 & n826 ;
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  assign n1501 = n1497 | n1500 ;
  assign n1502 = n1493 | n1501 ;
  assign n1503 = n1490 & ~n1502 ;
  assign n1504 = n1489 & n1503 ;
  assign n1505 = G42 & n826 ;
  buffer buf_n1506( .i (n1505), .o (n1506) );
  assign n1507 = G40 | G44 ;
  assign n1508 = ~n1452 & n1507 ;
  assign n1509 = n1506 | n1508 ;
  buffer buf_n1510( .i (n834), .o (n1510) );
  assign n1511 = G43 & ~n1510 ;
  buffer buf_n1512( .i (n817), .o (n1512) );
  assign n1513 = ~G14 & n1512 ;
  assign n1514 = n1511 | n1513 ;
  assign n1515 = n1509 | n1514 ;
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  assign n1518 = G39 & ~n1381 ;
  assign n1519 = G13 & ~G41 ;
  buffer buf_n1520( .i (n1519), .o (n1520) );
  assign n1521 = n1486 | n1520 ;
  assign n1522 = G4 & n1521 ;
  assign n1523 = ~n1518 & n1522 ;
  assign n1524 = ~n1517 & n1523 ;
  assign n1525 = n1504 | n1524 ;
  assign n1526 = ~n794 & n1525 ;
  assign n1527 = n767 & ~n1526 ;
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  assign n1531 = ~n1482 & n1530 ;
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  buffer buf_n1534( .i (n1533), .o (n1534) );
  buffer buf_n1535( .i (n1534), .o (n1535) );
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  assign n1543 = n717 | n1412 ;
  assign n1544 = ~n1236 & n1543 ;
  buffer buf_n1545( .i (n1544), .o (n1545) );
  assign n1546 = n1304 & ~n1545 ;
  assign n1547 = n1542 | n1546 ;
  assign n1548 = n1481 | n1547 ;
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  assign n1552 = n1028 & n1081 ;
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  assign n1554 = n1027 & n1053 ;
  buffer buf_n1555( .i (n1554), .o (n1555) );
  assign n1556 = n1074 | n1115 ;
  buffer buf_n1557( .i (n1556), .o (n1557) );
  assign n1558 = ~n1117 & n1557 ;
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  assign n1563 = ~n1555 & n1562 ;
  assign n1564 = n1553 | n1563 ;
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  assign n1572 = n1008 | n1112 ;
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  assign n1576 = n923 & n1027 ;
  assign n1577 = n1045 | n1576 ;
  assign n1578 = ~n1555 & n1577 ;
  buffer buf_n1579( .i (n1578), .o (n1579) );
  assign n1580 = n1575 | n1579 ;
  assign n1581 = n1575 & n1579 ;
  assign n1582 = n1580 & ~n1581 ;
  buffer buf_n1583( .i (n1582), .o (n1583) );
  assign n1584 = n1028 & ~n1093 ;
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  assign n1590 = n1583 | n1589 ;
  buffer buf_n1591( .i (n1590), .o (n1591) );
  assign n1592 = n725 | n1591 ;
  assign n1593 = ~n1244 & n1592 ;
  assign n1594 = n1571 & ~n1593 ;
  buffer buf_n1595( .i (n1594), .o (n1595) );
  assign n1596 = ~n725 & n1591 ;
  buffer buf_n1597( .i (n1596), .o (n1597) );
  assign n1598 = ~n1571 & n1597 ;
  assign n1599 = n925 & n1071 ;
  assign n1600 = n847 | n1369 ;
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  assign n1603 = n859 & n1602 ;
  assign n1604 = ~G14 & n829 ;
  assign n1605 = n867 & ~n1497 ;
  assign n1606 = ~n1604 & n1605 ;
  assign n1607 = G39 & ~n837 ;
  assign n1608 = G4 & n861 ;
  assign n1609 = ~n1607 & n1608 ;
  assign n1610 = n1606 & n1609 ;
  buffer buf_n1611( .i (n1610), .o (n1611) );
  assign n1612 = n1603 & n1611 ;
  assign n1613 = G16 & ~n1421 ;
  assign n1614 = G17 & ~n1510 ;
  assign n1615 = G22 & n1512 ;
  assign n1616 = n1614 | n1615 ;
  assign n1617 = n1613 | n1616 ;
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1621( .i (n856), .o (n1621) );
  assign n1622 = G21 & ~n1621 ;
  assign n1623 = G18 & n829 ;
  assign n1624 = n1349 | n1486 ;
  assign n1625 = ~n1623 & n1624 ;
  assign n1626 = ~n1622 & n1625 ;
  assign n1627 = ~n1495 & n1626 ;
  assign n1628 = ~n1620 & n1627 ;
  assign n1629 = n1612 | n1628 ;
  assign n1630 = ~n795 & n1629 ;
  buffer buf_n1631( .i (n767), .o (n1631) );
  assign n1632 = ~n1630 & n1631 ;
  buffer buf_n1633( .i (n1632), .o (n1633) );
  buffer buf_n1634( .i (n1633), .o (n1634) );
  assign n1635 = ~n1599 & n1634 ;
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n1637( .i (n1636), .o (n1637) );
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  assign n1654 = n1598 | n1653 ;
  assign n1655 = n1595 | n1654 ;
  buffer buf_n1656( .i (n1655), .o (n1656) );
  assign n1657 = n202 & n1059 ;
  buffer buf_n1658( .i (n1657), .o (n1658) );
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  assign n1662 = n263 | n1661 ;
  assign n1663 = n263 & n1661 ;
  assign n1664 = n1662 & ~n1663 ;
  buffer buf_n1665( .i (n1664), .o (n1665) );
  assign n1673 = n925 & n1665 ;
  assign n1674 = G18 | G22 ;
  buffer buf_n1675( .i (n1674), .o (n1675) );
  assign n1676 = ~n1437 & n1675 ;
  buffer buf_n1677( .i (n1676), .o (n1677) );
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  assign n1682 = G16 & ~n838 ;
  assign n1683 = G20 & ~n1621 ;
  assign n1684 = n1682 | n1683 ;
  assign n1685 = G17 & n827 ;
  assign n1686 = G15 | G19 ;
  assign n1687 = ~n1452 & n1686 ;
  assign n1688 = n1685 | n1687 ;
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  assign n1689 = G21 & n817 ;
  assign n1690 = n225 & ~n1689 ;
  buffer buf_n1691( .i (n1690), .o (n1691) );
  assign n1692 = ~n1688 & n1691 ;
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  assign n1695 = ~n1684 & n1694 ;
  assign n1696 = ~n1681 & n1695 ;
  assign n1697 = G5 & n1446 ;
  assign n1698 = G14 | n1418 ;
  assign n1699 = ~n1360 & n1698 ;
  assign n1700 = ~G13 & n1423 ;
  assign n1701 = n1439 & ~n1700 ;
  assign n1702 = n1699 & n1701 ;
  buffer buf_n1703( .i (n1421), .o (n1703) );
  assign n1704 = n948 | n1703 ;
  assign n1705 = n1449 & n1704 ;
  assign n1706 = n1702 & n1705 ;
  buffer buf_n1707( .i (n1706), .o (n1707) );
  assign n1708 = n1697 & n1707 ;
  assign n1709 = n1696 | n1708 ;
  buffer buf_n1710( .i (n794), .o (n1710) );
  assign n1711 = n1709 & ~n1710 ;
  assign n1712 = n1631 & ~n1711 ;
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  assign n1715 = ~n1673 & n1714 ;
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  assign n1734 = n1583 & n1589 ;
  buffer buf_n1735( .i (n1734), .o (n1735) );
  assign n1738 = ~n1565 & n1587 ;
  assign n1739 = n722 | n1738 ;
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  assign n1742 = n1735 | n1741 ;
  assign n1743 = ~n1244 & n1742 ;
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  assign n1744 = n1129 & ~n1672 ;
  assign n1745 = ~n1129 & n1672 ;
  assign n1746 = n1744 | n1745 ;
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  assign n1749 = n1553 & ~n1748 ;
  assign n1750 = ~n1553 & n1748 ;
  assign n1751 = n1749 | n1750 ;
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  assign n1758 = ~n1743 & n1757 ;
  assign n1759 = n1733 | n1758 ;
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  assign n1762 = n1597 & ~n1737 ;
  assign n1763 = n925 & n1036 ;
  assign n1764 = G39 & n1423 ;
  assign n1765 = G40 & ~n1418 ;
  assign n1766 = n1764 | n1765 ;
  assign n1767 = G10 & G14 ;
  assign n1768 = n806 | n1767 ;
  assign n1769 = ~n1451 & n1768 ;
  assign n1770 = ~n1766 & n1769 ;
  buffer buf_n1771( .i (n1770), .o (n1771) );
  assign n1772 = G12 | n1621 ;
  assign n1773 = n1520 | n1703 ;
  assign n1774 = G4 & n1773 ;
  assign n1775 = n1772 & n1774 ;
  assign n1776 = n1771 & n1775 ;
  assign n1777 = G17 & ~n1703 ;
  buffer buf_n1778( .i (n825), .o (n1778) );
  assign n1779 = G19 & n1778 ;
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  assign n1782 = n1454 | n1781 ;
  assign n1783 = n1777 | n1782 ;
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  assign n1784 = ~n1510 & n1675 ;
  assign n1785 = n275 | n1784 ;
  assign n1786 = ~G7 & n1512 ;
  assign n1787 = G20 & ~n1437 ;
  assign n1788 = n1786 | n1787 ;
  assign n1789 = n1785 | n1788 ;
  assign n1790 = n1449 & ~n1789 ;
  assign n1791 = ~n1783 & n1790 ;
  buffer buf_n1792( .i (n1791), .o (n1792) );
  assign n1793 = n1776 | n1792 ;
  buffer buf_n1794( .i (n793), .o (n1794) );
  assign n1795 = n1793 & ~n1794 ;
  buffer buf_n1796( .i (n766), .o (n1796) );
  assign n1797 = ~n1795 & n1796 ;
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  assign n1801 = ~n1763 & n1800 ;
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  buffer buf_n1813( .i (n1812), .o (n1813) );
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  assign n1816 = n1241 & ~n1583 ;
  assign n1817 = n1815 | n1816 ;
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  assign n1821 = n1762 | n1820 ;
  buffer buf_n1822( .i (n1821), .o (n1822) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  assign n1823 = n1656 | n1761 ;
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  assign n1825 = n1025 | n1822 ;
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  assign n1827 = n1409 | n1551 ;
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  assign n1829 = n906 & ~n1476 ;
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  assign n1836 = ~n1828 & n1835 ;
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  assign n1840 = ~n1826 & n1839 ;
  assign n1841 = ~n1824 & n1840 ;
  buffer buf_n1842( .i (n1841), .o (n1842) );
  inverter inv_n1895( .i (n1842), .o (n1895) );
  assign n1843 = G48 & ~n1824 ;
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  assign n1846 = G27 & ~n1842 ;
  assign n1847 = n1845 | ~n1846 ;
  assign n1848 = n1025 & n1822 ;
  buffer buf_n1849( .i (n1848), .o (n1849) );
  assign n1850 = n1826 & ~n1849 ;
  buffer buf_n1851( .i (n1850), .o (n1851) );
  assign n1852 = ~n906 & n1476 ;
  buffer buf_n1853( .i (n1852), .o (n1853) );
  assign n1854 = n1830 | n1853 ;
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1860( .i (n1859), .o (n1860) );
  assign n1861 = n1409 & n1551 ;
  buffer buf_n1862( .i (n1861), .o (n1862) );
  assign n1863 = n1828 & ~n1862 ;
  buffer buf_n1864( .i (n1863), .o (n1864) );
  assign n1865 = n1860 | n1864 ;
  assign n1866 = n1860 & n1864 ;
  assign n1867 = n1865 & ~n1866 ;
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  assign n1870 = n1851 & n1869 ;
  assign n1871 = n1851 | n1869 ;
  assign n1872 = ~n1870 & n1871 ;
  buffer buf_n1873( .i (n1872), .o (n1873) );
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n1875( .i (n1874), .o (n1875) );
  assign n1876 = n1656 & n1761 ;
  buffer buf_n1877( .i (n1876), .o (n1877) );
  assign n1878 = n1824 & ~n1877 ;
  buffer buf_n1879( .i (n1878), .o (n1879) );
  assign n1882 = G50 & n1879 ;
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  assign n1884 = G50 | n1879 ;
  assign n1885 = ~n651 & n1884 ;
  assign n1886 = ~n1883 & n1885 ;
  buffer buf_n1887( .i (n1886), .o (n1887) );
  assign n1888 = n1875 & n1887 ;
  assign n1889 = n1875 | n1887 ;
  assign n1890 = n1888 | ~n1889 ;
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1881( .i (n1880), .o (n1881) );
  assign n1891 = n1873 | n1881 ;
  assign n1892 = n1873 & n1881 ;
  assign n1893 = n1891 & ~n1892 ;
  assign G3519 = n57 ;
  assign G3520 = n60 ;
  assign G3521 = n97 ;
  assign G3522 = n124 ;
  assign G3523 = n149 ;
  assign G3524 = n577 ;
  assign G3525 = n607 ;
  assign G3526 = n689 ;
  assign G3527 = n755 ;
  assign G3528 = n1894 ;
  assign G3529 = n1018 ;
  assign G3530 = n1209 ;
  assign G3531 = n1409 ;
  assign G3532 = n1476 ;
  assign G3533 = n1549 ;
  assign G3534 = n1656 ;
  assign G3535 = n1760 ;
  assign G3536 = n1822 ;
  assign G3537 = n1895 ;
  assign G3538 = n1847 ;
  assign G3539 = n1890 ;
  assign G3540 = n1893 ;
endmodule
