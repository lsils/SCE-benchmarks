module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G158 , G159 , G16 , G160 , G161 , G162 , G163 , G164 , G165 , G166 , G167 , G168 , G169 , G17 , G170 , G171 , G172 , G173 , G174 , G175 , G176 , G177 , G178 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 , G5193 , G5194 , G5195 , G5196 , G5197 , G5198 , G5199 , G5200 , G5201 , G5202 , G5203 , G5204 , G5205 , G5206 , G5207 , G5208 , G5209 , G5210 , G5211 , G5212 , G5213 , G5214 , G5215 , G5216 , G5217 , G5218 , G5219 , G5220 , G5221 , G5222 , G5223 , G5224 , G5225 , G5226 , G5227 , G5228 , G5229 , G5230 , G5231 , G5232 , G5233 , G5234 , G5235 , G5236 , G5237 , G5238 , G5239 , G5240 , G5241 , G5242 , G5243 , G5244 , G5245 , G5246 , G5247 , G5248 , G5249 , G5250 , G5251 , G5252 , G5253 , G5254 , G5255 , G5256 , G5257 , G5258 , G5259 , G5260 , G5261 , G5262 , G5263 , G5264 , G5265 , G5266 , G5267 , G5268 , G5269 , G5270 , G5271 , G5272 , G5273 , G5274 , G5275 , G5276 , G5277 , G5278 , G5279 , G5280 , G5281 , G5282 , G5283 , G5284 , G5285 , G5286 , G5287 , G5288 , G5289 , G5290 , G5291 , G5292 , G5293 , G5294 , G5295 , G5296 , G5297 , G5298 , G5299 , G5300 , G5301 , G5302 , G5303 , G5304 , G5305 , G5306 , G5307 , G5308 , G5309 , G5310 , G5311 , G5312 , G5313 , G5314 , G5315 );
  input G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G158 , G159 , G16 , G160 , G161 , G162 , G163 , G164 , G165 , G166 , G167 , G168 , G169 , G17 , G170 , G171 , G172 , G173 , G174 , G175 , G176 , G177 , G178 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 ;
  output G5193 , G5194 , G5195 , G5196 , G5197 , G5198 , G5199 , G5200 , G5201 , G5202 , G5203 , G5204 , G5205 , G5206 , G5207 , G5208 , G5209 , G5210 , G5211 , G5212 , G5213 , G5214 , G5215 , G5216 , G5217 , G5218 , G5219 , G5220 , G5221 , G5222 , G5223 , G5224 , G5225 , G5226 , G5227 , G5228 , G5229 , G5230 , G5231 , G5232 , G5233 , G5234 , G5235 , G5236 , G5237 , G5238 , G5239 , G5240 , G5241 , G5242 , G5243 , G5244 , G5245 , G5246 , G5247 , G5248 , G5249 , G5250 , G5251 , G5252 , G5253 , G5254 , G5255 , G5256 , G5257 , G5258 , G5259 , G5260 , G5261 , G5262 , G5263 , G5264 , G5265 , G5266 , G5267 , G5268 , G5269 , G5270 , G5271 , G5272 , G5273 , G5274 , G5275 , G5276 , G5277 , G5278 , G5279 , G5280 , G5281 , G5282 , G5283 , G5284 , G5285 , G5286 , G5287 , G5288 , G5289 , G5290 , G5291 , G5292 , G5293 , G5294 , G5295 , G5296 , G5297 , G5298 , G5299 , G5300 , G5301 , G5302 , G5303 , G5304 , G5305 , G5306 , G5307 , G5308 , G5309 , G5310 , G5311 , G5312 , G5313 , G5314 , G5315 ;
  wire n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 ;
  assign n179 = G153 & G156 ;
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n187 = G66 & G67 ;
  buffer buf_n188( .i (n187), .o (n188) );
  assign n189 = G1 & G134 ;
  buffer buf_n190( .i (n189), .o (n190) );
  assign n191 = ~G165 & G63 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = G11 & ~G164 ;
  inverter inv_n194( .i (n193), .o (n194) );
  assign n195 = G136 & G154 ;
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  inverter inv_n203( .i (n202), .o (n203) );
  assign n204 = G11 & G12 ;
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  assign n211 = G65 & n208 ;
  inverter inv_n212( .i (n211), .o (n212) );
  buffer buf_n209( .i (n208), .o (n209) );
  inverter inv_n210( .i (n209), .o (n210) );
  assign n213 = G163 & G34 ;
  assign n214 = ~G163 & G33 ;
  assign n215 = n213 | n214 ;
  assign n216 = n208 & n215 ;
  inverter inv_n217( .i (n216), .o (n217) );
  assign n218 = G13 & G163 ;
  assign n219 = ~G163 & G35 ;
  assign n220 = n218 | n219 ;
  assign n221 = n207 & n220 ;
  buffer buf_n222( .i (n221), .o (n222) );
  inverter inv_n223( .i (n222), .o (n223) );
  assign n224 = G32 & n208 ;
  inverter inv_n225( .i (n224), .o (n225) );
  assign n226 = ~G163 & G9 ;
  assign n227 = G163 & G8 ;
  assign n228 = n206 & ~n227 ;
  assign n229 = ~n226 & n228 ;
  assign n230 = G66 & ~n229 ;
  buffer buf_n231( .i (n230), .o (n231) );
  assign n232 = ~G163 & G30 ;
  assign n233 = G10 & G163 ;
  assign n234 = n206 & ~n233 ;
  assign n235 = ~n232 & n234 ;
  assign n236 = G66 & ~n235 ;
  buffer buf_n237( .i (n236), .o (n237) );
  assign n238 = ~G163 & G7 ;
  assign n239 = G163 & G28 ;
  assign n240 = n206 & ~n239 ;
  assign n241 = ~n238 & n240 ;
  assign n242 = G66 & ~n241 ;
  buffer buf_n243( .i (n242), .o (n243) );
  assign n244 = ~G163 & G29 ;
  assign n245 = G163 & G31 ;
  buffer buf_n246( .i (n205), .o (n246) );
  assign n247 = ~n245 & n246 ;
  assign n248 = ~n244 & n247 ;
  assign n249 = G66 & ~n248 ;
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = G100 | G117 ;
  assign n252 = ~G101 & G117 ;
  assign n253 = n251 & ~n252 ;
  assign n254 = G145 & ~n253 ;
  assign n255 = G102 & G117 ;
  assign n256 = ~G117 & G98 ;
  assign n257 = n255 | n256 ;
  assign n258 = ~G145 & n257 ;
  assign n259 = n254 | n258 ;
  buffer buf_n260( .i (n259), .o (n260) );
  assign n270 = G100 | G119 ;
  assign n271 = ~G101 & G119 ;
  assign n272 = n270 & ~n271 ;
  assign n273 = G146 & ~n272 ;
  assign n274 = G102 & G119 ;
  assign n275 = ~G119 & G98 ;
  assign n276 = n274 | n275 ;
  assign n277 = ~G146 & n276 ;
  assign n278 = n273 | n277 ;
  buffer buf_n279( .i (n278), .o (n279) );
  assign n289 = n260 & n279 ;
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  assign n301 = G128 | G169 ;
  assign n302 = G128 & ~G168 ;
  assign n303 = n301 & ~n302 ;
  assign n304 = G150 & ~n303 ;
  assign n305 = G128 & G167 ;
  assign n306 = ~G128 & G166 ;
  assign n307 = n305 | n306 ;
  assign n308 = ~G150 & n307 ;
  assign n309 = n304 | n308 ;
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  assign n312 = G113 | G98 ;
  assign n313 = ~G102 & G113 ;
  assign n314 = n312 & ~n313 ;
  buffer buf_n315( .i (n314), .o (n315) );
  assign n331 = G100 | G115 ;
  assign n332 = ~G101 & G115 ;
  assign n333 = n331 & ~n332 ;
  buffer buf_n334( .i (n333), .o (n334) );
  assign n345 = n315 & ~n334 ;
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  assign n354 = G100 | G130 ;
  assign n355 = ~G101 & G130 ;
  assign n356 = n354 & ~n355 ;
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  assign n370 = ~G148 & G166 ;
  assign n371 = G148 & ~G169 ;
  assign n372 = n370 | n371 ;
  buffer buf_n373( .i (n372), .o (n373) );
  assign n374 = ~n367 & n373 ;
  assign n375 = n353 & n374 ;
  assign n376 = n311 & n375 ;
  assign n377 = G121 | G169 ;
  assign n378 = G121 & ~G168 ;
  assign n379 = n377 & ~n378 ;
  assign n380 = G147 & ~n379 ;
  assign n381 = G121 & G167 ;
  assign n382 = ~G121 & G166 ;
  assign n383 = n381 | n382 ;
  assign n384 = ~G147 & n383 ;
  assign n385 = n380 | n384 ;
  buffer buf_n386( .i (n385), .o (n386) );
  assign n387 = G126 | G169 ;
  assign n388 = G126 & ~G168 ;
  assign n389 = n387 & ~n388 ;
  assign n390 = G149 & ~n389 ;
  assign n391 = G126 & G167 ;
  assign n392 = ~G126 & G166 ;
  assign n393 = n391 | n392 ;
  assign n394 = ~G149 & n393 ;
  assign n395 = n390 | n394 ;
  buffer buf_n396( .i (n395), .o (n396) );
  assign n397 = n386 & n396 ;
  assign n398 = n376 & n397 ;
  assign n399 = n300 & n398 ;
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  assign n408 = G169 | G94 ;
  assign n409 = ~G168 & G94 ;
  assign n410 = n408 & ~n409 ;
  assign n411 = G140 & ~n410 ;
  assign n412 = G167 & G94 ;
  assign n413 = G166 & ~G94 ;
  assign n414 = n412 | n413 ;
  assign n415 = ~G140 & n414 ;
  assign n416 = n411 | n415 ;
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  assign n420 = G169 | G90 ;
  assign n421 = ~G168 & G90 ;
  assign n422 = n420 & ~n421 ;
  assign n423 = G143 & ~n422 ;
  assign n424 = G167 & G90 ;
  assign n425 = G166 & ~G90 ;
  assign n426 = n424 | n425 ;
  assign n427 = ~G143 & n426 ;
  assign n428 = n423 | n427 ;
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  assign n431 = G169 | G92 ;
  assign n432 = ~G168 & G92 ;
  assign n433 = n431 & ~n432 ;
  assign n434 = G144 & ~n433 ;
  assign n435 = G167 & G92 ;
  assign n436 = G166 & ~G92 ;
  assign n437 = n435 | n436 ;
  assign n438 = ~G144 & n437 ;
  assign n439 = n434 | n438 ;
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  assign n442 = n430 & n441 ;
  assign n443 = n419 & n442 ;
  assign n444 = G109 | G169 ;
  assign n445 = G109 & ~G168 ;
  assign n446 = n444 & ~n445 ;
  assign n447 = G135 & ~n446 ;
  assign n448 = G109 & G167 ;
  assign n449 = ~G109 & G166 ;
  assign n450 = n448 | n449 ;
  assign n451 = ~G135 & n450 ;
  assign n452 = n447 | n451 ;
  buffer buf_n453( .i (n452), .o (n453) );
  assign n454 = G169 | G96 ;
  assign n455 = ~G168 & G96 ;
  assign n456 = n454 & ~n455 ;
  assign n457 = G141 & ~n456 ;
  assign n458 = G167 & G96 ;
  assign n459 = G166 & ~G96 ;
  assign n460 = n458 | n459 ;
  assign n461 = ~G141 & n460 ;
  assign n462 = n457 | n461 ;
  buffer buf_n463( .i (n462), .o (n463) );
  assign n464 = n453 & n463 ;
  assign n465 = G107 | G169 ;
  assign n466 = G107 & ~G168 ;
  assign n467 = n465 & ~n466 ;
  assign n468 = G139 & ~n467 ;
  assign n469 = G107 & G167 ;
  assign n470 = ~G107 & G166 ;
  assign n471 = n469 | n470 ;
  assign n472 = ~G139 & n471 ;
  assign n473 = n468 | n472 ;
  buffer buf_n474( .i (n473), .o (n474) );
  assign n475 = G101 | G88 ;
  assign n476 = ~G100 & G88 ;
  assign n477 = n475 & ~n476 ;
  assign n478 = G142 & ~n477 ;
  assign n479 = G88 & G98 ;
  assign n480 = G102 & ~G88 ;
  assign n481 = n479 | n480 ;
  assign n482 = ~G142 & n481 ;
  assign n483 = n478 | n482 ;
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  assign n494 = n474 & n491 ;
  assign n495 = G103 | G169 ;
  assign n496 = G103 & ~G168 ;
  assign n497 = n495 & ~n496 ;
  assign n498 = G137 & ~n497 ;
  assign n499 = G103 & G167 ;
  assign n500 = ~G103 & G166 ;
  assign n501 = n499 | n500 ;
  assign n502 = ~G137 & n501 ;
  assign n503 = n498 | n502 ;
  buffer buf_n504( .i (n503), .o (n504) );
  assign n505 = G105 | G169 ;
  assign n506 = G105 & ~G168 ;
  assign n507 = n505 & ~n506 ;
  assign n508 = G138 & ~n507 ;
  assign n509 = G105 & G167 ;
  assign n510 = ~G105 & G166 ;
  assign n511 = n509 | n510 ;
  assign n512 = ~G138 & n511 ;
  assign n513 = n508 | n512 ;
  buffer buf_n514( .i (n513), .o (n514) );
  assign n515 = n504 & n514 ;
  assign n516 = n494 & n515 ;
  assign n517 = n464 & n516 ;
  assign n518 = n443 & n517 ;
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  assign n527 = G124 & G96 ;
  assign n528 = ~G124 & G97 ;
  assign n529 = n527 | n528 ;
  buffer buf_n530( .i (n529), .o (n530) );
  assign n548 = G141 & n530 ;
  buffer buf_n549( .i (n548), .o (n549) );
  assign n553 = G141 | n530 ;
  buffer buf_n554( .i (n553), .o (n554) );
  assign n557 = ~n549 & n554 ;
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  assign n566 = G109 & G124 ;
  assign n567 = G110 & ~G124 ;
  assign n568 = n566 | n567 ;
  buffer buf_n569( .i (n568), .o (n569) );
  assign n592 = G135 & n569 ;
  buffer buf_n593( .i (n592), .o (n593) );
  assign n605 = G135 | n569 ;
  buffer buf_n606( .i (n605), .o (n606) );
  assign n615 = ~n593 & n606 ;
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  assign n633 = G107 & G124 ;
  assign n634 = G108 & ~G124 ;
  assign n635 = n633 | n634 ;
  buffer buf_n636( .i (n635), .o (n636) );
  assign n659 = G139 | n636 ;
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  assign n669 = G139 & n636 ;
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  assign n686 = n661 & ~n671 ;
  buffer buf_n687( .i (n686), .o (n687) );
  assign n702 = n617 & n687 ;
  buffer buf_n703( .i (n702), .o (n703) );
  assign n707 = G105 & G124 ;
  assign n708 = G106 & ~G124 ;
  assign n709 = n707 | n708 ;
  buffer buf_n710( .i (n709), .o (n710) );
  assign n732 = G138 & n710 ;
  buffer buf_n733( .i (n732), .o (n733) );
  assign n734 = G138 | n710 ;
  buffer buf_n735( .i (n734), .o (n735) );
  assign n738 = ~n733 & n735 ;
  buffer buf_n739( .i (n738), .o (n739) );
  assign n754 = G103 & G124 ;
  assign n755 = G104 & ~G124 ;
  assign n756 = n754 | n755 ;
  buffer buf_n757( .i (n756), .o (n757) );
  assign n779 = G137 | n757 ;
  buffer buf_n780( .i (n779), .o (n780) );
  assign n786 = G137 & n757 ;
  buffer buf_n787( .i (n786), .o (n787) );
  assign n794 = n780 & ~n787 ;
  buffer buf_n795( .i (n794), .o (n795) );
  assign n810 = n739 & n795 ;
  buffer buf_n811( .i (n810), .o (n811) );
  assign n821 = n703 & n811 ;
  buffer buf_n822( .i (n821), .o (n822) );
  assign n833 = n561 & n822 ;
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  assign n844 = G124 & G88 ;
  assign n845 = ~G124 & G89 ;
  assign n846 = n844 | n845 ;
  buffer buf_n847( .i (n846), .o (n847) );
  assign n868 = G142 & n847 ;
  buffer buf_n869( .i (n868), .o (n869) );
  assign n889 = G142 | n847 ;
  buffer buf_n890( .i (n889), .o (n890) );
  assign n909 = ~n869 & n890 ;
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  assign n929 = G124 & G90 ;
  assign n930 = ~G124 & G91 ;
  assign n931 = n929 | n930 ;
  buffer buf_n932( .i (n931), .o (n932) );
  assign n956 = G143 & n932 ;
  buffer buf_n957( .i (n956), .o (n957) );
  assign n974 = G143 | n932 ;
  buffer buf_n975( .i (n974), .o (n975) );
  assign n984 = ~n957 & n975 ;
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  assign n1002 = G124 & G92 ;
  assign n1003 = ~G124 & G93 ;
  assign n1004 = n1002 | n1003 ;
  buffer buf_n1005( .i (n1004), .o (n1005) );
  assign n1031 = G144 & n1005 ;
  buffer buf_n1032( .i (n1031), .o (n1032) );
  assign n1035 = G144 | n1005 ;
  buffer buf_n1036( .i (n1035), .o (n1036) );
  assign n1037 = ~n1032 & n1036 ;
  buffer buf_n1038( .i (n1037), .o (n1038) );
  assign n1057 = G124 & G94 ;
  assign n1058 = ~G124 & G95 ;
  assign n1059 = n1057 | n1058 ;
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1083 = G140 & n1060 ;
  buffer buf_n1084( .i (n1083), .o (n1084) );
  assign n1102 = G140 | n1060 ;
  buffer buf_n1103( .i (n1102), .o (n1103) );
  assign n1121 = ~n1084 & n1103 ;
  buffer buf_n1122( .i (n1121), .o (n1122) );
  assign n1141 = n1038 & n1122 ;
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  assign n1156 = n998 & n1155 ;
  buffer buf_n1157( .i (n1156), .o (n1157) );
  assign n1158 = n925 & n1157 ;
  buffer buf_n1159( .i (n1158), .o (n1159) );
  assign n1160 = n843 & n1159 ;
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  assign n1173 = G123 | G125 ;
  buffer buf_n1174( .i (n1173), .o (n1174) );
  assign n1189 = G148 & n1174 ;
  buffer buf_n1190( .i (n1189), .o (n1190) );
  assign n1199 = G148 | n1174 ;
  buffer buf_n1200( .i (n1199), .o (n1200) );
  assign n1209 = ~n1190 & n1200 ;
  buffer buf_n1210( .i (n1209), .o (n1210) );
  assign n1221 = G123 & G128 ;
  assign n1222 = ~G123 & G129 ;
  assign n1223 = n1221 | n1222 ;
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  assign n1243 = G150 | n1226 ;
  buffer buf_n1244( .i (n1243), .o (n1244) );
  assign n1259 = G123 & G130 ;
  assign n1260 = ~G123 & G131 ;
  assign n1261 = n1259 | n1260 ;
  buffer buf_n1262( .i (n1261), .o (n1262) );
  assign n1282 = G150 & n1224 ;
  buffer buf_n1283( .i (n1282), .o (n1283) );
  assign n1300 = n1262 | n1283 ;
  buffer buf_n1301( .i (n1300), .o (n1301) );
  assign n1306 = n1244 & ~n1301 ;
  buffer buf_n1307( .i (n1306), .o (n1307) );
  assign n1322 = G123 & G126 ;
  assign n1323 = ~G123 & G127 ;
  assign n1324 = n1322 | n1323 ;
  buffer buf_n1325( .i (n1324), .o (n1325) );
  assign n1342 = G149 & n1325 ;
  buffer buf_n1343( .i (n1342), .o (n1343) );
  assign n1346 = G149 | n1325 ;
  buffer buf_n1347( .i (n1346), .o (n1347) );
  assign n1349 = ~n1343 & n1347 ;
  buffer buf_n1350( .i (n1349), .o (n1350) );
  assign n1365 = n1307 & n1350 ;
  buffer buf_n1366( .i (n1365), .o (n1366) );
  assign n1371 = n1210 & n1366 ;
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  assign n1386 = G117 & G123 ;
  assign n1387 = G118 & ~G123 ;
  assign n1388 = n1386 | n1387 ;
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  assign n1393 = G145 & n1390 ;
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  assign n1400 = G145 | n1391 ;
  buffer buf_n1401( .i (n1400), .o (n1401) );
  assign n1405 = ~n1395 & n1401 ;
  buffer buf_n1406( .i (n1405), .o (n1406) );
  assign n1411 = G119 & G123 ;
  assign n1412 = G120 & ~G123 ;
  assign n1413 = n1411 | n1412 ;
  buffer buf_n1414( .i (n1413), .o (n1414) );
  assign n1429 = G146 & n1414 ;
  buffer buf_n1430( .i (n1429), .o (n1430) );
  assign n1438 = G146 | n1414 ;
  buffer buf_n1439( .i (n1438), .o (n1439) );
  assign n1447 = ~n1430 & n1439 ;
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  assign n1457 = n1406 & n1452 ;
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  assign n1464 = G113 & G123 ;
  assign n1465 = G114 & ~G123 ;
  assign n1466 = n1464 | n1465 ;
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  assign n1482 = G115 & G123 ;
  assign n1483 = G116 & ~G123 ;
  assign n1484 = n1482 | n1483 ;
  buffer buf_n1485( .i (n1484), .o (n1485) );
  assign n1488 = n1475 | n1485 ;
  buffer buf_n1489( .i (n1488), .o (n1489) );
  assign n1490 = G122 | G123 ;
  buffer buf_n1491( .i (n1490), .o (n1491) );
  assign n1508 = ~G121 & G123 ;
  assign n1509 = n1491 & ~n1508 ;
  buffer buf_n1510( .i (n1509), .o (n1510) );
  assign n1525 = G147 & n1510 ;
  buffer buf_n1526( .i (n1525), .o (n1526) );
  assign n1534 = G147 | n1510 ;
  buffer buf_n1535( .i (n1534), .o (n1535) );
  assign n1542 = ~n1526 & n1535 ;
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n1556( .i (n1555), .o (n1556) );
  assign n1557 = ~n1489 & n1556 ;
  assign n1558 = n1463 & n1557 ;
  assign n1559 = n1385 & n1558 ;
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  assign n1569 = G113 | G115 ;
  assign n1570 = G113 & G115 ;
  assign n1571 = n1569 & ~n1570 ;
  buffer buf_n1572( .i (n1571), .o (n1572) );
  assign n1573 = G117 & ~G119 ;
  assign n1574 = ~G117 & G119 ;
  assign n1575 = n1573 | n1574 ;
  buffer buf_n1576( .i (n1575), .o (n1576) );
  assign n1577 = ~n1572 & n1576 ;
  assign n1578 = n1572 & ~n1576 ;
  assign n1579 = n1577 | n1578 ;
  buffer buf_n1580( .i (n1579), .o (n1580) );
  assign n1581 = G130 & ~G132 ;
  assign n1582 = ~G130 & G132 ;
  assign n1583 = n1581 | n1582 ;
  buffer buf_n1584( .i (n1583), .o (n1584) );
  assign n1585 = G121 & ~n1584 ;
  assign n1586 = ~G121 & n1584 ;
  assign n1587 = n1585 | n1586 ;
  buffer buf_n1588( .i (n1587), .o (n1588) );
  assign n1589 = G126 & ~G128 ;
  assign n1590 = ~G126 & G128 ;
  assign n1591 = n1589 | n1590 ;
  buffer buf_n1592( .i (n1591), .o (n1592) );
  assign n1593 = n1588 & ~n1592 ;
  assign n1594 = ~n1588 & n1592 ;
  assign n1595 = n1593 | n1594 ;
  buffer buf_n1596( .i (n1595), .o (n1596) );
  assign n1597 = n1580 | n1596 ;
  assign n1598 = n1580 & n1596 ;
  assign n1599 = n1597 & ~n1598 ;
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  inverter inv_n1605( .i (n1604), .o (n1605) );
  assign n1606 = G88 | G90 ;
  assign n1607 = G88 & G90 ;
  assign n1608 = n1606 & ~n1607 ;
  buffer buf_n1609( .i (n1608), .o (n1609) );
  assign n1610 = G92 & ~G94 ;
  assign n1611 = ~G92 & G94 ;
  assign n1612 = n1610 | n1611 ;
  buffer buf_n1613( .i (n1612), .o (n1613) );
  assign n1614 = ~n1609 & n1613 ;
  assign n1615 = n1609 & ~n1613 ;
  assign n1616 = n1614 | n1615 ;
  buffer buf_n1617( .i (n1616), .o (n1617) );
  assign n1618 = G103 | G96 ;
  assign n1619 = G103 & G96 ;
  assign n1620 = n1618 & ~n1619 ;
  buffer buf_n1621( .i (n1620), .o (n1621) );
  assign n1622 = G109 & ~G111 ;
  assign n1623 = ~G109 & G111 ;
  assign n1624 = n1622 | n1623 ;
  buffer buf_n1625( .i (n1624), .o (n1625) );
  assign n1626 = n1621 | n1625 ;
  assign n1627 = n1621 & n1625 ;
  assign n1628 = n1626 & ~n1627 ;
  buffer buf_n1629( .i (n1628), .o (n1629) );
  assign n1630 = G105 & ~G107 ;
  assign n1631 = ~G105 & G107 ;
  assign n1632 = n1630 | n1631 ;
  buffer buf_n1633( .i (n1632), .o (n1633) );
  assign n1634 = n1629 & ~n1633 ;
  assign n1635 = ~n1629 & n1633 ;
  assign n1636 = n1634 | n1635 ;
  buffer buf_n1637( .i (n1636), .o (n1637) );
  assign n1638 = n1617 & n1637 ;
  assign n1639 = n1617 | n1637 ;
  assign n1640 = ~n1638 & n1639 ;
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  inverter inv_n1645( .i (n1644), .o (n1645) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  assign n1646 = n593 & n660 ;
  buffer buf_n1647( .i (n1646), .o (n1647) );
  assign n1653 = n671 | n733 ;
  assign n1654 = n1647 | n1653 ;
  assign n1655 = n737 & n1654 ;
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n796( .i (n795), .o (n796) );
  assign n1666 = n558 & n796 ;
  assign n1667 = n1656 & n1666 ;
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  assign n1668 = n556 & n790 ;
  assign n1669 = n552 | n1668 ;
  assign n1670 = n1667 | n1669 ;
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  assign n1682 = n1159 & n1681 ;
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  assign n1683 = n1036 & n1084 ;
  buffer buf_n1684( .i (n1683), .o (n1684) );
  assign n1690 = n1034 | n1684 ;
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  assign n1706 = n979 & n1693 ;
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  assign n1718 = n973 | n1717 ;
  buffer buf_n1719( .i (n1718), .o (n1719) );
  assign n1720 = n908 & n1719 ;
  assign n1721 = n888 | n1720 ;
  assign n1722 = n1682 | n1721 ;
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  assign n1734 = ~n1475 & n1485 ;
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  inverter inv_n1747( .i (n1746), .o (n1747) );
  assign n1748 = G176 & ~G177 ;
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  assign n1758 = G60 & n1751 ;
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  assign n1759 = ~G21 & n1280 ;
  assign n1760 = G21 & ~n1280 ;
  assign n1761 = n1759 | n1760 ;
  buffer buf_n1762( .i (n1761), .o (n1762) );
  assign n1763 = ~G176 & n1762 ;
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  assign n1764 = G176 & ~n369 ;
  assign n1765 = G177 & ~n1764 ;
  assign n1766 = ~n1763 & n1765 ;
  assign n1767 = n1758 | n1766 ;
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  buffer buf_n1773( .i (n1772), .o (n1773) );
  inverter inv_n1774( .i (n1773), .o (n1774) );
  assign n1775 = G58 & n1750 ;
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n1247( .i (n1246), .o (n1247) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  assign n1776 = n1258 & ~n1299 ;
  assign n1777 = n1279 & ~n1776 ;
  assign n1778 = n1321 | n1777 ;
  buffer buf_n1779( .i (n1778), .o (n1779) );
  assign n1782 = G176 | n1779 ;
  assign n1783 = G176 & n310 ;
  assign n1784 = G177 & ~n1783 ;
  assign n1785 = n1782 & n1784 ;
  assign n1786 = n1775 | n1785 ;
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  inverter inv_n1794( .i (n1793), .o (n1794) );
  assign n1795 = G48 & n1751 ;
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  assign n1796 = G2 & n623 ;
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  assign n1806 = G2 | n632 ;
  assign n1807 = ~n1805 & n1806 ;
  buffer buf_n1808( .i (n1807), .o (n1808) );
  assign n1809 = G176 | n1808 ;
  assign n1810 = G176 & n453 ;
  assign n1811 = G177 & ~n1810 ;
  assign n1812 = n1809 & n1811 ;
  assign n1813 = n1795 | n1812 ;
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n1819( .i (n1818), .o (n1819) );
  inverter inv_n1820( .i (n1819), .o (n1820) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  assign n1821 = n1476 & n1486 ;
  assign n1822 = n1489 & ~n1821 ;
  buffer buf_n1823( .i (n1822), .o (n1823) );
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1825( .i (n1824), .o (n1825) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  assign n1834 = G173 | n1816 ;
  assign n1835 = G173 & ~n1769 ;
  assign n1836 = G172 & ~n1835 ;
  assign n1837 = n1834 & n1836 ;
  assign n1838 = ~G172 & G173 ;
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  assign n1841 = G3 & n1840 ;
  assign n1842 = G172 | G173 ;
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  assign n1845 = G22 & ~n1844 ;
  assign n1846 = n1841 | n1845 ;
  assign n1847 = n1837 | n1846 ;
  buffer buf_n1848( .i (n1847), .o (n1848) );
  assign n1849 = G19 & n1751 ;
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  assign n1850 = n1286 & n1348 ;
  assign n1851 = n1345 | n1850 ;
  buffer buf_n1852( .i (n1851), .o (n1852) );
  assign n1857 = n1192 | n1852 ;
  assign n1858 = n1203 & n1857 ;
  assign n1859 = n1372 | n1858 ;
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  assign n1869 = n1555 | n1868 ;
  assign n1870 = n1555 & n1868 ;
  assign n1871 = n1869 & ~n1870 ;
  buffer buf_n1872( .i (n1871), .o (n1872) );
  assign n1877 = ~G176 & n1872 ;
  assign n1878 = G176 & n386 ;
  assign n1879 = G177 & ~n1878 ;
  assign n1880 = ~n1877 & n1879 ;
  assign n1881 = n1849 | n1880 ;
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  inverter inv_n1888( .i (n1887), .o (n1888) );
  assign n1889 = G59 & n1749 ;
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  assign n1890 = n1370 | n1856 ;
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  assign n1896 = ~n1220 & n1895 ;
  assign n1897 = n1220 & ~n1895 ;
  assign n1898 = n1896 | n1897 ;
  buffer buf_n1899( .i (n1898), .o (n1899) );
  assign n1905 = ~G176 & n1899 ;
  assign n1906 = G176 & n373 ;
  assign n1907 = G177 & ~n1906 ;
  assign n1908 = ~n1905 & n1907 ;
  assign n1909 = n1889 | n1908 ;
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n1915( .i (n1914), .o (n1915) );
  buffer buf_n1916( .i (n1915), .o (n1916) );
  buffer buf_n1917( .i (n1916), .o (n1917) );
  inverter inv_n1918( .i (n1917), .o (n1918) );
  buffer buf_n1919( .i (n1750), .o (n1919) );
  assign n1920 = G50 & n1919 ;
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  assign n1921 = n1299 | n1319 ;
  buffer buf_n1922( .i (n1921), .o (n1922) );
  assign n1923 = n1364 | n1922 ;
  assign n1924 = n1364 & n1922 ;
  assign n1925 = n1923 & ~n1924 ;
  buffer buf_n1926( .i (n1925), .o (n1926) );
  assign n1929 = ~G176 & n1926 ;
  assign n1930 = G176 & n396 ;
  assign n1931 = G177 & ~n1930 ;
  assign n1932 = ~n1929 & n1931 ;
  assign n1933 = n1920 | n1932 ;
  buffer buf_n1934( .i (n1933), .o (n1934) );
  buffer buf_n1935( .i (n1934), .o (n1935) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  inverter inv_n1940( .i (n1939), .o (n1940) );
  assign n1941 = G174 | n1816 ;
  assign n1942 = G174 & ~n1769 ;
  assign n1943 = G175 & ~n1942 ;
  assign n1944 = n1941 & n1943 ;
  assign n1945 = G174 & ~G175 ;
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  assign n1948 = G3 & n1947 ;
  assign n1949 = G174 | G175 ;
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  assign n1952 = G22 & ~n1951 ;
  assign n1953 = n1948 | n1952 ;
  assign n1954 = n1944 | n1953 ;
  buffer buf_n1955( .i (n1954), .o (n1955) );
  assign n1956 = G53 & n1919 ;
  assign n1957 = G2 & n834 ;
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  buffer buf_n1960( .i (n1959), .o (n1960) );
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  assign n1967 = G2 & n832 ;
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  assign n1968 = n785 & n1657 ;
  assign n1969 = n793 | n1968 ;
  buffer buf_n1970( .i (n1969), .o (n1970) );
  buffer buf_n1971( .i (n1970), .o (n1971) );
  buffer buf_n1972( .i (n1971), .o (n1972) );
  assign n1973 = ~n565 & n1972 ;
  assign n1974 = n565 & ~n1972 ;
  assign n1975 = n1973 | n1974 ;
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  assign n1981 = n1967 | n1980 ;
  assign n1982 = ~n1966 & n1981 ;
  buffer buf_n1983( .i (n1982), .o (n1983) );
  assign n1987 = ~G176 & n1983 ;
  assign n1988 = G176 & n463 ;
  assign n1989 = G177 & ~n1988 ;
  assign n1990 = ~n1987 & n1989 ;
  assign n1991 = n1956 | n1990 ;
  buffer buf_n1992( .i (n1991), .o (n1992) );
  buffer buf_n1993( .i (n1992), .o (n1993) );
  buffer buf_n1994( .i (n1993), .o (n1994) );
  buffer buf_n1995( .i (n1994), .o (n1995) );
  buffer buf_n1996( .i (n1995), .o (n1996) );
  buffer buf_n1997( .i (n1996), .o (n1997) );
  inverter inv_n1998( .i (n1997), .o (n1998) );
  assign n1999 = G57 & n1750 ;
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n1658( .i (n1657), .o (n1658) );
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  assign n2000 = n706 & n744 ;
  assign n2001 = n1660 | n2000 ;
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n2003), .o (n2004) );
  buffer buf_n2005( .i (n2004), .o (n2005) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  assign n2007 = G2 | n1665 ;
  assign n2008 = n2006 & n2007 ;
  buffer buf_n2009( .i (n2008), .o (n2009) );
  assign n2010 = ~n809 & n2009 ;
  assign n2011 = n809 & ~n2009 ;
  assign n2012 = n2010 | n2011 ;
  buffer buf_n2013( .i (n2012), .o (n2013) );
  assign n2016 = ~G176 & n2013 ;
  assign n2017 = G176 & n504 ;
  assign n2018 = G177 & ~n2017 ;
  assign n2019 = ~n2016 & n2018 ;
  assign n2020 = n1999 | n2019 ;
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  inverter inv_n2028( .i (n2027), .o (n2028) );
  buffer buf_n2029( .i (n1749), .o (n2029) );
  assign n2030 = G56 & n2029 ;
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  assign n2031 = n604 | n1797 ;
  buffer buf_n2032( .i (n2031), .o (n2032) );
  assign n2037 = n697 & n2032 ;
  buffer buf_n2038( .i (n2037), .o (n2038) );
  assign n2042 = n685 | n2038 ;
  buffer buf_n2043( .i (n2042), .o (n2043) );
  assign n2044 = n753 | n2043 ;
  assign n2045 = n753 & n2043 ;
  assign n2046 = n2044 & ~n2045 ;
  buffer buf_n2047( .i (n2046), .o (n2047) );
  assign n2051 = ~G176 & n2047 ;
  assign n2052 = G176 & n514 ;
  assign n2053 = G177 & ~n2052 ;
  assign n2054 = ~n2051 & n2053 ;
  assign n2055 = n2030 | n2054 ;
  buffer buf_n2056( .i (n2055), .o (n2056) );
  buffer buf_n2057( .i (n2056), .o (n2057) );
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  inverter inv_n2063( .i (n2062), .o (n2063) );
  assign n2064 = G55 & n2029 ;
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n2033( .i (n2032), .o (n2033) );
  buffer buf_n2034( .i (n2033), .o (n2034) );
  buffer buf_n2035( .i (n2034), .o (n2035) );
  buffer buf_n2036( .i (n2035), .o (n2036) );
  assign n2065 = n701 | n2036 ;
  assign n2066 = ~n2041 & n2065 ;
  buffer buf_n2067( .i (n2066), .o (n2067) );
  assign n2069 = ~G176 & n2067 ;
  assign n2070 = G176 & n474 ;
  assign n2071 = G177 & ~n2070 ;
  assign n2072 = ~n2069 & n2071 ;
  assign n2073 = n2064 | n2072 ;
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n2075( .i (n2074), .o (n2075) );
  buffer buf_n2076( .i (n2075), .o (n2076) );
  buffer buf_n2077( .i (n2076), .o (n2077) );
  buffer buf_n2078( .i (n2077), .o (n2078) );
  buffer buf_n2079( .i (n2078), .o (n2079) );
  buffer buf_n2080( .i (n2079), .o (n2080) );
  inverter inv_n2081( .i (n2080), .o (n2081) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  assign n2082 = n1392 & n1468 ;
  assign n2083 = n1392 | n1468 ;
  assign n2084 = ~n2082 & n2083 ;
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2089( .i (n2088), .o (n2089) );
  buffer buf_n2090( .i (n2089), .o (n2090) );
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  assign n2095 = n1428 & n1487 ;
  assign n2096 = n1428 | n1487 ;
  assign n2097 = ~n2095 & n2096 ;
  buffer buf_n2098( .i (n2097), .o (n2098) );
  assign n2099 = ~n2094 & n2098 ;
  assign n2100 = n2094 & ~n2098 ;
  assign n2101 = n2099 | n2100 ;
  buffer buf_n2102( .i (n2101), .o (n2102) );
  assign n2103 = G123 & G132 ;
  assign n2104 = ~G123 & G133 ;
  assign n2105 = n2103 | n2104 ;
  buffer buf_n2106( .i (n2105), .o (n2106) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  assign n2107 = n1242 | n1341 ;
  assign n2108 = n1242 & n1341 ;
  assign n2109 = n2107 & ~n2108 ;
  buffer buf_n2110( .i (n2109), .o (n2110) );
  assign n2111 = n2106 | n2110 ;
  assign n2112 = n2106 & n2110 ;
  assign n2113 = n2111 & ~n2112 ;
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n1522( .i (n1521), .o (n1522) );
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  assign n2115 = n1188 & n1524 ;
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  assign n2116 = G125 | n1507 ;
  assign n2117 = ~n2115 & n2116 ;
  buffer buf_n2118( .i (n2117), .o (n2118) );
  assign n2119 = ~n1281 & n2118 ;
  assign n2120 = n1281 & ~n2118 ;
  assign n2121 = n2119 | n2120 ;
  buffer buf_n2122( .i (n2121), .o (n2122) );
  assign n2123 = n2114 & ~n2122 ;
  assign n2124 = ~n2114 & n2122 ;
  assign n2125 = n2123 | n2124 ;
  buffer buf_n2126( .i (n2125), .o (n2126) );
  assign n2127 = ~n2102 & n2126 ;
  assign n2128 = n2102 & ~n2126 ;
  assign n2129 = n2127 | n2128 ;
  buffer buf_n2130( .i (n2129), .o (n2130) );
  buffer buf_n2131( .i (n2130), .o (n2131) );
  buffer buf_n2132( .i (n2131), .o (n2132) );
  inverter inv_n2133( .i (n2132), .o (n2133) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  assign n2134 = n731 & n778 ;
  assign n2135 = n731 | n778 ;
  assign n2136 = ~n2134 & n2135 ;
  buffer buf_n2137( .i (n2136), .o (n2137) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  assign n2138 = ~n591 & n658 ;
  assign n2139 = n591 & ~n658 ;
  assign n2140 = n2138 | n2139 ;
  buffer buf_n2141( .i (n2140), .o (n2141) );
  assign n2142 = n2137 | n2141 ;
  assign n2143 = n2137 & n2141 ;
  assign n2144 = n2142 & ~n2143 ;
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  assign n2146 = n955 & n1030 ;
  assign n2147 = n955 | n1030 ;
  assign n2148 = ~n2146 & n2147 ;
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  assign n2150 = G111 & G124 ;
  assign n2151 = G112 & ~G124 ;
  assign n2152 = n2150 | n2151 ;
  buffer buf_n2153( .i (n2152), .o (n2153) );
  assign n2154 = n1082 & ~n2153 ;
  assign n2155 = ~n1082 & n2153 ;
  assign n2156 = n2154 | n2155 ;
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  assign n2158 = ~n547 & n867 ;
  assign n2159 = n547 & ~n867 ;
  assign n2160 = n2158 | n2159 ;
  buffer buf_n2161( .i (n2160), .o (n2161) );
  assign n2162 = ~n2157 & n2161 ;
  assign n2163 = n2157 & ~n2161 ;
  assign n2164 = n2162 | n2163 ;
  buffer buf_n2165( .i (n2164), .o (n2165) );
  assign n2166 = ~n2149 & n2165 ;
  assign n2167 = n2149 & ~n2165 ;
  assign n2168 = n2166 | n2167 ;
  buffer buf_n2169( .i (n2168), .o (n2169) );
  assign n2170 = ~n2145 & n2169 ;
  assign n2171 = n2145 & ~n2169 ;
  assign n2172 = n2170 | n2171 ;
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n2174( .i (n2173), .o (n2174) );
  inverter inv_n2175( .i (n2174), .o (n2175) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  assign n2176 = n1674 | n1958 ;
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n2177), .o (n2178) );
  buffer buf_n2179( .i (n2178), .o (n2179) );
  buffer buf_n2180( .i (n2179), .o (n2180) );
  assign n2182 = n1157 & n2180 ;
  assign n2183 = n1719 | n2182 ;
  buffer buf_n2184( .i (n2183), .o (n2184) );
  assign n2185 = n928 | n2184 ;
  assign n2186 = n928 & n2184 ;
  assign n2187 = n2185 & ~n2186 ;
  buffer buf_n2188( .i (n2187), .o (n2188) );
  buffer buf_n2189( .i (n2188), .o (n2189) );
  buffer buf_n2190( .i (n2189), .o (n2190) );
  buffer buf_n2191( .i (n2190), .o (n2191) );
  buffer buf_n2192( .i (n2191), .o (n2192) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  assign n2193 = n1140 | n2181 ;
  assign n2194 = n1140 & n2181 ;
  assign n2195 = n2193 & ~n2194 ;
  buffer buf_n2196( .i (n2195), .o (n2196) );
  buffer buf_n2197( .i (n2196), .o (n2197) );
  buffer buf_n2198( .i (n2197), .o (n2198) );
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n2200( .i (n2199), .o (n2200) );
  buffer buf_n2201( .i (n2200), .o (n2201) );
  buffer buf_n1984( .i (n1983), .o (n1984) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n1986( .i (n1985), .o (n1986) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2014( .i (n2013), .o (n2014) );
  buffer buf_n2015( .i (n2014), .o (n2015) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  assign n2202 = ~n1808 & n2068 ;
  assign n2203 = n2015 & n2202 ;
  assign n2204 = n2050 & n2203 ;
  assign n2205 = n1986 & n2204 ;
  assign n2206 = ~n2201 & n2205 ;
  assign n2207 = n2192 & n2206 ;
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  assign n2208 = n1155 & n2178 ;
  assign n2209 = n1705 | n2208 ;
  buffer buf_n2210( .i (n2209), .o (n2210) );
  assign n2211 = ~n1001 & n2210 ;
  assign n2212 = n1001 & ~n2210 ;
  assign n2213 = n2211 | n2212 ;
  buffer buf_n2214( .i (n2213), .o (n2214) );
  buffer buf_n2215( .i (n2214), .o (n2215) );
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  assign n2221 = n1120 & n2178 ;
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  assign n2222 = n1101 | n2178 ;
  assign n2223 = ~n2221 & n2222 ;
  buffer buf_n2224( .i (n2223), .o (n2224) );
  assign n2225 = n1056 | n2224 ;
  assign n2226 = n1056 & n2224 ;
  assign n2227 = n2225 & ~n2226 ;
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  buffer buf_n2231( .i (n2230), .o (n2231) );
  buffer buf_n2232( .i (n2231), .o (n2232) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  assign n2235 = n2220 & ~n2234 ;
  assign n2236 = n2207 & n2235 ;
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  assign n2240 = n1541 & n1860 ;
  assign n2241 = n1533 | n2240 ;
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  assign n2247 = n1446 & n2243 ;
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  assign n2248 = n1437 | n2243 ;
  assign n2249 = ~n2247 & n2248 ;
  buffer buf_n2250( .i (n2249), .o (n2250) );
  assign n2251 = n1410 & n2250 ;
  assign n2252 = n1410 | n2250 ;
  assign n2253 = ~n2251 & n2252 ;
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  assign n2263 = n1404 & n1437 ;
  assign n2264 = n1399 | n2263 ;
  buffer buf_n2244( .i (n2243), .o (n2244) );
  assign n2265 = n1458 & n2244 ;
  assign n2266 = n2264 | n2265 ;
  buffer buf_n2267( .i (n2266), .o (n2267) );
  assign n2268 = n1486 | n2267 ;
  assign n2269 = n1486 & n2267 ;
  assign n2270 = n2268 & ~n2269 ;
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2273( .i (n2272), .o (n2273) );
  buffer buf_n2274( .i (n2273), .o (n2274) );
  buffer buf_n2275( .i (n2274), .o (n2275) );
  buffer buf_n2276( .i (n2275), .o (n2276) );
  buffer buf_n2277( .i (n2276), .o (n2277) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  buffer buf_n1455( .i (n1454), .o (n1455) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n2246( .i (n2245), .o (n2246) );
  assign n2278 = n1456 & n2246 ;
  assign n2279 = n1456 | n2246 ;
  assign n2280 = ~n2278 & n2279 ;
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n1873( .i (n1872), .o (n1873) );
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  assign n2288 = n1762 & n1823 ;
  assign n2289 = ~n1781 & n2288 ;
  assign n2290 = n1928 & n2289 ;
  assign n2291 = n1904 & n2290 ;
  assign n2292 = n1876 & n2291 ;
  assign n2293 = ~n2287 & n2292 ;
  assign n2294 = ~n2277 & n2293 ;
  assign n2295 = ~n2262 & n2294 ;
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n2297( .i (n2296), .o (n2297) );
  assign n2298 = G158 | n1815 ;
  assign n2299 = G158 & ~n1768 ;
  assign n2300 = G159 & ~n2299 ;
  assign n2301 = n2298 & n2300 ;
  assign n2302 = G158 | G159 ;
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  assign n2305 = G81 & ~n2304 ;
  assign n2306 = G158 & ~G159 ;
  buffer buf_n2307( .i (n2306), .o (n2307) );
  buffer buf_n2308( .i (n2307), .o (n2308) );
  assign n2309 = G80 & n2308 ;
  assign n2310 = n2305 | n2309 ;
  assign n2311 = n2301 | n2310 ;
  assign n2312 = G64 & n2311 ;
  buffer buf_n2313( .i (n2312), .o (n2313) );
  assign n2314 = G160 | n1815 ;
  assign n2315 = G160 & ~n1768 ;
  assign n2316 = G161 & ~n2315 ;
  assign n2317 = n2314 & n2316 ;
  assign n2318 = G160 | G161 ;
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  assign n2321 = G81 & ~n2320 ;
  assign n2322 = G160 & ~G161 ;
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  assign n2325 = G80 & n2324 ;
  assign n2326 = n2321 | n2325 ;
  assign n2327 = n2317 | n2326 ;
  assign n2328 = G64 & n2327 ;
  buffer buf_n2329( .i (n2328), .o (n2329) );
  assign n2330 = G173 | n1994 ;
  assign n2331 = G173 & ~n1883 ;
  assign n2332 = G172 & ~n2331 ;
  assign n2333 = n2330 & n2332 ;
  assign n2334 = G16 & n1840 ;
  assign n2335 = G14 & ~n1844 ;
  assign n2336 = n2334 | n2335 ;
  assign n2337 = n2333 | n2336 ;
  buffer buf_n2338( .i (n2337), .o (n2338) );
  assign n2339 = G173 | n2024 ;
  assign n2340 = G173 & ~n1913 ;
  assign n2341 = G172 & ~n2340 ;
  assign n2342 = n2339 & n2341 ;
  assign n2343 = G6 & ~n1844 ;
  assign n2344 = G27 & n1840 ;
  assign n2345 = n2343 | n2344 ;
  assign n2346 = n2342 | n2345 ;
  buffer buf_n2347( .i (n2346), .o (n2347) );
  assign n2348 = G173 | n2059 ;
  assign n2349 = G173 & ~n1935 ;
  assign n2350 = G172 & ~n2349 ;
  assign n2351 = n2348 & n2350 ;
  assign n2352 = G26 & n1840 ;
  assign n2353 = G5 & ~n1844 ;
  assign n2354 = n2352 | n2353 ;
  assign n2355 = n2351 | n2354 ;
  buffer buf_n2356( .i (n2355), .o (n2356) );
  assign n2357 = G173 | n2077 ;
  assign n2358 = G173 & ~n1789 ;
  assign n2359 = G172 & ~n2358 ;
  assign n2360 = n2357 & n2359 ;
  buffer buf_n2361( .i (n1839), .o (n2361) );
  assign n2362 = G24 & n2361 ;
  buffer buf_n2363( .i (n1843), .o (n2363) );
  assign n2364 = G25 & ~n2363 ;
  assign n2365 = n2362 | n2364 ;
  assign n2366 = n2360 | n2365 ;
  buffer buf_n2367( .i (n2366), .o (n2367) );
  assign n2368 = G174 | n1994 ;
  assign n2369 = G174 & ~n1883 ;
  assign n2370 = G175 & ~n2369 ;
  assign n2371 = n2368 & n2370 ;
  assign n2372 = G14 & ~n1951 ;
  assign n2373 = G16 & n1947 ;
  assign n2374 = n2372 | n2373 ;
  assign n2375 = n2371 | n2374 ;
  buffer buf_n2376( .i (n2375), .o (n2376) );
  assign n2377 = G174 | n2024 ;
  assign n2378 = G174 & ~n1913 ;
  assign n2379 = G175 & ~n2378 ;
  assign n2380 = n2377 & n2379 ;
  assign n2381 = G27 & n1947 ;
  assign n2382 = G6 & ~n1951 ;
  assign n2383 = n2381 | n2382 ;
  assign n2384 = n2380 | n2383 ;
  buffer buf_n2385( .i (n2384), .o (n2385) );
  assign n2386 = G174 | n2059 ;
  assign n2387 = G174 & ~n1935 ;
  assign n2388 = G175 & ~n2387 ;
  assign n2389 = n2386 & n2388 ;
  assign n2390 = G5 & ~n1951 ;
  assign n2391 = G26 & n1947 ;
  assign n2392 = n2390 | n2391 ;
  assign n2393 = n2389 | n2392 ;
  buffer buf_n2394( .i (n2393), .o (n2394) );
  assign n2395 = G174 | n2077 ;
  assign n2396 = G174 & ~n1789 ;
  assign n2397 = G175 & ~n2396 ;
  assign n2398 = n2395 & n2397 ;
  buffer buf_n2399( .i (n1946), .o (n2399) );
  assign n2400 = G24 & n2399 ;
  buffer buf_n2401( .i (n1950), .o (n2401) );
  assign n2402 = G25 & ~n2401 ;
  assign n2403 = n2400 | n2402 ;
  assign n2404 = n2398 | n2403 ;
  buffer buf_n2405( .i (n2404), .o (n2405) );
  assign n2406 = G158 | n1993 ;
  assign n2407 = G158 & ~n1882 ;
  assign n2408 = G159 & ~n2407 ;
  assign n2409 = n2406 & n2408 ;
  assign n2410 = G76 & ~n2304 ;
  assign n2411 = G86 & n2308 ;
  assign n2412 = n2410 | n2411 ;
  assign n2413 = n2409 | n2412 ;
  assign n2414 = G64 & n2413 ;
  buffer buf_n2415( .i (n2414), .o (n2415) );
  assign n2416 = G158 | n2076 ;
  assign n2417 = G158 & ~n1788 ;
  assign n2418 = G159 & ~n2417 ;
  assign n2419 = n2416 & n2418 ;
  assign n2420 = G72 & ~n2304 ;
  assign n2421 = G82 & n2308 ;
  assign n2422 = n2420 | n2421 ;
  assign n2423 = n2419 | n2422 ;
  assign n2424 = G64 & n2423 ;
  buffer buf_n2425( .i (n2424), .o (n2425) );
  assign n2426 = G158 | n2058 ;
  assign n2427 = G158 & ~n1934 ;
  assign n2428 = G159 & ~n2427 ;
  assign n2429 = n2426 & n2428 ;
  assign n2430 = G70 & ~n2304 ;
  assign n2431 = G71 & n2308 ;
  assign n2432 = n2430 | n2431 ;
  assign n2433 = n2429 | n2432 ;
  assign n2434 = G64 & n2433 ;
  buffer buf_n2435( .i (n2434), .o (n2435) );
  assign n2436 = G158 | n2023 ;
  assign n2437 = G158 & ~n1912 ;
  assign n2438 = G159 & ~n2437 ;
  assign n2439 = n2436 & n2438 ;
  buffer buf_n2440( .i (n2303), .o (n2440) );
  assign n2441 = G68 & ~n2440 ;
  buffer buf_n2442( .i (n2307), .o (n2442) );
  assign n2443 = G69 & n2442 ;
  assign n2444 = n2441 | n2443 ;
  assign n2445 = n2439 | n2444 ;
  assign n2446 = G64 & n2445 ;
  buffer buf_n2447( .i (n2446), .o (n2447) );
  assign n2448 = G160 | n1993 ;
  assign n2449 = G160 & ~n1882 ;
  assign n2450 = G161 & ~n2449 ;
  assign n2451 = n2448 & n2450 ;
  assign n2452 = G76 & ~n2320 ;
  assign n2453 = G86 & n2324 ;
  assign n2454 = n2452 | n2453 ;
  assign n2455 = n2451 | n2454 ;
  assign n2456 = G64 & n2455 ;
  buffer buf_n2457( .i (n2456), .o (n2457) );
  assign n2458 = G160 | n2076 ;
  assign n2459 = G160 & ~n1788 ;
  assign n2460 = G161 & ~n2459 ;
  assign n2461 = n2458 & n2460 ;
  assign n2462 = G72 & ~n2320 ;
  assign n2463 = G82 & n2324 ;
  assign n2464 = n2462 | n2463 ;
  assign n2465 = n2461 | n2464 ;
  assign n2466 = G64 & n2465 ;
  buffer buf_n2467( .i (n2466), .o (n2467) );
  assign n2468 = G160 | n2058 ;
  assign n2469 = G160 & ~n1934 ;
  assign n2470 = G161 & ~n2469 ;
  assign n2471 = n2468 & n2470 ;
  assign n2472 = G70 & ~n2320 ;
  assign n2473 = G71 & n2324 ;
  assign n2474 = n2472 | n2473 ;
  assign n2475 = n2471 | n2474 ;
  assign n2476 = G64 & n2475 ;
  buffer buf_n2477( .i (n2476), .o (n2477) );
  assign n2478 = G160 | n2023 ;
  assign n2479 = G160 & ~n1912 ;
  assign n2480 = G161 & ~n2479 ;
  assign n2481 = n2478 & n2480 ;
  buffer buf_n2482( .i (n2319), .o (n2482) );
  assign n2483 = G68 & ~n2482 ;
  buffer buf_n2484( .i (n2323), .o (n2484) );
  assign n2485 = G69 & n2484 ;
  assign n2486 = n2483 | n2485 ;
  assign n2487 = n2481 | n2486 ;
  assign n2488 = G64 & n2487 ;
  buffer buf_n2489( .i (n2488), .o (n2489) );
  assign n2490 = G170 & n1828 ;
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  assign n2491 = ~G61 & n1481 ;
  assign n2492 = G61 & ~n1481 ;
  assign n2493 = n2491 | n2492 ;
  buffer buf_n2494( .i (n2493), .o (n2494) );
  assign n2497 = G170 | n2494 ;
  assign n2498 = ~n2490 & n2497 ;
  assign n2499 = G171 & ~n2498 ;
  assign n2500 = G178 & G62 ;
  assign n2501 = G170 & ~G54 ;
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  assign n2502 = G170 | n330 ;
  assign n2503 = ~n2501 & n2502 ;
  assign n2504 = G171 | n2503 ;
  assign n2505 = ~n2500 & n2504 ;
  assign n2506 = ~n2499 & n2505 ;
  buffer buf_n2507( .i (n2506), .o (n2507) );
  buffer buf_n2495( .i (n2494), .o (n2495) );
  buffer buf_n2496( .i (n2495), .o (n2496) );
  assign n2508 = n1830 & n2496 ;
  assign n2509 = n1830 | n2496 ;
  assign n2510 = ~n2508 & n2509 ;
  inverter inv_n2511( .i (n2510), .o (n2511) );
  assign n2512 = G54 & n1919 ;
  assign n2513 = ~G176 & n1823 ;
  assign n2514 = G176 & ~n325 ;
  assign n2515 = G177 & ~n2514 ;
  assign n2516 = ~n2513 & n2515 ;
  assign n2517 = n2512 | n2516 ;
  buffer buf_n2518( .i (n2517), .o (n2518) );
  buffer buf_n2519( .i (n2518), .o (n2519) );
  buffer buf_n2520( .i (n2519), .o (n2520) );
  buffer buf_n2521( .i (n2520), .o (n2521) );
  buffer buf_n2522( .i (n2521), .o (n2522) );
  buffer buf_n2523( .i (n2522), .o (n2523) );
  inverter inv_n2524( .i (n2523), .o (n2524) );
  assign n2525 = G52 & n1919 ;
  assign n2526 = G176 | n2271 ;
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  assign n2527 = G176 & ~n344 ;
  assign n2528 = G177 & ~n2527 ;
  assign n2529 = n2526 & n2528 ;
  assign n2530 = n2525 | n2529 ;
  buffer buf_n2531( .i (n2530), .o (n2531) );
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n2532), .o (n2533) );
  buffer buf_n2534( .i (n2533), .o (n2534) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  buffer buf_n2536( .i (n2535), .o (n2536) );
  inverter inv_n2537( .i (n2536), .o (n2537) );
  assign n2538 = G47 & n2029 ;
  assign n2539 = G176 | n2254 ;
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  assign n2540 = G176 & n269 ;
  assign n2541 = G177 & ~n2540 ;
  assign n2542 = n2539 & n2541 ;
  assign n2543 = n2538 | n2542 ;
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  inverter inv_n2551( .i (n2550), .o (n2551) );
  assign n2552 = G43 & n2029 ;
  assign n2553 = G176 | n2281 ;
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  assign n2554 = G176 & n288 ;
  assign n2555 = G177 & ~n2554 ;
  assign n2556 = n2553 & n2555 ;
  assign n2557 = n2552 | n2556 ;
  buffer buf_n2558( .i (n2557), .o (n2558) );
  buffer buf_n2559( .i (n2558), .o (n2559) );
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  buffer buf_n2563( .i (n2562), .o (n2563) );
  buffer buf_n2564( .i (n2563), .o (n2564) );
  inverter inv_n2565( .i (n2564), .o (n2565) );
  assign n2566 = G155 & G99 ;
  assign n2567 = n196 & n2566 ;
  assign n2568 = n180 & n2567 ;
  assign n2569 = ~n1600 & n2568 ;
  assign n2570 = ~n1641 & n2569 ;
  assign n2571 = ~n2130 & n2570 ;
  assign n2572 = ~n2173 & n2571 ;
  buffer buf_n2573( .i (n2572), .o (n2573) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  assign n2574 = G46 & n1752 ;
  assign n2575 = ~G176 & n2188 ;
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  assign n2576 = G176 & n493 ;
  assign n2577 = G177 & ~n2576 ;
  assign n2578 = ~n2575 & n2577 ;
  assign n2579 = n2574 | n2578 ;
  buffer buf_n2580( .i (n2579), .o (n2580) );
  buffer buf_n2581( .i (n2580), .o (n2581) );
  buffer buf_n2582( .i (n2581), .o (n2582) );
  buffer buf_n2583( .i (n2582), .o (n2583) );
  buffer buf_n2584( .i (n2583), .o (n2584) );
  inverter inv_n2585( .i (n2584), .o (n2585) );
  buffer buf_n2586( .i (n1749), .o (n2586) );
  assign n2587 = G45 & n2586 ;
  assign n2588 = ~G176 & n2214 ;
  assign n2589 = G176 & n429 ;
  assign n2590 = G177 & ~n2589 ;
  assign n2591 = ~n2588 & n2590 ;
  assign n2592 = n2587 | n2591 ;
  buffer buf_n2593( .i (n2592), .o (n2593) );
  buffer buf_n2594( .i (n2593), .o (n2594) );
  buffer buf_n2595( .i (n2594), .o (n2595) );
  buffer buf_n2596( .i (n2595), .o (n2596) );
  buffer buf_n2597( .i (n2596), .o (n2597) );
  buffer buf_n2598( .i (n2597), .o (n2598) );
  buffer buf_n2599( .i (n2598), .o (n2599) );
  inverter inv_n2600( .i (n2599), .o (n2600) );
  assign n2601 = G20 & n2586 ;
  assign n2602 = G176 | n2228 ;
  assign n2603 = G176 & n440 ;
  assign n2604 = G177 & ~n2603 ;
  assign n2605 = n2602 & n2604 ;
  assign n2606 = n2601 | n2605 ;
  buffer buf_n2607( .i (n2606), .o (n2607) );
  buffer buf_n2608( .i (n2607), .o (n2608) );
  buffer buf_n2609( .i (n2608), .o (n2609) );
  buffer buf_n2610( .i (n2609), .o (n2610) );
  buffer buf_n2611( .i (n2610), .o (n2611) );
  buffer buf_n2612( .i (n2611), .o (n2612) );
  buffer buf_n2613( .i (n2612), .o (n2613) );
  inverter inv_n2614( .i (n2613), .o (n2614) );
  assign n2615 = G44 & n2586 ;
  assign n2616 = G176 | n2196 ;
  assign n2617 = G176 & n417 ;
  assign n2618 = G177 & ~n2617 ;
  assign n2619 = n2616 & n2618 ;
  assign n2620 = n2615 | n2619 ;
  buffer buf_n2621( .i (n2620), .o (n2621) );
  buffer buf_n2622( .i (n2621), .o (n2622) );
  buffer buf_n2623( .i (n2622), .o (n2623) );
  buffer buf_n2624( .i (n2623), .o (n2624) );
  buffer buf_n2625( .i (n2624), .o (n2625) );
  buffer buf_n2626( .i (n2625), .o (n2626) );
  buffer buf_n2627( .i (n2626), .o (n2627) );
  inverter inv_n2628( .i (n2627), .o (n2628) );
  assign n2629 = G174 | n2581 ;
  assign n2630 = G174 & ~n2519 ;
  assign n2631 = G175 & ~n2630 ;
  assign n2632 = n2629 & n2631 ;
  assign n2633 = G41 & ~n2401 ;
  assign n2634 = G42 & n2399 ;
  assign n2635 = n2633 | n2634 ;
  assign n2636 = n2632 | n2635 ;
  buffer buf_n2637( .i (n2636), .o (n2637) );
  assign n2638 = G173 | n2581 ;
  assign n2639 = G173 & ~n2519 ;
  assign n2640 = G172 & ~n2639 ;
  assign n2641 = n2638 & n2640 ;
  assign n2642 = G41 & ~n2363 ;
  assign n2643 = G42 & n2361 ;
  assign n2644 = n2642 | n2643 ;
  assign n2645 = n2641 | n2644 ;
  buffer buf_n2646( .i (n2645), .o (n2646) );
  assign n2647 = G173 & ~n2533 ;
  assign n2648 = G173 | n2595 ;
  assign n2649 = G172 & n2648 ;
  assign n2650 = ~n2647 & n2649 ;
  assign n2651 = G17 & n2361 ;
  assign n2652 = G18 & ~n2363 ;
  assign n2653 = n2651 | n2652 ;
  assign n2654 = n2650 | n2653 ;
  buffer buf_n2655( .i (n2654), .o (n2655) );
  assign n2656 = G173 & ~n2547 ;
  assign n2657 = G173 | n2609 ;
  assign n2658 = G172 & n2657 ;
  assign n2659 = ~n2656 & n2658 ;
  assign n2660 = G39 & n2361 ;
  assign n2661 = G40 & ~n2363 ;
  assign n2662 = n2660 | n2661 ;
  assign n2663 = n2659 | n2662 ;
  buffer buf_n2664( .i (n2663), .o (n2664) );
  assign n2665 = G173 & ~n2561 ;
  assign n2666 = G173 | n2623 ;
  assign n2667 = G172 & n2666 ;
  assign n2668 = ~n2665 & n2667 ;
  buffer buf_n2669( .i (n1839), .o (n2669) );
  assign n2670 = G36 & n2669 ;
  buffer buf_n2671( .i (n1843), .o (n2671) );
  assign n2672 = G15 & ~n2671 ;
  assign n2673 = n2670 | n2672 ;
  assign n2674 = n2668 | n2673 ;
  buffer buf_n2675( .i (n2674), .o (n2675) );
  assign n2676 = G174 | n2596 ;
  assign n2677 = G174 & ~n2532 ;
  assign n2678 = G175 & ~n2677 ;
  assign n2679 = n2676 & n2678 ;
  assign n2680 = G17 & n2399 ;
  assign n2681 = G18 & ~n2401 ;
  assign n2682 = n2680 | n2681 ;
  assign n2683 = n2679 | n2682 ;
  buffer buf_n2684( .i (n2683), .o (n2684) );
  assign n2685 = G174 | n2610 ;
  assign n2686 = G174 & ~n2546 ;
  assign n2687 = G175 & ~n2686 ;
  assign n2688 = n2685 & n2687 ;
  assign n2689 = G39 & n2399 ;
  assign n2690 = G40 & ~n2401 ;
  assign n2691 = n2689 | n2690 ;
  assign n2692 = n2688 | n2691 ;
  buffer buf_n2693( .i (n2692), .o (n2693) );
  assign n2694 = G174 | n2624 ;
  assign n2695 = G174 & ~n2560 ;
  assign n2696 = G175 & ~n2695 ;
  assign n2697 = n2694 & n2696 ;
  buffer buf_n2698( .i (n1946), .o (n2698) );
  assign n2699 = G36 & n2698 ;
  buffer buf_n2700( .i (n1950), .o (n2700) );
  assign n2701 = G15 & ~n2700 ;
  assign n2702 = n2699 | n2701 ;
  assign n2703 = n2697 | n2702 ;
  buffer buf_n2704( .i (n2703), .o (n2704) );
  assign n2705 = G158 & ~n2560 ;
  assign n2706 = G158 | n2622 ;
  assign n2707 = G159 & n2706 ;
  assign n2708 = ~n2705 & n2707 ;
  assign n2709 = G77 & ~n2440 ;
  assign n2710 = G87 & n2442 ;
  assign n2711 = n2709 | n2710 ;
  assign n2712 = n2708 | n2711 ;
  assign n2713 = G64 & n2712 ;
  buffer buf_n2714( .i (n2713), .o (n2714) );
  assign n2715 = G158 & ~n2546 ;
  assign n2716 = G158 | n2608 ;
  assign n2717 = G159 & n2716 ;
  assign n2718 = ~n2715 & n2717 ;
  assign n2719 = G75 & ~n2440 ;
  assign n2720 = G85 & n2442 ;
  assign n2721 = n2719 | n2720 ;
  assign n2722 = n2718 | n2721 ;
  assign n2723 = G64 & n2722 ;
  buffer buf_n2724( .i (n2723), .o (n2724) );
  assign n2725 = G158 & ~n2532 ;
  assign n2726 = G158 | n2594 ;
  assign n2727 = G159 & n2726 ;
  assign n2728 = ~n2725 & n2727 ;
  assign n2729 = G84 & n2442 ;
  assign n2730 = G74 & ~n2440 ;
  assign n2731 = n2729 | n2730 ;
  assign n2732 = n2728 | n2731 ;
  assign n2733 = G64 & n2732 ;
  buffer buf_n2734( .i (n2733), .o (n2734) );
  assign n2735 = G158 | n2580 ;
  assign n2736 = G158 & ~n2518 ;
  assign n2737 = G159 & ~n2736 ;
  assign n2738 = n2735 & n2737 ;
  buffer buf_n2739( .i (n2303), .o (n2739) );
  assign n2740 = G73 & ~n2739 ;
  buffer buf_n2741( .i (n2307), .o (n2741) );
  assign n2742 = G83 & n2741 ;
  assign n2743 = n2740 | n2742 ;
  assign n2744 = n2738 | n2743 ;
  assign n2745 = G64 & n2744 ;
  buffer buf_n2746( .i (n2745), .o (n2746) );
  assign n2747 = G160 | n2623 ;
  assign n2748 = G160 & ~n2559 ;
  assign n2749 = G161 & ~n2748 ;
  assign n2750 = n2747 & n2749 ;
  assign n2751 = G77 & ~n2482 ;
  assign n2752 = G87 & n2484 ;
  assign n2753 = n2751 | n2752 ;
  assign n2754 = n2750 | n2753 ;
  assign n2755 = G64 & n2754 ;
  buffer buf_n2756( .i (n2755), .o (n2756) );
  assign n2757 = G160 | n2609 ;
  assign n2758 = G160 & ~n2545 ;
  assign n2759 = G161 & ~n2758 ;
  assign n2760 = n2757 & n2759 ;
  assign n2761 = G85 & n2484 ;
  assign n2762 = G75 & ~n2482 ;
  assign n2763 = n2761 | n2762 ;
  assign n2764 = n2760 | n2763 ;
  assign n2765 = G64 & n2764 ;
  buffer buf_n2766( .i (n2765), .o (n2766) );
  assign n2767 = G160 & ~n2532 ;
  assign n2768 = G160 | n2594 ;
  assign n2769 = G161 & n2768 ;
  assign n2770 = ~n2767 & n2769 ;
  assign n2771 = G74 & ~n2482 ;
  assign n2772 = G84 & n2484 ;
  assign n2773 = n2771 | n2772 ;
  assign n2774 = n2770 | n2773 ;
  assign n2775 = G64 & n2774 ;
  buffer buf_n2776( .i (n2775), .o (n2776) );
  assign n2777 = G160 | n2580 ;
  assign n2778 = G160 & ~n2518 ;
  assign n2779 = G161 & ~n2778 ;
  assign n2780 = n2777 & n2779 ;
  buffer buf_n2781( .i (n2319), .o (n2781) );
  assign n2782 = G73 & ~n2781 ;
  buffer buf_n2783( .i (n2323), .o (n2783) );
  assign n2784 = G83 & n2783 ;
  assign n2785 = n2782 | n2784 ;
  assign n2786 = n2780 | n2785 ;
  assign n2787 = G64 & n2786 ;
  buffer buf_n2788( .i (n2787), .o (n2788) );
  assign n2789 = ~G145 & n1389 ;
  buffer buf_n2790( .i (n2789), .o (n2790) );
  buffer buf_n2791( .i (n2790), .o (n2791) );
  assign n2792 = n1433 & ~n2791 ;
  assign n2793 = G145 & ~n1440 ;
  assign n2794 = n2790 | n2793 ;
  assign n2795 = n1391 & ~n1448 ;
  assign n2796 = n2794 & ~n2795 ;
  assign n2797 = n2792 | n2796 ;
  buffer buf_n2798( .i (n2797), .o (n2798) );
  assign n2799 = n2085 & n2798 ;
  assign n2800 = n2085 | n2798 ;
  assign n2801 = ~n2799 & n2800 ;
  assign n2802 = n2244 & ~n2801 ;
  assign n2803 = ~n1394 & n1433 ;
  assign n2804 = n1401 & ~n2803 ;
  buffer buf_n2805( .i (n2804), .o (n2805) );
  assign n2806 = ~n1442 & n1468 ;
  buffer buf_n2807( .i (n1467), .o (n2807) );
  assign n2808 = n1442 & ~n2807 ;
  assign n2809 = n2806 | n2808 ;
  buffer buf_n2810( .i (n2809), .o (n2810) );
  assign n2811 = n2805 & n2810 ;
  assign n2812 = n2805 | n2810 ;
  assign n2813 = ~n2811 & n2812 ;
  assign n2814 = n2244 | n2813 ;
  assign n2815 = ~n2802 & n2814 ;
  buffer buf_n2816( .i (n2815), .o (n2816) );
  buffer buf_n2817( .i (n2816), .o (n2817) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  assign n2818 = n1198 & ~n1891 ;
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  assign n2819 = ~n1208 & n1891 ;
  assign n2820 = n2818 | n2819 ;
  buffer buf_n2821( .i (n2820), .o (n2821) );
  assign n2822 = G162 & n1267 ;
  assign n2823 = n1248 & n2822 ;
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  assign n2824 = G162 | n1247 ;
  assign n2825 = n1305 & n2824 ;
  assign n2826 = ~n2823 & n2825 ;
  buffer buf_n2827( .i (n2826), .o (n2827) );
  assign n2828 = ~n1210 & n1543 ;
  assign n2829 = n1210 & ~n1543 ;
  assign n2830 = n2828 | n2829 ;
  buffer buf_n2831( .i (n2830), .o (n2831) );
  assign n2832 = n2827 & n2831 ;
  assign n2833 = n2827 | n2831 ;
  assign n2834 = ~n2832 & n2833 ;
  buffer buf_n2835( .i (n2834), .o (n2835) );
  assign n2836 = ~n1358 & n2835 ;
  assign n2837 = n1358 & ~n2835 ;
  assign n2838 = n2836 | n2837 ;
  buffer buf_n2839( .i (n2838), .o (n2839) );
  assign n2840 = n2821 & ~n2839 ;
  assign n2841 = ~n2821 & n2839 ;
  assign n2842 = n2840 | n2841 ;
  buffer buf_n2843( .i (n2842), .o (n2843) );
  buffer buf_n2844( .i (n2843), .o (n2844) );
  assign n2845 = n2817 | n2844 ;
  assign n2846 = n2816 & n2843 ;
  assign n2847 = G176 | n2846 ;
  assign n2848 = n2845 & ~n2847 ;
  assign n2849 = ~G148 & G98 ;
  assign n2850 = ~G100 & G148 ;
  assign n2851 = n2849 | n2850 ;
  buffer buf_n2852( .i (n2851), .o (n2852) );
  assign n2853 = ~n357 & n2852 ;
  assign n2854 = n357 & ~n2852 ;
  assign n2855 = n2853 | n2854 ;
  buffer buf_n2856( .i (n2855), .o (n2856) );
  assign n2857 = G100 | G121 ;
  assign n2858 = ~G101 & G121 ;
  assign n2859 = n2857 & ~n2858 ;
  assign n2860 = G147 & ~n2859 ;
  assign n2861 = G102 & G121 ;
  assign n2862 = ~G121 & G98 ;
  assign n2863 = n2861 | n2862 ;
  assign n2864 = ~G147 & n2863 ;
  assign n2865 = n2860 | n2864 ;
  buffer buf_n2866( .i (n2865), .o (n2866) );
  assign n2867 = n2856 | n2866 ;
  assign n2868 = n2856 & n2866 ;
  assign n2869 = n2867 & ~n2868 ;
  buffer buf_n2870( .i (n2869), .o (n2870) );
  assign n2871 = G100 | G128 ;
  assign n2872 = ~G101 & G128 ;
  assign n2873 = n2871 & ~n2872 ;
  assign n2874 = G150 & ~n2873 ;
  assign n2875 = G102 & G128 ;
  assign n2876 = ~G128 & G98 ;
  assign n2877 = n2875 | n2876 ;
  assign n2878 = ~G150 & n2877 ;
  assign n2879 = n2874 | n2878 ;
  buffer buf_n2880( .i (n2879), .o (n2880) );
  assign n2881 = G100 | G126 ;
  assign n2882 = ~G101 & G126 ;
  assign n2883 = n2881 & ~n2882 ;
  assign n2884 = G149 & ~n2883 ;
  assign n2885 = G102 & G126 ;
  assign n2886 = ~G126 & G98 ;
  assign n2887 = n2885 | n2886 ;
  assign n2888 = ~G149 & n2887 ;
  assign n2889 = n2884 | n2888 ;
  buffer buf_n2890( .i (n2889), .o (n2890) );
  assign n2891 = n2880 | n2890 ;
  assign n2892 = n2880 & n2890 ;
  assign n2893 = n2891 & ~n2892 ;
  buffer buf_n2894( .i (n2893), .o (n2894) );
  assign n2895 = n2870 | n2894 ;
  assign n2896 = n2870 & n2894 ;
  assign n2897 = n2895 & ~n2896 ;
  buffer buf_n2898( .i (n2897), .o (n2898) );
  buffer buf_n2899( .i (n2898), .o (n2899) );
  assign n2900 = n261 | n280 ;
  assign n2901 = ~n290 & n2900 ;
  buffer buf_n2902( .i (n2901), .o (n2902) );
  assign n2903 = ~n316 & n335 ;
  assign n2904 = n346 | n2903 ;
  buffer buf_n2905( .i (n2904), .o (n2905) );
  assign n2906 = n2902 | n2905 ;
  assign n2907 = n2902 & n2905 ;
  assign n2908 = n2906 & ~n2907 ;
  buffer buf_n2909( .i (n2908), .o (n2909) );
  buffer buf_n2910( .i (n2909), .o (n2910) );
  assign n2911 = n2899 | n2910 ;
  assign n2912 = n2898 & n2909 ;
  assign n2913 = G176 & ~n2912 ;
  assign n2914 = n2911 & n2913 ;
  assign n2915 = G177 & ~n2914 ;
  assign n2916 = ~n2848 & n2915 ;
  buffer buf_n2917( .i (n2916), .o (n2917) );
  buffer buf_n2918( .i (n2917), .o (n2918) );
  buffer buf_n2919( .i (n2918), .o (n2919) );
  buffer buf_n2920( .i (n2919), .o (n2920) );
  buffer buf_n2921( .i (n2920), .o (n2921) );
  buffer buf_n2922( .i (n2921), .o (n2922) );
  buffer buf_n2923( .i (n2922), .o (n2923) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  assign n2924 = ~G51 & n1757 ;
  assign n2925 = n2923 | n2924 ;
  inverter inv_n2926( .i (n2925), .o (n2926) );
  assign n2927 = n622 & n678 ;
  assign n2928 = n619 | n689 ;
  assign n2929 = ~n704 & n2928 ;
  buffer buf_n2930( .i (n2929), .o (n2930) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  assign n2931 = n599 | n676 ;
  assign n2932 = ~n1652 & n2931 ;
  assign n2933 = n2930 | n2932 ;
  assign n2934 = ~n2927 & n2933 ;
  buffer buf_n2935( .i (n2934), .o (n2935) );
  assign n2936 = n1662 & ~n2935 ;
  assign n2937 = ~n1662 & n2935 ;
  assign n2938 = n2936 | n2937 ;
  buffer buf_n2939( .i (n2938), .o (n2939) );
  buffer buf_n2940( .i (n2939), .o (n2940) );
  assign n2941 = n1977 | n2940 ;
  assign n2942 = n1976 & n2939 ;
  assign n2943 = G157 | n2942 ;
  assign n2944 = n2941 & ~n2943 ;
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  assign n2945 = n614 & n668 ;
  assign n2946 = n614 | n678 ;
  assign n2947 = ~n2945 & n2946 ;
  buffer buf_n2948( .i (n2947), .o (n2948) );
  assign n2949 = n2002 & ~n2948 ;
  assign n2950 = ~n2002 & n2948 ;
  assign n2951 = n2949 | n2950 ;
  buffer buf_n2952( .i (n2951), .o (n2952) );
  buffer buf_n2953( .i (n2952), .o (n2953) );
  assign n2954 = n562 | n2930 ;
  assign n2955 = n562 & n2930 ;
  assign n2956 = n2954 & ~n2955 ;
  buffer buf_n2957( .i (n2956), .o (n2957) );
  assign n2958 = n824 | n1970 ;
  buffer buf_n2959( .i (n2958), .o (n2959) );
  assign n2960 = n2957 & ~n2959 ;
  assign n2961 = ~n2957 & n2959 ;
  assign n2962 = n2960 | n2961 ;
  buffer buf_n2963( .i (n2962), .o (n2963) );
  buffer buf_n2964( .i (n2963), .o (n2964) );
  assign n2965 = n2953 & n2964 ;
  assign n2966 = n2952 | n2963 ;
  assign n2967 = G157 & n2966 ;
  assign n2968 = ~n2965 & n2967 ;
  assign n2969 = n2944 | n2968 ;
  buffer buf_n2970( .i (n2969), .o (n2970) );
  buffer buf_n2971( .i (n2970), .o (n2971) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  assign n2972 = n1142 | n1691 ;
  buffer buf_n2973( .i (n2972), .o (n2973) );
  buffer buf_n2974( .i (n2973), .o (n2974) );
  buffer buf_n2975( .i (n2974), .o (n2975) );
  buffer buf_n2976( .i (n2975), .o (n2976) );
  assign n2977 = ~n964 & n2976 ;
  assign n2978 = n983 & ~n2977 ;
  buffer buf_n2979( .i (n2978), .o (n2979) );
  assign n2980 = n910 | n1040 ;
  assign n2981 = n910 & n1040 ;
  assign n2982 = n2980 & ~n2981 ;
  buffer buf_n2983( .i (n2982), .o (n2983) );
  buffer buf_n2984( .i (n2983), .o (n2984) );
  buffer buf_n2985( .i (n2984), .o (n2985) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1689( .i (n1688), .o (n1689) );
  assign n2986 = n1090 | n2973 ;
  assign n2987 = ~n1689 & n2986 ;
  buffer buf_n2988( .i (n2987), .o (n2988) );
  assign n2989 = n2985 & n2988 ;
  assign n2990 = n2985 | n2988 ;
  assign n2991 = ~n2989 & n2990 ;
  buffer buf_n2992( .i (n2991), .o (n2992) );
  assign n2993 = n2979 & n2992 ;
  assign n2994 = n2979 | n2992 ;
  assign n2995 = ~n2993 & n2994 ;
  buffer buf_n2996( .i (n2995), .o (n2996) );
  assign n2997 = n1675 & n2996 ;
  assign n2998 = n962 | n1694 ;
  assign n2999 = ~n1707 & n2998 ;
  buffer buf_n3000( .i (n2999), .o (n3000) );
  buffer buf_n3001( .i (n3000), .o (n3001) );
  assign n3002 = ~n985 & n1107 ;
  assign n3003 = n985 & ~n1107 ;
  assign n3004 = n3002 | n3003 ;
  buffer buf_n3005( .i (n3004), .o (n3005) );
  assign n3006 = n2983 & ~n3005 ;
  assign n3007 = ~n2983 & n3005 ;
  assign n3008 = n3006 | n3007 ;
  buffer buf_n3009( .i (n3008), .o (n3009) );
  buffer buf_n3010( .i (n3009), .o (n3010) );
  assign n3011 = n3001 | n3010 ;
  assign n3012 = n3000 & n3009 ;
  assign n3013 = n1671 | n3012 ;
  assign n3014 = n3011 & ~n3013 ;
  buffer buf_n3015( .i (n3014), .o (n3015) );
  buffer buf_n3016( .i (n3015), .o (n3016) );
  assign n3017 = G157 | n3016 ;
  assign n3018 = n2997 | n3017 ;
  assign n3019 = n836 | n1674 ;
  assign n3020 = n2996 & n3019 ;
  assign n3021 = ~n836 & n3015 ;
  assign n3022 = G157 & ~n3021 ;
  assign n3023 = ~n3020 & n3022 ;
  assign n3024 = n3018 & ~n3023 ;
  buffer buf_n3025( .i (n3024), .o (n3025) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  assign n3026 = n749 | n805 ;
  assign n3027 = ~n820 & n3026 ;
  buffer buf_n3028( .i (n3027), .o (n3028) );
  assign n3029 = n3025 & ~n3028 ;
  assign n3030 = ~n3025 & n3028 ;
  assign n3031 = n3029 | n3030 ;
  buffer buf_n3032( .i (n3031), .o (n3032) );
  buffer buf_n3033( .i (n3032), .o (n3033) );
  assign n3034 = ~n2971 & n3033 ;
  assign n3035 = n2970 & ~n3032 ;
  assign n3036 = G176 | n3035 ;
  assign n3037 = n3034 | n3036 ;
  assign n3038 = G100 | G90 ;
  assign n3039 = ~G101 & G90 ;
  assign n3040 = n3038 & ~n3039 ;
  assign n3041 = G143 & ~n3040 ;
  assign n3042 = G102 & G90 ;
  assign n3043 = ~G90 & G98 ;
  assign n3044 = n3042 | n3043 ;
  assign n3045 = ~G143 & n3044 ;
  assign n3046 = n3041 | n3045 ;
  buffer buf_n3047( .i (n3046), .o (n3047) );
  assign n3048 = G100 | G92 ;
  assign n3049 = ~G101 & G92 ;
  assign n3050 = n3048 & ~n3049 ;
  assign n3051 = G144 & ~n3050 ;
  assign n3052 = G102 & G92 ;
  assign n3053 = ~G92 & G98 ;
  assign n3054 = n3052 | n3053 ;
  assign n3055 = ~G144 & n3054 ;
  assign n3056 = n3051 | n3055 ;
  buffer buf_n3057( .i (n3056), .o (n3057) );
  assign n3058 = n3047 & ~n3057 ;
  assign n3059 = ~n3047 & n3057 ;
  assign n3060 = n3058 | n3059 ;
  buffer buf_n3061( .i (n3060), .o (n3061) );
  assign n3062 = G100 | G94 ;
  assign n3063 = ~G101 & G94 ;
  assign n3064 = n3062 & ~n3063 ;
  assign n3065 = G140 & ~n3064 ;
  assign n3066 = G102 & G94 ;
  assign n3067 = ~G94 & G98 ;
  assign n3068 = n3066 | n3067 ;
  assign n3069 = ~G140 & n3068 ;
  assign n3070 = n3065 | n3069 ;
  buffer buf_n3071( .i (n3070), .o (n3071) );
  assign n3072 = n484 & n3071 ;
  assign n3073 = n484 | n3071 ;
  assign n3074 = ~n3072 & n3073 ;
  buffer buf_n3075( .i (n3074), .o (n3075) );
  assign n3076 = ~n3061 & n3075 ;
  assign n3077 = n3061 & ~n3075 ;
  assign n3078 = n3076 | n3077 ;
  buffer buf_n3079( .i (n3078), .o (n3079) );
  buffer buf_n3080( .i (n3079), .o (n3080) );
  assign n3081 = G100 | G107 ;
  assign n3082 = ~G101 & G107 ;
  assign n3083 = n3081 & ~n3082 ;
  assign n3084 = G139 & ~n3083 ;
  assign n3085 = G102 & G107 ;
  assign n3086 = ~G107 & G98 ;
  assign n3087 = n3085 | n3086 ;
  assign n3088 = ~G139 & n3087 ;
  assign n3089 = n3084 | n3088 ;
  buffer buf_n3090( .i (n3089), .o (n3090) );
  assign n3091 = G100 | G105 ;
  assign n3092 = ~G101 & G105 ;
  assign n3093 = n3091 & ~n3092 ;
  assign n3094 = G138 & ~n3093 ;
  assign n3095 = G102 & G105 ;
  assign n3096 = ~G105 & G98 ;
  assign n3097 = n3095 | n3096 ;
  assign n3098 = ~G138 & n3097 ;
  assign n3099 = n3094 | n3098 ;
  buffer buf_n3100( .i (n3099), .o (n3100) );
  assign n3101 = n3090 & n3100 ;
  assign n3102 = n3090 | n3100 ;
  assign n3103 = ~n3101 & n3102 ;
  buffer buf_n3104( .i (n3103), .o (n3104) );
  assign n3105 = G100 | G96 ;
  assign n3106 = ~G101 & G96 ;
  assign n3107 = n3105 & ~n3106 ;
  assign n3108 = G141 & ~n3107 ;
  assign n3109 = G102 & G96 ;
  assign n3110 = ~G96 & G98 ;
  assign n3111 = n3109 | n3110 ;
  assign n3112 = ~G141 & n3111 ;
  assign n3113 = n3108 | n3112 ;
  buffer buf_n3114( .i (n3113), .o (n3114) );
  assign n3115 = G100 | G109 ;
  assign n3116 = ~G101 & G109 ;
  assign n3117 = n3115 & ~n3116 ;
  assign n3118 = G135 & ~n3117 ;
  assign n3119 = G102 & G109 ;
  assign n3120 = ~G109 & G98 ;
  assign n3121 = n3119 | n3120 ;
  assign n3122 = ~G135 & n3121 ;
  assign n3123 = n3118 | n3122 ;
  buffer buf_n3124( .i (n3123), .o (n3124) );
  assign n3125 = G100 | G103 ;
  assign n3126 = ~G101 & G103 ;
  assign n3127 = n3125 & ~n3126 ;
  assign n3128 = G137 & ~n3127 ;
  assign n3129 = G102 & G103 ;
  assign n3130 = ~G103 & G98 ;
  assign n3131 = n3129 | n3130 ;
  assign n3132 = ~G137 & n3131 ;
  assign n3133 = n3128 | n3132 ;
  buffer buf_n3134( .i (n3133), .o (n3134) );
  assign n3135 = n3124 & n3134 ;
  assign n3136 = n3124 | n3134 ;
  assign n3137 = ~n3135 & n3136 ;
  buffer buf_n3138( .i (n3137), .o (n3138) );
  assign n3139 = n3114 & ~n3138 ;
  assign n3140 = ~n3114 & n3138 ;
  assign n3141 = n3139 | n3140 ;
  buffer buf_n3142( .i (n3141), .o (n3142) );
  assign n3143 = ~n3104 & n3142 ;
  assign n3144 = n3104 & ~n3142 ;
  assign n3145 = n3143 | n3144 ;
  buffer buf_n3146( .i (n3145), .o (n3146) );
  buffer buf_n3147( .i (n3146), .o (n3147) );
  assign n3148 = ~n3080 & n3147 ;
  assign n3149 = n3079 & ~n3146 ;
  assign n3150 = G176 & ~n3149 ;
  assign n3151 = ~n3148 & n3150 ;
  assign n3152 = G177 & ~n3151 ;
  assign n3153 = n3037 & n3152 ;
  buffer buf_n3154( .i (n3153), .o (n3154) );
  buffer buf_n3155( .i (n3154), .o (n3155) );
  buffer buf_n3156( .i (n3155), .o (n3156) );
  buffer buf_n3157( .i (n3156), .o (n3157) );
  buffer buf_n3158( .i (n3157), .o (n3158) );
  buffer buf_n3159( .i (n3158), .o (n3159) );
  assign n3160 = ~G49 & n1757 ;
  assign n3161 = n3159 | n3160 ;
  inverter inv_n3162( .i (n3161), .o (n3162) );
  assign n3163 = ~G177 & G38 ;
  assign n3164 = n3154 | n3163 ;
  buffer buf_n3165( .i (n3164), .o (n3165) );
  buffer buf_n3166( .i (n3165), .o (n3166) );
  assign n3167 = G173 | n3166 ;
  assign n3168 = ~G177 & G37 ;
  assign n3169 = n2917 | n3168 ;
  buffer buf_n3170( .i (n3169), .o (n3170) );
  buffer buf_n3171( .i (n3170), .o (n3171) );
  assign n3172 = G173 & ~n3171 ;
  assign n3173 = G172 & ~n3172 ;
  assign n3174 = n3167 & n3173 ;
  assign n3175 = G23 & ~n2671 ;
  assign n3176 = G4 & n2669 ;
  assign n3177 = n3175 | n3176 ;
  assign n3178 = n3174 | n3177 ;
  buffer buf_n3179( .i (n3178), .o (n3179) );
  assign n3180 = G174 | n3166 ;
  assign n3181 = G174 & ~n3171 ;
  assign n3182 = G175 & ~n3181 ;
  assign n3183 = n3180 & n3182 ;
  assign n3184 = G23 & ~n2700 ;
  assign n3185 = G4 & n2698 ;
  assign n3186 = n3184 | n3185 ;
  assign n3187 = n3183 | n3186 ;
  buffer buf_n3188( .i (n3187), .o (n3188) );
  assign n3189 = G158 | n3165 ;
  assign n3190 = G158 & ~n3170 ;
  assign n3191 = G159 & ~n3190 ;
  assign n3192 = n3189 & n3191 ;
  assign n3193 = G79 & ~n2739 ;
  assign n3194 = G78 & n2741 ;
  assign n3195 = n3193 | n3194 ;
  assign n3196 = n3192 | n3195 ;
  assign n3197 = G64 & n3196 ;
  inverter inv_n3198( .i (n3197), .o (n3198) );
  assign n3199 = G160 | n3165 ;
  assign n3200 = G160 & ~n3170 ;
  assign n3201 = G161 & ~n3200 ;
  assign n3202 = n3199 & n3201 ;
  assign n3203 = G79 & ~n2781 ;
  assign n3204 = G78 & n2783 ;
  assign n3205 = n3203 | n3204 ;
  assign n3206 = n3202 | n3205 ;
  assign n3207 = G64 & n3206 ;
  inverter inv_n3208( .i (n3207), .o (n3208) );
  assign G5193 = ~G66 ;
  assign G5194 = ~G113 ;
  assign G5195 = ~G165 ;
  assign G5196 = ~G151 ;
  assign G5197 = ~G127 ;
  assign G5198 = ~G131 ;
  assign G5199 = n186 ;
  assign G5200 = ~G152 ;
  assign G5201 = ~G151 ;
  assign G5202 = ~G151 ;
  assign G5203 = ~G125 ;
  assign G5204 = ~G129 ;
  assign G5205 = n188 ;
  assign G5206 = ~G99 ;
  assign G5207 = ~G153 ;
  assign G5208 = ~G156 ;
  assign G5209 = ~G155 ;
  assign G5210 = n190 ;
  assign G5211 = n192 ;
  assign G5212 = n194 ;
  assign G5213 = n203 ;
  assign G5214 = G64 ;
  assign G5215 = G66 ;
  assign G5216 = G1 ;
  assign G5217 = G152 ;
  assign G5218 = G114 ;
  assign G5219 = G152 ;
  assign G5220 = n212 ;
  assign G5221 = n210 ;
  assign G5222 = ~G1 ;
  assign G5223 = ~G1 ;
  assign G5224 = ~G1 ;
  assign G5225 = ~G1 ;
  assign G5226 = ~G114 ;
  assign G5227 = ~G114 ;
  assign G5228 = n217 ;
  assign G5229 = n223 ;
  assign G5230 = n223 ;
  assign G5231 = n225 ;
  assign G5232 = n231 ;
  assign G5233 = n237 ;
  assign G5234 = n243 ;
  assign G5235 = n250 ;
  assign G5236 = n407 ;
  assign G5237 = n526 ;
  assign G5238 = n1172 ;
  assign G5239 = n1568 ;
  assign G5240 = n1568 ;
  assign G5241 = n1172 ;
  assign G5242 = n1605 ;
  assign G5243 = n1645 ;
  assign G5244 = n1733 ;
  assign G5245 = n1747 ;
  assign G5246 = n1733 ;
  assign G5247 = n1747 ;
  assign G5248 = n1774 ;
  assign G5249 = n1794 ;
  assign G5250 = n1820 ;
  assign G5251 = n1833 ;
  assign G5252 = n1848 ;
  assign G5253 = n1888 ;
  assign G5254 = n1918 ;
  assign G5255 = n1940 ;
  assign G5256 = n1955 ;
  assign G5257 = n1998 ;
  assign G5258 = n2028 ;
  assign G5259 = n2063 ;
  assign G5260 = n2081 ;
  assign G5261 = n2133 ;
  assign G5262 = n2175 ;
  assign G5263 = n2239 ;
  assign G5264 = n2297 ;
  assign G5265 = n2313 ;
  assign G5266 = n2329 ;
  assign G5267 = n2338 ;
  assign G5268 = n2347 ;
  assign G5269 = n2356 ;
  assign G5270 = n2367 ;
  assign G5271 = n2376 ;
  assign G5272 = n2385 ;
  assign G5273 = n2394 ;
  assign G5274 = n2405 ;
  assign G5275 = n2415 ;
  assign G5276 = n2425 ;
  assign G5277 = n2435 ;
  assign G5278 = n2447 ;
  assign G5279 = n2457 ;
  assign G5280 = n2467 ;
  assign G5281 = n2477 ;
  assign G5282 = n2489 ;
  assign G5283 = n2507 ;
  assign G5284 = n2511 ;
  assign G5285 = n2524 ;
  assign G5286 = n2537 ;
  assign G5287 = n2551 ;
  assign G5288 = n2565 ;
  assign G5289 = n2573 ;
  assign G5290 = n2585 ;
  assign G5291 = n2600 ;
  assign G5292 = n2614 ;
  assign G5293 = n2628 ;
  assign G5294 = n2637 ;
  assign G5295 = n2646 ;
  assign G5296 = n2655 ;
  assign G5297 = n2664 ;
  assign G5298 = n2675 ;
  assign G5299 = n2684 ;
  assign G5300 = n2693 ;
  assign G5301 = n2704 ;
  assign G5302 = n2714 ;
  assign G5303 = n2724 ;
  assign G5304 = n2734 ;
  assign G5305 = n2746 ;
  assign G5306 = n2756 ;
  assign G5307 = n2766 ;
  assign G5308 = n2776 ;
  assign G5309 = n2788 ;
  assign G5310 = n2926 ;
  assign G5311 = n3162 ;
  assign G5312 = n3179 ;
  assign G5313 = n3188 ;
  assign G5314 = n3198 ;
  assign G5315 = n3208 ;
endmodule
