module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 , y1 , y2 , y3 , y4 , y5 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 , y1 , y2 , y3 , y4 , y5 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n51 , n52 , n53 , n54 , n55 , n56 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 ;
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n13( .i (x1), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n51( .i (x5), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n58( .i (x6), .o (n58) );
  buffer buf_n66( .i (x7), .o (n66) );
  assign n83 = n58 & n66 ;
  buffer buf_n84( .i (n83), .o (n84) );
  assign n91 = n53 & ~n84 ;
  buffer buf_n92( .i (n91), .o (n92) );
  assign n95 = n17 & ~n92 ;
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n39( .i (x4), .o (n39) );
  assign n98 = n39 & n51 ;
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n22( .i (x2), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n30( .i (x3), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  assign n106 = n23 & n31 ;
  buffer buf_n107( .i (n106), .o (n107) );
  assign n111 = n100 & n107 ;
  buffer buf_n112( .i (n111), .o (n112) );
  assign n113 = n7 | n112 ;
  assign n114 = ( n8 & n96 ) | ( n8 & n113 ) | ( n96 & n113 ) ;
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  assign n121 = n14 & ~n23 ;
  buffer buf_n122( .i (n121), .o (n122) );
  assign n127 = n3 & n23 ;
  buffer buf_n128( .i (n127), .o (n128) );
  assign n131 = n122 | n128 ;
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n32( .i (n31), .o (n32) );
  assign n134 = n32 & n53 ;
  buffer buf_n135( .i (n134), .o (n135) );
  assign n138 = ~n4 & n15 ;
  buffer buf_n139( .i (n138), .o (n139) );
  assign n140 = ~n135 & n139 ;
  assign n141 = n132 | n140 ;
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n59( .i (n58), .o (n59) );
  assign n143 = n40 & n59 ;
  buffer buf_n144( .i (n143), .o (n144) );
  assign n148 = n69 & n144 ;
  assign n149 = n139 & ~n148 ;
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  assign n152 = n142 | n151 ;
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  assign n153 = n5 | n25 ;
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  assign n156 = n18 | n102 ;
  assign n157 = n155 & n156 ;
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n85( .i (n84), .o (n85) );
  assign n158 = n85 & n100 ;
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  assign n161 = n36 | n160 ;
  assign n162 = n157 | n161 ;
  assign n163 = n152 & n162 ;
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  assign n168 = ~n13 & n30 ;
  buffer buf_n169( .i (n168), .o (n169) );
  assign n171 = n22 | n39 ;
  buffer buf_n172( .i (n171), .o (n172) );
  assign n176 = n169 & ~n172 ;
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n54( .i (n53), .o (n54) );
  assign n179 = n58 | n66 ;
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  assign n184 = n54 & n181 ;
  assign n185 = n177 & ~n184 ;
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  assign n191 = ~n25 & n33 ;
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  assign n195 = n27 | n102 ;
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n19( .i (n18), .o (n19) );
  assign n197 = n19 | n193 ;
  assign n198 = ( n194 & n196 ) | ( n194 & n197 ) | ( n196 & n197 ) ;
  assign n199 = n10 & n198 ;
  buffer buf_n200( .i (n22), .o (n200) );
  assign n201 = n14 | n200 ;
  buffer buf_n202( .i (n201), .o (n202) );
  assign n207 = ~n33 & n202 ;
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  assign n211 = ~n4 & n24 ;
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n216 = n3 & ~n200 ;
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  assign n222 = n102 | n219 ;
  assign n223 = n214 | n222 ;
  assign n224 = n210 & ~n223 ;
  buffer buf_n225( .i (n224), .o (n225) );
  assign n226 = n199 | n225 ;
  assign n227 = ~n190 & n226 ;
  assign n228 = n4 & n53 ;
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n74( .i (x8), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  assign n231 = n67 & n75 ;
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  assign n236 = n230 & n234 ;
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  assign n237 = n54 | n181 ;
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n240( .i (n3), .o (n240) );
  assign n241 = n76 | n240 ;
  buffer buf_n242( .i (n241), .o (n242) );
  assign n244 = n43 & n242 ;
  assign n245 = ( n44 & n238 ) | ( n44 & n244 ) | ( n238 & n244 ) ;
  assign n246 = n236 | n245 ;
  buffer buf_n247( .i (n246), .o (n247) );
  assign n248 = n15 & ~n32 ;
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = n16 & n25 ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n253 = n250 | n252 ;
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n60( .i (n59), .o (n60) );
  assign n255 = n41 | n60 ;
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  assign n259 = ~n160 & n258 ;
  assign n260 = n254 & n259 ;
  assign n261 = n247 & n260 ;
  assign n262 = n22 & ~n30 ;
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  assign n266 = ~n144 & n264 ;
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n52), .o (n268) );
  assign n269 = n263 & ~n268 ;
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  assign n273 = n267 | n271 ;
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n170( .i (n169), .o (n170) );
  assign n276 = n144 & ~n170 ;
  buffer buf_n277( .i (n276), .o (n277) );
  assign n278 = ~n208 & n277 ;
  buffer buf_n279( .i (n278), .o (n279) );
  assign n280 = n215 & ~n279 ;
  assign n281 = ~n275 & n280 ;
  assign n282 = n261 | n281 ;
  buffer buf_n283( .i (n282), .o (n283) );
  assign n284 = n227 | n283 ;
  buffer buf_n285( .i (n284), .o (n285) );
  assign n286 = n254 | n274 ;
  assign n287 = n32 & n41 ;
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n136( .i (n135), .o (n136) );
  assign n291 = ~n136 & n252 ;
  assign n292 = ~n290 & n291 ;
  assign n293 = n24 & n41 ;
  buffer buf_n294( .i (n293), .o (n294) );
  assign n297 = n6 & ~n294 ;
  buffer buf_n298( .i (n297), .o (n298) );
  assign n299 = n159 | n230 ;
  assign n300 = n298 | n299 ;
  assign n301 = n292 | n300 ;
  assign n302 = n286 & ~n301 ;
  assign n313 = n250 & ~n257 ;
  assign n314 = n186 | n313 ;
  assign n315 = n9 & n314 ;
  buffer buf_n303( .i (n31), .o (n303) );
  buffer buf_n304( .i (n40), .o (n304) );
  assign n305 = n303 | n304 ;
  buffer buf_n306( .i (n305), .o (n306) );
  assign n309 = ~n288 & n306 ;
  buffer buf_n310( .i (n309), .o (n310) );
  assign n311 = n27 & n238 ;
  assign n312 = ~n310 & n311 ;
  assign n316 = n279 | n312 ;
  assign n317 = ( n10 & n315 ) | ( n10 & n316 ) | ( n315 & n316 ) ;
  assign n318 = n302 | n317 ;
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n320( .i (n101), .o (n320) );
  assign n321 = n192 & n320 ;
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  assign n324 = n62 | n233 ;
  buffer buf_n325( .i (n324), .o (n325) );
  assign n326 = n136 | n289 ;
  assign n327 = ( n290 & n325 ) | ( n290 & n326 ) | ( n325 & n326 ) ;
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  assign n329 = n206 & ~n322 ;
  assign n330 = ( n323 & n328 ) | ( n323 & ~n329 ) | ( n328 & ~n329 ) ;
  assign n331 = ~n11 & n330 ;
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  assign n332 = ~n14 & n200 ;
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  assign n335 = ~n78 & n334 ;
  buffer buf_n336( .i (n335), .o (n336) );
  assign n337 = n209 & ~n336 ;
  buffer buf_n338( .i (n337), .o (n338) );
  assign n339 = ~n247 & n338 ;
  buffer buf_n20( .i (n19), .o (n20) );
  assign n340 = n31 | n200 ;
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  assign n346 = ( n9 & ~n20 ) | ( n9 & n345 ) | ( ~n20 & n345 ) ;
  assign n347 = ( n20 & n196 ) | ( n20 & ~n345 ) | ( n196 & ~n345 ) ;
  assign n348 = n346 & n347 ;
  assign n349 = n339 | n348 ;
  assign n350 = n331 | n349 ;
  assign n351 = n319 | n350 ;
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  assign n353 = ~n308 & n336 ;
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  assign n358 = ~n319 & n357 ;
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n455( .i (n5), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  assign n457 = ~n183 & n456 ;
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  assign n459 = n56 & ~n307 ;
  assign n460 = ~n133 & n459 ;
  assign n461 = ~n458 & n460 ;
  buffer buf_n178( .i (n177), .o (n178) );
  assign n363 = n15 | n60 ;
  buffer buf_n364( .i (n363), .o (n364) );
  assign n462 = n242 | n364 ;
  assign n463 = n178 & ~n462 ;
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n384( .i (n13), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  assign n389 = ~n268 & n385 ;
  buffer buf_n390( .i (n389), .o (n390) );
  assign n465 = n108 & n390 ;
  buffer buf_n466( .i (n465), .o (n466) );
  assign n467 = n235 & n466 ;
  assign n468 = n464 | n467 ;
  assign n469 = n461 | n468 ;
  buffer buf_n470( .i (n52), .o (n470) );
  assign n471 = n68 & n470 ;
  buffer buf_n472( .i (n471), .o (n472) );
  assign n474 = ~n42 & n122 ;
  assign n475 = n472 & n474 ;
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n79( .i (n78), .o (n79) );
  assign n477 = ~n5 & n61 ;
  buffer buf_n478( .i (n477), .o (n478) );
  assign n479 = n34 & n78 ;
  assign n480 = ( n79 & n478 ) | ( n79 & n479 ) | ( n478 & n479 ) ;
  assign n481 = n476 & n480 ;
  buffer buf_n482( .i (n51), .o (n482) );
  assign n483 = n75 & n482 ;
  buffer buf_n484( .i (n483), .o (n484) );
  assign n486 = n16 & ~n484 ;
  buffer buf_n404( .i (n30), .o (n404) );
  assign n405 = n384 | n404 ;
  buffer buf_n406( .i (n405), .o (n406) );
  assign n487 = ~n406 & n484 ;
  assign n488 = n486 | n487 ;
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  assign n490 = ~n175 & n456 ;
  assign n491 = n489 & n490 ;
  assign n492 = n481 | n491 ;
  buffer buf_n493( .i (n492), .o (n493) );
  assign n494 = n469 | n493 ;
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n109( .i (n108), .o (n109) );
  assign n428 = ~n203 & n288 ;
  assign n429 = n109 | n428 ;
  assign n430 = n298 & n429 ;
  buffer buf_n431( .i (n430), .o (n431) );
  assign n432 = n240 & ~n268 ;
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  assign n435 = n267 & ~n434 ;
  buffer buf_n436( .i (n435), .o (n436) );
  assign n437 = n89 & n436 ;
  assign n438 = ( n90 & n431 ) | ( n90 & n437 ) | ( n431 & n437 ) ;
  buffer buf_n265( .i (n264), .o (n265) );
  assign n439 = n139 & n265 ;
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  assign n442 = n7 & n35 ;
  assign n443 = ~n18 & n56 ;
  assign n444 = ( ~n19 & n442 ) | ( ~n19 & n443 ) | ( n442 & n443 ) ;
  assign n445 = n441 | n444 ;
  assign n446 = n76 & ~n268 ;
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  assign n450 = ~n192 & n234 ;
  assign n451 = n449 | n450 ;
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  assign n452 = n64 & ~n296 ;
  assign n453 = n451 & n452 ;
  assign n454 = n445 & n453 ;
  assign n495 = n438 | n454 ;
  assign n496 = n494 | n495 ;
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n37( .i (n36), .o (n37) );
  assign n367 = n52 & n59 ;
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  assign n371 = n252 & n370 ;
  assign n372 = ~n36 & n371 ;
  assign n359 = ~n54 & n333 ;
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n365( .i (n364), .o (n365) );
  assign n366 = n230 | n365 ;
  assign n373 = ~n361 & n366 ;
  assign n374 = ( n37 & ~n372 ) | ( n37 & n373 ) | ( ~n372 & n373 ) ;
  buffer buf_n97( .i (n96), .o (n97) );
  assign n375 = ~n109 & n343 ;
  assign n376 = n8 | n375 ;
  assign n377 = n97 | n376 ;
  assign n378 = n374 & n377 ;
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  assign n379 = n76 | n303 ;
  buffer buf_n380( .i (n379), .o (n380) );
  assign n382 = ~n6 & n380 ;
  assign n383 = n238 | n382 ;
  assign n386 = n240 & n385 ;
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  assign n392 = ~n212 & n390 ;
  assign n393 = n388 | n392 ;
  assign n394 = n383 & ~n393 ;
  assign n395 = n221 | n394 ;
  assign n396 = ~n204 & n230 ;
  assign n397 = ~n27 & n63 ;
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n398( .i (n26), .o (n398) );
  assign n399 = ( n63 & n391 ) | ( n63 & ~n398 ) | ( n391 & ~n398 ) ;
  assign n400 = ( n396 & ~n397 ) | ( n396 & n399 ) | ( ~n397 & n399 ) ;
  assign n401 = n37 & n400 ;
  assign n402 = n395 & ~n401 ;
  assign n403 = n378 & n402 ;
  assign n497 = n49 & n403 ;
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  assign n410 = ~n6 & n86 ;
  buffer buf_n411( .i (n410), .o (n411) );
  assign n412 = n370 & ~n408 ;
  assign n413 = ( ~n409 & n411 ) | ( ~n409 & n412 ) | ( n411 & n412 ) ;
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  assign n416 = n33 & n368 ;
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  assign n419 = n7 & ~n87 ;
  assign n420 = n418 | n419 ;
  assign n421 = n126 & n420 ;
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n422( .i (n229), .o (n422) );
  assign n423 = n391 | n422 ;
  assign n424 = n110 & n423 ;
  assign n425 = n187 | n424 ;
  assign n426 = n421 | n425 ;
  assign n427 = n415 | n426 ;
  assign n498 = n49 | n427 ;
  assign n499 = ( n496 & ~n497 ) | ( n496 & n498 ) | ( ~n497 & n498 ) ;
  assign n500 = n358 | n499 ;
  assign n539 = n20 | n464 ;
  buffer buf_n540( .i (n539), .o (n540) );
  assign n541 = n86 & n447 ;
  buffer buf_n542( .i (n541), .o (n542) );
  assign n543 = n310 & n542 ;
  buffer buf_n544( .i (n543), .o (n544) );
  assign n545 = ~n304 & n470 ;
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  assign n549 = n88 & n548 ;
  assign n550 = n215 & ~n549 ;
  assign n551 = ~n544 & n550 ;
  assign n552 = n540 & ~n551 ;
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n556( .i (n303), .o (n556) );
  buffer buf_n561( .i (n470), .o (n561) );
  assign n562 = n556 & ~n561 ;
  buffer buf_n563( .i (n562), .o (n563) );
  assign n564 = n473 | n563 ;
  assign n565 = n220 & n564 ;
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  assign n553 = n72 & n310 ;
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  assign n554 = ~n147 & n258 ;
  assign n555 = ~n553 & n554 ;
  assign n568 = n82 & n555 ;
  assign n557 = n69 & n556 ;
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  assign n560 = n147 & ~n559 ;
  assign n569 = ~n81 & n560 ;
  buffer buf_n570( .i (n569), .o (n570) );
  assign n571 = ( n567 & n568 ) | ( n567 & n570 ) | ( n568 & n570 ) ;
  assign n572 = n552 | n571 ;
  assign n577 = n71 | n257 ;
  assign n581 = n150 & n577 ;
  assign n573 = ~n181 & n217 ;
  buffer buf_n574( .i (n573), .o (n574) );
  assign n575 = n43 & n387 ;
  assign n576 = ( n388 & n574 ) | ( n388 & n575 ) | ( n574 & n575 ) ;
  assign n578 = n249 & n369 ;
  assign n579 = ~n265 & n390 ;
  assign n580 = n578 | n579 ;
  assign n582 = n576 | n580 ;
  assign n583 = n581 | n582 ;
  assign n584 = n108 | n212 ;
  buffer buf_n585( .i (n584), .o (n585) );
  assign n586 = n258 & n585 ;
  assign n525 = n39 | n51 ;
  buffer buf_n526( .i (n525), .o (n526) );
  assign n528 = ~n99 & n526 ;
  buffer buf_n529( .i (n528), .o (n529) );
  assign n531 = ~n455 & n529 ;
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n587( .i (n86), .o (n587) );
  assign n588 = ~n381 & n587 ;
  assign n589 = n532 & n588 ;
  assign n590 = n586 | n589 ;
  assign n591 = n583 & ~n590 ;
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  assign n521 = n108 | n270 ;
  buffer buf_n522( .i (n521), .o (n522) );
  assign n533 = n522 | n532 ;
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  assign n501 = n63 | n343 ;
  assign n502 = n71 & ~n154 ;
  assign n503 = ( n72 & ~n501 ) | ( n72 & n502 ) | ( ~n501 & n502 ) ;
  buffer buf_n504( .i (n62), .o (n504) );
  assign n505 = n192 & n504 ;
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  assign n506 = n87 & n130 ;
  assign n507 = n505 | n506 ;
  assign n508 = n503 | n507 ;
  assign n536 = n105 & n508 ;
  assign n509 = ~n145 & n433 ;
  buffer buf_n510( .i (n509), .o (n510) );
  assign n511 = n44 | n87 ;
  assign n512 = n510 & n511 ;
  assign n513 = n59 & ~n404 ;
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  assign n518 = ( n44 & ~n398 ) | ( n44 & n456 ) | ( ~n398 & n456 ) ;
  assign n519 = n517 | n518 ;
  assign n520 = ~n512 & n519 ;
  assign n537 = n520 | n534 ;
  assign n538 = ( n535 & ~n536 ) | ( n535 & n537 ) | ( ~n536 & n537 ) ;
  assign n594 = n538 | n592 ;
  assign n595 = ( ~n572 & n593 ) | ( ~n572 & n594 ) | ( n593 & n594 ) ;
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  assign n596 = n94 | n542 ;
  assign n597 = n16 & ~n341 ;
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n240), .o (n600) );
  buffer buf_n601( .i (n385), .o (n601) );
  assign n602 = n600 | n601 ;
  buffer buf_n603( .i (n602), .o (n603) );
  assign n604 = n109 & ~n603 ;
  assign n605 = n599 | n604 ;
  assign n606 = n596 & n605 ;
  buffer buf_n607( .i (n180), .o (n607) );
  assign n608 = n77 | n607 ;
  buffer buf_n609( .i (n608), .o (n609) );
  assign n610 = n112 & n609 ;
  assign n611 = ~n96 & n610 ;
  assign n612 = ~n325 & n476 ;
  assign n613 = n611 | n612 ;
  assign n614 = n606 | n613 ;
  assign n615 = ~n69 & n514 ;
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n530( .i (n529), .o (n530) );
  assign n618 = n204 | n530 ;
  assign n619 = n617 & ~n618 ;
  assign n620 = n130 & n417 ;
  assign n621 = n277 & n360 ;
  assign n622 = n620 | n621 ;
  assign n623 = n619 | n622 ;
  assign n624 = n547 & n574 ;
  assign n625 = ~n489 & n624 ;
  assign n626 = n67 | n75 ;
  buffer buf_n627( .i (n626), .o (n627) );
  assign n629 = ~n232 & n627 ;
  buffer buf_n630( .i (n629), .o (n630) );
  assign n631 = n146 | n630 ;
  assign n632 = n422 & n598 ;
  assign n633 = n631 & n632 ;
  assign n634 = n625 | n633 ;
  assign n635 = n623 | n634 ;
  assign n636 = n614 | n635 ;
  buffer buf_n239( .i (n238), .o (n239) );
  assign n637 = n18 & n381 ;
  assign n638 = n239 | n637 ;
  assign n639 = n55 | n387 ;
  assign n640 = n234 & n639 ;
  buffer buf_n243( .i (n242), .o (n243) );
  assign n641 = ~n243 & n558 ;
  assign n642 = n640 | n641 ;
  assign n643 = n638 & ~n642 ;
  assign n644 = ~n64 & n585 ;
  assign n645 = n142 & n644 ;
  assign n646 = ~n643 & n645 ;
  assign n647 = n290 & n510 ;
  assign n648 = n182 & ~n455 ;
  buffer buf_n649( .i (n648), .o (n649) );
  assign n650 = ~n295 & n563 ;
  assign n651 = n649 & n650 ;
  assign n652 = n647 | n651 ;
  buffer buf_n28( .i (n27), .o (n28) );
  assign n658 = n28 | n258 ;
  buffer buf_n628( .i (n627), .o (n628) );
  assign n653 = n62 & n628 ;
  buffer buf_n654( .i (n653), .o (n654) );
  assign n659 = n28 & n654 ;
  assign n660 = ( n20 & n658 ) | ( n20 & n659 ) | ( n658 & n659 ) ;
  assign n661 = n652 & n660 ;
  assign n662 = n646 | n661 ;
  assign n663 = n636 | n662 ;
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n527( .i (n526), .o (n527) );
  assign n664 = n264 & ~n527 ;
  buffer buf_n665( .i (n664), .o (n665) );
  assign n666 = ~n456 & n665 ;
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n362( .i (n361), .o (n362) );
  assign n669 = n362 | n667 ;
  assign n670 = ( n431 & n668 ) | ( n431 & n669 ) | ( n668 & n669 ) ;
  assign n671 = ~n657 & n670 ;
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n672( .i (n257), .o (n672) );
  assign n673 = ~n411 & n672 ;
  buffer buf_n485( .i (n484), .o (n485) );
  assign n674 = n407 & ~n485 ;
  buffer buf_n675( .i (n674), .o (n675) );
  assign n676 = n71 | n478 ;
  assign n677 = ~n675 & n676 ;
  assign n678 = n673 & n677 ;
  assign n679 = n524 & n678 ;
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n272( .i (n271), .o (n272) );
  assign n680 = n137 | n272 ;
  buffer buf_n681( .i (n107), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  assign n683 = n504 & ~n682 ;
  assign n684 = ~n603 & n630 ;
  assign n685 = ~n683 & n684 ;
  assign n686 = n680 & n685 ;
  buffer buf_n687( .i (n256), .o (n687) );
  assign n688 = ~n183 & n687 ;
  assign n689 = n466 & n688 ;
  assign n690 = ~n609 & n665 ;
  assign n691 = n17 & n546 ;
  assign n692 = n616 & n691 ;
  assign n693 = n690 | n692 ;
  assign n694 = n689 | n693 ;
  assign n695 = n686 | n694 ;
  assign n696 = n679 | n695 ;
  assign n697 = n671 | n696 ;
  assign n698 = n663 | n697 ;
  assign n699 = n595 & ~n698 ;
  assign y0 = n120 ;
  assign y1 = n167 ;
  assign y2 = n285 ;
  assign y3 = n352 ;
  assign y4 = n500 ;
  assign y5 = ~n699 ;
endmodule
