module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( in_18_ , in_1_ , in_7_ , in_109_ , in_13_ , in_106_ , in_54_ , in_118_ , in_101_ , in_3_ , in_0_ , in_113_ , in_56_ , in_30_ , in_89_ , in_35_ , in_70_ , in_38_ , in_100_ , in_105_ , in_28_ , in_10_ , in_9_ , in_78_ , in_29_ , in_60_ , in_94_ , in_108_ , in_117_ , in_103_ , in_67_ , in_44_ , in_57_ , in_76_ , in_47_ , in_20_ , in_84_ , in_17_ , in_72_ , in_116_ , in_16_ , in_120_ , in_104_ , in_64_ , in_125_ , in_58_ , in_42_ , in_40_ , in_81_ , in_115_ , in_88_ , in_24_ , in_33_ , in_123_ , in_61_ , in_79_ , in_31_ , in_36_ , in_82_ , in_111_ , in_68_ , in_2_ , in_87_ , in_74_ , in_114_ , in_53_ , in_83_ , in_86_ , in_65_ , in_102_ , in_6_ , in_75_ , in_4_ , in_93_ , in_45_ , in_90_ , in_80_ , in_73_ , in_46_ , in_25_ , in_107_ , in_37_ , in_85_ , in_49_ , in_39_ , in_63_ , in_12_ , in_112_ , in_32_ , in_119_ , in_77_ , in_34_ , in_41_ , in_122_ , in_124_ , in_48_ , in_92_ , in_15_ , in_55_ , in_50_ , in_5_ , in_127_ , in_96_ , in_22_ , in_43_ , in_52_ , in_51_ , in_21_ , in_95_ , in_59_ , in_69_ , in_121_ , in_97_ , in_11_ , in_98_ , in_126_ , in_14_ , in_91_ , in_26_ , in_99_ , in_27_ , in_71_ , in_8_ , in_23_ , in_110_ , in_62_ , in_66_ , in_19_ , out_3_ , out_2_ , out_5_ , out_1_ , out_0_ , out_7_ , out_4_ , out_6_ );
  input in_18_ , in_1_ , in_7_ , in_109_ , in_13_ , in_106_ , in_54_ , in_118_ , in_101_ , in_3_ , in_0_ , in_113_ , in_56_ , in_30_ , in_89_ , in_35_ , in_70_ , in_38_ , in_100_ , in_105_ , in_28_ , in_10_ , in_9_ , in_78_ , in_29_ , in_60_ , in_94_ , in_108_ , in_117_ , in_103_ , in_67_ , in_44_ , in_57_ , in_76_ , in_47_ , in_20_ , in_84_ , in_17_ , in_72_ , in_116_ , in_16_ , in_120_ , in_104_ , in_64_ , in_125_ , in_58_ , in_42_ , in_40_ , in_81_ , in_115_ , in_88_ , in_24_ , in_33_ , in_123_ , in_61_ , in_79_ , in_31_ , in_36_ , in_82_ , in_111_ , in_68_ , in_2_ , in_87_ , in_74_ , in_114_ , in_53_ , in_83_ , in_86_ , in_65_ , in_102_ , in_6_ , in_75_ , in_4_ , in_93_ , in_45_ , in_90_ , in_80_ , in_73_ , in_46_ , in_25_ , in_107_ , in_37_ , in_85_ , in_49_ , in_39_ , in_63_ , in_12_ , in_112_ , in_32_ , in_119_ , in_77_ , in_34_ , in_41_ , in_122_ , in_124_ , in_48_ , in_92_ , in_15_ , in_55_ , in_50_ , in_5_ , in_127_ , in_96_ , in_22_ , in_43_ , in_52_ , in_51_ , in_21_ , in_95_ , in_59_ , in_69_ , in_121_ , in_97_ , in_11_ , in_98_ , in_126_ , in_14_ , in_91_ , in_26_ , in_99_ , in_27_ , in_71_ , in_8_ , in_23_ , in_110_ , in_62_ , in_66_ , in_19_ ;
  output out_3_ , out_2_ , out_5_ , out_1_ , out_0_ , out_7_ , out_4_ , out_6_ ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 ;
  assign n129 = in_127_ & in_126_ ;
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  assign n139 = in_125_ | in_124_ ;
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  assign n147 = in_117_ | in_116_ ;
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  assign n151 = in_113_ | in_112_ ;
  buffer buf_n152( .i (n151), .o (n152) );
  assign n153 = in_115_ & in_114_ ;
  buffer buf_n154( .i (n153), .o (n154) );
  assign n155 = ( n148 & n152 ) | ( n148 & n154 ) | ( n152 & n154 ) ;
  buffer buf_n156( .i (n155), .o (n156) );
  assign n161 = ( ~n148 & n152 ) | ( ~n148 & n154 ) | ( n152 & n154 ) ;
  buffer buf_n162( .i (n161), .o (n162) );
  assign n163 = ( n150 & ~n156 ) | ( n150 & n162 ) | ( ~n156 & n162 ) ;
  buffer buf_n164( .i (n163), .o (n164) );
  assign n165 = in_123_ & in_122_ ;
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = in_118_ & in_119_ ;
  buffer buf_n170( .i (n169), .o (n170) );
  assign n171 = in_120_ | in_121_ ;
  buffer buf_n172( .i (n171), .o (n172) );
  assign n173 = ( n166 & n170 ) | ( n166 & n172 ) | ( n170 & n172 ) ;
  buffer buf_n174( .i (n173), .o (n174) );
  assign n179 = ( ~n166 & n170 ) | ( ~n166 & n172 ) | ( n170 & n172 ) ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = ( n168 & ~n174 ) | ( n168 & n180 ) | ( ~n174 & n180 ) ;
  buffer buf_n182( .i (n181), .o (n182) );
  assign n183 = ( n144 & n164 ) | ( n144 & n182 ) | ( n164 & n182 ) ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n187 = ( ~n144 & n164 ) | ( ~n144 & n182 ) | ( n164 & n182 ) ;
  buffer buf_n188( .i (n187), .o (n188) );
  assign n189 = ( n146 & ~n184 ) | ( n146 & n188 ) | ( ~n184 & n188 ) ;
  buffer buf_n190( .i (n189), .o (n190) );
  assign n191 = n138 & n190 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = n138 | n190 ;
  buffer buf_n194( .i (n193), .o (n194) );
  assign n195 = ~n192 & n194 ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n197 = in_111_ & in_110_ ;
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  assign n207 = in_109_ | in_108_ ;
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n215 = in_101_ | in_100_ ;
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  assign n219 = in_96_ | in_97_ ;
  buffer buf_n220( .i (n219), .o (n220) );
  assign n221 = in_98_ & in_99_ ;
  buffer buf_n222( .i (n221), .o (n222) );
  assign n223 = ( ~n216 & n220 ) | ( ~n216 & n222 ) | ( n220 & n222 ) ;
  buffer buf_n224( .i (n223), .o (n224) );
  assign n225 = ( n216 & n220 ) | ( n216 & n222 ) | ( n220 & n222 ) ;
  buffer buf_n226( .i (n225), .o (n226) );
  assign n231 = ( n218 & n224 ) | ( n218 & ~n226 ) | ( n224 & ~n226 ) ;
  buffer buf_n232( .i (n231), .o (n232) );
  assign n233 = in_106_ & in_107_ ;
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  assign n237 = in_103_ & in_102_ ;
  buffer buf_n238( .i (n237), .o (n238) );
  assign n239 = in_105_ | in_104_ ;
  buffer buf_n240( .i (n239), .o (n240) );
  assign n241 = ( n234 & n238 ) | ( n234 & n240 ) | ( n238 & n240 ) ;
  buffer buf_n242( .i (n241), .o (n242) );
  assign n247 = ( ~n234 & n238 ) | ( ~n234 & n240 ) | ( n238 & n240 ) ;
  buffer buf_n248( .i (n247), .o (n248) );
  assign n249 = ( n236 & ~n242 ) | ( n236 & n248 ) | ( ~n242 & n248 ) ;
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = ( n212 & n232 ) | ( n212 & n250 ) | ( n232 & n250 ) ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n255 = ( ~n212 & n232 ) | ( ~n212 & n250 ) | ( n232 & n250 ) ;
  buffer buf_n256( .i (n255), .o (n256) );
  assign n257 = ( n214 & ~n252 ) | ( n214 & n256 ) | ( ~n252 & n256 ) ;
  buffer buf_n258( .i (n257), .o (n258) );
  assign n259 = n206 & n258 ;
  buffer buf_n260( .i (n259), .o (n260) );
  assign n261 = n206 | n258 ;
  buffer buf_n262( .i (n261), .o (n262) );
  assign n263 = ~n260 & n262 ;
  buffer buf_n264( .i (n263), .o (n264) );
  assign n265 = n196 & n264 ;
  buffer buf_n266( .i (n265), .o (n266) );
  assign n270 = n196 | n264 ;
  buffer buf_n271( .i (n270), .o (n271) );
  assign n272 = ~n266 & n271 ;
  buffer buf_n273( .i (n272), .o (n273) );
  assign n274 = in_94_ & in_95_ ;
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  assign n284 = in_93_ | in_92_ ;
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  assign n292 = in_84_ | in_85_ ;
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = in_81_ | in_80_ ;
  buffer buf_n297( .i (n296), .o (n297) );
  assign n298 = in_82_ & in_83_ ;
  buffer buf_n299( .i (n298), .o (n299) );
  assign n300 = ( n293 & n297 ) | ( n293 & n299 ) | ( n297 & n299 ) ;
  buffer buf_n301( .i (n300), .o (n301) );
  assign n306 = ( ~n293 & n297 ) | ( ~n293 & n299 ) | ( n297 & n299 ) ;
  buffer buf_n307( .i (n306), .o (n307) );
  assign n308 = ( n295 & ~n301 ) | ( n295 & n307 ) | ( ~n301 & n307 ) ;
  buffer buf_n309( .i (n308), .o (n309) );
  assign n310 = in_90_ & in_91_ ;
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  assign n314 = in_87_ & in_86_ ;
  buffer buf_n315( .i (n314), .o (n315) );
  assign n316 = in_89_ | in_88_ ;
  buffer buf_n317( .i (n316), .o (n317) );
  assign n318 = ( n311 & n315 ) | ( n311 & n317 ) | ( n315 & n317 ) ;
  buffer buf_n319( .i (n318), .o (n319) );
  assign n324 = ( ~n311 & n315 ) | ( ~n311 & n317 ) | ( n315 & n317 ) ;
  buffer buf_n325( .i (n324), .o (n325) );
  assign n326 = ( n313 & ~n319 ) | ( n313 & n325 ) | ( ~n319 & n325 ) ;
  buffer buf_n327( .i (n326), .o (n327) );
  assign n328 = ( n289 & n309 ) | ( n289 & n327 ) | ( n309 & n327 ) ;
  buffer buf_n329( .i (n328), .o (n329) );
  assign n332 = ( ~n289 & n309 ) | ( ~n289 & n327 ) | ( n309 & n327 ) ;
  buffer buf_n333( .i (n332), .o (n333) );
  assign n334 = ( n291 & ~n329 ) | ( n291 & n333 ) | ( ~n329 & n333 ) ;
  buffer buf_n335( .i (n334), .o (n335) );
  assign n336 = n283 & n335 ;
  buffer buf_n337( .i (n336), .o (n337) );
  assign n338 = n283 | n335 ;
  buffer buf_n339( .i (n338), .o (n339) );
  assign n340 = ~n337 & n339 ;
  buffer buf_n341( .i (n340), .o (n341) );
  assign n342 = in_78_ & in_79_ ;
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  assign n352 = in_76_ | in_77_ ;
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  assign n360 = in_68_ | in_69_ ;
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  assign n364 = in_64_ | in_65_ ;
  buffer buf_n365( .i (n364), .o (n365) );
  assign n366 = in_67_ & in_66_ ;
  buffer buf_n367( .i (n366), .o (n367) );
  assign n368 = ( n361 & n365 ) | ( n361 & n367 ) | ( n365 & n367 ) ;
  buffer buf_n369( .i (n368), .o (n369) );
  assign n374 = ( ~n361 & n365 ) | ( ~n361 & n367 ) | ( n365 & n367 ) ;
  buffer buf_n375( .i (n374), .o (n375) );
  assign n376 = ( n363 & ~n369 ) | ( n363 & n375 ) | ( ~n369 & n375 ) ;
  buffer buf_n377( .i (n376), .o (n377) );
  assign n378 = in_74_ & in_75_ ;
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  assign n382 = in_70_ & in_71_ ;
  buffer buf_n383( .i (n382), .o (n383) );
  assign n384 = in_72_ | in_73_ ;
  buffer buf_n385( .i (n384), .o (n385) );
  assign n386 = ( n379 & n383 ) | ( n379 & n385 ) | ( n383 & n385 ) ;
  buffer buf_n387( .i (n386), .o (n387) );
  assign n392 = ( ~n379 & n383 ) | ( ~n379 & n385 ) | ( n383 & n385 ) ;
  buffer buf_n393( .i (n392), .o (n393) );
  assign n394 = ( n381 & ~n387 ) | ( n381 & n393 ) | ( ~n387 & n393 ) ;
  buffer buf_n395( .i (n394), .o (n395) );
  assign n396 = ( n357 & n377 ) | ( n357 & n395 ) | ( n377 & n395 ) ;
  buffer buf_n397( .i (n396), .o (n397) );
  assign n400 = ( ~n357 & n377 ) | ( ~n357 & n395 ) | ( n377 & n395 ) ;
  buffer buf_n401( .i (n400), .o (n401) );
  assign n402 = ( n359 & ~n397 ) | ( n359 & n401 ) | ( ~n397 & n401 ) ;
  buffer buf_n403( .i (n402), .o (n403) );
  assign n404 = n351 & n403 ;
  buffer buf_n405( .i (n404), .o (n405) );
  assign n406 = n351 | n403 ;
  buffer buf_n407( .i (n406), .o (n407) );
  assign n408 = ~n405 & n407 ;
  buffer buf_n409( .i (n408), .o (n409) );
  assign n410 = n341 & n409 ;
  buffer buf_n411( .i (n410), .o (n411) );
  assign n415 = n341 | n409 ;
  buffer buf_n416( .i (n415), .o (n416) );
  assign n417 = ~n411 & n416 ;
  buffer buf_n418( .i (n417), .o (n418) );
  assign n419 = n273 & n418 ;
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  assign n426 = ( n160 & n178 ) | ( n160 & n184 ) | ( n178 & n184 ) ;
  buffer buf_n427( .i (n426), .o (n427) );
  assign n432 = ( n160 & n178 ) | ( n160 & ~n184 ) | ( n178 & ~n184 ) ;
  buffer buf_n433( .i (n432), .o (n433) );
  assign n434 = ( n186 & ~n427 ) | ( n186 & n433 ) | ( ~n427 & n433 ) ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n436 = n192 & n435 ;
  buffer buf_n437( .i (n436), .o (n437) );
  assign n438 = n192 | n435 ;
  buffer buf_n439( .i (n438), .o (n439) );
  assign n440 = ~n437 & n439 ;
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  assign n442 = ( n230 & n246 ) | ( n230 & n252 ) | ( n246 & n252 ) ;
  buffer buf_n443( .i (n442), .o (n443) );
  assign n448 = ( n230 & n246 ) | ( n230 & ~n252 ) | ( n246 & ~n252 ) ;
  buffer buf_n449( .i (n448), .o (n449) );
  assign n450 = ( n254 & ~n443 ) | ( n254 & n449 ) | ( ~n443 & n449 ) ;
  buffer buf_n451( .i (n450), .o (n451) );
  assign n452 = n260 & n451 ;
  buffer buf_n453( .i (n452), .o (n453) );
  assign n454 = n260 | n451 ;
  buffer buf_n455( .i (n454), .o (n455) );
  assign n456 = ~n453 & n455 ;
  buffer buf_n457( .i (n456), .o (n457) );
  assign n458 = n441 & n457 ;
  assign n459 = n441 | n457 ;
  assign n460 = ~n458 & n459 ;
  buffer buf_n461( .i (n460), .o (n461) );
  assign n462 = n269 & n461 ;
  assign n463 = n269 | n461 ;
  assign n464 = ~n462 & n463 ;
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  assign n466 = ( n305 & n323 ) | ( n305 & n329 ) | ( n323 & n329 ) ;
  buffer buf_n467( .i (n466), .o (n467) );
  assign n472 = ( n305 & n323 ) | ( n305 & ~n329 ) | ( n323 & ~n329 ) ;
  buffer buf_n473( .i (n472), .o (n473) );
  assign n474 = ( n331 & ~n467 ) | ( n331 & n473 ) | ( ~n467 & n473 ) ;
  buffer buf_n475( .i (n474), .o (n475) );
  assign n476 = n337 & n475 ;
  buffer buf_n477( .i (n476), .o (n477) );
  assign n478 = n337 | n475 ;
  buffer buf_n479( .i (n478), .o (n479) );
  assign n480 = ~n477 & n479 ;
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  assign n482 = ( n373 & n391 ) | ( n373 & n397 ) | ( n391 & n397 ) ;
  buffer buf_n483( .i (n482), .o (n483) );
  assign n488 = ( n373 & n391 ) | ( n373 & ~n397 ) | ( n391 & ~n397 ) ;
  buffer buf_n489( .i (n488), .o (n489) );
  assign n490 = ( n399 & ~n483 ) | ( n399 & n489 ) | ( ~n483 & n489 ) ;
  buffer buf_n491( .i (n490), .o (n491) );
  assign n492 = n405 & n491 ;
  buffer buf_n493( .i (n492), .o (n493) );
  assign n494 = n405 | n491 ;
  buffer buf_n495( .i (n494), .o (n495) );
  assign n496 = ~n493 & n495 ;
  buffer buf_n497( .i (n496), .o (n497) );
  assign n498 = n481 & n497 ;
  assign n499 = n481 | n497 ;
  assign n500 = ~n498 & n499 ;
  buffer buf_n501( .i (n500), .o (n501) );
  assign n502 = n414 & n501 ;
  assign n503 = n414 | n501 ;
  assign n504 = ~n502 & n503 ;
  buffer buf_n505( .i (n504), .o (n505) );
  assign n506 = n465 & n505 ;
  assign n507 = n465 | n505 ;
  assign n508 = ~n506 & n507 ;
  buffer buf_n509( .i (n508), .o (n509) );
  assign n510 = n425 & n509 ;
  assign n511 = n425 | n509 ;
  assign n512 = ~n510 & n511 ;
  buffer buf_n513( .i (n512), .o (n513) );
  assign n514 = n273 | n418 ;
  buffer buf_n515( .i (n514), .o (n515) );
  assign n516 = ~n420 & n515 ;
  buffer buf_n517( .i (n516), .o (n517) );
  assign n518 = in_30_ & in_31_ ;
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  assign n528 = in_28_ | in_29_ ;
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  assign n536 = in_26_ & in_27_ ;
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  assign n540 = in_22_ & in_23_ ;
  buffer buf_n541( .i (n540), .o (n541) );
  assign n542 = in_24_ | in_25_ ;
  buffer buf_n543( .i (n542), .o (n543) );
  assign n544 = ( n537 & n541 ) | ( n537 & n543 ) | ( n541 & n543 ) ;
  buffer buf_n545( .i (n544), .o (n545) );
  assign n550 = ( ~n537 & n541 ) | ( ~n537 & n543 ) | ( n541 & n543 ) ;
  buffer buf_n551( .i (n550), .o (n551) );
  assign n552 = ( n539 & ~n545 ) | ( n539 & n551 ) | ( ~n545 & n551 ) ;
  buffer buf_n553( .i (n552), .o (n553) );
  assign n554 = in_20_ | in_21_ ;
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  assign n558 = in_17_ | in_16_ ;
  buffer buf_n559( .i (n558), .o (n559) );
  assign n560 = in_18_ & in_19_ ;
  buffer buf_n561( .i (n560), .o (n561) );
  assign n562 = ( n555 & n559 ) | ( n555 & n561 ) | ( n559 & n561 ) ;
  buffer buf_n563( .i (n562), .o (n563) );
  assign n568 = ( ~n555 & n559 ) | ( ~n555 & n561 ) | ( n559 & n561 ) ;
  buffer buf_n569( .i (n568), .o (n569) );
  assign n570 = ( n557 & ~n563 ) | ( n557 & n569 ) | ( ~n563 & n569 ) ;
  buffer buf_n571( .i (n570), .o (n571) );
  assign n572 = ( n533 & n553 ) | ( n533 & n571 ) | ( n553 & n571 ) ;
  buffer buf_n573( .i (n572), .o (n573) );
  assign n576 = ( ~n533 & n553 ) | ( ~n533 & n571 ) | ( n553 & n571 ) ;
  buffer buf_n577( .i (n576), .o (n577) );
  assign n578 = ( n535 & ~n573 ) | ( n535 & n577 ) | ( ~n573 & n577 ) ;
  buffer buf_n579( .i (n578), .o (n579) );
  assign n580 = n527 & n579 ;
  buffer buf_n581( .i (n580), .o (n581) );
  assign n582 = n527 | n579 ;
  buffer buf_n583( .i (n582), .o (n583) );
  assign n584 = ~n581 & n583 ;
  buffer buf_n585( .i (n584), .o (n585) );
  assign n586 = in_15_ & in_14_ ;
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  assign n596 = in_13_ | in_12_ ;
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  assign n604 = in_4_ | in_5_ ;
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  assign n608 = in_1_ | in_0_ ;
  buffer buf_n609( .i (n608), .o (n609) );
  assign n610 = in_3_ & in_2_ ;
  buffer buf_n611( .i (n610), .o (n611) );
  assign n612 = ( n605 & n609 ) | ( n605 & n611 ) | ( n609 & n611 ) ;
  buffer buf_n613( .i (n612), .o (n613) );
  assign n618 = ( ~n605 & n609 ) | ( ~n605 & n611 ) | ( n609 & n611 ) ;
  buffer buf_n619( .i (n618), .o (n619) );
  assign n620 = ( n607 & ~n613 ) | ( n607 & n619 ) | ( ~n613 & n619 ) ;
  buffer buf_n621( .i (n620), .o (n621) );
  assign n622 = in_10_ & in_11_ ;
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  assign n626 = in_7_ & in_6_ ;
  buffer buf_n627( .i (n626), .o (n627) );
  assign n628 = in_9_ | in_8_ ;
  buffer buf_n629( .i (n628), .o (n629) );
  assign n630 = ( n623 & n627 ) | ( n623 & n629 ) | ( n627 & n629 ) ;
  buffer buf_n631( .i (n630), .o (n631) );
  assign n636 = ( ~n623 & n627 ) | ( ~n623 & n629 ) | ( n627 & n629 ) ;
  buffer buf_n637( .i (n636), .o (n637) );
  assign n638 = ( n625 & ~n631 ) | ( n625 & n637 ) | ( ~n631 & n637 ) ;
  buffer buf_n639( .i (n638), .o (n639) );
  assign n640 = ( n601 & n621 ) | ( n601 & n639 ) | ( n621 & n639 ) ;
  buffer buf_n641( .i (n640), .o (n641) );
  assign n644 = ( ~n601 & n621 ) | ( ~n601 & n639 ) | ( n621 & n639 ) ;
  buffer buf_n645( .i (n644), .o (n645) );
  assign n646 = ( n603 & ~n641 ) | ( n603 & n645 ) | ( ~n641 & n645 ) ;
  buffer buf_n647( .i (n646), .o (n647) );
  assign n648 = n595 & n647 ;
  buffer buf_n649( .i (n648), .o (n649) );
  assign n650 = n595 | n647 ;
  buffer buf_n651( .i (n650), .o (n651) );
  assign n652 = ~n649 & n651 ;
  buffer buf_n653( .i (n652), .o (n653) );
  assign n654 = n585 & n653 ;
  buffer buf_n655( .i (n654), .o (n655) );
  assign n659 = n585 | n653 ;
  buffer buf_n660( .i (n659), .o (n660) );
  assign n661 = ~n655 & n660 ;
  buffer buf_n662( .i (n661), .o (n662) );
  assign n663 = in_47_ & in_46_ ;
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  assign n673 = in_44_ | in_45_ ;
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  assign n681 = in_36_ | in_37_ ;
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  assign n685 = in_33_ | in_32_ ;
  buffer buf_n686( .i (n685), .o (n686) );
  assign n687 = in_35_ & in_34_ ;
  buffer buf_n688( .i (n687), .o (n688) );
  assign n689 = ( n682 & n686 ) | ( n682 & n688 ) | ( n686 & n688 ) ;
  buffer buf_n690( .i (n689), .o (n690) );
  assign n695 = ( ~n682 & n686 ) | ( ~n682 & n688 ) | ( n686 & n688 ) ;
  buffer buf_n696( .i (n695), .o (n696) );
  assign n697 = ( n684 & ~n690 ) | ( n684 & n696 ) | ( ~n690 & n696 ) ;
  buffer buf_n698( .i (n697), .o (n698) );
  assign n699 = in_42_ & in_43_ ;
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  assign n703 = in_38_ & in_39_ ;
  buffer buf_n704( .i (n703), .o (n704) );
  assign n705 = in_40_ | in_41_ ;
  buffer buf_n706( .i (n705), .o (n706) );
  assign n707 = ( n700 & n704 ) | ( n700 & n706 ) | ( n704 & n706 ) ;
  buffer buf_n708( .i (n707), .o (n708) );
  assign n713 = ( ~n700 & n704 ) | ( ~n700 & n706 ) | ( n704 & n706 ) ;
  buffer buf_n714( .i (n713), .o (n714) );
  assign n715 = ( n702 & ~n708 ) | ( n702 & n714 ) | ( ~n708 & n714 ) ;
  buffer buf_n716( .i (n715), .o (n716) );
  assign n717 = ( n678 & n698 ) | ( n678 & n716 ) | ( n698 & n716 ) ;
  buffer buf_n718( .i (n717), .o (n718) );
  assign n721 = ( ~n678 & n698 ) | ( ~n678 & n716 ) | ( n698 & n716 ) ;
  buffer buf_n722( .i (n721), .o (n722) );
  assign n723 = ( n680 & ~n718 ) | ( n680 & n722 ) | ( ~n718 & n722 ) ;
  buffer buf_n724( .i (n723), .o (n724) );
  assign n725 = n672 & n724 ;
  buffer buf_n726( .i (n725), .o (n726) );
  assign n727 = n672 | n724 ;
  buffer buf_n728( .i (n727), .o (n728) );
  assign n729 = ~n726 & n728 ;
  buffer buf_n730( .i (n729), .o (n730) );
  assign n731 = in_63_ & in_62_ ;
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  assign n741 = in_60_ | in_61_ ;
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  assign n749 = in_58_ & in_59_ ;
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  assign n753 = in_54_ & in_55_ ;
  buffer buf_n754( .i (n753), .o (n754) );
  assign n755 = in_56_ | in_57_ ;
  buffer buf_n756( .i (n755), .o (n756) );
  assign n757 = ( n750 & n754 ) | ( n750 & n756 ) | ( n754 & n756 ) ;
  buffer buf_n758( .i (n757), .o (n758) );
  assign n763 = ( ~n750 & n754 ) | ( ~n750 & n756 ) | ( n754 & n756 ) ;
  buffer buf_n764( .i (n763), .o (n764) );
  assign n765 = ( n752 & ~n758 ) | ( n752 & n764 ) | ( ~n758 & n764 ) ;
  buffer buf_n766( .i (n765), .o (n766) );
  assign n767 = in_53_ | in_52_ ;
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  assign n771 = in_49_ | in_48_ ;
  buffer buf_n772( .i (n771), .o (n772) );
  assign n773 = in_50_ & in_51_ ;
  buffer buf_n774( .i (n773), .o (n774) );
  assign n775 = ( n768 & n772 ) | ( n768 & n774 ) | ( n772 & n774 ) ;
  buffer buf_n776( .i (n775), .o (n776) );
  assign n781 = ( ~n768 & n772 ) | ( ~n768 & n774 ) | ( n772 & n774 ) ;
  buffer buf_n782( .i (n781), .o (n782) );
  assign n783 = ( n770 & ~n776 ) | ( n770 & n782 ) | ( ~n776 & n782 ) ;
  buffer buf_n784( .i (n783), .o (n784) );
  assign n785 = ( n746 & n766 ) | ( n746 & n784 ) | ( n766 & n784 ) ;
  buffer buf_n786( .i (n785), .o (n786) );
  assign n789 = ( ~n746 & n766 ) | ( ~n746 & n784 ) | ( n766 & n784 ) ;
  buffer buf_n790( .i (n789), .o (n790) );
  assign n791 = ( n748 & ~n786 ) | ( n748 & n790 ) | ( ~n786 & n790 ) ;
  buffer buf_n792( .i (n791), .o (n792) );
  assign n793 = n740 & n792 ;
  buffer buf_n794( .i (n793), .o (n794) );
  assign n795 = n740 | n792 ;
  buffer buf_n796( .i (n795), .o (n796) );
  assign n797 = ~n794 & n796 ;
  buffer buf_n798( .i (n797), .o (n798) );
  assign n799 = n730 | n798 ;
  buffer buf_n800( .i (n799), .o (n800) );
  assign n801 = n730 & n798 ;
  buffer buf_n802( .i (n801), .o (n802) );
  assign n806 = n800 & ~n802 ;
  buffer buf_n807( .i (n806), .o (n807) );
  assign n808 = n662 & n807 ;
  buffer buf_n809( .i (n808), .o (n809) );
  assign n815 = n662 | n807 ;
  buffer buf_n816( .i (n815), .o (n816) );
  assign n817 = ~n809 & n816 ;
  buffer buf_n818( .i (n817), .o (n818) );
  assign n819 = n517 & n818 ;
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  assign n828 = ( n549 & n567 ) | ( n549 & n573 ) | ( n567 & n573 ) ;
  buffer buf_n829( .i (n828), .o (n829) );
  assign n834 = ( n549 & n567 ) | ( n549 & ~n573 ) | ( n567 & ~n573 ) ;
  buffer buf_n835( .i (n834), .o (n835) );
  assign n836 = ( n575 & ~n829 ) | ( n575 & n835 ) | ( ~n829 & n835 ) ;
  buffer buf_n837( .i (n836), .o (n837) );
  assign n838 = n581 | n837 ;
  buffer buf_n839( .i (n838), .o (n839) );
  assign n840 = n581 & n837 ;
  buffer buf_n841( .i (n840), .o (n841) );
  assign n842 = n839 & ~n841 ;
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  assign n844 = ( n617 & n635 ) | ( n617 & n641 ) | ( n635 & n641 ) ;
  buffer buf_n845( .i (n844), .o (n845) );
  assign n850 = ( n617 & n635 ) | ( n617 & ~n641 ) | ( n635 & ~n641 ) ;
  buffer buf_n851( .i (n850), .o (n851) );
  assign n852 = ( n643 & ~n845 ) | ( n643 & n851 ) | ( ~n845 & n851 ) ;
  buffer buf_n853( .i (n852), .o (n853) );
  assign n854 = n649 & n853 ;
  buffer buf_n855( .i (n854), .o (n855) );
  assign n856 = n649 | n853 ;
  buffer buf_n857( .i (n856), .o (n857) );
  assign n858 = ~n855 & n857 ;
  buffer buf_n859( .i (n858), .o (n859) );
  assign n860 = n843 & n859 ;
  assign n861 = n843 | n859 ;
  assign n862 = ~n860 & n861 ;
  buffer buf_n863( .i (n862), .o (n863) );
  assign n864 = n658 & n863 ;
  assign n865 = n658 | n863 ;
  assign n866 = ~n864 & n865 ;
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  assign n868 = ( n762 & n780 ) | ( n762 & n786 ) | ( n780 & n786 ) ;
  buffer buf_n869( .i (n868), .o (n869) );
  assign n874 = ( n762 & n780 ) | ( n762 & ~n786 ) | ( n780 & ~n786 ) ;
  buffer buf_n875( .i (n874), .o (n875) );
  assign n876 = ( n788 & ~n869 ) | ( n788 & n875 ) | ( ~n869 & n875 ) ;
  buffer buf_n877( .i (n876), .o (n877) );
  assign n878 = n794 & n877 ;
  buffer buf_n879( .i (n878), .o (n879) );
  assign n880 = n794 | n877 ;
  buffer buf_n881( .i (n880), .o (n881) );
  assign n882 = ~n879 & n881 ;
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  assign n884 = ( n694 & n712 ) | ( n694 & n718 ) | ( n712 & n718 ) ;
  buffer buf_n885( .i (n884), .o (n885) );
  assign n890 = ( n694 & n712 ) | ( n694 & ~n718 ) | ( n712 & ~n718 ) ;
  buffer buf_n891( .i (n890), .o (n891) );
  assign n892 = ( n720 & ~n885 ) | ( n720 & n891 ) | ( ~n885 & n891 ) ;
  buffer buf_n893( .i (n892), .o (n893) );
  assign n894 = n726 & n893 ;
  buffer buf_n895( .i (n894), .o (n895) );
  assign n896 = n726 | n893 ;
  buffer buf_n897( .i (n896), .o (n897) );
  assign n898 = ~n895 & n897 ;
  buffer buf_n899( .i (n898), .o (n899) );
  assign n900 = n883 & n899 ;
  assign n901 = n883 | n899 ;
  assign n902 = ~n900 & n901 ;
  buffer buf_n903( .i (n902), .o (n903) );
  assign n904 = n805 & n903 ;
  assign n905 = n805 | n903 ;
  assign n906 = ~n904 & n905 ;
  buffer buf_n907( .i (n906), .o (n907) );
  assign n908 = n867 & n907 ;
  assign n909 = n867 | n907 ;
  assign n910 = ~n908 & n909 ;
  buffer buf_n911( .i (n910), .o (n911) );
  assign n912 = n814 & n911 ;
  assign n913 = n814 | n911 ;
  assign n914 = ~n912 & n913 ;
  buffer buf_n915( .i (n914), .o (n915) );
  assign n916 = ( n513 & n824 ) | ( n513 & n915 ) | ( n824 & n915 ) ;
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  assign n921 = ( n811 & n867 ) | ( n811 & n907 ) | ( n867 & n907 ) ;
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  assign n926 = ( n655 & n843 ) | ( n655 & n859 ) | ( n843 & n859 ) ;
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  assign n931 = n833 & n841 ;
  buffer buf_n932( .i (n931), .o (n932) );
  assign n937 = n833 | n841 ;
  buffer buf_n938( .i (n937), .o (n938) );
  assign n939 = ~n932 & n938 ;
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  assign n941 = n849 & n855 ;
  buffer buf_n942( .i (n941), .o (n942) );
  assign n947 = n849 | n855 ;
  buffer buf_n948( .i (n947), .o (n948) );
  assign n949 = ~n942 & n948 ;
  buffer buf_n950( .i (n949), .o (n950) );
  assign n951 = n940 & n950 ;
  assign n952 = n940 | n950 ;
  assign n953 = ~n951 & n952 ;
  buffer buf_n954( .i (n953), .o (n954) );
  assign n955 = n930 & n954 ;
  assign n956 = n930 | n954 ;
  assign n957 = ~n955 & n956 ;
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  assign n959 = n889 & n895 ;
  buffer buf_n960( .i (n959), .o (n960) );
  assign n965 = n889 | n895 ;
  buffer buf_n966( .i (n965), .o (n966) );
  assign n967 = ~n960 & n966 ;
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  assign n969 = n873 & n879 ;
  buffer buf_n970( .i (n969), .o (n970) );
  assign n975 = n873 | n879 ;
  buffer buf_n976( .i (n975), .o (n976) );
  assign n977 = ~n970 & n976 ;
  buffer buf_n978( .i (n977), .o (n978) );
  assign n979 = n968 & n978 ;
  assign n980 = n968 | n978 ;
  assign n981 = ~n979 & n980 ;
  buffer buf_n982( .i (n981), .o (n982) );
  assign n983 = ( n802 & n883 ) | ( n802 & n899 ) | ( n883 & n899 ) ;
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  assign n988 = n982 & n987 ;
  assign n989 = n982 | n987 ;
  assign n990 = ~n988 & n989 ;
  buffer buf_n991( .i (n990), .o (n991) );
  assign n992 = n958 & n991 ;
  assign n993 = n958 | n991 ;
  assign n994 = ~n992 & n993 ;
  buffer buf_n995( .i (n994), .o (n995) );
  assign n996 = n925 & n995 ;
  assign n997 = n925 | n995 ;
  assign n998 = ~n996 & n997 ;
  buffer buf_n999( .i (n998), .o (n999) );
  assign n1000 = ( n422 & n465 ) | ( n422 & n505 ) | ( n465 & n505 ) ;
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  assign n1005 = ( n266 & n441 ) | ( n266 & n457 ) | ( n441 & n457 ) ;
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  assign n1010 = n431 & n437 ;
  buffer buf_n1011( .i (n1010), .o (n1011) );
  assign n1016 = n431 | n437 ;
  buffer buf_n1017( .i (n1016), .o (n1017) );
  assign n1018 = ~n1011 & n1017 ;
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  assign n1020 = n447 & n453 ;
  buffer buf_n1021( .i (n1020), .o (n1021) );
  assign n1026 = n447 | n453 ;
  buffer buf_n1027( .i (n1026), .o (n1027) );
  assign n1028 = ~n1021 & n1027 ;
  buffer buf_n1029( .i (n1028), .o (n1029) );
  assign n1030 = n1019 & n1029 ;
  assign n1031 = n1019 | n1029 ;
  assign n1032 = ~n1030 & n1031 ;
  buffer buf_n1033( .i (n1032), .o (n1033) );
  assign n1034 = n1009 & n1033 ;
  assign n1035 = n1009 | n1033 ;
  assign n1036 = ~n1034 & n1035 ;
  buffer buf_n1037( .i (n1036), .o (n1037) );
  assign n1038 = ( n411 & n481 ) | ( n411 & n497 ) | ( n481 & n497 ) ;
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  assign n1043 = n471 & n477 ;
  buffer buf_n1044( .i (n1043), .o (n1044) );
  assign n1049 = n471 | n477 ;
  buffer buf_n1050( .i (n1049), .o (n1050) );
  assign n1051 = ~n1044 & n1050 ;
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  assign n1053 = n487 & n493 ;
  buffer buf_n1054( .i (n1053), .o (n1054) );
  assign n1059 = n487 | n493 ;
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1061 = ~n1054 & n1060 ;
  buffer buf_n1062( .i (n1061), .o (n1062) );
  assign n1063 = n1052 & n1062 ;
  assign n1064 = n1052 | n1062 ;
  assign n1065 = ~n1063 & n1064 ;
  buffer buf_n1066( .i (n1065), .o (n1066) );
  assign n1067 = n1042 & n1066 ;
  assign n1068 = n1042 | n1066 ;
  assign n1069 = ~n1067 & n1068 ;
  buffer buf_n1070( .i (n1069), .o (n1070) );
  assign n1071 = n1037 & n1070 ;
  assign n1072 = n1037 | n1070 ;
  assign n1073 = ~n1071 & n1072 ;
  buffer buf_n1074( .i (n1073), .o (n1074) );
  assign n1075 = n1004 & n1074 ;
  assign n1076 = n1004 | n1074 ;
  assign n1077 = ~n1075 & n1076 ;
  buffer buf_n1078( .i (n1077), .o (n1078) );
  assign n1079 = n999 & n1078 ;
  assign n1080 = n999 | n1078 ;
  assign n1081 = ~n1079 & n1080 ;
  buffer buf_n1082( .i (n1081), .o (n1082) );
  assign n1083 = n920 & n1082 ;
  assign n1084 = n920 | n1082 ;
  assign n1085 = ~n1083 & n1084 ;
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  assign n1086 = n513 & n915 ;
  assign n1087 = n513 | n915 ;
  assign n1088 = ~n1086 & n1087 ;
  buffer buf_n1089( .i (n1088), .o (n1089) );
  assign n1090 = n827 & n1089 ;
  assign n1091 = n827 | n1089 ;
  assign n1092 = ~n1090 & n1091 ;
  assign n1093 = ( n922 & n958 ) | ( n922 & n991 ) | ( n958 & n991 ) ;
  buffer buf_n1094( .i (n1093), .o (n1094) );
  assign n1095 = n932 & n942 ;
  assign n1096 = n932 | n942 ;
  assign n1097 = ~n1095 & n1096 ;
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  assign n1100 = ( n927 & n940 ) | ( n927 & n950 ) | ( n940 & n950 ) ;
  buffer buf_n1101( .i (n1100), .o (n1101) );
  assign n1102 = n1099 & n1101 ;
  assign n1103 = n1099 | n1101 ;
  assign n1104 = ~n1102 & n1103 ;
  buffer buf_n1105( .i (n1104), .o (n1105) );
  assign n1109 = n960 & n970 ;
  assign n1110 = n960 | n970 ;
  assign n1111 = ~n1109 & n1110 ;
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  assign n1114 = ( n968 & n978 ) | ( n968 & n984 ) | ( n978 & n984 ) ;
  buffer buf_n1115( .i (n1114), .o (n1115) );
  assign n1116 = n1113 & n1115 ;
  assign n1117 = n1113 | n1115 ;
  assign n1118 = ~n1116 & n1117 ;
  buffer buf_n1119( .i (n1118), .o (n1119) );
  assign n1123 = n1105 & n1119 ;
  assign n1124 = n1105 | n1119 ;
  assign n1125 = ~n1123 & n1124 ;
  buffer buf_n1126( .i (n1125), .o (n1126) );
  assign n1127 = n1094 & n1126 ;
  assign n1128 = n1094 | n1126 ;
  assign n1129 = ~n1127 & n1128 ;
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  assign n1134 = ( n917 & n999 ) | ( n917 & n1078 ) | ( n999 & n1078 ) ;
  buffer buf_n1135( .i (n1134), .o (n1135) );
  assign n1136 = n1011 & n1021 ;
  assign n1137 = n1011 | n1021 ;
  assign n1138 = ~n1136 & n1137 ;
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  assign n1141 = ( n1006 & n1019 ) | ( n1006 & n1029 ) | ( n1019 & n1029 ) ;
  buffer buf_n1142( .i (n1141), .o (n1142) );
  assign n1143 = n1140 & n1142 ;
  assign n1144 = n1140 | n1142 ;
  assign n1145 = ~n1143 & n1144 ;
  buffer buf_n1146( .i (n1145), .o (n1146) );
  assign n1150 = n1044 & n1054 ;
  assign n1151 = n1044 | n1054 ;
  assign n1152 = ~n1150 & n1151 ;
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  assign n1155 = ( n1039 & n1052 ) | ( n1039 & n1062 ) | ( n1052 & n1062 ) ;
  buffer buf_n1156( .i (n1155), .o (n1156) );
  assign n1157 = n1154 & n1156 ;
  assign n1158 = n1154 | n1156 ;
  assign n1159 = ~n1157 & n1158 ;
  buffer buf_n1160( .i (n1159), .o (n1160) );
  assign n1164 = n1146 & n1160 ;
  assign n1165 = n1146 | n1160 ;
  assign n1166 = ~n1164 & n1165 ;
  buffer buf_n1167( .i (n1166), .o (n1167) );
  assign n1168 = ( n1001 & n1037 ) | ( n1001 & n1070 ) | ( n1037 & n1070 ) ;
  buffer buf_n1169( .i (n1168), .o (n1169) );
  assign n1170 = n1167 & n1169 ;
  assign n1171 = n1167 | n1169 ;
  assign n1172 = ~n1170 & n1171 ;
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  assign n1177 = ( n1133 & n1135 ) | ( n1133 & n1176 ) | ( n1135 & n1176 ) ;
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  assign n1179 = ( n1094 & n1108 ) | ( n1094 & n1122 ) | ( n1108 & n1122 ) ;
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  assign n1181 = ( n936 & n946 ) | ( n936 & n1101 ) | ( n946 & n1101 ) ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  assign n1189 = ( n964 & n974 ) | ( n964 & n1115 ) | ( n974 & n1115 ) ;
  buffer buf_n1190( .i (n1189), .o (n1190) );
  assign n1197 = n1182 & n1190 ;
  assign n1198 = n1182 | n1190 ;
  assign n1199 = ~n1197 & n1198 ;
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  assign n1204 = n1180 & n1203 ;
  assign n1205 = n1180 | n1203 ;
  assign n1206 = ~n1204 & n1205 ;
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  assign n1211 = ( n1015 & n1025 ) | ( n1015 & n1142 ) | ( n1025 & n1142 ) ;
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  assign n1219 = ( n1048 & n1058 ) | ( n1048 & n1156 ) | ( n1058 & n1156 ) ;
  buffer buf_n1220( .i (n1219), .o (n1220) );
  assign n1227 = n1212 & n1220 ;
  assign n1228 = n1212 | n1220 ;
  assign n1229 = ~n1227 & n1228 ;
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  assign n1234 = ( n1149 & n1163 ) | ( n1149 & n1169 ) | ( n1163 & n1169 ) ;
  buffer buf_n1235( .i (n1234), .o (n1235) );
  assign n1236 = n1233 & n1235 ;
  assign n1237 = n1233 | n1235 ;
  assign n1238 = ~n1236 & n1237 ;
  buffer buf_n1239( .i (n1238), .o (n1239) );
  assign n1243 = n1207 & n1239 ;
  assign n1244 = n1207 | n1239 ;
  assign n1245 = ~n1243 & n1244 ;
  buffer buf_n1246( .i (n1245), .o (n1246) );
  assign n1247 = n1178 & n1246 ;
  assign n1248 = n1178 | n1246 ;
  assign n1249 = ~n1247 & n1248 ;
  assign n1250 = n517 | n818 ;
  buffer buf_n1251( .i (n1250), .o (n1251) );
  assign n1252 = ~n820 & n1251 ;
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  assign n1253 = ( n1180 & n1188 ) | ( n1180 & n1196 ) | ( n1188 & n1196 ) ;
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  assign n1261 = ( n1178 & n1210 ) | ( n1178 & n1242 ) | ( n1210 & n1242 ) ;
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  assign n1263 = ( n1218 & n1226 ) | ( n1218 & n1235 ) | ( n1226 & n1235 ) ;
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  assign n1271 = ( n1260 & n1262 ) | ( n1260 & n1270 ) | ( n1262 & n1270 ) ;
  assign n1272 = n1130 & n1173 ;
  assign n1273 = n1130 | n1173 ;
  assign n1274 = ~n1272 & n1273 ;
  buffer buf_n1275( .i (n1274), .o (n1275) );
  assign n1276 = n1135 & n1275 ;
  assign n1277 = n1135 | n1275 ;
  assign n1278 = ~n1276 & n1277 ;
  assign n1279 = n1254 & n1264 ;
  assign n1280 = n1254 | n1264 ;
  assign n1281 = ~n1279 & n1280 ;
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  assign n1286 = n1262 & n1285 ;
  assign n1287 = n1262 | n1285 ;
  assign n1288 = ~n1286 & n1287 ;
  assign out_3_ = n1085 ;
  assign out_2_ = n1092 ;
  assign out_5_ = n1249 ;
  assign out_1_ = n1252 ;
  assign out_0_ = 1'b0 ;
  assign out_7_ = n1271 ;
  assign out_4_ = n1278 ;
  assign out_6_ = n1288 ;
endmodule
