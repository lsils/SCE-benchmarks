module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 ;
  buffer buf_n9( .i (x0), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  inverter inv_n30( .i (n29), .o (n30) );
  buffer buf_n52( .i (x2), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n71( .i (x3), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  assign n158 = n59 | n78 ;
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n31( .i (x1), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n90( .i (x4), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n108( .i (x5), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n125( .i (x6), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n142( .i (x7), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  assign n167 = n135 & n152 ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n171 = ~n120 & n168 ;
  buffer buf_n172( .i (n171), .o (n172) );
  assign n173 = n104 & n172 ;
  assign n174 = ~n46 & n173 ;
  assign n175 = ~n166 & n174 ;
  assign n176 = n99 & n117 ;
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n79( .i (n78), .o (n79) );
  assign n182 = n39 | n79 ;
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  assign n192 = ( n66 & ~n180 ) | ( n66 & n187 ) | ( ~n180 & n187 ) ;
  assign n193 = n181 | n192 ;
  assign n194 = ~n25 & n193 ;
  assign n195 = ( ~n26 & n175 ) | ( ~n26 & n194 ) | ( n175 & n194 ) ;
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  assign n199 = ~n134 & n151 ;
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  assign n206 = n67 & n123 ;
  assign n207 = ( n106 & n205 ) | ( n106 & n206 ) | ( n205 & n206 ) ;
  assign n208 = ~n107 & n207 ;
  assign n209 = n132 & ~n149 ;
  buffer buf_n210( .i (n209), .o (n210) );
  assign n212 = ~n117 & n210 ;
  buffer buf_n213( .i (n212), .o (n213) );
  assign n216 = ( n63 & n101 ) | ( n63 & n213 ) | ( n101 & n213 ) ;
  assign n217 = ~n64 & n216 ;
  assign n218 = ~n84 & n217 ;
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  assign n223 = ( ~n89 & n208 ) | ( ~n89 & n222 ) | ( n208 & n222 ) ;
  assign n224 = ( ~n28 & n50 ) | ( ~n28 & n223 ) | ( n50 & n223 ) ;
  assign n225 = ( ~n40 & n80 ) | ( ~n40 & n99 ) | ( n80 & n99 ) ;
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  assign n229 = n65 & ~n228 ;
  assign n230 = ( n44 & ~n65 ) | ( n44 & n228 ) | ( ~n65 & n228 ) ;
  assign n231 = ( ~n45 & n229 ) | ( ~n45 & n230 ) | ( n229 & n230 ) ;
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  assign n235 = ( n61 & n99 ) | ( n61 & ~n117 ) | ( n99 & ~n117 ) ;
  assign n236 = ( n62 & ~n135 ) | ( n62 & n235 ) | ( ~n135 & n235 ) ;
  buffer buf_n237( .i (n236), .o (n237) );
  assign n240 = n64 & ~n237 ;
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  assign n243 = n239 | n241 ;
  assign n244 = ( ~n67 & n242 ) | ( ~n67 & n243 ) | ( n242 & n243 ) ;
  assign n245 = ( n47 & n232 ) | ( n47 & ~n244 ) | ( n232 & ~n244 ) ;
  assign n246 = ~n88 & n245 ;
  assign n247 = ( n89 & n234 ) | ( n89 & n246 ) | ( n234 & n246 ) ;
  assign n248 = n28 | n247 ;
  assign n249 = ( ~n51 & n224 ) | ( ~n51 & ~n248 ) | ( n224 & ~n248 ) ;
  assign n250 = n81 | n118 ;
  buffer buf_n251( .i (n98), .o (n251) );
  assign n252 = n80 & n251 ;
  buffer buf_n253( .i (n252), .o (n253) );
  assign n255 = n100 & ~n118 ;
  assign n256 = ( n250 & ~n253 ) | ( n250 & n255 ) | ( ~n253 & n255 ) ;
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  assign n259 = n65 & ~n257 ;
  assign n260 = ( n45 & ~n258 ) | ( n45 & n259 ) | ( ~n258 & n259 ) ;
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  assign n263 = ( ~n43 & n83 ) | ( ~n43 & n120 ) | ( n83 & n120 ) ;
  buffer buf_n264( .i (n263), .o (n264) );
  assign n265 = ( n104 & n122 ) | ( n104 & ~n264 ) | ( n122 & ~n264 ) ;
  assign n266 = ( ~n85 & n104 ) | ( ~n85 & n264 ) | ( n104 & n264 ) ;
  assign n267 = n265 & ~n266 ;
  assign n268 = ~n81 & n118 ;
  buffer buf_n269( .i (n268), .o (n269) );
  assign n270 = ~n102 & n269 ;
  assign n271 = ~n44 & n270 ;
  assign n272 = ~n66 & n271 ;
  assign n273 = ( n84 & n103 ) | ( n84 & ~n228 ) | ( n103 & ~n228 ) ;
  assign n274 = n64 & n227 ;
  assign n275 = ( n44 & n228 ) | ( n44 & n274 ) | ( n228 & n274 ) ;
  assign n276 = n273 & ~n275 ;
  assign n277 = n272 | n276 ;
  assign n278 = ( ~n261 & n267 ) | ( ~n261 & n277 ) | ( n267 & n277 ) ;
  assign n279 = n262 | n278 ;
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  assign n282 = ( n59 & n78 ) | ( n59 & ~n115 ) | ( n78 & ~n115 ) ;
  buffer buf_n283( .i (n282), .o (n283) );
  assign n288 = ( n61 & n251 ) | ( n61 & ~n283 ) | ( n251 & ~n283 ) ;
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  assign n293 = ( ~n82 & n119 ) | ( ~n82 & n289 ) | ( n119 & n289 ) ;
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  assign n296 = n287 | n294 ;
  assign n297 = ( ~n292 & n295 ) | ( ~n292 & n296 ) | ( n295 & n296 ) ;
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  assign n300 = ( ~n47 & n141 ) | ( ~n47 & n298 ) | ( n141 & n298 ) ;
  buffer buf_n301( .i (n116), .o (n301) );
  assign n302 = n134 | n301 ;
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n103), .o (n308) );
  assign n309 = ~n164 & n308 ;
  assign n310 = ~n307 & n309 ;
  assign n311 = ~n47 & n310 ;
  assign n312 = ( ~n299 & n300 ) | ( ~n299 & n311 ) | ( n300 & n311 ) ;
  assign n313 = ( n60 & n116 ) | ( n60 & n133 ) | ( n116 & n133 ) ;
  assign n314 = ( n134 & ~n251 ) | ( n134 & n313 ) | ( ~n251 & n313 ) ;
  buffer buf_n315( .i (n314), .o (n315) );
  assign n318 = n136 & ~n315 ;
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  assign n321 = n317 | n319 ;
  assign n322 = ( ~n139 & n320 ) | ( ~n139 & n321 ) | ( n320 & n321 ) ;
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  assign n325 = n46 | n157 ;
  assign n326 = ( n87 & n323 ) | ( n87 & n325 ) | ( n323 & n325 ) ;
  assign n327 = n324 & ~n326 ;
  assign n328 = ( ~n27 & n312 ) | ( ~n27 & n327 ) | ( n312 & n327 ) ;
  assign n329 = ~n280 & n328 ;
  assign n330 = ( ~n29 & n281 ) | ( ~n29 & n329 ) | ( n281 & n329 ) ;
  buffer buf_n331( .i (n301), .o (n331) );
  assign n332 = ( n81 & n135 ) | ( n81 & n331 ) | ( n135 & n331 ) ;
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  assign n335 = n84 & n334 ;
  buffer buf_n336( .i (n63), .o (n336) );
  assign n337 = ( ~n83 & n333 ) | ( ~n83 & n336 ) | ( n333 & n336 ) ;
  assign n338 = ~n334 & n337 ;
  assign n339 = n335 | n338 ;
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n46), .o (n342) );
  assign n343 = n340 & ~n342 ;
  buffer buf_n344( .i (n336), .o (n344) );
  assign n345 = n305 | n344 ;
  assign n346 = ( ~n45 & n85 ) | ( ~n45 & n345 ) | ( n85 & n345 ) ;
  buffer buf_n347( .i (n43), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  assign n350 = n346 | n349 ;
  assign n351 = ( n61 & ~n80 ) | ( n61 & n301 ) | ( ~n80 & n301 ) ;
  buffer buf_n352( .i (n60), .o (n352) );
  buffer buf_n353( .i (n79), .o (n353) );
  buffer buf_n354( .i (n133), .o (n354) );
  assign n355 = ( n352 & n353 ) | ( n352 & ~n354 ) | ( n353 & ~n354 ) ;
  assign n356 = n351 | n355 ;
  assign n357 = ( n82 & ~n119 ) | ( n82 & n356 ) | ( ~n119 & n356 ) ;
  assign n358 = n102 | n357 ;
  assign n359 = ~n352 & n353 ;
  buffer buf_n360( .i (n359), .o (n360) );
  assign n365 = n301 & n354 ;
  buffer buf_n366( .i (n365), .o (n366) );
  assign n370 = n360 & n366 ;
  assign n371 = n102 & ~n370 ;
  assign n372 = n358 & ~n371 ;
  assign n373 = n348 | n372 ;
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  assign n374 = n101 | n303 ;
  buffer buf_n375( .i (n374), .o (n375) );
  assign n376 = n362 & ~n375 ;
  assign n377 = n348 & ~n376 ;
  assign n378 = n373 & ~n377 ;
  assign n379 = n350 & ~n378 ;
  assign n380 = ( ~n341 & n343 ) | ( ~n341 & n379 ) | ( n343 & n379 ) ;
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n124( .i (n123), .o (n124) );
  assign n383 = ( n103 & n344 ) | ( n103 & n347 ) | ( n344 & n347 ) ;
  assign n384 = ( n85 & n139 ) | ( n85 & n383 ) | ( n139 & n383 ) ;
  buffer buf_n385( .i (n384), .o (n385) );
  assign n386 = ( n124 & ~n141 ) | ( n124 & n385 ) | ( ~n141 & n385 ) ;
  assign n387 = ( n87 & n124 ) | ( n87 & ~n385 ) | ( n124 & ~n385 ) ;
  assign n388 = n386 & ~n387 ;
  assign n389 = ~n62 & n100 ;
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n83), .o (n392) );
  assign n393 = n391 & n392 ;
  assign n394 = n121 & n202 ;
  assign n395 = n393 & n394 ;
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  assign n398 = ( ~n95 & n130 ) | ( ~n95 & n147 ) | ( n130 & n147 ) ;
  buffer buf_n399( .i (n398), .o (n399) );
  assign n404 = ( n59 & ~n132 ) | ( n59 & n399 ) | ( ~n132 & n399 ) ;
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  assign n409 = ( n151 & ~n251 ) | ( n151 & n405 ) | ( ~n251 & n405 ) ;
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  assign n412 = ~n403 & n410 ;
  assign n413 = ( ~n408 & n411 ) | ( ~n408 & n412 ) | ( n411 & n412 ) ;
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n392), .o (n416) );
  assign n417 = ( ~n122 & n414 ) | ( ~n122 & n416 ) | ( n414 & n416 ) ;
  assign n418 = ( n219 & n415 ) | ( n219 & ~n417 ) | ( n415 & ~n417 ) ;
  assign n419 = n43 & ~n162 ;
  assign n420 = ( ~n179 & n202 ) | ( ~n179 & n419 ) | ( n202 & n419 ) ;
  assign n421 = n180 & n420 ;
  buffer buf_n422( .i (n421), .o (n422) );
  assign n423 = ( ~n396 & n418 ) | ( ~n396 & n422 ) | ( n418 & n422 ) ;
  assign n424 = n342 & ~n422 ;
  assign n425 = ( n397 & n423 ) | ( n397 & ~n424 ) | ( n423 & ~n424 ) ;
  assign n426 = ( ~n27 & n388 ) | ( ~n27 & n425 ) | ( n388 & n425 ) ;
  assign n427 = n381 & n426 ;
  assign n428 = ( ~n29 & ~n382 ) | ( ~n29 & n427 ) | ( ~n382 & n427 ) ;
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  assign n429 = n79 & n116 ;
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n115), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  assign n437 = ~n151 & n436 ;
  assign n438 = ( n41 & n430 ) | ( n41 & n437 ) | ( n430 & n437 ) ;
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n42), .o (n442) );
  assign n443 = ( n154 & n439 ) | ( n154 & ~n442 ) | ( n439 & ~n442 ) ;
  assign n444 = ( ~n121 & n433 ) | ( ~n121 & n443 ) | ( n433 & n443 ) ;
  assign n445 = ( ~n434 & n441 ) | ( ~n434 & n444 ) | ( n441 & n444 ) ;
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n446( .i (n353), .o (n446) );
  assign n447 = n211 & ~n446 ;
  assign n448 = ( n42 & ~n119 ) | ( n42 & n447 ) | ( ~n119 & n447 ) ;
  assign n449 = ~n442 & n448 ;
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  assign n452 = n139 & ~n450 ;
  assign n453 = ( n445 & n451 ) | ( n445 & ~n452 ) | ( n451 & ~n452 ) ;
  assign n454 = n106 & ~n453 ;
  assign n455 = ( n78 & n132 ) | ( n78 & n149 ) | ( n132 & n149 ) ;
  buffer buf_n456( .i (n455), .o (n456) );
  assign n461 = ( ~n353 & n436 ) | ( ~n353 & n456 ) | ( n436 & n456 ) ;
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  assign n466 = ( n136 & n153 ) | ( n136 & n462 ) | ( n153 & n462 ) ;
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  assign n469 = ~n460 & n467 ;
  assign n470 = ( ~n465 & n468 ) | ( ~n465 & n469 ) | ( n468 & n469 ) ;
  assign n471 = ~n349 & n470 ;
  assign n472 = n106 | n471 ;
  assign n473 = ~n454 & n472 ;
  assign n474 = n70 | n473 ;
  buffer buf_n475( .i (n150), .o (n475) );
  assign n476 = ( ~n354 & n436 ) | ( ~n354 & n475 ) | ( n436 & n475 ) ;
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  assign n481 = ~n153 & n477 ;
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n101), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  assign n486 = ( ~n121 & n482 ) | ( ~n121 & n485 ) | ( n482 & n485 ) ;
  assign n487 = ( n480 & n483 ) | ( n480 & n486 ) | ( n483 & n486 ) ;
  assign n488 = n86 | n487 ;
  assign n489 = n172 & ~n308 ;
  assign n490 = n86 & ~n489 ;
  assign n491 = n488 & ~n490 ;
  assign n492 = ~n48 & n491 ;
  assign n493 = n70 & ~n492 ;
  assign n494 = n474 & ~n493 ;
  assign n495 = ( ~n41 & n62 ) | ( ~n41 & n160 ) | ( n62 & n160 ) ;
  buffer buf_n496( .i (n352), .o (n496) );
  assign n497 = ( n41 & ~n160 ) | ( n41 & n496 ) | ( ~n160 & n496 ) ;
  assign n498 = ( ~n63 & n495 ) | ( ~n63 & n497 ) | ( n495 & n497 ) ;
  assign n499 = ( n120 & n137 ) | ( n120 & n498 ) | ( n137 & n498 ) ;
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n138), .o (n501) );
  assign n502 = ( n308 & n500 ) | ( n308 & ~n501 ) | ( n500 & ~n501 ) ;
  assign n503 = ( n122 & n308 ) | ( n122 & ~n500 ) | ( n308 & ~n500 ) ;
  assign n504 = n502 & ~n503 ;
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n40), .o (n507) );
  assign n508 = n496 & ~n507 ;
  buffer buf_n509( .i (n508), .o (n509) );
  assign n514 = n100 & ~n507 ;
  buffer buf_n515( .i (n514), .o (n515) );
  assign n517 = ( n390 & n509 ) | ( n390 & ~n515 ) | ( n509 & ~n515 ) ;
  assign n518 = ( n138 & ~n392 ) | ( n138 & n517 ) | ( ~n392 & n517 ) ;
  buffer buf_n519( .i (n518), .o (n519) );
  assign n520 = ( n123 & ~n140 ) | ( n123 & n519 ) | ( ~n140 & n519 ) ;
  assign n521 = ( n86 & ~n123 ) | ( n86 & n519 ) | ( ~n123 & n519 ) ;
  assign n522 = n520 & n521 ;
  assign n523 = ~n496 & n507 ;
  assign n524 = n160 | n507 ;
  assign n525 = ( ~n42 & n523 ) | ( ~n42 & n524 ) | ( n523 & n524 ) ;
  assign n526 = ( ~n137 & n484 ) | ( ~n137 & n525 ) | ( n484 & n525 ) ;
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n331), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  assign n532 = ( n501 & n527 ) | ( n501 & ~n531 ) | ( n527 & ~n531 ) ;
  buffer buf_n533( .i (n485), .o (n533) );
  assign n534 = ( n527 & n531 ) | ( n527 & ~n533 ) | ( n531 & ~n533 ) ;
  assign n535 = n532 | n534 ;
  assign n536 = n137 | n484 ;
  buffer buf_n537( .i (n98), .o (n537) );
  assign n538 = ( ~n352 & n354 ) | ( ~n352 & n537 ) | ( n354 & n537 ) ;
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n537), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  assign n543 = ( n82 & n539 ) | ( n82 & n542 ) | ( n539 & n542 ) ;
  assign n544 = n540 & n543 ;
  assign n545 = n536 & ~n544 ;
  assign n546 = n348 & ~n545 ;
  buffer buf_n547( .i (n446), .o (n547) );
  assign n548 = ~n136 & n547 ;
  buffer buf_n549( .i (n133), .o (n549) );
  assign n550 = n537 & ~n549 ;
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n549), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  assign n554 = ( ~n528 & n551 ) | ( ~n528 & n553 ) | ( n551 & n553 ) ;
  assign n555 = ( ~n528 & n547 ) | ( ~n528 & n551 ) | ( n547 & n551 ) ;
  assign n556 = ( n548 & n554 ) | ( n548 & ~n555 ) | ( n554 & ~n555 ) ;
  assign n557 = n344 & n556 ;
  buffer buf_n558( .i (n347), .o (n558) );
  assign n559 = n557 | n558 ;
  assign n560 = ~n546 & n559 ;
  assign n561 = n535 & ~n560 ;
  assign n562 = ( n505 & ~n522 ) | ( n505 & n561 ) | ( ~n522 & n561 ) ;
  assign n563 = ~n506 & n562 ;
  assign n564 = n28 | n563 ;
  assign n565 = ( ~n29 & n494 ) | ( ~n29 & ~n564 ) | ( n494 & ~n564 ) ;
  assign n566 = ( ~n19 & n183 ) | ( ~n19 & n496 ) | ( n183 & n496 ) ;
  assign n567 = n20 | n566 ;
  assign n568 = n529 | n567 ;
  assign n569 = ( n138 & ~n485 ) | ( n138 & n568 ) | ( ~n485 & n568 ) ;
  assign n570 = n533 | n569 ;
  assign n571 = n157 | n570 ;
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  inverter inv_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n553), .o (n577) );
  assign n578 = n529 & ~n577 ;
  assign n579 = ~n155 & n578 ;
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n531), .o (n582) );
  assign n583 = n580 | n582 ;
  assign n584 = n542 | n547 ;
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  assign n589 = ( ~n581 & n583 ) | ( ~n581 & n588 ) | ( n583 & n588 ) ;
  assign n590 = n48 | n589 ;
  assign n591 = ( ~n27 & n70 ) | ( ~n27 & n590 ) | ( n70 & n590 ) ;
  buffer buf_n592( .i (n26), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  assign n594 = n591 | n593 ;
  inverter inv_n595( .i (n594), .o (n595) );
  assign n596 = ( n484 & ~n529 ) | ( n484 & n577 ) | ( ~n529 & n577 ) ;
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  assign n599 = ( ~n105 & n582 ) | ( ~n105 & n598 ) | ( n582 & n598 ) ;
  assign n600 = n156 & ~n597 ;
  assign n601 = ( n140 & ~n598 ) | ( n140 & n600 ) | ( ~n598 & n600 ) ;
  assign n602 = n599 & ~n601 ;
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  assign n605 = ( n70 & n191 ) | ( n70 & ~n603 ) | ( n191 & ~n603 ) ;
  assign n606 = n604 | n605 ;
  buffer buf_n607( .i (n593), .o (n607) );
  assign n608 = ~n606 & ~n607 ;
  assign n609 = ( n76 & n113 ) | ( n76 & ~n147 ) | ( n113 & ~n147 ) ;
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n615( .i (n77), .o (n615) );
  assign n616 = ( n97 & ~n610 ) | ( n97 & n615 ) | ( ~n610 & n615 ) ;
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  assign n621 = ( ~n436 & n475 ) | ( ~n436 & n617 ) | ( n475 & n617 ) ;
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  assign n624 = n614 | n622 ;
  assign n625 = ( ~n620 & n623 ) | ( ~n620 & n624 ) | ( n623 & n624 ) ;
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  assign n628 = n501 & ~n626 ;
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  assign n629 = n215 & ~n585 ;
  buffer buf_n630( .i (n615), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n435), .o (n632) );
  assign n633 = ( n537 & ~n631 ) | ( n537 & n632 ) | ( ~n631 & n632 ) ;
  assign n634 = n446 & ~n633 ;
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  assign n637 = ( n269 & n577 ) | ( n269 & n635 ) | ( n577 & n635 ) ;
  assign n638 = n636 | n637 ;
  assign n639 = n629 | n638 ;
  assign n640 = ( n627 & n628 ) | ( n627 & ~n639 ) | ( n628 & ~n639 ) ;
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  assign n643 = n25 | n68 ;
  assign n644 = ( n48 & ~n641 ) | ( n48 & n643 ) | ( ~n641 & n643 ) ;
  assign n645 = n642 | n644 ;
  buffer buf_n646( .i (n645), .o (n646) );
  inverter inv_n647( .i (n646), .o (n647) );
  assign n648 = ~n331 & n552 ;
  buffer buf_n649( .i (n648), .o (n649) );
  assign n652 = n577 & ~n649 ;
  buffer buf_n653( .i (n652), .o (n653) );
  assign n654 = n533 & n653 ;
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  assign n655 = ( n416 & n651 ) | ( n416 & ~n653 ) | ( n651 & ~n653 ) ;
  assign n656 = ( n582 & ~n654 ) | ( n582 & n655 ) | ( ~n654 & n655 ) ;
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n131), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  assign n661 = ( ~n435 & n630 ) | ( ~n435 & n660 ) | ( n630 & n660 ) ;
  assign n662 = ( ~n475 & n631 ) | ( ~n475 & n661 ) | ( n631 & n661 ) ;
  buffer buf_n663( .i (n662), .o (n663) );
  assign n666 = n547 & ~n663 ;
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  assign n669 = n665 | n667 ;
  assign n670 = ( ~n416 & n668 ) | ( ~n416 & n669 ) | ( n668 & n669 ) ;
  assign n671 = n105 & ~n670 ;
  assign n672 = ( n152 & n331 ) | ( n152 & n552 ) | ( n331 & n552 ) ;
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n553), .o (n675) );
  assign n676 = n673 & ~n675 ;
  assign n677 = ( ~n530 & n674 ) | ( ~n530 & n676 ) | ( n674 & n676 ) ;
  assign n678 = ~n416 & n677 ;
  assign n679 = n105 | n678 ;
  assign n680 = ~n671 & n679 ;
  buffer buf_n681( .i (n392), .o (n681) );
  assign n682 = n66 & ~n681 ;
  assign n683 = n528 & ~n542 ;
  buffer buf_n684( .i (n446), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n542), .o (n686) );
  assign n687 = ( n683 & n685 ) | ( n683 & n686 ) | ( n685 & n686 ) ;
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n344), .o (n690) );
  assign n691 = ( n681 & n688 ) | ( n681 & ~n690 ) | ( n688 & ~n690 ) ;
  assign n692 = ( n682 & ~n689 ) | ( n682 & n691 ) | ( ~n689 & n691 ) ;
  buffer buf_n693( .i (n692), .o (n693) );
  assign n694 = ( n657 & n680 ) | ( n657 & n693 ) | ( n680 & n693 ) ;
  assign n695 = n69 & ~n693 ;
  assign n696 = ( n658 & ~n694 ) | ( n658 & n695 ) | ( ~n694 & n695 ) ;
  assign n697 = n50 | n696 ;
  assign n698 = ~n607 & ~n697 ;
  assign n699 = ( n77 & ~n96 ) | ( n77 & n131 ) | ( ~n96 & n131 ) ;
  buffer buf_n700( .i (n699), .o (n700) );
  assign n705 = ( ~n150 & n630 ) | ( ~n150 & n700 ) | ( n630 & n700 ) ;
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n709( .i (n631), .o (n709) );
  assign n710 = ~n706 & n709 ;
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  assign n713 = n708 | n711 ;
  buffer buf_n714( .i (n685), .o (n714) );
  assign n715 = ( n712 & n713 ) | ( n712 & ~n714 ) | ( n713 & ~n714 ) ;
  assign n716 = n531 & ~n715 ;
  buffer buf_n717( .i (n541), .o (n717) );
  assign n718 = ( n153 & n551 ) | ( n153 & n717 ) | ( n551 & n717 ) ;
  buffer buf_n719( .i (n152), .o (n719) );
  assign n720 = ( n551 & ~n717 ) | ( n551 & n719 ) | ( ~n717 & n719 ) ;
  assign n721 = ( n686 & ~n718 ) | ( n686 & n720 ) | ( ~n718 & n720 ) ;
  assign n722 = n714 | n721 ;
  buffer buf_n723( .i (n530), .o (n723) );
  assign n724 = n722 & ~n723 ;
  assign n725 = n716 | n724 ;
  assign n726 = ~n68 & n725 ;
  assign n727 = n580 & ~n587 ;
  assign n728 = n68 & ~n727 ;
  assign n729 = n726 | n728 ;
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  assign n732 = ( n50 & n593 ) | ( n50 & ~n730 ) | ( n593 & ~n730 ) ;
  assign n733 = ( n37 & ~n77 ) | ( n37 & n114 ) | ( ~n77 & n114 ) ;
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n739( .i (n60), .o (n739) );
  assign n740 = ( ~n632 & n735 ) | ( ~n632 & n739 ) | ( n735 & n739 ) ;
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n746( .i (n40), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n632), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  assign n750 = ( n741 & ~n747 ) | ( n741 & n749 ) | ( ~n747 & n749 ) ;
  assign n751 = ~n738 & n750 ;
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  assign n754 = n690 & ~n752 ;
  assign n755 = ( n745 & n753 ) | ( n745 & ~n754 ) | ( n753 & ~n754 ) ;
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = n107 & n756 ;
  assign n759 = n533 & n690 ;
  buffer buf_n760( .i (n681), .o (n760) );
  assign n761 = ( n349 & n759 ) | ( n349 & n760 ) | ( n759 & n760 ) ;
  assign n762 = ~n342 & n761 ;
  assign n763 = n553 & n717 ;
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n675), .o (n766) );
  assign n767 = n347 & ~n766 ;
  buffer buf_n768( .i (n442), .o (n768) );
  assign n769 = n585 & n768 ;
  assign n770 = ( n765 & n767 ) | ( n765 & ~n769 ) | ( n767 & ~n769 ) ;
  assign n771 = n582 & n770 ;
  buffer buf_n772( .i (n67), .o (n772) );
  assign n773 = n771 & ~n772 ;
  assign n774 = n762 | n773 ;
  assign n775 = ( n757 & ~n758 ) | ( n757 & n774 ) | ( ~n758 & n774 ) ;
  assign n776 = ~n593 & n775 ;
  assign n777 = ( ~n731 & ~n732 ) | ( ~n731 & n776 ) | ( ~n732 & n776 ) ;
  assign n778 = ( n530 & ~n766 ) | ( n530 & n768 ) | ( ~n766 & n768 ) ;
  assign n779 = ( n485 & ~n650 ) | ( n485 & n768 ) | ( ~n650 & n768 ) ;
  assign n780 = ~n778 & n779 ;
  buffer buf_n781( .i (n690), .o (n781) );
  assign n782 = ( n760 & n780 ) | ( n760 & ~n781 ) | ( n780 & ~n781 ) ;
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n783( .i (n749), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  assign n785 = ( n516 & n764 ) | ( n516 & ~n784 ) | ( n764 & ~n784 ) ;
  assign n786 = ( ~n516 & n766 ) | ( ~n516 & n784 ) | ( n766 & n784 ) ;
  assign n787 = ( ~n501 & n785 ) | ( ~n501 & n786 ) | ( n785 & n786 ) ;
  assign n788 = ( n760 & n781 ) | ( n760 & ~n787 ) | ( n781 & ~n787 ) ;
  assign n789 = n782 & ~n788 ;
  buffer buf_n790( .i (n739), .o (n790) );
  assign n791 = n746 | n790 ;
  assign n792 = ~n183 & n790 ;
  buffer buf_n793( .i (n790), .o (n793) );
  assign n794 = ( n791 & n792 ) | ( n791 & ~n793 ) | ( n792 & ~n793 ) ;
  assign n795 = ( n675 & n686 ) | ( n675 & n794 ) | ( n686 & n794 ) ;
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n766), .o (n797) );
  assign n798 = ( n723 & n796 ) | ( n723 & ~n797 ) | ( n796 & ~n797 ) ;
  buffer buf_n799( .i (n686), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  assign n801 = ( n723 & ~n796 ) | ( n723 & n800 ) | ( ~n796 & n800 ) ;
  assign n802 = n798 & ~n801 ;
  assign n803 = ( n98 & n435 ) | ( n98 & ~n734 ) | ( n435 & ~n734 ) ;
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  assign n808 = ( n709 & ~n746 ) | ( n709 & n804 ) | ( ~n746 & n804 ) ;
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  assign n811 = n738 | n809 ;
  assign n812 = ( ~n807 & n810 ) | ( ~n807 & n811 ) | ( n810 & n811 ) ;
  buffer buf_n813( .i (n336), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  assign n815 = n812 & ~n814 ;
  buffer buf_n816( .i (n97), .o (n816) );
  assign n817 = n630 & ~n816 ;
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  assign n822 = ~n768 & n821 ;
  assign n823 = n814 & ~n822 ;
  assign n824 = n815 | n823 ;
  assign n825 = ~n802 & n824 ;
  assign n826 = ~n789 & n825 ;
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  assign n829 = ( n34 & n74 ) | ( n34 & ~n145 ) | ( n74 & ~n145 ) ;
  buffer buf_n830( .i (n829), .o (n830) );
  assign n835 = ( n36 & n130 ) | ( n36 & ~n830 ) | ( n130 & ~n830 ) ;
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  assign n840 = ( n149 & ~n615 ) | ( n149 & n836 ) | ( ~n615 & n836 ) ;
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  assign n843 = n834 | n841 ;
  assign n844 = ( ~n839 & n842 ) | ( ~n839 & n843 ) | ( n842 & n843 ) ;
  assign n845 = n717 & ~n844 ;
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n552), .o (n848) );
  assign n849 = ( ~n684 & n719 ) | ( ~n684 & n848 ) | ( n719 & n848 ) ;
  buffer buf_n850( .i (n541), .o (n850) );
  assign n851 = ( n719 & n848 ) | ( n719 & n850 ) | ( n848 & n850 ) ;
  assign n852 = n849 & ~n851 ;
  assign n853 = n846 | n852 ;
  assign n854 = ( ~n558 & n847 ) | ( ~n558 & n853 ) | ( n847 & n853 ) ;
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  assign n857 = ( ~n124 & n772 ) | ( ~n124 & n855 ) | ( n772 & n855 ) ;
  assign n858 = ~n748 & n818 ;
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  assign n862 = ( n203 & n558 ) | ( n203 & n861 ) | ( n558 & n861 ) ;
  assign n863 = ~n349 & n862 ;
  assign n864 = ~n772 & n863 ;
  assign n865 = ( n856 & ~n857 ) | ( n856 & n864 ) | ( ~n857 & n864 ) ;
  assign n866 = n541 & ~n709 ;
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  assign n869 = ( ~n155 & n784 ) | ( ~n155 & n868 ) | ( n784 & n868 ) ;
  buffer buf_n870( .i (n850), .o (n870) );
  assign n871 = ( n783 & ~n867 ) | ( n783 & n870 ) | ( ~n867 & n870 ) ;
  assign n872 = ( n155 & n714 ) | ( n155 & ~n871 ) | ( n714 & ~n871 ) ;
  assign n873 = n869 | n872 ;
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  assign n876 = ( ~n141 & n513 ) | ( ~n141 & n874 ) | ( n513 & n874 ) ;
  assign n877 = ~n875 & n876 ;
  assign n878 = ( ~n592 & n865 ) | ( ~n592 & n877 ) | ( n865 & n877 ) ;
  assign n879 = n827 & n878 ;
  assign n880 = ( ~n607 & ~n828 ) | ( ~n607 & n879 ) | ( ~n828 & n879 ) ;
  buffer buf_n881( .i (n154), .o (n881) );
  assign n882 = ( ~n799 & n813 ) | ( ~n799 & n881 ) | ( n813 & n881 ) ;
  assign n883 = ~n684 & n848 ;
  assign n884 = ( n269 & n649 ) | ( n269 & ~n883 ) | ( n649 & ~n883 ) ;
  assign n885 = n154 | n336 ;
  assign n886 = ( ~n799 & n884 ) | ( ~n799 & n885 ) | ( n884 & n885 ) ;
  assign n887 = ~n882 & n886 ;
  buffer buf_n888( .i (n793), .o (n888) );
  assign n889 = ( n201 & n859 ) | ( n201 & n888 ) | ( n859 & n888 ) ;
  assign n890 = ~n813 & n889 ;
  buffer buf_n891( .i (n675), .o (n891) );
  assign n892 = n881 | n891 ;
  buffer buf_n254( .i (n253), .o (n254) );
  assign n893 = n793 & ~n850 ;
  assign n894 = n748 & ~n790 ;
  assign n895 = n684 & ~n894 ;
  assign n896 = ( n254 & n893 ) | ( n254 & ~n895 ) | ( n893 & ~n895 ) ;
  assign n897 = ( n881 & n891 ) | ( n881 & ~n896 ) | ( n891 & ~n896 ) ;
  assign n898 = ( n890 & n892 ) | ( n890 & ~n897 ) | ( n892 & ~n897 ) ;
  assign n899 = n887 | n898 ;
  assign n900 = n342 | n899 ;
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  assign n901 = n170 & n180 ;
  assign n902 = n364 & n901 ;
  buffer buf_n903( .i (n558), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  assign n905 = ~n902 & n904 ;
  assign n906 = n900 & ~n905 ;
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n909( .i (n848), .o (n909) );
  assign n910 = ( ~n704 & n783 ) | ( ~n704 & n909 ) | ( n783 & n909 ) ;
  assign n911 = ( ~n685 & n704 ) | ( ~n685 & n783 ) | ( n704 & n783 ) ;
  assign n912 = n910 & ~n911 ;
  assign n913 = n814 & ~n912 ;
  assign n914 = n375 | n714 ;
  assign n915 = ~n814 & n914 ;
  assign n916 = n913 | n915 ;
  assign n917 = ~n904 & n916 ;
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  assign n918 = n369 & ~n800 ;
  assign n919 = ~n165 & n918 ;
  assign n920 = n904 & ~n919 ;
  assign n921 = n917 | n920 ;
  buffer buf_n922( .i (n719), .o (n922) );
  assign n923 = ( n178 & n685 ) | ( n178 & n922 ) | ( n685 & n922 ) ;
  buffer buf_n924( .i (n709), .o (n924) );
  buffer buf_n925( .i (n475), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  assign n927 = ( ~n177 & n924 ) | ( ~n177 & n926 ) | ( n924 & n926 ) ;
  buffer buf_n928( .i (n749), .o (n928) );
  assign n929 = ( n870 & n927 ) | ( n870 & n928 ) | ( n927 & n928 ) ;
  assign n930 = ~n923 & n929 ;
  buffer buf_n931( .i (n813), .o (n931) );
  assign n932 = n930 | n931 ;
  assign n933 = ~n749 & n926 ;
  assign n934 = n870 & n933 ;
  buffer buf_n935( .i (n924), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  assign n937 = n934 & n936 ;
  assign n938 = n931 & ~n937 ;
  assign n939 = n932 & ~n938 ;
  assign n940 = n511 & n861 ;
  buffer buf_n941( .i (n940), .o (n941) );
  assign n942 = ( ~n904 & n939 ) | ( ~n904 & n941 ) | ( n939 & n941 ) ;
  assign n943 = n800 | n931 ;
  assign n944 = ( ~n760 & n781 ) | ( ~n760 & n943 ) | ( n781 & n943 ) ;
  buffer buf_n945( .i (n903), .o (n945) );
  assign n946 = ( n941 & n944 ) | ( n941 & n945 ) | ( n944 & n945 ) ;
  assign n947 = n942 | n946 ;
  assign n948 = ( n592 & n921 ) | ( n592 & ~n947 ) | ( n921 & ~n947 ) ;
  assign n949 = n907 | n948 ;
  assign n950 = ( ~n607 & n908 ) | ( ~n607 & ~n949 ) | ( n908 & ~n949 ) ;
  assign y0 = n30 ;
  assign y1 = n30 ;
  assign y2 = n30 ;
  assign y3 = n198 ;
  assign y4 = n249 ;
  assign y5 = n330 ;
  assign y6 = n428 ;
  assign y7 = n565 ;
  assign y8 = n576 ;
  assign y9 = n595 ;
  assign y10 = n608 ;
  assign y11 = n647 ;
  assign y12 = n698 ;
  assign y13 = n777 ;
  assign y14 = n880 ;
  assign y15 = n950 ;
endmodule
