module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 ;
  buffer buf_n66( .i (x2), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n124( .i (x4), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n94( .i (x3), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n154( .i (x5), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n212( .i (x7), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n240( .i (x8), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  assign n268 = n220 & ~n248 ;
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  assign n286 = ~n167 & n272 ;
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  assign n297 = ~n118 & n296 ;
  assign n298 = ( n91 & ~n149 ) | ( n91 & n297 ) | ( ~n149 & n297 ) ;
  assign n299 = ~n92 & n298 ;
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n10( .i (x0), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n38( .i (x1), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  assign n302 = n46 | n74 ;
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  assign n318 = n113 | n312 ;
  buffer buf_n319( .i (n318), .o (n319) );
  assign n320 = n31 & n319 ;
  assign n321 = n31 | n319 ;
  assign n322 = ~n320 & n321 ;
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  assign n325 = n220 | n248 ;
  buffer buf_n326( .i (n325), .o (n326) );
  assign n341 = ( ~n222 & n269 ) | ( ~n222 & n326 ) | ( n269 & n326 ) ;
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  assign n361 = ~n130 & n160 ;
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  assign n379 = ~n113 & n373 ;
  buffer buf_n380( .i (n379), .o (n380) );
  assign n387 = ~n31 & n380 ;
  assign n388 = ~n315 & n387 ;
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  assign n389 = ~n103 & n133 ;
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  assign n404 = ~n83 & n396 ;
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n30), .o (n408) );
  assign n409 = n407 & ~n408 ;
  assign n410 = ~n60 & n409 ;
  assign n411 = ( n353 & n388 ) | ( n353 & n410 ) | ( n388 & n410 ) ;
  assign n412 = ~n323 & n411 ;
  assign n413 = ( n324 & n355 ) | ( n324 & n412 ) | ( n355 & n412 ) ;
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  assign n417 = ( n37 & n65 ) | ( n37 & ~n414 ) | ( n65 & ~n414 ) ;
  assign n418 = n300 & n417 ;
  assign n419 = ( n301 & n416 ) | ( n301 & ~n418 ) | ( n416 & ~n418 ) ;
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  assign n421 = n77 & n105 ;
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  assign n435 = ~n103 & n163 ;
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  assign n447 = n162 | n248 ;
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  assign n460 = n84 & n456 ;
  assign n461 = ( n428 & n444 ) | ( n428 & ~n460 ) | ( n444 & ~n460 ) ;
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  assign n464 = n58 | n232 ;
  assign n465 = ( n145 & n462 ) | ( n145 & n464 ) | ( n462 & n464 ) ;
  assign n466 = n463 & ~n465 ;
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  assign n469 = ( n76 & ~n164 ) | ( n76 & n222 ) | ( ~n164 & n222 ) ;
  buffer buf_n470( .i (n469), .o (n470) );
  assign n478 = ( ~n136 & n224 ) | ( ~n136 & n470 ) | ( n224 & n470 ) ;
  buffer buf_n479( .i (n478), .o (n479) );
  assign n482 = n226 & ~n479 ;
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  assign n485 = n481 | n483 ;
  assign n486 = ( ~n229 & n484 ) | ( ~n229 & n485 ) | ( n484 & n485 ) ;
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n182( .i (x6), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  assign n489 = ~n194 & n252 ;
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  assign n505 = ( n57 & ~n487 ) | ( n57 & n495 ) | ( ~n487 & n495 ) ;
  assign n506 = n488 & n505 ;
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n195( .i (n194), .o (n195) );
  assign n509 = ~n167 & n195 ;
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  assign n522 = n79 | n137 ;
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  assign n530 = n514 & ~n527 ;
  assign n531 = ( n58 & ~n336 ) | ( n58 & n530 ) | ( ~n336 & n530 ) ;
  assign n532 = ~n59 & n531 ;
  assign n533 = ~n50 & n78 ;
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  assign n545 = n193 | n327 ;
  buffer buf_n546( .i (n545), .o (n546) );
  assign n554 = n167 & ~n546 ;
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  assign n560 = n107 & ~n137 ;
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  assign n573 = n559 & n565 ;
  assign n574 = n540 & n573 ;
  buffer buf_n575( .i (n574), .o (n575) );
  assign n576 = ( ~n507 & n532 ) | ( ~n507 & n575 ) | ( n532 & n575 ) ;
  assign n577 = n116 & ~n575 ;
  assign n578 = ( n508 & n576 ) | ( n508 & ~n577 ) | ( n576 & ~n577 ) ;
  assign n579 = n75 | n103 ;
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  assign n592 = n140 & ~n170 ;
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  assign n602 = n222 & n250 ;
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  assign n613 = n58 & n611 ;
  assign n614 = ( n590 & n596 ) | ( n590 & n613 ) | ( n596 & n613 ) ;
  assign n615 = ~n591 & n614 ;
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  assign n616 = ( n49 & n77 ) | ( n49 & ~n223 ) | ( n77 & ~n223 ) ;
  buffer buf_n617( .i (n616), .o (n617) );
  assign n628 = n225 | n617 ;
  assign n629 = ~n49 & n105 ;
  buffer buf_n630( .i (n629), .o (n630) );
  assign n638 = ( ~n79 & n617 ) | ( ~n79 & n630 ) | ( n617 & n630 ) ;
  assign n639 = ( ~n52 & n628 ) | ( ~n52 & n638 ) | ( n628 & n638 ) ;
  assign n640 = n255 & n639 ;
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  assign n643 = ( n81 & n109 ) | ( n81 & ~n227 ) | ( n109 & ~n227 ) ;
  assign n644 = ( n81 & n109 ) | ( n81 & n255 ) | ( n109 & n255 ) ;
  assign n645 = n643 & ~n644 ;
  assign n646 = n641 | n645 ;
  assign n647 = ( ~n56 & n642 ) | ( ~n56 & n646 ) | ( n642 & n646 ) ;
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  assign n651 = n135 & ~n223 ;
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  assign n662 = n51 & n225 ;
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n256( .i (n255), .o (n256) );
  assign n668 = ~n140 & n256 ;
  buffer buf_n669( .i (n668), .o (n669) );
  assign n672 = n56 & ~n669 ;
  assign n673 = ( n658 & n667 ) | ( n658 & ~n672 ) | ( n667 & ~n672 ) ;
  assign n674 = ( ~n86 & n648 ) | ( ~n86 & n673 ) | ( n648 & n673 ) ;
  assign n675 = n115 | n674 ;
  assign n676 = ( ~n116 & n650 ) | ( ~n116 & n675 ) | ( n650 & n675 ) ;
  assign n677 = n615 | n676 ;
  assign n678 = ( ~n467 & n578 ) | ( ~n467 & n677 ) | ( n578 & n677 ) ;
  assign n679 = n468 | n678 ;
  assign n680 = ~n36 & n679 ;
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  assign n683 = n106 | n136 ;
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  assign n696 = n520 & ~n695 ;
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  assign n697 = n87 & n400 ;
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  assign n700 = n23 & ~n51 ;
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  assign n711 = ~n587 & n704 ;
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  assign n721 = ( n432 & ~n698 ) | ( n432 & n715 ) | ( ~n698 & n715 ) ;
  assign n722 = ~n22 & n50 ;
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  assign n734 = n715 | n732 ;
  assign n735 = ( n699 & n721 ) | ( n699 & n734 ) | ( n721 & n734 ) ;
  buffer buf_n736( .i (n735), .o (n736) );
  assign n737 = ( ~n385 & n696 ) | ( ~n385 & n736 ) | ( n696 & n736 ) ;
  assign n738 = n49 & n77 ;
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  assign n750 = ~n26 & n742 ;
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  assign n761 = n736 | n759 ;
  assign n762 = ( n386 & n737 ) | ( n386 & n761 ) | ( n737 & n761 ) ;
  assign n763 = n681 | n762 ;
  assign n764 = ( n359 & n682 ) | ( n359 & n763 ) | ( n682 & n763 ) ;
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  assign n766 = ( n130 & n160 ) | ( n130 & ~n188 ) | ( n160 & ~n188 ) ;
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  assign n783 = ( ~n117 & n205 ) | ( ~n117 & n782 ) | ( n205 & n782 ) ;
  assign n784 = ( n117 & ~n147 ) | ( n117 & n782 ) | ( ~n147 & n782 ) ;
  assign n785 = n783 | n784 ;
  assign n786 = n91 & ~n785 ;
  assign n787 = ( n36 & n64 ) | ( n36 & n786 ) | ( n64 & n786 ) ;
  assign n788 = ~n37 & n787 ;
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  assign n791 = n134 & n164 ;
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  assign n806 = n112 & n798 ;
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  assign n816 = n22 & ~n106 ;
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n825( .i (n48), .o (n825) );
  assign n826 = ~n105 & n825 ;
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  assign n838 = ( n723 & n817 ) | ( n723 & ~n828 ) | ( n817 & ~n828 ) ;
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  assign n847 = ( n382 & ~n402 ) | ( n382 & n846 ) | ( ~n402 & n846 ) ;
  assign n848 = n732 | n846 ;
  assign n849 = ( n403 & n847 ) | ( n403 & n848 ) | ( n847 & n848 ) ;
  assign n850 = ~n91 & n849 ;
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n760( .i (n759), .o (n760) );
  assign n853 = n760 | n851 ;
  assign n854 = ( n815 & n852 ) | ( n815 & n853 ) | ( n852 & n853 ) ;
  buffer buf_n855( .i (n102), .o (n855) );
  assign n856 = ~n221 & n855 ;
  buffer buf_n857( .i (n856), .o (n857) );
  assign n863 = n163 & ~n221 ;
  buffer buf_n864( .i (n863), .o (n864) );
  assign n876 = ( n436 & n857 ) | ( n436 & ~n864 ) | ( n857 & ~n864 ) ;
  buffer buf_n877( .i (n876), .o (n877) );
  assign n882 = n253 & n877 ;
  assign n883 = n80 & ~n882 ;
  assign n884 = n164 | n326 ;
  buffer buf_n885( .i (n884), .o (n885) );
  assign n892 = n106 & ~n885 ;
  assign n893 = n79 | n892 ;
  buffer buf_n894( .i (n893), .o (n894) );
  assign n900 = ~n883 & n894 ;
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  assign n903 = ( ~n141 & n199 ) | ( ~n141 & n901 ) | ( n199 & n901 ) ;
  assign n904 = n196 & n439 ;
  assign n905 = ( n81 & n606 ) | ( n81 & n904 ) | ( n606 & n904 ) ;
  assign n906 = ~n82 & n905 ;
  assign n907 = n141 & n906 ;
  assign n908 = ( n902 & ~n903 ) | ( n902 & n907 ) | ( ~n903 & n907 ) ;
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  assign n912 = n83 & ~n687 ;
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  assign n917 = ~n223 & n251 ;
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  assign n931 = ( n909 & n914 ) | ( n909 & n925 ) | ( n914 & n925 ) ;
  assign n932 = n516 & ~n931 ;
  assign n933 = ( n517 & n911 ) | ( n517 & ~n932 ) | ( n911 & ~n932 ) ;
  assign n934 = n61 & ~n933 ;
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n935( .i (n104), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  assign n937 = ( n194 & n252 ) | ( n194 & n936 ) | ( n252 & n936 ) ;
  buffer buf_n938( .i (n937), .o (n938) );
  assign n944 = ( ~n226 & n254 ) | ( ~n226 & n938 ) | ( n254 & n938 ) ;
  buffer buf_n945( .i (n944), .o (n945) );
  assign n948 = n256 & ~n945 ;
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  assign n951 = n947 | n949 ;
  assign n952 = ( ~n259 & n950 ) | ( ~n259 & n951 ) | ( n950 & n951 ) ;
  buffer buf_n953( .i (n80), .o (n953) );
  assign n954 = ~n169 & n953 ;
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  assign n961 = n84 & ~n956 ;
  buffer buf_n962( .i (n961), .o (n962) );
  assign n963 = n952 & n962 ;
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  assign n964 = ( n101 & n189 ) | ( n101 & ~n219 ) | ( n189 & ~n219 ) ;
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  assign n976 = ~n943 & n975 ;
  assign n977 = ( ~n958 & n962 ) | ( ~n958 & n976 ) | ( n962 & n976 ) ;
  assign n978 = ( ~n175 & n963 ) | ( ~n175 & n977 ) | ( n963 & n977 ) ;
  assign n979 = ~n146 & n978 ;
  assign n980 = n61 | n979 ;
  assign n981 = ~n934 & n980 ;
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  assign n984 = ( ~n52 & n168 ) | ( ~n52 & n226 ) | ( n168 & n226 ) ;
  assign n985 = ( n169 & n953 ) | ( n169 & n984 ) | ( n953 & n984 ) ;
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  assign n989 = ( n55 & ~n83 ) | ( n55 & n986 ) | ( ~n83 & n986 ) ;
  assign n990 = ~n230 & n989 ;
  assign n991 = ( ~n173 & n988 ) | ( ~n173 & n990 ) | ( n988 & n990 ) ;
  assign n992 = n144 | n991 ;
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  assign n993 = ~n163 & n221 ;
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  assign n1004 = n745 & n1002 ;
  assign n1005 = n144 & ~n1004 ;
  assign n1006 = n992 & ~n1005 ;
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  assign n1009 = ( n117 & ~n263 ) | ( n117 & n1007 ) | ( ~n263 & n1007 ) ;
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n1010( .i (n166), .o (n1010) );
  assign n1011 = ~n329 & n1010 ;
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  assign n1019 = ( n59 & ~n529 ) | ( n59 & n1018 ) | ( ~n529 & n1018 ) ;
  assign n1020 = ~n60 & n1019 ;
  buffer buf_n1021( .i (n116), .o (n1021) );
  assign n1022 = n1020 & ~n1021 ;
  assign n1023 = ( n1008 & ~n1009 ) | ( n1008 & n1022 ) | ( ~n1009 & n1022 ) ;
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  assign n1024 = ( n50 & n136 ) | ( n50 & ~n252 ) | ( n136 & ~n252 ) ;
  buffer buf_n1025( .i (n1024), .o (n1025) );
  assign n1030 = ( n80 & n254 ) | ( n80 & n1025 ) | ( n254 & n1025 ) ;
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  assign n1035 = ( n54 & n140 ) | ( n54 & n1031 ) | ( n140 & n1031 ) ;
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  assign n1038 = n1029 & ~n1036 ;
  assign n1039 = ( n1034 & ~n1037 ) | ( n1034 & n1038 ) | ( ~n1037 & n1038 ) ;
  assign n1040 = n114 | n1039 ;
  assign n1041 = n134 & n250 ;
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  assign n1049 = ( n84 & n142 ) | ( n84 & n1048 ) | ( n142 & n1048 ) ;
  assign n1050 = ~n57 & n1049 ;
  assign n1051 = n114 & ~n1050 ;
  assign n1052 = n1040 & ~n1051 ;
  assign n1053 = n107 & n137 ;
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  assign n1063 = ( n85 & ~n259 ) | ( n85 & n312 ) | ( ~n259 & n312 ) ;
  assign n1064 = ( n85 & n259 ) | ( n85 & ~n312 ) | ( n259 & ~n312 ) ;
  assign n1065 = ( ~n86 & n1063 ) | ( ~n86 & n1064 ) | ( n1063 & n1064 ) ;
  assign n1066 = ( n115 & n145 ) | ( n115 & n1065 ) | ( n145 & n1065 ) ;
  assign n1067 = ( n1052 & ~n1061 ) | ( n1052 & n1066 ) | ( ~n1061 & n1066 ) ;
  assign n1068 = n235 | n1067 ;
  buffer buf_n1069( .i (n82), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  assign n1071 = ( n56 & n112 ) | ( n56 & ~n1070 ) | ( n112 & ~n1070 ) ;
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n57), .o (n1073) );
  assign n1074 = ~n1072 & n1073 ;
  buffer buf_n1075( .i (n78), .o (n1075) );
  buffer buf_n1076( .i (n135), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  assign n1078 = n1075 & n1077 ;
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  assign n1087 = ( ~n114 & n1072 ) | ( ~n114 & n1084 ) | ( n1072 & n1084 ) ;
  assign n1088 = ( n87 & ~n1074 ) | ( n87 & n1087 ) | ( ~n1074 & n1087 ) ;
  assign n1089 = n262 & ~n1088 ;
  assign n1090 = n235 & ~n1089 ;
  assign n1091 = n1068 & ~n1090 ;
  assign n1092 = ( ~n35 & n1023 ) | ( ~n35 & n1091 ) | ( n1023 & n1091 ) ;
  assign n1093 = ~n982 & n1092 ;
  assign n1094 = ( ~n37 & n983 ) | ( ~n37 & n1093 ) | ( n983 & n1093 ) ;
  buffer buf_n1095( .i (n1094), .o (n1095) );
  assign n1096 = ( ~n789 & n854 ) | ( ~n789 & n1095 ) | ( n854 & n1095 ) ;
  assign n1097 = n359 | n1095 ;
  assign n1098 = ( n790 & n1096 ) | ( n790 & n1097 ) | ( n1096 & n1097 ) ;
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n1099( .i (n220), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  assign n1102 = ( n165 & n935 ) | ( n165 & ~n1101 ) | ( n935 & ~n1101 ) ;
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  assign n1108 = n168 & ~n1104 ;
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  assign n1111 = ( ~n228 & n256 ) | ( ~n228 & n1109 ) | ( n256 & n1109 ) ;
  assign n1112 = ( ~n1107 & n1110 ) | ( ~n1107 & n1111 ) | ( n1110 & n1111 ) ;
  assign n1113 = n1070 & n1112 ;
  buffer buf_n1114( .i (n219), .o (n1114) );
  buffer buf_n1115( .i (n247), .o (n1115) );
  assign n1116 = ( n102 & ~n1114 ) | ( n102 & n1115 ) | ( ~n1114 & n1115 ) ;
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  assign n1127 = ( ~n165 & n251 ) | ( ~n165 & n1118 ) | ( n251 & n1118 ) ;
  buffer buf_n1128( .i (n1127), .o (n1128) );
  assign n1131 = n253 & ~n1128 ;
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n1134 = n1130 | n1132 ;
  buffer buf_n1135( .i (n255), .o (n1135) );
  assign n1136 = ( n1133 & n1134 ) | ( n1133 & ~n1135 ) | ( n1134 & ~n1135 ) ;
  buffer buf_n1137( .i (n1136), .o (n1137) );
  assign n1138 = n1070 | n1137 ;
  assign n1139 = ( ~n85 & n1113 ) | ( ~n85 & n1138 ) | ( n1113 & n1138 ) ;
  assign n1140 = n1073 & ~n1139 ;
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  assign n1141 = n170 & n275 ;
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  assign n1145 = n72 & ~n100 ;
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  assign n1158 = n1143 & n1157 ;
  assign n1159 = n1073 | n1158 ;
  assign n1160 = ~n1140 & n1159 ;
  assign n1161 = n146 & ~n1160 ;
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n1162( .i (n162), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  assign n1164 = ( n104 & n1100 ) | ( n104 & n1163 ) | ( n1100 & n1163 ) ;
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  assign n1173 = ( n111 & n257 ) | ( n111 & ~n1170 ) | ( n257 & ~n1170 ) ;
  assign n1174 = ( ~n225 & n253 ) | ( ~n225 & n1166 ) | ( n253 & n1166 ) ;
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  assign n1179 = ~n1173 & n1178 ;
  buffer buf_n1180( .i (n1070), .o (n1180) );
  assign n1181 = ~n1179 & n1180 ;
  assign n1182 = n899 & ~n1181 ;
  assign n1183 = ~n59 & n1182 ;
  assign n1184 = n146 | n1183 ;
  assign n1185 = ~n1161 & n1184 ;
  assign n1186 = n206 & ~n1185 ;
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  assign n1187 = n135 | n1101 ;
  buffer buf_n1188( .i (n1187), .o (n1188) );
  assign n1194 = ( n652 & ~n1077 ) | ( n652 & n1188 ) | ( ~n1077 & n1188 ) ;
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1207( .i (n254), .o (n1207) );
  assign n1208 = n1195 | n1207 ;
  assign n1209 = n170 | n1208 ;
  assign n1210 = n1069 & n1209 ;
  assign n1211 = n168 & n605 ;
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1222( .i (n139), .o (n1222) );
  assign n1223 = n1212 & n1222 ;
  assign n1224 = n1069 | n1223 ;
  assign n1225 = ~n1210 & n1224 ;
  assign n1226 = n113 & n1225 ;
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  assign n1229 = n293 | n1227 ;
  assign n1230 = ( n916 & n1228 ) | ( n916 & n1229 ) | ( n1228 & n1229 ) ;
  assign n1231 = n61 & n1230 ;
  assign n1232 = n206 | n1231 ;
  assign n1233 = ~n1186 & n1232 ;
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  assign n1236 = n37 & n1234 ;
  assign n1237 = n196 & n273 ;
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n1247( .i (n1246), .o (n1247) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  assign n1249 = n377 & n715 ;
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  assign n1252 = n1248 & n1251 ;
  assign n1253 = n561 & n953 ;
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  assign n1258 = n26 & n54 ;
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1262( .i (n55), .o (n1262) );
  assign n1263 = ~n1259 & n1262 ;
  buffer buf_n1264( .i (n1263), .o (n1264) );
  assign n1265 = n1257 & n1264 ;
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  assign n1266 = ( n406 & ~n1261 ) | ( n406 & n1264 ) | ( ~n1261 & n1264 ) ;
  assign n1267 = ( n408 & n1265 ) | ( n408 & n1266 ) | ( n1265 & n1266 ) ;
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  assign n1272 = ~n355 & n1270 ;
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  assign n1273 = ( n112 & ~n172 ) | ( n112 & n258 ) | ( ~n172 & n258 ) ;
  assign n1274 = n1126 & ~n1273 ;
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  assign n1277 = ( ~n249 & n855 ) | ( ~n249 & n1099 ) | ( n855 & n1099 ) ;
  assign n1278 = ( n134 & ~n250 ) | ( n134 & n1277 ) | ( ~n250 & n1277 ) ;
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1282( .i (n251), .o (n1282) );
  assign n1283 = n1279 & n1282 ;
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  assign n1286 = n1281 & ~n1284 ;
  assign n1287 = ( n1207 & ~n1285 ) | ( n1207 & n1286 ) | ( ~n1285 & n1286 ) ;
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  assign n1290 = ( ~n171 & n1069 ) | ( ~n171 & n1288 ) | ( n1069 & n1288 ) ;
  assign n1291 = n139 & n274 ;
  assign n1292 = ~n585 & n1291 ;
  assign n1293 = ~n171 & n1292 ;
  assign n1294 = ( ~n1289 & n1290 ) | ( ~n1289 & n1293 ) | ( n1290 & n1293 ) ;
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  assign n1298 = ( n86 & n144 ) | ( n86 & ~n1295 ) | ( n144 & ~n1295 ) ;
  assign n1299 = n1275 & n1298 ;
  assign n1300 = ( n1276 & n1297 ) | ( n1276 & ~n1299 ) | ( n1297 & ~n1299 ) ;
  buffer buf_n1301( .i (n60), .o (n1301) );
  assign n1302 = ( ~n33 & n1300 ) | ( ~n33 & n1301 ) | ( n1300 & n1301 ) ;
  assign n1303 = n918 & n1010 ;
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  assign n1311 = ~n1075 & n1077 ;
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  assign n1319 = n141 & ~n1314 ;
  buffer buf_n1320( .i (n1319), .o (n1320) );
  assign n1321 = n1308 & n1320 ;
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  assign n1322 = ( n291 & ~n1316 ) | ( n291 & n1320 ) | ( ~n1316 & n1320 ) ;
  buffer buf_n1323( .i (n1180), .o (n1323) );
  assign n1324 = ( n1321 & n1322 ) | ( n1321 & ~n1323 ) | ( n1322 & ~n1323 ) ;
  assign n1325 = n115 | n1324 ;
  assign n1326 = ( n224 & n1076 ) | ( n224 & n1282 ) | ( n1076 & n1282 ) ;
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1332( .i (n1010), .o (n1332) );
  buffer buf_n1333( .i (n1282), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  assign n1335 = ( n1327 & n1332 ) | ( n1327 & ~n1334 ) | ( n1332 & ~n1334 ) ;
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  assign n1340 = ( n228 & n1222 ) | ( n228 & n1336 ) | ( n1222 & n1336 ) ;
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  assign n1343 = ~n1331 & n1341 ;
  assign n1344 = ( ~n1339 & n1342 ) | ( ~n1339 & n1343 ) | ( n1342 & n1343 ) ;
  assign n1345 = ~n1323 & n1344 ;
  buffer buf_n1346( .i (n111), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  assign n1350 = ~n1345 & n1349 ;
  assign n1351 = n1325 & ~n1350 ;
  assign n1352 = ( n33 & n1301 ) | ( n33 & ~n1351 ) | ( n1301 & ~n1351 ) ;
  assign n1353 = n1302 & ~n1352 ;
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  assign n1354 = ( n110 & n1135 ) | ( n110 & n1191 ) | ( n1135 & n1191 ) ;
  buffer buf_n1355( .i (n1354), .o (n1355) );
  assign n1356 = n230 & ~n1355 ;
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  assign n1357 = ( ~n142 & n1193 ) | ( ~n142 & n1355 ) | ( n1193 & n1355 ) ;
  assign n1358 = ( ~n231 & n1356 ) | ( ~n231 & n1357 ) | ( n1356 & n1357 ) ;
  assign n1359 = ( ~n1073 & n1323 ) | ( ~n1073 & n1358 ) | ( n1323 & n1358 ) ;
  assign n1360 = ~n936 & n1282 ;
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  assign n1370 = ( ~n142 & n230 ) | ( ~n142 & n1365 ) | ( n230 & n1365 ) ;
  buffer buf_n1371( .i (n1222), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  assign n1373 = ( ~n258 & n1365 ) | ( ~n258 & n1372 ) | ( n1365 & n1372 ) ;
  assign n1374 = ( n1347 & n1370 ) | ( n1347 & n1373 ) | ( n1370 & n1373 ) ;
  buffer buf_n1375( .i (n1262), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  assign n1377 = ( n1323 & ~n1374 ) | ( n1323 & n1376 ) | ( ~n1374 & n1376 ) ;
  assign n1378 = n1359 & ~n1377 ;
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n1075), .o (n1381) );
  assign n1382 = n1334 | n1381 ;
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  assign n1389 = ( n143 & ~n231 ) | ( n143 & n1386 ) | ( ~n231 & n1386 ) ;
  assign n1390 = ( n143 & n1180 ) | ( n143 & ~n1386 ) | ( n1180 & ~n1386 ) ;
  assign n1391 = ( n260 & ~n1389 ) | ( n260 & n1390 ) | ( ~n1389 & n1390 ) ;
  buffer buf_n1392( .i (n1376), .o (n1392) );
  assign n1393 = ( ~n1349 & n1391 ) | ( ~n1349 & n1392 ) | ( n1391 & n1392 ) ;
  buffer buf_n1394( .i (n1180), .o (n1394) );
  assign n1395 = ( n336 & n528 ) | ( n336 & ~n1394 ) | ( n528 & ~n1394 ) ;
  assign n1396 = ( n1349 & n1392 ) | ( n1349 & ~n1395 ) | ( n1392 & ~n1395 ) ;
  assign n1397 = n1393 & n1396 ;
  buffer buf_n926( .i (n925), .o (n926) );
  assign n1398 = n26 & ~n309 ;
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  assign n1407 = ~n689 & n1400 ;
  buffer buf_n1408( .i (n1407), .o (n1408) );
  assign n1412 = n926 & n1408 ;
  buffer buf_n1413( .i (n1412), .o (n1413) );
  assign n1414 = ( ~n1379 & n1397 ) | ( ~n1379 & n1413 ) | ( n1397 & n1413 ) ;
  assign n1415 = n33 & ~n1413 ;
  assign n1416 = ( n1380 & n1414 ) | ( n1380 & ~n1415 ) | ( n1414 & ~n1415 ) ;
  assign n1417 = n1353 | n1416 ;
  assign n1418 = ( n1271 & ~n1272 ) | ( n1271 & n1417 ) | ( ~n1272 & n1417 ) ;
  assign n1419 = n1252 | n1418 ;
  assign n1420 = ( n1235 & ~n1236 ) | ( n1235 & n1419 ) | ( ~n1236 & n1419 ) ;
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  assign n1423 = n132 & ~n190 ;
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n207( .i (n206), .o (n207) );
  assign n1445 = ~n171 & n608 ;
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n249), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  assign n1453 = ( n166 & ~n936 ) | ( n166 & n1452 ) | ( ~n936 & n1452 ) ;
  buffer buf_n1454( .i (n1453), .o (n1454) );
  assign n1455 = ( n138 & ~n1334 ) | ( n138 & n1454 ) | ( ~n1334 & n1454 ) ;
  assign n1456 = ( n138 & n1332 ) | ( n138 & ~n1454 ) | ( n1332 & ~n1454 ) ;
  assign n1457 = n1455 & ~n1456 ;
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  assign n1460 = ( ~n55 & n229 ) | ( ~n55 & n1458 ) | ( n229 & n1458 ) ;
  buffer buf_n631( .i (n630), .o (n631) );
  assign n1461 = n138 & n631 ;
  assign n1462 = ( n169 & n1207 ) | ( n169 & n1461 ) | ( n1207 & n1461 ) ;
  assign n1463 = ~n1135 & n1462 ;
  assign n1464 = ~n229 & n1463 ;
  assign n1465 = ( n1459 & ~n1460 ) | ( n1459 & n1464 ) | ( ~n1460 & n1464 ) ;
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n566( .i (n565), .o (n566) );
  assign n1469 = ( n566 & ~n1376 ) | ( n566 & n1466 ) | ( ~n1376 & n1466 ) ;
  assign n1470 = n1448 & ~n1469 ;
  assign n1471 = ( n1449 & n1468 ) | ( n1449 & ~n1470 ) | ( n1468 & ~n1470 ) ;
  assign n1472 = n89 & ~n1471 ;
  assign n1473 = ( n110 & n228 ) | ( n110 & n1222 ) | ( n228 & n1222 ) ;
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  assign n1477 = ( n107 & n1077 ) | ( n107 & ~n1333 ) | ( n1077 & ~n1333 ) ;
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  assign n1484 = n1476 & ~n1483 ;
  assign n1485 = n175 & n1484 ;
  buffer buf_n1486( .i (n1392), .o (n1486) );
  assign n1487 = n1485 & ~n1486 ;
  assign n1488 = n89 | n1487 ;
  assign n1489 = ~n1472 & n1488 ;
  assign n1490 = ( ~n35 & n207 ) | ( ~n35 & n1489 ) | ( n207 & n1489 ) ;
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n1491( .i (n1076), .o (n1491) );
  assign n1492 = ~n51 & n1491 ;
  buffer buf_n1493( .i (n1492), .o (n1493) );
  assign n1498 = n139 & ~n1493 ;
  buffer buf_n1499( .i (n1498), .o (n1499) );
  assign n1500 = n881 & n1499 ;
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  assign n1501 = n166 | n224 ;
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1505( .i (n1504), .o (n1505) );
  assign n1513 = ( n1495 & ~n1499 ) | ( n1495 & n1505 ) | ( ~n1499 & n1505 ) ;
  assign n1514 = ( n1262 & ~n1500 ) | ( n1262 & n1513 ) | ( ~n1500 & n1513 ) ;
  buffer buf_n1515( .i (n82), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  assign n1518 = n1514 & ~n1517 ;
  assign n1519 = ( n48 & n104 ) | ( n48 & n1163 ) | ( n104 & n1163 ) ;
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1525( .i (n1101), .o (n1525) );
  assign n1526 = ( ~n936 & n1520 ) | ( ~n936 & n1525 ) | ( n1520 & n1525 ) ;
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  assign n1531 = ( n52 & n1332 ) | ( n52 & n1527 ) | ( n1332 & n1527 ) ;
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n1522( .i (n1521), .o (n1522) );
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  assign n1534 = n1524 & ~n1532 ;
  assign n1535 = ( n1530 & ~n1533 ) | ( n1530 & n1534 ) | ( ~n1533 & n1534 ) ;
  assign n1536 = ~n1372 & n1535 ;
  assign n1537 = n1517 & ~n1536 ;
  assign n1538 = n1518 | n1537 ;
  assign n1539 = n261 | n1538 ;
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  assign n1542 = ~n110 & n1212 ;
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n145), .o (n1548) );
  assign n1549 = n1547 & ~n1548 ;
  assign n1550 = n1540 & ~n1549 ;
  assign n1551 = ( n62 & n1541 ) | ( n62 & n1550 ) | ( n1541 & n1550 ) ;
  assign n1552 = ( n35 & n207 ) | ( n35 & n1551 ) | ( n207 & n1551 ) ;
  assign n1553 = n1490 & ~n1552 ;
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n1556( .i (n935), .o (n1556) );
  buffer buf_n1557( .i (n165), .o (n1557) );
  assign n1558 = n1556 | n1557 ;
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  assign n1565 = n143 | n1564 ;
  buffer buf_n1566( .i (n1565), .o (n1566) );
  assign n1569 = n23 & n1075 ;
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  assign n1577 = n29 & ~n1574 ;
  buffer buf_n1578( .i (n1577), .o (n1578) );
  assign n1579 = ~n1566 & n1578 ;
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  assign n1580 = ( n808 & ~n1576 ) | ( n808 & n1578 ) | ( ~n1576 & n1578 ) ;
  assign n1581 = ( n88 & n1579 ) | ( n88 & n1580 ) | ( n1579 & n1580 ) ;
  assign n1582 = n1301 | n1581 ;
  buffer buf_n1583( .i (n1491), .o (n1583) );
  assign n1584 = ( ~n1332 & n1381 ) | ( ~n1332 & n1583 ) | ( n1381 & n1583 ) ;
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  assign n1591 = n172 | n1587 ;
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  assign n1594 = ( n1348 & n1394 ) | ( n1348 & ~n1592 ) | ( n1394 & ~n1592 ) ;
  assign n1595 = ( n1590 & n1593 ) | ( n1590 & ~n1594 ) | ( n1593 & ~n1594 ) ;
  assign n1596 = n32 | n1595 ;
  assign n1597 = n1301 & n1596 ;
  assign n1598 = n1582 & ~n1597 ;
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  assign n1601 = ~n238 & n1599 ;
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  assign n1602 = n757 & ~n1512 ;
  assign n1603 = ~n695 & n1602 ;
  buffer buf_n1604( .i (n133), .o (n1604) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  assign n1606 = n1101 & n1605 ;
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  assign n1615 = ( n257 & ~n1314 ) | ( n257 & n1371 ) | ( ~n1314 & n1371 ) ;
  buffer buf_n1616( .i (n227), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  assign n1618 = ( ~n257 & n1314 ) | ( ~n257 & n1617 ) | ( n1314 & n1617 ) ;
  assign n1619 = ( ~n1612 & n1615 ) | ( ~n1612 & n1618 ) | ( n1615 & n1618 ) ;
  assign n1620 = n173 & n1619 ;
  buffer buf_n1621( .i (n1525), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  assign n1623 = ( n1334 & ~n1381 ) | ( n1334 & n1622 ) | ( ~n1381 & n1622 ) ;
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  assign n1629 = ~n1616 & n1624 ;
  assign n1630 = ( n1515 & n1625 ) | ( n1515 & n1629 ) | ( n1625 & n1629 ) ;
  assign n1631 = n1372 & n1630 ;
  assign n1632 = n173 | n1631 ;
  assign n1633 = ~n1620 & n1632 ;
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  assign n1634 = ( n367 & n652 ) | ( n367 & ~n866 ) | ( n652 & ~n866 ) ;
  buffer buf_n1635( .i (n1634), .o (n1635) );
  assign n1638 = ( n953 & n1207 ) | ( n953 & n1635 ) | ( n1207 & n1635 ) ;
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1135), .o (n1640) );
  assign n1641 = ( n27 & n1639 ) | ( n27 & ~n1640 ) | ( n1639 & ~n1640 ) ;
  assign n1642 = ( n27 & n1515 ) | ( n27 & ~n1639 ) | ( n1515 & ~n1639 ) ;
  assign n1643 = n1641 & ~n1642 ;
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  assign n1646 = n30 & ~n1644 ;
  assign n1647 = ( n1633 & n1645 ) | ( n1633 & ~n1646 ) | ( n1645 & ~n1646 ) ;
  buffer buf_n1648( .i (n1349), .o (n1648) );
  assign n1649 = n1647 | n1648 ;
  assign n1650 = n525 & n1640 ;
  assign n1651 = ( n609 & n657 ) | ( n609 & ~n1650 ) | ( n657 & ~n1650 ) ;
  buffer buf_n1652( .i (n172), .o (n1652) );
  assign n1653 = n1651 | n1652 ;
  assign n1654 = n334 | n526 ;
  assign n1655 = n1652 & n1654 ;
  assign n1656 = n1653 & ~n1655 ;
  assign n1657 = ~n408 & n1656 ;
  assign n1658 = n1648 & ~n1657 ;
  assign n1659 = n1649 & ~n1658 ;
  assign n1660 = n62 | n1659 ;
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  assign n1661 = n915 & ~n1310 ;
  assign n1662 = ( ~n76 & n1163 ) | ( ~n76 & n1604 ) | ( n1163 & n1604 ) ;
  buffer buf_n1663( .i (n1662), .o (n1663) );
  assign n1669 = ( n78 & ~n1525 ) | ( n78 & n1663 ) | ( ~n1525 & n1663 ) ;
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1010), .o (n1674) );
  assign n1675 = ( n1583 & n1670 ) | ( n1583 & n1674 ) | ( n1670 & n1674 ) ;
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  assign n1678 = ~n1667 & n1676 ;
  assign n1679 = ( ~n1673 & n1677 ) | ( ~n1673 & n1678 ) | ( n1677 & n1678 ) ;
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n258), .o (n1682) );
  assign n1683 = ( ~n1347 & n1680 ) | ( ~n1347 & n1682 ) | ( n1680 & n1682 ) ;
  assign n1684 = ~n580 & n1605 ;
  buffer buf_n1685( .i (n1684), .o (n1685) );
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  assign n1692 = ~n1506 & n1690 ;
  assign n1693 = ~n1682 & n1692 ;
  assign n1694 = ( n1681 & ~n1683 ) | ( n1681 & n1693 ) | ( ~n1683 & n1693 ) ;
  assign n1695 = ~n1081 & n1515 ;
  buffer buf_n1696( .i (n1695), .o (n1696) );
  assign n1697 = n1446 & n1696 ;
  assign n1698 = ( n1016 & ~n1083 ) | ( n1016 & n1696 ) | ( ~n1083 & n1696 ) ;
  buffer buf_n1699( .i (n1372), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  assign n1701 = ( n1697 & n1698 ) | ( n1697 & n1700 ) | ( n1698 & n1700 ) ;
  assign n1702 = n1694 | n1701 ;
  assign n1703 = ( n916 & ~n1661 ) | ( n916 & n1702 ) | ( ~n1661 & n1702 ) ;
  buffer buf_n1704( .i (n32), .o (n1704) );
  assign n1705 = n1703 & ~n1704 ;
  assign n1706 = n62 & ~n1705 ;
  assign n1707 = n1660 & ~n1706 ;
  assign n1708 = n1603 | n1707 ;
  assign n1709 = ( n1600 & ~n1601 ) | ( n1600 & n1708 ) | ( ~n1601 & n1708 ) ;
  assign n1710 = n132 | n190 ;
  buffer buf_n1711( .i (n1710), .o (n1711) );
  assign n1730 = ( n1424 & ~n1604 ) | ( n1424 & n1711 ) | ( ~n1604 & n1711 ) ;
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1381), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  assign n1744 = n1640 & ~n1743 ;
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  assign n1748 = ( n1348 & n1739 ) | ( n1348 & ~n1746 ) | ( n1739 & ~n1746 ) ;
  assign n1749 = n1740 & ~n1748 ;
  assign n1750 = n1486 | n1749 ;
  assign n1751 = n194 | n1452 ;
  buffer buf_n1752( .i (n1751), .o (n1752) );
  assign n1760 = n1583 & ~n1752 ;
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  assign n1767 = n430 & n1766 ;
  assign n1768 = n1486 & ~n1767 ;
  assign n1769 = n1750 & ~n1768 ;
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n867( .i (n866), .o (n867) );
  assign n1772 = ( n867 & n1502 ) | ( n867 & ~n1674 ) | ( n1502 & ~n1674 ) ;
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n34), .o (n1783) );
  assign n1784 = ( n1770 & ~n1782 ) | ( n1770 & n1783 ) | ( ~n1782 & n1783 ) ;
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  assign n1785 = n260 & n399 ;
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  assign n1788 = ( n205 & n1404 ) | ( n205 & n1787 ) | ( n1404 & n1787 ) ;
  assign n1789 = ~n206 & n1788 ;
  assign n1790 = n1782 & n1789 ;
  assign n1791 = ( n1771 & ~n1784 ) | ( n1771 & n1790 ) | ( ~n1784 & n1790 ) ;
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  assign n1792 = ~n130 & n188 ;
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  assign n1811 = n930 & n1810 ;
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n1812( .i (n1333), .o (n1812) );
  buffer buf_n1813( .i (n1812), .o (n1813) );
  assign n1814 = ( n53 & n1741 ) | ( n53 & ~n1813 ) | ( n1741 & ~n1813 ) ;
  assign n1815 = n620 & ~n1814 ;
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  assign n1819 = ( n277 & ~n311 ) | ( n277 & n1816 ) | ( ~n311 & n1816 ) ;
  assign n1820 = n1347 & ~n1819 ;
  assign n1821 = ( n1348 & n1818 ) | ( n1348 & ~n1820 ) | ( n1818 & ~n1820 ) ;
  buffer buf_n1822( .i (n1583), .o (n1822) );
  assign n1823 = n197 & n1822 ;
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1825( .i (n1824), .o (n1825) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  assign n1829 = n201 & ~n1826 ;
  buffer buf_n1830( .i (n1829), .o (n1830) );
  assign n1831 = n1821 & n1830 ;
  buffer buf_n1827( .i (n1826), .o (n1827) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1832( .i (n76), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  assign n1836 = ( n108 & ~n1812 ) | ( n108 & n1835 ) | ( ~n1812 & n1835 ) ;
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n109), .o (n1841) );
  assign n1842 = n1837 & ~n1841 ;
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  assign n1845 = ( n1262 & n1516 ) | ( n1262 & ~n1843 ) | ( n1516 & ~n1843 ) ;
  assign n1846 = ( n1840 & n1844 ) | ( n1840 & ~n1845 ) | ( n1844 & ~n1845 ) ;
  assign n1847 = n231 | n1817 ;
  assign n1848 = ( n1818 & n1846 ) | ( n1818 & n1847 ) | ( n1846 & n1847 ) ;
  assign n1849 = ( ~n1828 & n1830 ) | ( ~n1828 & n1848 ) | ( n1830 & n1848 ) ;
  assign n1850 = ( n1548 & n1831 ) | ( n1548 & n1849 ) | ( n1831 & n1849 ) ;
  assign n1851 = ~n1704 & n1850 ;
  buffer buf_n1852( .i (n1851), .o (n1852) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  assign n1854 = n717 | n1852 ;
  assign n1855 = ( n1811 & n1853 ) | ( n1811 & n1854 ) | ( n1853 & n1854 ) ;
  assign n1856 = n1791 | n1855 ;
  assign n1857 = ( ~n1554 & n1709 ) | ( ~n1554 & n1856 ) | ( n1709 & n1856 ) ;
  assign n1858 = n1555 | n1857 ;
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n1859( .i (n75), .o (n1859) );
  assign n1860 = ( n1100 & ~n1450 ) | ( n1100 & n1859 ) | ( ~n1450 & n1859 ) ;
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  buffer buf_n1872( .i (n1871), .o (n1872) );
  assign n1873 = ( n1100 & n1163 ) | ( n1100 & n1450 ) | ( n1163 & n1450 ) ;
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  buffer buf_n1879( .i (n1878), .o (n1879) );
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  assign n1886 = ~n1872 & n1885 ;
  buffer buf_n1887( .i (n1674), .o (n1887) );
  buffer buf_n1888( .i (n1887), .o (n1888) );
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  assign n1891 = ( n348 & n1516 ) | ( n348 & n1890 ) | ( n1516 & n1890 ) ;
  buffer buf_n1892( .i (n1891), .o (n1892) );
  assign n1893 = ( n30 & ~n174 ) | ( n30 & n1892 ) | ( ~n174 & n1892 ) ;
  buffer buf_n1894( .i (n29), .o (n1894) );
  assign n1895 = ( n1394 & ~n1892 ) | ( n1394 & n1894 ) | ( ~n1892 & n1894 ) ;
  assign n1896 = n1893 & ~n1895 ;
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  assign n1899 = n1704 & ~n1897 ;
  assign n1900 = ( n1886 & n1898 ) | ( n1886 & ~n1899 ) | ( n1898 & ~n1899 ) ;
  assign n1901 = n63 | n1900 ;
  assign n1902 = ( n1617 & ~n1625 ) | ( n1617 & n1889 ) | ( ~n1625 & n1889 ) ;
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1907( .i (n1906), .o (n1907) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1908( .i (n1617), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  assign n1910 = ( n1682 & n1903 ) | ( n1682 & ~n1909 ) | ( n1903 & ~n1909 ) ;
  assign n1911 = n1628 & n1910 ;
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n176( .i (n175), .o (n176) );
  assign n1914 = n176 & ~n1912 ;
  assign n1915 = ( n1907 & n1913 ) | ( n1907 & ~n1914 ) | ( n1913 & ~n1914 ) ;
  assign n1916 = ~n34 & n1915 ;
  assign n1917 = n63 & ~n1916 ;
  assign n1918 = n1901 & ~n1917 ;
  assign n1919 = n121 | n1918 ;
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  assign n1920 = ( n53 & n1741 ) | ( n53 & n1813 ) | ( n1741 & n1813 ) ;
  buffer buf_n1921( .i (n1920), .o (n1921) );
  assign n1926 = ( n1617 & ~n1640 ) | ( n1617 & n1921 ) | ( ~n1640 & n1921 ) ;
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  buffer buf_n1930( .i (n1929), .o (n1930) );
  assign n1931 = ( n1375 & n1517 ) | ( n1375 & n1927 ) | ( n1517 & n1927 ) ;
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  assign n1934 = n1925 & ~n1932 ;
  assign n1935 = ( n1930 & ~n1933 ) | ( n1930 & n1934 ) | ( ~n1933 & n1934 ) ;
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n825), .o (n1938) );
  assign n1939 = ~n1833 & n1938 ;
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  assign n1951 = n1936 | n1950 ;
  assign n1952 = ( n1221 & n1937 ) | ( n1221 & n1951 ) | ( n1937 & n1951 ) ;
  assign n1953 = ~n36 & n1952 ;
  assign n1954 = n121 & ~n1953 ;
  assign n1955 = n1919 & ~n1954 ;
  assign n1956 = ( n153 & ~n211 ) | ( n153 & n1955 ) | ( ~n211 & n1955 ) ;
  assign n1957 = ( ~n1444 & n1858 ) | ( ~n1444 & n1956 ) | ( n1858 & n1956 ) ;
  buffer buf_n177( .i (n176), .o (n177) );
  assign n1958 = ( n27 & ~n1371 ) | ( n27 & n1889 ) | ( ~n1371 & n1889 ) ;
  assign n1959 = ( ~n1346 & n1890 ) | ( ~n1346 & n1958 ) | ( n1890 & n1958 ) ;
  buffer buf_n1960( .i (n1959), .o (n1960) );
  assign n1963 = n174 & ~n1960 ;
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  assign n1966 = n1962 | n1964 ;
  assign n1967 = ( ~n177 & n1965 ) | ( ~n177 & n1966 ) | ( n1965 & n1966 ) ;
  assign n1968 = n90 | n1967 ;
  buffer buf_n1969( .i (n1822), .o (n1969) );
  assign n1970 = ( n1841 & n1888 ) | ( n1841 & ~n1969 ) | ( n1888 & ~n1969 ) ;
  buffer buf_n1971( .i (n1970), .o (n1971) );
  buffer buf_n1972( .i (n1971), .o (n1972) );
  buffer buf_n1973( .i (n1972), .o (n1973) );
  buffer buf_n1974( .i (n1973), .o (n1974) );
  assign n1975 = n203 | n1974 ;
  assign n1976 = ( ~n175 & n203 ) | ( ~n175 & n1974 ) | ( n203 & n1974 ) ;
  assign n1977 = ( n176 & ~n1975 ) | ( n176 & n1976 ) | ( ~n1975 & n1976 ) ;
  assign n1978 = ~n1704 & n1977 ;
  assign n1979 = n90 & ~n1978 ;
  assign n1980 = n1968 & ~n1979 ;
  assign n1981 = n64 | n1980 ;
  buffer buf_n1982( .i (n108), .o (n1982) );
  assign n1983 = ( ~n1741 & n1887 ) | ( ~n1741 & n1982 ) | ( n1887 & n1982 ) ;
  buffer buf_n1984( .i (n1983), .o (n1984) );
  assign n1989 = ( ~n1371 & n1743 ) | ( ~n1371 & n1984 ) | ( n1743 & n1984 ) ;
  buffer buf_n1990( .i (n1989), .o (n1990) );
  buffer buf_n1991( .i (n1990), .o (n1991) );
  buffer buf_n1992( .i (n1991), .o (n1992) );
  buffer buf_n1993( .i (n1992), .o (n1993) );
  buffer buf_n1994( .i (n1346), .o (n1994) );
  assign n1995 = ( n1652 & n1990 ) | ( n1652 & n1994 ) | ( n1990 & n1994 ) ;
  buffer buf_n1996( .i (n1995), .o (n1996) );
  buffer buf_n1997( .i (n1996), .o (n1997) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n1986( .i (n1985), .o (n1986) );
  buffer buf_n1987( .i (n1986), .o (n1987) );
  buffer buf_n1988( .i (n1987), .o (n1988) );
  assign n1998 = ~n1988 & n1996 ;
  assign n1999 = ( ~n1993 & n1997 ) | ( ~n1993 & n1998 ) | ( n1997 & n1998 ) ;
  assign n2000 = n205 & ~n1999 ;
  assign n2001 = ~n1491 & n1834 ;
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n2003), .o (n2004) );
  buffer buf_n2005( .i (n2004), .o (n2005) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n2007( .i (n2006), .o (n2007) );
  buffer buf_n2008( .i (n2007), .o (n2008) );
  buffer buf_n2012( .i (n1700), .o (n2012) );
  assign n2013 = ( ~n400 & n2008 ) | ( ~n400 & n2012 ) | ( n2008 & n2012 ) ;
  assign n2014 = n176 | n2013 ;
  buffer buf_n2015( .i (n204), .o (n2015) );
  assign n2016 = n2014 & ~n2015 ;
  assign n2017 = n2000 | n2016 ;
  assign n2018 = n1783 | n2017 ;
  assign n2019 = n64 & n2018 ;
  assign n2020 = n1981 & ~n2019 ;
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  assign n2023 = n359 & n2021 ;
  assign n2024 = ~n200 & n1775 ;
  buffer buf_n2025( .i (n1969), .o (n2025) );
  assign n2026 = ~n1081 & n2025 ;
  buffer buf_n2027( .i (n2026), .o (n2027) );
  assign n2028 = n2024 & n2027 ;
  assign n2029 = ~n191 & n1099 ;
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n2047( .i (n1162), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  assign n2049 = n2030 & ~n2048 ;
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  buffer buf_n2055( .i (n2054), .o (n2055) );
  assign n2057 = n196 & n867 ;
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  assign n2061 = n2055 | n2060 ;
  assign n2062 = ( ~n1083 & n2027 ) | ( ~n1083 & n2061 ) | ( n2027 & n2061 ) ;
  assign n2063 = ( n1394 & n2028 ) | ( n1394 & n2062 ) | ( n2028 & n2062 ) ;
  assign n2064 = n1392 & ~n2063 ;
  buffer buf_n2065( .i (n1099), .o (n2065) );
  assign n2066 = ( n1604 & n2047 ) | ( n1604 & ~n2065 ) | ( n2047 & ~n2065 ) ;
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n2073( .i (n2072), .o (n2073) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  assign n2075 = n1969 & ~n2071 ;
  buffer buf_n2076( .i (n2075), .o (n2076) );
  buffer buf_n2077( .i (n2076), .o (n2077) );
  assign n2078 = ( n200 & n1890 ) | ( n200 & n2076 ) | ( n1890 & n2076 ) ;
  assign n2079 = ( ~n2074 & n2077 ) | ( ~n2074 & n2078 ) | ( n2077 & n2078 ) ;
  buffer buf_n2080( .i (n1517), .o (n2080) );
  assign n2081 = n2079 & ~n2080 ;
  buffer buf_n2082( .i (n1376), .o (n2082) );
  assign n2083 = n2081 | n2082 ;
  assign n2084 = ~n2064 & n2083 ;
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  assign n2087 = ( n34 & ~n118 ) | ( n34 & n2085 ) | ( ~n118 & n2085 ) ;
  buffer buf_n2088( .i (n2065), .o (n2088) );
  assign n2089 = n193 | n2088 ;
  buffer buf_n2090( .i (n2089), .o (n2090) );
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n2099( .i (n2098), .o (n2099) );
  assign n2103 = ~n590 & n596 ;
  assign n2104 = ( n1486 & ~n2099 ) | ( n1486 & n2103 ) | ( ~n2099 & n2103 ) ;
  buffer buf_n2105( .i (n2082), .o (n2105) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  assign n2107 = n2104 & ~n2106 ;
  buffer buf_n2108( .i (n32), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  assign n2110 = n2107 & ~n2109 ;
  assign n2111 = ( n2086 & ~n2087 ) | ( n2086 & n2110 ) | ( ~n2087 & n2110 ) ;
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  assign n2114 = n192 & n2065 ;
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  buffer buf_n2119( .i (n2118), .o (n2119) );
  buffer buf_n2120( .i (n2119), .o (n2120) );
  buffer buf_n2121( .i (n2120), .o (n2121) );
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  assign n2129 = n717 & n2128 ;
  assign n2130 = n601 & n2129 ;
  buffer buf_n2131( .i (n195), .o (n2131) );
  assign n2132 = n919 & n2131 ;
  buffer buf_n2133( .i (n2132), .o (n2133) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  buffer buf_n2137( .i (n2136), .o (n2137) );
  buffer buf_n2138( .i (n2137), .o (n2138) );
  buffer buf_n2139( .i (n2138), .o (n2139) );
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n632( .i (n631), .o (n632) );
  assign n2143 = ~n44 & n160 ;
  buffer buf_n2144( .i (n2143), .o (n2144) );
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  assign n2158 = ( n632 & n1153 ) | ( n632 & ~n2151 ) | ( n1153 & ~n2151 ) ;
  assign n2159 = ( n1154 & ~n1742 ) | ( n1154 & n2158 ) | ( ~n1742 & n2158 ) ;
  assign n2160 = ~n2025 & n2159 ;
  assign n2161 = ~n28 & n2160 ;
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n2163( .i (n2162), .o (n2163) );
  buffer buf_n2164( .i (n2163), .o (n2164) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n2165( .i (n1994), .o (n2165) );
  assign n2166 = ( n800 & n2162 ) | ( n800 & ~n2165 ) | ( n2162 & ~n2165 ) ;
  assign n2167 = n1402 & ~n2166 ;
  assign n2168 = ( n1403 & n2164 ) | ( n1403 & ~n2167 ) | ( n2164 & ~n2167 ) ;
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  assign n2171 = ~n192 & n269 ;
  buffer buf_n2172( .i (n2171), .o (n2172) );
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n2175( .i (n2174), .o (n2175) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n2177), .o (n2178) );
  buffer buf_n2179( .i (n2178), .o (n2179) );
  buffer buf_n2180( .i (n2179), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  buffer buf_n2182( .i (n2181), .o (n2182) );
  buffer buf_n2183( .i (n2182), .o (n2183) );
  buffer buf_n2184( .i (n2183), .o (n2184) );
  assign n2185 = n2169 & n2184 ;
  assign n2186 = ( n2142 & n2170 ) | ( n2142 & n2185 ) | ( n2170 & n2185 ) ;
  assign n2187 = n162 | n190 ;
  buffer buf_n2188( .i (n2187), .o (n2188) );
  buffer buf_n2189( .i (n2188), .o (n2189) );
  buffer buf_n2190( .i (n2189), .o (n2190) );
  buffer buf_n2191( .i (n2190), .o (n2191) );
  buffer buf_n2192( .i (n2191), .o (n2192) );
  buffer buf_n2193( .i (n2192), .o (n2193) );
  buffer buf_n2194( .i (n2193), .o (n2194) );
  buffer buf_n2195( .i (n2194), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  buffer buf_n2197( .i (n2196), .o (n2197) );
  buffer buf_n2198( .i (n2197), .o (n2198) );
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n2200( .i (n2199), .o (n2200) );
  buffer buf_n2201( .i (n2200), .o (n2201) );
  assign n2203 = ( n195 & n1333 ) | ( n195 & n1834 ) | ( n1333 & n1834 ) ;
  assign n2204 = n1452 & n1557 ;
  buffer buf_n2205( .i (n2204), .o (n2205) );
  assign n2211 = ( ~n2131 & n2203 ) | ( ~n2131 & n2205 ) | ( n2203 & n2205 ) ;
  buffer buf_n2212( .i (n2211), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  assign n2214 = ( ~n72 & n188 ) | ( ~n72 & n218 ) | ( n188 & n218 ) ;
  buffer buf_n2215( .i (n2214), .o (n2215) );
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  assign n2219 = n74 & n2215 ;
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n2221( .i (n2220), .o (n2221) );
  assign n2222 = ( n192 & n2047 ) | ( n192 & ~n2220 ) | ( n2047 & ~n2220 ) ;
  assign n2223 = ( n2218 & n2221 ) | ( n2218 & ~n2222 ) | ( n2221 & ~n2222 ) ;
  assign n2224 = ( n1076 & ~n1452 ) | ( n1076 & n2223 ) | ( ~n1452 & n2223 ) ;
  buffer buf_n2225( .i (n159), .o (n2225) );
  buffer buf_n2226( .i (n187), .o (n2226) );
  assign n2227 = n2225 & n2226 ;
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  assign n2247 = n189 & ~n219 ;
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  assign n2259 = ( ~n1859 & n2230 ) | ( ~n1859 & n2249 ) | ( n2230 & n2249 ) ;
  assign n2260 = ( ~n1859 & n2065 ) | ( ~n1859 & n2230 ) | ( n2065 & n2230 ) ;
  assign n2261 = ( n2088 & n2259 ) | ( n2088 & ~n2260 ) | ( n2259 & ~n2260 ) ;
  buffer buf_n2262( .i (n1605), .o (n2262) );
  buffer buf_n2263( .i (n1451), .o (n2263) );
  assign n2264 = ( ~n2261 & n2262 ) | ( ~n2261 & n2263 ) | ( n2262 & n2263 ) ;
  assign n2265 = n2224 & ~n2264 ;
  buffer buf_n2266( .i (n2265), .o (n2266) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  assign n2269 = ( n227 & n1822 ) | ( n227 & ~n2266 ) | ( n1822 & ~n2266 ) ;
  assign n2270 = n2212 & n2269 ;
  assign n2271 = ( n2213 & n2268 ) | ( n2213 & ~n2270 ) | ( n2268 & ~n2270 ) ;
  assign n2272 = ( ~n28 & n1346 ) | ( ~n28 & n2271 ) | ( n1346 & n2271 ) ;
  buffer buf_n2273( .i (n218), .o (n2273) );
  assign n2274 = ( n161 & n247 ) | ( n161 & ~n2273 ) | ( n247 & ~n2273 ) ;
  buffer buf_n2275( .i (n2274), .o (n2275) );
  buffer buf_n2285( .i (n1114), .o (n2285) );
  assign n2286 = ( n75 & n2275 ) | ( n75 & n2285 ) | ( n2275 & n2285 ) ;
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n2289( .i (n2288), .o (n2289) );
  buffer buf_n2276( .i (n2275), .o (n2276) );
  buffer buf_n2277( .i (n2276), .o (n2277) );
  buffer buf_n2278( .i (n2277), .o (n2278) );
  assign n2290 = ( n1451 & n2088 ) | ( n1451 & ~n2287 ) | ( n2088 & ~n2287 ) ;
  assign n2291 = n2278 & n2290 ;
  assign n2292 = ( n1834 & ~n2289 ) | ( n1834 & n2291 ) | ( ~n2289 & n2291 ) ;
  assign n2293 = n2131 | n2292 ;
  assign n2294 = ~n246 & n2225 ;
  buffer buf_n2295( .i (n2294), .o (n2295) );
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n2297( .i (n2296), .o (n2297) );
  assign n2305 = ( n448 & ~n2047 ) | ( n448 & n2297 ) | ( ~n2047 & n2297 ) ;
  buffer buf_n2306( .i (n2305), .o (n2306) );
  assign n2321 = n1525 & n2306 ;
  buffer buf_n2322( .i (n1833), .o (n2322) );
  assign n2323 = n2321 & n2322 ;
  assign n2324 = n2131 & ~n2323 ;
  assign n2325 = n2293 & ~n2324 ;
  assign n2326 = n1969 | n2325 ;
  buffer buf_n2327( .i (n161), .o (n2327) );
  buffer buf_n2328( .i (n189), .o (n2328) );
  assign n2329 = ( ~n1115 & n2327 ) | ( ~n1115 & n2328 ) | ( n2327 & n2328 ) ;
  buffer buf_n2330( .i (n2329), .o (n2330) );
  buffer buf_n2334( .i (n1162), .o (n2334) );
  assign n2335 = ( n1859 & n2330 ) | ( n1859 & ~n2334 ) | ( n2330 & ~n2334 ) ;
  buffer buf_n2336( .i (n2335), .o (n2336) );
  buffer buf_n2337( .i (n2336), .o (n2337) );
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2331( .i (n2330), .o (n2331) );
  buffer buf_n2332( .i (n2331), .o (n2332) );
  buffer buf_n2333( .i (n2332), .o (n2333) );
  assign n2339 = ( n1557 & n2263 ) | ( n1557 & n2336 ) | ( n2263 & n2336 ) ;
  assign n2340 = n2333 & ~n2339 ;
  assign n2341 = ( n1835 & ~n2338 ) | ( n1835 & n2340 ) | ( ~n2338 & n2340 ) ;
  buffer buf_n2342( .i (n1622), .o (n2342) );
  assign n2343 = n2341 & n2342 ;
  buffer buf_n2344( .i (n1822), .o (n2344) );
  assign n2345 = ~n2343 & n2344 ;
  assign n2346 = n2326 & ~n2345 ;
  buffer buf_n2347( .i (n111), .o (n2347) );
  assign n2348 = ( n28 & ~n2346 ) | ( n28 & n2347 ) | ( ~n2346 & n2347 ) ;
  assign n2349 = n2272 & ~n2348 ;
  buffer buf_n2350( .i (n2349), .o (n2350) );
  buffer buf_n2351( .i (n2350), .o (n2351) );
  buffer buf_n2352( .i (n2351), .o (n2352) );
  assign n2353 = n684 | n1835 ;
  buffer buf_n2354( .i (n2353), .o (n2354) );
  buffer buf_n2355( .i (n2354), .o (n2355) );
  buffer buf_n2356( .i (n2355), .o (n2356) );
  buffer buf_n2357( .i (n2356), .o (n2357) );
  buffer buf_n2358( .i (n2357), .o (n2358) );
  assign n2359 = n1894 & ~n2358 ;
  assign n2360 = ( n926 & n2350 ) | ( n926 & n2359 ) | ( n2350 & n2359 ) ;
  assign n2361 = n2200 | n2360 ;
  assign n2362 = ( ~n2201 & n2352 ) | ( ~n2201 & n2361 ) | ( n2352 & n2361 ) ;
  buffer buf_n2363( .i (n2106), .o (n2363) );
  assign n2364 = n2362 | n2363 ;
  assign n2365 = ( n133 & n191 ) | ( n133 & ~n1162 ) | ( n191 & ~n1162 ) ;
  buffer buf_n2366( .i (n2365), .o (n2366) );
  assign n2372 = ( n2048 & ~n2088 ) | ( n2048 & n2366 ) | ( ~n2088 & n2366 ) ;
  buffer buf_n2373( .i (n2372), .o (n2373) );
  buffer buf_n2374( .i (n2373), .o (n2374) );
  buffer buf_n2375( .i (n2374), .o (n2375) );
  buffer buf_n2376( .i (n2375), .o (n2376) );
  buffer buf_n2377( .i (n193), .o (n2377) );
  buffer buf_n2378( .i (n2377), .o (n2378) );
  assign n2379 = ( n1491 & n2373 ) | ( n1491 & n2378 ) | ( n2373 & n2378 ) ;
  buffer buf_n2380( .i (n2379), .o (n2380) );
  buffer buf_n2381( .i (n2380), .o (n2381) );
  buffer buf_n2367( .i (n2366), .o (n2367) );
  buffer buf_n2368( .i (n2367), .o (n2368) );
  buffer buf_n2369( .i (n2368), .o (n2369) );
  buffer buf_n2370( .i (n2369), .o (n2370) );
  assign n2382 = n2370 & ~n2380 ;
  assign n2383 = ( n2376 & ~n2381 ) | ( n2376 & n2382 ) | ( ~n2381 & n2382 ) ;
  buffer buf_n2384( .i (n1841), .o (n2384) );
  assign n2385 = n2383 & n2384 ;
  buffer buf_n2386( .i (n132), .o (n2386) );
  buffer buf_n2387( .i (n2386), .o (n2387) );
  buffer buf_n2388( .i (n191), .o (n2388) );
  assign n2389 = ( n2334 & n2387 ) | ( n2334 & n2388 ) | ( n2387 & n2388 ) ;
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2391( .i (n2390), .o (n2391) );
  buffer buf_n2392( .i (n2391), .o (n2392) );
  buffer buf_n2393( .i (n2392), .o (n2393) );
  buffer buf_n2394( .i (n2393), .o (n2394) );
  buffer buf_n2231( .i (n2230), .o (n2231) );
  buffer buf_n2232( .i (n2231), .o (n2232) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  buffer buf_n2235( .i (n2234), .o (n2235) );
  buffer buf_n2395( .i (n2262), .o (n2395) );
  buffer buf_n2396( .i (n2395), .o (n2396) );
  buffer buf_n2397( .i (n2396), .o (n2397) );
  assign n2398 = ( n2235 & ~n2342 ) | ( n2235 & n2397 ) | ( ~n2342 & n2397 ) ;
  assign n2399 = n2394 & ~n2398 ;
  assign n2400 = n2384 | n2399 ;
  assign n2401 = ( ~n2347 & n2385 ) | ( ~n2347 & n2400 ) | ( n2385 & n2400 ) ;
  assign n2402 = n1682 | n2401 ;
  buffer buf_n2403( .i (n2285), .o (n2403) );
  buffer buf_n2404( .i (n2403), .o (n2404) );
  buffer buf_n2405( .i (n2404), .o (n2405) );
  assign n2406 = ( n2377 & ~n2390 ) | ( n2377 & n2405 ) | ( ~n2390 & n2405 ) ;
  buffer buf_n2407( .i (n2406), .o (n2407) );
  buffer buf_n2408( .i (n2407), .o (n2408) );
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  assign n2411 = ( n1674 & n2396 ) | ( n1674 & ~n2407 ) | ( n2396 & ~n2407 ) ;
  buffer buf_n2412( .i (n2411), .o (n2412) );
  buffer buf_n2413( .i (n2412), .o (n2413) );
  assign n2414 = ~n2394 & n2412 ;
  assign n2415 = ( n2410 & n2413 ) | ( n2410 & n2414 ) | ( n2413 & n2414 ) ;
  assign n2416 = ~n2347 & n2415 ;
  buffer buf_n2417( .i (n1813), .o (n2417) );
  buffer buf_n2418( .i (n2417), .o (n2418) );
  buffer buf_n2419( .i (n2418), .o (n2419) );
  buffer buf_n2420( .i (n2419), .o (n2420) );
  assign n2421 = ~n2416 & n2420 ;
  assign n2422 = n2402 & ~n2421 ;
  assign n2423 = n1056 & n1743 ;
  buffer buf_n2424( .i (n2423), .o (n2424) );
  assign n2429 = n288 & ~n2354 ;
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  assign n2432 = n1307 | n2430 ;
  assign n2433 = ( n2424 & n2431 ) | ( n2424 & n2432 ) | ( n2431 & n2432 ) ;
  buffer buf_n2434( .i (n2433), .o (n2434) );
  assign n2435 = ( n87 & n2422 ) | ( n87 & n2434 ) | ( n2422 & n2434 ) ;
  buffer buf_n2436( .i (n855), .o (n2436) );
  assign n2437 = ( n2387 & n2388 ) | ( n2387 & ~n2436 ) | ( n2388 & ~n2436 ) ;
  buffer buf_n2438( .i (n2437), .o (n2438) );
  assign n2443 = ( n2262 & n2405 ) | ( n2262 & ~n2438 ) | ( n2405 & ~n2438 ) ;
  buffer buf_n2444( .i (n2443), .o (n2444) );
  buffer buf_n2445( .i (n2444), .o (n2445) );
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n2448( .i (n2378), .o (n2448) );
  assign n2449 = ( n108 & n2444 ) | ( n108 & ~n2448 ) | ( n2444 & ~n2448 ) ;
  buffer buf_n2450( .i (n2449), .o (n2450) );
  buffer buf_n2451( .i (n2450), .o (n2451) );
  buffer buf_n2439( .i (n2438), .o (n2439) );
  buffer buf_n2440( .i (n2439), .o (n2440) );
  buffer buf_n2441( .i (n2440), .o (n2441) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  assign n2452 = n2442 & n2450 ;
  assign n2453 = ( ~n2447 & n2451 ) | ( ~n2447 & n2452 ) | ( n2451 & n2452 ) ;
  assign n2454 = n2419 | n2453 ;
  assign n2455 = ( n561 & n1982 ) | ( n561 & n2342 ) | ( n1982 & n2342 ) ;
  assign n2456 = ( n561 & ~n1982 ) | ( n561 & n2342 ) | ( ~n1982 & n2342 ) ;
  assign n2457 = ( n1841 & ~n2455 ) | ( n1841 & n2456 ) | ( ~n2455 & n2456 ) ;
  assign n2458 = n199 & n2457 ;
  assign n2459 = n2419 & ~n2458 ;
  assign n2460 = n2454 & ~n2459 ;
  assign n2461 = n1556 & ~n1557 ;
  buffer buf_n2462( .i (n2461), .o (n2462) );
  buffer buf_n2463( .i (n2462), .o (n2463) );
  buffer buf_n2464( .i (n2463), .o (n2464) );
  assign n2470 = ( n2176 & n2344 ) | ( n2176 & n2464 ) | ( n2344 & n2464 ) ;
  assign n2471 = ~n2025 & n2470 ;
  buffer buf_n2472( .i (n2471), .o (n2472) );
  buffer buf_n2473( .i (n2472), .o (n2473) );
  assign n2474 = n1652 | n2472 ;
  assign n2475 = ( n2460 & n2473 ) | ( n2460 & n2474 ) | ( n2473 & n2474 ) ;
  buffer buf_n2476( .i (n2080), .o (n2476) );
  assign n2477 = ( n2434 & n2475 ) | ( n2434 & ~n2476 ) | ( n2475 & ~n2476 ) ;
  assign n2478 = n2435 | n2477 ;
  assign n2479 = ~n2108 & n2478 ;
  assign n2480 = n2363 & ~n2479 ;
  assign n2481 = n2364 & ~n2480 ;
  assign n2482 = n2186 | n2481 ;
  assign n2483 = ( ~n2112 & n2130 ) | ( ~n2112 & n2482 ) | ( n2130 & n2482 ) ;
  assign n2484 = n2113 | n2483 ;
  assign n2485 = ( n200 & n1516 ) | ( n200 & ~n2419 ) | ( n1516 & ~n2419 ) ;
  buffer buf_n2486( .i (n2485), .o (n2486) );
  assign n2487 = ( n1700 & ~n2080 ) | ( n1700 & n2486 ) | ( ~n2080 & n2486 ) ;
  assign n2488 = ( n260 & ~n1700 ) | ( n260 & n2486 ) | ( ~n1700 & n2486 ) ;
  assign n2489 = n2487 & n2488 ;
  buffer buf_n2490( .i (n2489), .o (n2490) );
  buffer buf_n2491( .i (n2490), .o (n2491) );
  assign n2492 = ~n1451 & n1605 ;
  buffer buf_n2493( .i (n2492), .o (n2493) );
  assign n2501 = ( n23 & n2322 ) | ( n23 & n2493 ) | ( n2322 & n2493 ) ;
  buffer buf_n2502( .i (n2501), .o (n2502) );
  buffer buf_n2503( .i (n2502), .o (n2503) );
  buffer buf_n2504( .i (n2503), .o (n2504) );
  buffer buf_n2505( .i (n1835), .o (n2505) );
  assign n2506 = ( n2397 & ~n2502 ) | ( n2397 & n2505 ) | ( ~n2502 & n2505 ) ;
  buffer buf_n2507( .i (n25), .o (n2507) );
  assign n2508 = ( ~n2417 & n2506 ) | ( ~n2417 & n2507 ) | ( n2506 & n2507 ) ;
  assign n2509 = ~n2504 & n2508 ;
  buffer buf_n2510( .i (n2509), .o (n2510) );
  buffer buf_n2511( .i (n2510), .o (n2511) );
  buffer buf_n2512( .i (n1890), .o (n2512) );
  assign n2513 = ( n201 & n2510 ) | ( n201 & ~n2512 ) | ( n2510 & ~n2512 ) ;
  buffer buf_n2514( .i (n2048), .o (n2514) );
  assign n2515 = n2263 & ~n2514 ;
  buffer buf_n2516( .i (n2515), .o (n2516) );
  buffer buf_n2517( .i (n2516), .o (n2517) );
  buffer buf_n2518( .i (n2517), .o (n2518) );
  assign n2523 = n2344 & n2518 ;
  buffer buf_n2524( .i (n2507), .o (n2524) );
  assign n2525 = ( n1743 & n2523 ) | ( n1743 & n2524 ) | ( n2523 & n2524 ) ;
  buffer buf_n2526( .i (n2524), .o (n2526) );
  assign n2527 = n2525 & ~n2526 ;
  assign n2528 = ~n201 & n2527 ;
  assign n2529 = ( n2511 & ~n2513 ) | ( n2511 & n2528 ) | ( ~n2513 & n2528 ) ;
  buffer buf_n2530( .i (n2529), .o (n2530) );
  buffer buf_n2531( .i (n2530), .o (n2531) );
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n408), .o (n2533) );
  buffer buf_n2534( .i (n174), .o (n2534) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  assign n2536 = ( ~n2530 & n2533 ) | ( ~n2530 & n2535 ) | ( n2533 & n2535 ) ;
  assign n2537 = n2490 & n2536 ;
  assign n2538 = ( n2491 & n2532 ) | ( n2491 & ~n2537 ) | ( n2532 & ~n2537 ) ;
  assign n2539 = n119 | n2538 ;
  buffer buf_n2540( .i (n2388), .o (n2540) );
  assign n2541 = ( ~n1832 & n2048 ) | ( ~n1832 & n2540 ) | ( n2048 & n2540 ) ;
  buffer buf_n2542( .i (n2541), .o (n2542) );
  buffer buf_n2543( .i (n2542), .o (n2543) );
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  buffer buf_n2551( .i (n1742), .o (n2551) );
  assign n2552 = ( n2025 & n2546 ) | ( n2025 & n2551 ) | ( n2546 & n2551 ) ;
  buffer buf_n2553( .i (n2552), .o (n2553) );
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2555( .i (n2554), .o (n2555) );
  buffer buf_n2556( .i (n2555), .o (n2556) );
  buffer buf_n2557( .i (n199), .o (n2557) );
  buffer buf_n2558( .i (n2557), .o (n2558) );
  assign n2559 = ( n2512 & n2553 ) | ( n2512 & n2558 ) | ( n2553 & n2558 ) ;
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  assign n2562 = n2550 & ~n2560 ;
  assign n2563 = ( n2556 & ~n2561 ) | ( n2556 & n2562 ) | ( ~n2561 & n2562 ) ;
  assign n2564 = ~n263 & n2563 ;
  assign n2565 = ~n2109 & n2564 ;
  assign n2566 = n119 & ~n2565 ;
  assign n2567 = n2539 & ~n2566 ;
  assign n2568 = n65 | n2567 ;
  buffer buf_n178( .i (n177), .o (n178) );
  assign n2569 = n1742 & ~n2417 ;
  buffer buf_n2570( .i (n2569), .o (n2570) );
  buffer buf_n2573( .i (n2551), .o (n2573) );
  assign n2574 = ~n2570 & n2573 ;
  buffer buf_n2575( .i (n2574), .o (n2575) );
  buffer buf_n2576( .i (n1699), .o (n2576) );
  assign n2577 = n2575 & n2576 ;
  buffer buf_n2571( .i (n2570), .o (n2571) );
  buffer buf_n2572( .i (n2571), .o (n2572) );
  assign n2578 = ( n202 & ~n2572 ) | ( n202 & n2575 ) | ( ~n2572 & n2575 ) ;
  assign n2579 = ( ~n261 & n2577 ) | ( ~n261 & n2578 ) | ( n2577 & n2578 ) ;
  assign n2580 = n1648 & n2579 ;
  buffer buf_n2581( .i (n131), .o (n2581) );
  assign n2582 = ( n74 & n1115 ) | ( n74 & n2581 ) | ( n1115 & n2581 ) ;
  buffer buf_n2583( .i (n2582), .o (n2583) );
  buffer buf_n2584( .i (n2583), .o (n2584) );
  buffer buf_n2585( .i (n2584), .o (n2585) );
  buffer buf_n2586( .i (n2585), .o (n2586) );
  buffer buf_n2587( .i (n2586), .o (n2587) );
  buffer buf_n2588( .i (n2587), .o (n2588) );
  buffer buf_n2589( .i (n2588), .o (n2589) );
  assign n2590 = ( ~n198 & n2344 ) | ( ~n198 & n2589 ) | ( n2344 & n2589 ) ;
  buffer buf_n2591( .i (n2590), .o (n2591) );
  buffer buf_n2594( .i (n2397), .o (n2594) );
  buffer buf_n2595( .i (n2594), .o (n2595) );
  buffer buf_n2596( .i (n2595), .o (n2596) );
  assign n2597 = ~n2591 & n2596 ;
  buffer buf_n2598( .i (n2597), .o (n2598) );
  buffer buf_n2599( .i (n2598), .o (n2599) );
  buffer buf_n2592( .i (n2591), .o (n2592) );
  buffer buf_n2593( .i (n2592), .o (n2593) );
  assign n2600 = n2593 | n2598 ;
  assign n2601 = ( ~n2012 & n2599 ) | ( ~n2012 & n2600 ) | ( n2599 & n2600 ) ;
  assign n2602 = n1648 | n2601 ;
  assign n2603 = ( ~n1021 & n2580 ) | ( ~n1021 & n2602 ) | ( n2580 & n2602 ) ;
  assign n2604 = n178 | n2603 ;
  buffer buf_n2425( .i (n2424), .o (n2425) );
  buffer buf_n2426( .i (n2425), .o (n2426) );
  buffer buf_n2427( .i (n2426), .o (n2427) );
  buffer buf_n2428( .i (n2427), .o (n2428) );
  assign n2605 = ~n2263 & n2377 ;
  buffer buf_n2606( .i (n2605), .o (n2606) );
  buffer buf_n2607( .i (n2606), .o (n2607) );
  buffer buf_n2608( .i (n2607), .o (n2608) );
  buffer buf_n2609( .i (n2608), .o (n2609) );
  buffer buf_n2610( .i (n2609), .o (n2610) );
  buffer buf_n2611( .i (n2610), .o (n2611) );
  buffer buf_n2612( .i (n2611), .o (n2612) );
  buffer buf_n2613( .i (n2612), .o (n2613) );
  buffer buf_n2614( .i (n2613), .o (n2614) );
  buffer buf_n2615( .i (n2614), .o (n2615) );
  assign n2616 = n2428 & n2615 ;
  assign n2617 = n178 & ~n2616 ;
  assign n2618 = n2604 & ~n2617 ;
  buffer buf_n2619( .i (n1783), .o (n2619) );
  assign n2620 = n2618 & ~n2619 ;
  assign n2621 = n65 & ~n2620 ;
  assign n2622 = n2568 & ~n2621 ;
  assign n2623 = n2484 | n2622 ;
  assign n2624 = ( n2022 & ~n2023 ) | ( n2022 & n2623 ) | ( ~n2023 & n2623 ) ;
  buffer buf_n2625( .i (n2334), .o (n2625) );
  assign n2626 = n2404 & n2625 ;
  buffer buf_n2627( .i (n2626), .o (n2627) );
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  buffer buf_n2631( .i (n2630), .o (n2631) );
  buffer buf_n2632( .i (n2631), .o (n2632) );
  buffer buf_n2633( .i (n2632), .o (n2633) );
  buffer buf_n2634( .i (n2633), .o (n2634) );
  buffer buf_n2635( .i (n2634), .o (n2635) );
  buffer buf_n2636( .i (n2635), .o (n2636) );
  buffer buf_n2637( .i (n2636), .o (n2637) );
  assign n2638 = ( ~n177 & n402 ) | ( ~n177 & n2637 ) | ( n402 & n2637 ) ;
  assign n2639 = ~n2363 & n2638 ;
  buffer buf_n2640( .i (n90), .o (n2640) );
  assign n2641 = n2639 & ~n2640 ;
  assign n2642 = n2619 & n2641 ;
  buffer buf_n2643( .i (n54), .o (n2643) );
  buffer buf_n2644( .i (n1616), .o (n2644) );
  assign n2645 = ( n2551 & ~n2643 ) | ( n2551 & n2644 ) | ( ~n2643 & n2644 ) ;
  buffer buf_n2646( .i (n2645), .o (n2646) );
  buffer buf_n2647( .i (n2646), .o (n2647) );
  buffer buf_n2648( .i (n2647), .o (n2648) );
  buffer buf_n2649( .i (n2648), .o (n2649) );
  buffer buf_n2650( .i (n2573), .o (n2650) );
  assign n2651 = n2646 & ~n2650 ;
  buffer buf_n2652( .i (n2651), .o (n2652) );
  buffer buf_n2653( .i (n2652), .o (n2653) );
  assign n2654 = ( n2082 & ~n2534 ) | ( n2082 & n2652 ) | ( ~n2534 & n2652 ) ;
  assign n2655 = ( n2649 & n2653 ) | ( n2649 & n2654 ) | ( n2653 & n2654 ) ;
  assign n2656 = ( n147 & ~n1021 ) | ( n147 & n2655 ) | ( ~n1021 & n2655 ) ;
  assign n2657 = ( n1889 & ~n2551 ) | ( n1889 & n2643 ) | ( ~n2551 & n2643 ) ;
  buffer buf_n2658( .i (n2657), .o (n2658) );
  buffer buf_n2659( .i (n2658), .o (n2659) );
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2660), .o (n2661) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  assign n2662 = n477 & ~n2658 ;
  buffer buf_n2663( .i (n2662), .o (n2663) );
  buffer buf_n2664( .i (n2663), .o (n2664) );
  assign n2665 = n233 & ~n2663 ;
  assign n2666 = ( n2661 & n2664 ) | ( n2661 & ~n2665 ) | ( n2664 & ~n2665 ) ;
  assign n2667 = ( n147 & n1021 ) | ( n147 & n2666 ) | ( n1021 & n2666 ) ;
  assign n2668 = n2656 & ~n2667 ;
  assign n2669 = ( ~n793 & n866 ) | ( ~n793 & n1188 ) | ( n866 & n1188 ) ;
  buffer buf_n2670( .i (n2669), .o (n2670) );
  buffer buf_n2671( .i (n2670), .o (n2671) );
  buffer buf_n2672( .i (n2671), .o (n2672) );
  buffer buf_n2673( .i (n2672), .o (n2673) );
  buffer buf_n2674( .i (n2673), .o (n2674) );
  buffer buf_n2675( .i (n2674), .o (n2675) );
  buffer buf_n2676( .i (n2675), .o (n2676) );
  buffer buf_n2685( .i (n2165), .o (n2685) );
  assign n2686 = ( n2476 & ~n2676 ) | ( n2476 & n2685 ) | ( ~n2676 & n2685 ) ;
  buffer buf_n2687( .i (n2686), .o (n2687) );
  buffer buf_n2688( .i (n2685), .o (n2688) );
  buffer buf_n2689( .i (n2688), .o (n2689) );
  assign n2690 = ( n2106 & n2687 ) | ( n2106 & ~n2689 ) | ( n2687 & ~n2689 ) ;
  assign n2691 = ( n89 & n2106 ) | ( n89 & ~n2687 ) | ( n2106 & ~n2687 ) ;
  assign n2692 = n2690 & ~n2691 ;
  assign n2693 = n2668 | n2692 ;
  assign n2694 = ~n2619 & n2693 ;
  assign n2695 = n2642 | n2694 ;
  buffer buf_n2696( .i (n2695), .o (n2696) );
  buffer buf_n2697( .i (n2696), .o (n2697) );
  assign n2698 = ( n1752 & ~n2448 ) | ( n1752 & n2606 ) | ( ~n2448 & n2606 ) ;
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n2700( .i (n2699), .o (n2700) );
  buffer buf_n2701( .i (n2700), .o (n2701) );
  buffer buf_n2702( .i (n2701), .o (n2702) );
  buffer buf_n2703( .i (n2702), .o (n2703) );
  buffer buf_n2704( .i (n2703), .o (n2704) );
  buffer buf_n2705( .i (n2704), .o (n2705) );
  buffer buf_n2706( .i (n2705), .o (n2706) );
  buffer buf_n2707( .i (n2706), .o (n2707) );
  buffer buf_n2708( .i (n2707), .o (n2708) );
  buffer buf_n2709( .i (n2708), .o (n2709) );
  buffer buf_n2710( .i (n2709), .o (n2710) );
  buffer buf_n2711( .i (n2710), .o (n2711) );
  buffer buf_n2712( .i (n2711), .o (n2712) );
  assign n2714 = n2696 & n2712 ;
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n2715( .i (n2514), .o (n2715) );
  assign n2716 = n2395 | n2715 ;
  buffer buf_n2717( .i (n2716), .o (n2717) );
  buffer buf_n2718( .i (n2717), .o (n2718) );
  buffer buf_n2719( .i (n2718), .o (n2719) );
  buffer buf_n2720( .i (n2719), .o (n2720) );
  buffer buf_n2721( .i (n2720), .o (n2721) );
  assign n2726 = ( n1994 & n2650 ) | ( n1994 & n2721 ) | ( n2650 & n2721 ) ;
  assign n2727 = ( n1982 & n2505 ) | ( n1982 & ~n2717 ) | ( n2505 & ~n2717 ) ;
  buffer buf_n2728( .i (n2727), .o (n2728) );
  buffer buf_n2729( .i (n2728), .o (n2729) );
  buffer buf_n2730( .i (n2729), .o (n2730) );
  assign n2731 = ( n1699 & n2512 ) | ( n1699 & n2730 ) | ( n2512 & n2730 ) ;
  assign n2732 = n2726 & ~n2731 ;
  assign n2733 = n2082 & n2732 ;
  buffer buf_n2734( .i (n1888), .o (n2734) );
  buffer buf_n2735( .i (n2734), .o (n2735) );
  assign n2736 = n2573 | n2735 ;
  buffer buf_n2737( .i (n2736), .o (n2737) );
  assign n2738 = ( n566 & n2080 ) | ( n566 & ~n2737 ) | ( n2080 & ~n2737 ) ;
  buffer buf_n2739( .i (n1375), .o (n2739) );
  buffer buf_n2740( .i (n2739), .o (n2740) );
  assign n2741 = n2738 | n2740 ;
  assign n2742 = ( ~n2105 & n2733 ) | ( ~n2105 & n2741 ) | ( n2733 & n2741 ) ;
  assign n2743 = ( n235 & ~n2108 ) | ( n235 & n2742 ) | ( ~n2108 & n2742 ) ;
  buffer buf_n2744( .i (n2505), .o (n2744) );
  buffer buf_n2745( .i (n2744), .o (n2745) );
  assign n2746 = n442 | n2745 ;
  buffer buf_n2747( .i (n2746), .o (n2747) );
  buffer buf_n2748( .i (n2747), .o (n2748) );
  assign n2749 = ( n443 & n2573 ) | ( n443 & ~n2596 ) | ( n2573 & ~n2596 ) ;
  assign n2750 = n2747 & ~n2749 ;
  buffer buf_n2751( .i (n2650), .o (n2751) );
  assign n2752 = ( n2748 & n2750 ) | ( n2748 & ~n2751 ) | ( n2750 & ~n2751 ) ;
  assign n2753 = n2740 | n2752 ;
  assign n2754 = n807 & n2751 ;
  assign n2755 = n2740 & ~n2754 ;
  assign n2756 = n2753 & ~n2755 ;
  buffer buf_n2757( .i (n234), .o (n2757) );
  assign n2758 = ( n2108 & ~n2756 ) | ( n2108 & n2757 ) | ( ~n2756 & n2757 ) ;
  assign n2759 = n2743 & ~n2758 ;
  assign n2760 = ~n2387 & n2403 ;
  buffer buf_n2761( .i (n2760), .o (n2761) );
  buffer buf_n2762( .i (n2761), .o (n2762) );
  buffer buf_n2763( .i (n2762), .o (n2763) );
  buffer buf_n2764( .i (n2763), .o (n2764) );
  buffer buf_n2765( .i (n2764), .o (n2765) );
  buffer buf_n2766( .i (n2765), .o (n2766) );
  buffer buf_n2767( .i (n2766), .o (n2767) );
  buffer buf_n2768( .i (n2767), .o (n2768) );
  buffer buf_n2769( .i (n2768), .o (n2769) );
  buffer buf_n2770( .i (n2769), .o (n2770) );
  buffer buf_n2771( .i (n2770), .o (n2771) );
  buffer buf_n2772( .i (n2771), .o (n2772) );
  buffer buf_n2773( .i (n2772), .o (n2773) );
  assign n2774 = n1888 & n2744 ;
  buffer buf_n2775( .i (n2774), .o (n2775) );
  buffer buf_n2776( .i (n2775), .o (n2776) );
  assign n2777 = ( ~n728 & n1994 ) | ( ~n728 & n2776 ) | ( n1994 & n2776 ) ;
  assign n2778 = n729 & n2777 ;
  buffer buf_n2779( .i (n1556), .o (n2779) );
  buffer buf_n2780( .i (n2779), .o (n2780) );
  buffer buf_n2781( .i (n2780), .o (n2781) );
  assign n2782 = n701 & ~n2781 ;
  buffer buf_n2783( .i (n2782), .o (n2783) );
  buffer buf_n2784( .i (n2783), .o (n2784) );
  buffer buf_n2785( .i (n2784), .o (n2785) );
  assign n2786 = ( ~n2512 & n2650 ) | ( ~n2512 & n2785 ) | ( n2650 & n2785 ) ;
  assign n2787 = ~n2751 & n2786 ;
  assign n2788 = n2778 | n2787 ;
  buffer buf_n2789( .i (n2788), .o (n2789) );
  buffer buf_n2790( .i (n2789), .o (n2790) );
  buffer buf_n2791( .i (n1548), .o (n2791) );
  assign n2792 = ( n2757 & n2789 ) | ( n2757 & ~n2791 ) | ( n2789 & ~n2791 ) ;
  assign n2793 = ( n2773 & n2790 ) | ( n2773 & ~n2792 ) | ( n2790 & ~n2792 ) ;
  assign n2794 = n2759 | n2793 ;
  buffer buf_n2795( .i (n2794), .o (n2795) );
  buffer buf_n2796( .i (n2795), .o (n2796) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  assign n2797 = ( ~n209 & n267 ) | ( ~n209 & n2795 ) | ( n267 & n2795 ) ;
  assign n2798 = ( n504 & n2796 ) | ( n504 & ~n2797 ) | ( n2796 & ~n2797 ) ;
  assign n2799 = ( n1556 & n1833 ) | ( n1556 & n2405 ) | ( n1833 & n2405 ) ;
  buffer buf_n2800( .i (n2799), .o (n2800) );
  buffer buf_n2806( .i (n2715), .o (n2806) );
  assign n2807 = ( n1622 & n2800 ) | ( n1622 & ~n2806 ) | ( n2800 & ~n2806 ) ;
  buffer buf_n2808( .i (n2807), .o (n2808) );
  assign n2812 = n1616 & ~n2808 ;
  buffer buf_n2813( .i (n2812), .o (n2813) );
  buffer buf_n2814( .i (n2813), .o (n2814) );
  buffer buf_n2809( .i (n2808), .o (n2809) );
  buffer buf_n2810( .i (n2809), .o (n2810) );
  assign n2815 = n2810 | n2813 ;
  assign n2816 = ( ~n1909 & n2814 ) | ( ~n1909 & n2815 ) | ( n2814 & n2815 ) ;
  buffer buf_n2817( .i (n2816), .o (n2817) );
  buffer buf_n2818( .i (n2817), .o (n2818) );
  assign n2819 = ( n203 & n2740 ) | ( n203 & ~n2817 ) | ( n2740 & ~n2817 ) ;
  buffer buf_n2820( .i (n2347), .o (n2820) );
  assign n2821 = n539 & n2820 ;
  assign n2822 = ~n1508 & n2821 ;
  buffer buf_n2823( .i (n202), .o (n2823) );
  assign n2824 = n2822 & n2823 ;
  assign n2825 = ( n2818 & n2819 ) | ( n2818 & n2824 ) | ( n2819 & n2824 ) ;
  buffer buf_n2826( .i (n2825), .o (n2826) );
  buffer buf_n2827( .i (n2826), .o (n2827) );
  assign n2828 = n2199 | n2685 ;
  assign n2829 = ( n88 & n2105 ) | ( n88 & ~n2828 ) | ( n2105 & ~n2828 ) ;
  buffer buf_n2830( .i (n2105), .o (n2830) );
  assign n2831 = n2829 & ~n2830 ;
  assign n2832 = ~n2091 & n2806 ;
  buffer buf_n2833( .i (n2832), .o (n2833) );
  buffer buf_n2834( .i (n2833), .o (n2834) );
  buffer buf_n2835( .i (n2834), .o (n2835) );
  assign n2838 = ~n73 & n161 ;
  buffer buf_n2839( .i (n2838), .o (n2839) );
  assign n2848 = ( ~n855 & n2386 ) | ( ~n855 & n2839 ) | ( n2386 & n2839 ) ;
  buffer buf_n2849( .i (n2848), .o (n2849) );
  buffer buf_n2850( .i (n2849), .o (n2850) );
  buffer buf_n2851( .i (n2850), .o (n2851) );
  assign n2852 = ( n935 & n1832 ) | ( n935 & n2849 ) | ( n1832 & n2849 ) ;
  assign n2853 = ( n2262 & n2514 ) | ( n2262 & ~n2852 ) | ( n2514 & ~n2852 ) ;
  assign n2854 = ~n2851 & n2853 ;
  assign n2855 = n1147 & n2386 ;
  buffer buf_n2856( .i (n2855), .o (n2856) );
  assign n2863 = n994 & n2856 ;
  buffer buf_n2864( .i (n2863), .o (n2864) );
  buffer buf_n2865( .i (n2864), .o (n2865) );
  assign n2866 = n1621 & ~n2864 ;
  assign n2867 = ( n2854 & n2865 ) | ( n2854 & ~n2866 ) | ( n2865 & ~n2866 ) ;
  assign n2868 = n197 & n2867 ;
  buffer buf_n2869( .i (n2868), .o (n2869) );
  buffer buf_n2870( .i (n2869), .o (n2870) );
  assign n2871 = n1254 | n2869 ;
  assign n2872 = ( n2835 & n2870 ) | ( n2835 & n2871 ) | ( n2870 & n2871 ) ;
  assign n2873 = n2420 & n2872 ;
  assign n2874 = n2225 & ~n2226 ;
  buffer buf_n2875( .i (n2874), .o (n2875) );
  assign n2884 = ( ~n362 & n1793 ) | ( ~n362 & n2875 ) | ( n1793 & n2875 ) ;
  buffer buf_n2885( .i (n73), .o (n2885) );
  buffer buf_n2886( .i (n2885), .o (n2886) );
  assign n2887 = ( n2285 & n2884 ) | ( n2285 & ~n2886 ) | ( n2884 & ~n2886 ) ;
  buffer buf_n2888( .i (n2887), .o (n2888) );
  buffer buf_n2889( .i (n2888), .o (n2889) );
  buffer buf_n2890( .i (n2889), .o (n2890) );
  buffer buf_n2891( .i (n2890), .o (n2891) );
  assign n2892 = ~n2404 & n2888 ;
  buffer buf_n2893( .i (n2892), .o (n2893) );
  buffer buf_n2894( .i (n2893), .o (n2894) );
  assign n2895 = ( n2322 & n2779 ) | ( n2322 & n2893 ) | ( n2779 & n2893 ) ;
  assign n2896 = ( n2891 & n2894 ) | ( n2891 & n2895 ) | ( n2894 & n2895 ) ;
  buffer buf_n2897( .i (n2896), .o (n2897) );
  buffer buf_n2898( .i (n2897), .o (n2898) );
  buffer buf_n2899( .i (n2898), .o (n2899) );
  assign n2900 = ( n390 & n1832 ) | ( n390 & ~n2625 ) | ( n1832 & ~n2625 ) ;
  buffer buf_n2901( .i (n2900), .o (n2901) );
  buffer buf_n2902( .i (n2901), .o (n2902) );
  buffer buf_n2903( .i (n2902), .o (n2903) );
  buffer buf_n2904( .i (n102), .o (n2904) );
  buffer buf_n2905( .i (n2327), .o (n2905) );
  assign n2906 = ( n2886 & n2904 ) | ( n2886 & ~n2905 ) | ( n2904 & ~n2905 ) ;
  buffer buf_n2907( .i (n2906), .o (n2907) );
  buffer buf_n2908( .i (n2907), .o (n2908) );
  buffer buf_n2909( .i (n2908), .o (n2909) );
  buffer buf_n2910( .i (n2909), .o (n2910) );
  assign n2911 = ( n2395 & ~n2779 ) | ( n2395 & n2901 ) | ( ~n2779 & n2901 ) ;
  assign n2912 = ( n393 & n2910 ) | ( n393 & ~n2911 ) | ( n2910 & ~n2911 ) ;
  assign n2913 = n2903 & ~n2912 ;
  assign n2914 = ( ~n198 & n2897 ) | ( ~n198 & n2913 ) | ( n2897 & n2913 ) ;
  assign n2915 = n2644 | n2914 ;
  assign n2916 = ( ~n1908 & n2899 ) | ( ~n1908 & n2915 ) | ( n2899 & n2915 ) ;
  assign n2917 = n2420 | n2916 ;
  buffer buf_n2918( .i (n2420), .o (n2918) );
  assign n2919 = ( n2873 & n2917 ) | ( n2873 & ~n2918 ) | ( n2917 & ~n2918 ) ;
  buffer buf_n2920( .i (n2739), .o (n2920) );
  assign n2921 = n2919 & n2920 ;
  buffer buf_n2922( .i (n2886), .o (n2922) );
  buffer buf_n2923( .i (n2922), .o (n2923) );
  buffer buf_n2924( .i (n2923), .o (n2924) );
  buffer buf_n2925( .i (n2436), .o (n2925) );
  buffer buf_n2926( .i (n2925), .o (n2926) );
  assign n2927 = ~n2924 & n2926 ;
  buffer buf_n2928( .i (n2927), .o (n2928) );
  buffer buf_n2929( .i (n2928), .o (n2929) );
  buffer buf_n2840( .i (n2839), .o (n2840) );
  buffer buf_n2841( .i (n2840), .o (n2841) );
  buffer buf_n2842( .i (n2841), .o (n2842) );
  buffer buf_n2843( .i (n2842), .o (n2843) );
  buffer buf_n2844( .i (n2843), .o (n2844) );
  buffer buf_n2936( .i (n2322), .o (n2936) );
  assign n2937 = ( n1622 & n2844 ) | ( n1622 & n2936 ) | ( n2844 & n2936 ) ;
  buffer buf_n2938( .i (n1621), .o (n2938) );
  assign n2939 = ( n2780 & n2844 ) | ( n2780 & n2938 ) | ( n2844 & n2938 ) ;
  assign n2940 = ( n2929 & n2937 ) | ( n2929 & ~n2939 ) | ( n2937 & ~n2939 ) ;
  assign n2941 = ~n582 & n2050 ;
  buffer buf_n2942( .i (n2941), .o (n2942) );
  buffer buf_n2943( .i (n2942), .o (n2943) );
  assign n2944 = n197 | n2942 ;
  assign n2945 = ( n2940 & n2943 ) | ( n2940 & n2944 ) | ( n2943 & n2944 ) ;
  buffer buf_n2946( .i (n2945), .o (n2946) );
  buffer buf_n2947( .i (n2946), .o (n2947) );
  buffer buf_n2948( .i (n2418), .o (n2948) );
  assign n2949 = ( n2596 & n2946 ) | ( n2596 & ~n2948 ) | ( n2946 & ~n2948 ) ;
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  assign n2950 = ~n549 & n2744 ;
  assign n2951 = n442 & n2950 ;
  assign n2952 = ~n2596 & n2951 ;
  assign n2953 = ( n2947 & ~n2949 ) | ( n2947 & n2952 ) | ( ~n2949 & n2952 ) ;
  assign n2954 = ( ~n2276 & n2334 ) | ( ~n2276 & n2388 ) | ( n2334 & n2388 ) ;
  buffer buf_n2955( .i (n2954), .o (n2955) );
  buffer buf_n2956( .i (n2955), .o (n2956) );
  buffer buf_n2957( .i (n2956), .o (n2957) );
  buffer buf_n2958( .i (n2957), .o (n2958) );
  buffer buf_n2959( .i (n1450), .o (n2959) );
  buffer buf_n2960( .i (n2959), .o (n2960) );
  assign n2961 = ( n2405 & n2955 ) | ( n2405 & ~n2960 ) | ( n2955 & ~n2960 ) ;
  buffer buf_n2962( .i (n2961), .o (n2962) );
  buffer buf_n2963( .i (n2962), .o (n2963) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  buffer buf_n2280( .i (n2279), .o (n2280) );
  assign n2964 = n2280 & n2962 ;
  assign n2965 = ( ~n2958 & n2963 ) | ( ~n2958 & n2964 ) | ( n2963 & n2964 ) ;
  assign n2966 = n2744 & n2965 ;
  buffer buf_n2967( .i (n2960), .o (n2967) );
  assign n2968 = ( n1621 & ~n2378 ) | ( n1621 & n2967 ) | ( ~n2378 & n2967 ) ;
  assign n2969 = ( n2448 & n2806 ) | ( n2448 & ~n2968 ) | ( n2806 & ~n2968 ) ;
  buffer buf_n2970( .i (n2448), .o (n2970) );
  assign n2971 = ( n2517 & n2969 ) | ( n2517 & ~n2970 ) | ( n2969 & ~n2970 ) ;
  buffer buf_n2972( .i (n2505), .o (n2972) );
  assign n2973 = n2971 | n2972 ;
  assign n2974 = ( ~n2745 & n2966 ) | ( ~n2745 & n2973 ) | ( n2966 & n2973 ) ;
  buffer buf_n2975( .i (n2384), .o (n2975) );
  buffer buf_n2976( .i (n2595), .o (n2976) );
  assign n2977 = ( n2974 & ~n2975 ) | ( n2974 & n2976 ) | ( ~n2975 & n2976 ) ;
  buffer buf_n2978( .i (n2404), .o (n2978) );
  assign n2979 = ( n2377 & n2960 ) | ( n2377 & ~n2978 ) | ( n2960 & ~n2978 ) ;
  buffer buf_n2980( .i (n2979), .o (n2980) );
  assign n2981 = ( ~n1812 & n2936 ) | ( ~n1812 & n2980 ) | ( n2936 & n2980 ) ;
  buffer buf_n2982( .i (n2378), .o (n2982) );
  assign n2983 = ( n2936 & ~n2980 ) | ( n2936 & n2982 ) | ( ~n2980 & n2982 ) ;
  assign n2984 = n2981 & ~n2983 ;
  buffer buf_n2985( .i (n1887), .o (n2985) );
  assign n2986 = ~n2984 & n2985 ;
  buffer buf_n2987( .i (n2936), .o (n2987) );
  assign n2988 = n606 & ~n2987 ;
  assign n2989 = n2985 | n2988 ;
  assign n2990 = ~n2986 & n2989 ;
  assign n2991 = ( n2975 & n2976 ) | ( n2975 & n2990 ) | ( n2976 & n2990 ) ;
  assign n2992 = n2977 & n2991 ;
  assign n2993 = n2953 | n2992 ;
  assign n2994 = ~n2920 & n2993 ;
  assign n2995 = n2921 | n2994 ;
  buffer buf_n2996( .i (n2995), .o (n2996) );
  assign n2997 = ( ~n2826 & n2831 ) | ( ~n2826 & n2996 ) | ( n2831 & n2996 ) ;
  assign n2998 = n249 | n2386 ;
  buffer buf_n2999( .i (n2998), .o (n2999) );
  buffer buf_n3000( .i (n2999), .o (n3000) );
  buffer buf_n3001( .i (n3000), .o (n3001) );
  assign n3005 = ( ~n2395 & n2493 ) | ( ~n2395 & n3001 ) | ( n2493 & n3001 ) ;
  buffer buf_n3006( .i (n3005), .o (n3006) );
  buffer buf_n3007( .i (n3006), .o (n3007) );
  buffer buf_n3008( .i (n3007), .o (n3008) );
  buffer buf_n3009( .i (n3008), .o (n3009) );
  buffer buf_n3010( .i (n3009), .o (n3010) );
  buffer buf_n3011( .i (n3010), .o (n3011) );
  buffer buf_n3012( .i (n3011), .o (n3012) );
  buffer buf_n3013( .i (n3012), .o (n3013) );
  buffer buf_n3014( .i (n3013), .o (n3014) );
  buffer buf_n3015( .i (n3014), .o (n3015) );
  assign n3016 = n2996 | n3015 ;
  assign n3017 = ( n2827 & n2997 ) | ( n2827 & n3016 ) | ( n2997 & n3016 ) ;
  buffer buf_n3018( .i (n3017), .o (n3018) );
  buffer buf_n3019( .i (n3018), .o (n3019) );
  buffer buf_n3020( .i (n2619), .o (n3020) );
  assign n3021 = n3018 & n3020 ;
  buffer buf_n3022( .i (n2540), .o (n3022) );
  assign n3023 = n603 & ~n3022 ;
  buffer buf_n3024( .i (n3023), .o (n3024) );
  buffer buf_n3025( .i (n3024), .o (n3025) );
  buffer buf_n3026( .i (n3025), .o (n3026) );
  buffer buf_n3027( .i (n3026), .o (n3027) );
  buffer buf_n3028( .i (n3027), .o (n3028) );
  buffer buf_n3029( .i (n3028), .o (n3029) );
  buffer buf_n3030( .i (n3029), .o (n3030) );
  buffer buf_n3031( .i (n3030), .o (n3031) );
  buffer buf_n3032( .i (n3031), .o (n3032) );
  buffer buf_n3033( .i (n3032), .o (n3033) );
  buffer buf_n3034( .i (n3033), .o (n3034) );
  buffer buf_n3035( .i (n3034), .o (n3035) );
  assign n3036 = n1250 & n3035 ;
  buffer buf_n3037( .i (n3036), .o (n3037) );
  assign n3038 = n22 & n2514 ;
  buffer buf_n3039( .i (n3022), .o (n3039) );
  assign n3040 = ( n2779 & n3038 ) | ( n2779 & ~n3039 ) | ( n3038 & ~n3039 ) ;
  buffer buf_n3041( .i (n3040), .o (n3041) );
  buffer buf_n3042( .i (n3041), .o (n3042) );
  buffer buf_n3043( .i (n3042), .o (n3043) );
  assign n3044 = ( n25 & n2781 ) | ( n25 & ~n3041 ) | ( n2781 & ~n3041 ) ;
  assign n3045 = ( ~n198 & n2985 ) | ( ~n198 & n3044 ) | ( n2985 & n3044 ) ;
  assign n3046 = ~n3043 & n3045 ;
  assign n3047 = ~n1908 & n3046 ;
  assign n3048 = n1375 | n3047 ;
  assign n3049 = ( ~n1562 & n2120 ) | ( ~n1562 & n2384 ) | ( n2120 & n2384 ) ;
  assign n3050 = ~n2526 & n3049 ;
  buffer buf_n3051( .i (n2643), .o (n3051) );
  buffer buf_n3052( .i (n3051), .o (n3052) );
  assign n3053 = ~n3050 & n3052 ;
  assign n3054 = n3048 & ~n3053 ;
  assign n3055 = n2476 | n3054 ;
  buffer buf_n3056( .i (n2328), .o (n3056) );
  assign n3057 = ( n47 & n2905 ) | ( n47 & n3056 ) | ( n2905 & n3056 ) ;
  buffer buf_n3058( .i (n3057), .o (n3058) );
  buffer buf_n3059( .i (n3058), .o (n3059) );
  buffer buf_n3060( .i (n3059), .o (n3060) );
  buffer buf_n3065( .i (n1938), .o (n3065) );
  buffer buf_n3066( .i (n2926), .o (n3066) );
  assign n3067 = ( n3060 & ~n3065 ) | ( n3060 & n3066 ) | ( ~n3065 & n3066 ) ;
  buffer buf_n3068( .i (n3067), .o (n3068) );
  buffer buf_n3069( .i (n3068), .o (n3069) );
  buffer buf_n3070( .i (n3069), .o (n3070) );
  buffer buf_n3071( .i (n3070), .o (n3071) );
  assign n3072 = ( n1887 & n2970 ) | ( n1887 & n3068 ) | ( n2970 & n3068 ) ;
  buffer buf_n3073( .i (n3072), .o (n3073) );
  buffer buf_n3074( .i (n3073), .o (n3074) );
  buffer buf_n3061( .i (n3060), .o (n3061) );
  buffer buf_n3062( .i (n3061), .o (n3062) );
  buffer buf_n3063( .i (n3062), .o (n3063) );
  buffer buf_n3064( .i (n3063), .o (n3064) );
  assign n3075 = ~n3064 & n3073 ;
  assign n3076 = ( ~n3071 & n3074 ) | ( ~n3071 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3077 = n1909 & n3076 ;
  assign n3078 = ~n1894 & n3077 ;
  assign n3079 = n2476 & ~n3078 ;
  assign n3080 = n3055 & ~n3079 ;
  assign n3081 = ~n2791 & n3080 ;
  buffer buf_n3082( .i (n3081), .o (n3082) );
  buffer buf_n3083( .i (n3082), .o (n3083) );
  buffer buf_n3084( .i (n2745), .o (n3084) );
  buffer buf_n3085( .i (n3084), .o (n3085) );
  assign n3086 = ( ~n1909 & n2558 ) | ( ~n1909 & n3085 ) | ( n2558 & n3085 ) ;
  buffer buf_n3087( .i (n3086), .o (n3087) );
  buffer buf_n3089( .i (n2735), .o (n3089) );
  buffer buf_n3090( .i (n3089), .o (n3090) );
  assign n3091 = ( n202 & n2751 ) | ( n202 & ~n3090 ) | ( n2751 & ~n3090 ) ;
  assign n3092 = ~n3087 & n3091 ;
  buffer buf_n3093( .i (n3092), .o (n3093) );
  buffer buf_n3094( .i (n3093), .o (n3094) );
  assign n3095 = n53 & n2397 ;
  buffer buf_n3096( .i (n3095), .o (n3096) );
  buffer buf_n3097( .i (n3096), .o (n3097) );
  buffer buf_n3098( .i (n3097), .o (n3098) );
  buffer buf_n3099( .i (n3098), .o (n3099) );
  buffer buf_n3100( .i (n3099), .o (n3100) );
  buffer buf_n3101( .i (n3100), .o (n3101) );
  buffer buf_n3102( .i (n3101), .o (n3102) );
  assign n3103 = ( n2689 & ~n3093 ) | ( n2689 & n3102 ) | ( ~n3093 & n3102 ) ;
  assign n3104 = n3094 & n3103 ;
  assign n3105 = n3082 | n3104 ;
  buffer buf_n3106( .i (n1783), .o (n3106) );
  assign n3107 = ( n3083 & n3105 ) | ( n3083 & ~n3106 ) | ( n3105 & ~n3106 ) ;
  assign n3108 = n3037 | n3107 ;
  assign n3109 = ( n3019 & ~n3021 ) | ( n3019 & n3108 ) | ( ~n3021 & n3108 ) ;
  assign n3110 = n2798 | n3109 ;
  assign n3111 = ( n2697 & ~n2714 ) | ( n2697 & n3110 ) | ( ~n2714 & n3110 ) ;
  buffer buf_n2713( .i (n2712), .o (n2713) );
  assign n3112 = n2960 & n3022 ;
  buffer buf_n3113( .i (n3112), .o (n3113) );
  buffer buf_n3114( .i (n3113), .o (n3114) );
  buffer buf_n3115( .i (n3114), .o (n3115) );
  buffer buf_n3116( .i (n3115), .o (n3116) );
  buffer buf_n3117( .i (n3116), .o (n3117) );
  buffer buf_n3118( .i (n3117), .o (n3118) );
  buffer buf_n3119( .i (n3118), .o (n3119) );
  buffer buf_n3120( .i (n3119), .o (n3120) );
  buffer buf_n3121( .i (n3120), .o (n3121) );
  buffer buf_n3122( .i (n3121), .o (n3122) );
  buffer buf_n3123( .i (n3122), .o (n3123) );
  buffer buf_n3124( .i (n3123), .o (n3124) );
  buffer buf_n3125( .i (n3124), .o (n3125) );
  buffer buf_n3126( .i (n3125), .o (n3126) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  buffer buf_n3127( .i (n2387), .o (n3127) );
  buffer buf_n3128( .i (n3127), .o (n3128) );
  buffer buf_n3129( .i (n3128), .o (n3129) );
  assign n3130 = n3065 & ~n3129 ;
  buffer buf_n3131( .i (n3130), .o (n3131) );
  buffer buf_n3132( .i (n3131), .o (n3132) );
  buffer buf_n3133( .i (n3132), .o (n3133) );
  buffer buf_n3135( .i (n2781), .o (n3135) );
  buffer buf_n3136( .i (n3135), .o (n3136) );
  assign n3137 = n3133 & n3136 ;
  buffer buf_n3138( .i (n3065), .o (n3138) );
  buffer buf_n3139( .i (n3138), .o (n3139) );
  buffer buf_n3140( .i (n3139), .o (n3140) );
  assign n3141 = ( n2972 & n3132 ) | ( n2972 & ~n3140 ) | ( n3132 & ~n3140 ) ;
  assign n3142 = ( n1943 & ~n3136 ) | ( n1943 & n3141 ) | ( ~n3136 & n3141 ) ;
  assign n3143 = ( n2975 & ~n3137 ) | ( n2975 & n3142 ) | ( ~n3137 & n3142 ) ;
  buffer buf_n3144( .i (n2581), .o (n3144) );
  buffer buf_n3145( .i (n3144), .o (n3145) );
  assign n3146 = ( n48 & n2922 ) | ( n48 & ~n3145 ) | ( n2922 & ~n3145 ) ;
  assign n3147 = ( n825 & ~n2625 ) | ( n825 & n3146 ) | ( ~n2625 & n3146 ) ;
  buffer buf_n3148( .i (n3147), .o (n3148) );
  assign n3151 = n3065 & ~n3148 ;
  buffer buf_n3152( .i (n3151), .o (n3152) );
  buffer buf_n3153( .i (n3152), .o (n3153) );
  buffer buf_n3149( .i (n3148), .o (n3149) );
  buffer buf_n3150( .i (n3149), .o (n3150) );
  assign n3154 = n3150 | n3152 ;
  assign n3155 = ( ~n3140 & n3153 ) | ( ~n3140 & n3154 ) | ( n3153 & n3154 ) ;
  buffer buf_n3156( .i (n3155), .o (n3156) );
  buffer buf_n3157( .i (n3156), .o (n3157) );
  assign n3158 = n2735 & ~n3156 ;
  assign n3159 = ( n3143 & ~n3157 ) | ( n3143 & n3158 ) | ( ~n3157 & n3158 ) ;
  assign n3160 = n2918 & ~n3159 ;
  assign n3161 = ( n396 & ~n955 ) | ( n396 & n2728 ) | ( ~n955 & n2728 ) ;
  assign n3162 = n3051 | n3161 ;
  assign n3163 = n369 & n2781 ;
  buffer buf_n3164( .i (n3163), .o (n3164) );
  assign n3171 = n2745 & n3164 ;
  assign n3172 = n3051 & ~n3171 ;
  assign n3173 = n3162 & ~n3172 ;
  assign n3174 = n2918 | n3173 ;
  assign n3175 = ( ~n261 & n3160 ) | ( ~n261 & n3174 ) | ( n3160 & n3174 ) ;
  assign n3176 = ( n204 & ~n2533 ) | ( n204 & n3175 ) | ( ~n2533 & n3175 ) ;
  buffer buf_n3177( .i (n2972), .o (n3177) );
  assign n3178 = ( n2418 & n3136 ) | ( n2418 & ~n3177 ) | ( n3136 & ~n3177 ) ;
  assign n3179 = n1985 & ~n3178 ;
  buffer buf_n3180( .i (n3179), .o (n3180) );
  buffer buf_n3181( .i (n3180), .o (n3181) );
  buffer buf_n3182( .i (n2924), .o (n3182) );
  assign n3183 = ( ~n422 & n3066 ) | ( ~n422 & n3182 ) | ( n3066 & n3182 ) ;
  assign n3184 = ( ~n2396 & n3138 ) | ( ~n2396 & n3183 ) | ( n3138 & n3183 ) ;
  assign n3185 = ~n424 & n3184 ;
  assign n3186 = ( n2417 & ~n2985 ) | ( n2417 & n3185 ) | ( ~n2985 & n3185 ) ;
  buffer buf_n3187( .i (n101), .o (n3187) );
  assign n3188 = ( n46 & n2581 ) | ( n46 & n3187 ) | ( n2581 & n3187 ) ;
  buffer buf_n3189( .i (n3188), .o (n3189) );
  assign n3201 = ( ~n2922 & n3145 ) | ( ~n2922 & n3189 ) | ( n3145 & n3189 ) ;
  buffer buf_n3202( .i (n3201), .o (n3202) );
  assign n3205 = n3128 & ~n3202 ;
  buffer buf_n3206( .i (n3205), .o (n3206) );
  buffer buf_n3207( .i (n3206), .o (n3207) );
  buffer buf_n3203( .i (n3202), .o (n3203) );
  buffer buf_n3204( .i (n3203), .o (n3204) );
  assign n3208 = n3204 | n3206 ;
  buffer buf_n3209( .i (n2396), .o (n3209) );
  assign n3210 = ( n3207 & n3208 ) | ( n3207 & ~n3209 ) | ( n3208 & ~n3209 ) ;
  buffer buf_n3211( .i (n2806), .o (n3211) );
  buffer buf_n3212( .i (n3211), .o (n3212) );
  buffer buf_n3213( .i (n1813), .o (n3213) );
  assign n3214 = ( n3210 & n3212 ) | ( n3210 & n3213 ) | ( n3212 & n3213 ) ;
  assign n3215 = n3186 & n3214 ;
  buffer buf_n3216( .i (n3215), .o (n3216) );
  buffer buf_n3217( .i (n3216), .o (n3217) );
  buffer buf_n3218( .i (n3217), .o (n3218) );
  assign n3219 = ( ~n1699 & n3052 ) | ( ~n1699 & n3216 ) | ( n3052 & n3216 ) ;
  assign n3220 = n3180 & ~n3219 ;
  assign n3221 = ( n3181 & n3218 ) | ( n3181 & ~n3220 ) | ( n3218 & ~n3220 ) ;
  assign n3222 = ( n204 & n2533 ) | ( n204 & ~n3221 ) | ( n2533 & ~n3221 ) ;
  assign n3223 = n3176 & ~n3222 ;
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  assign n3224 = n1368 & ~n2012 ;
  buffer buf_n3225( .i (n2959), .o (n3225) );
  assign n3226 = ( n1938 & ~n3128 ) | ( n1938 & n3225 ) | ( ~n3128 & n3225 ) ;
  buffer buf_n3227( .i (n3226), .o (n3227) );
  buffer buf_n3228( .i (n3227), .o (n3228) );
  buffer buf_n3229( .i (n3228), .o (n3229) );
  buffer buf_n3230( .i (n3229), .o (n3230) );
  assign n3231 = n1812 & ~n3227 ;
  buffer buf_n3232( .i (n3231), .o (n3232) );
  buffer buf_n3233( .i (n3232), .o (n3233) );
  assign n3234 = ( n2972 & n3140 ) | ( n2972 & n3232 ) | ( n3140 & n3232 ) ;
  assign n3235 = ( ~n3230 & n3233 ) | ( ~n3230 & n3234 ) | ( n3233 & n3234 ) ;
  assign n3236 = n2975 & n3235 ;
  assign n3237 = ~n29 & n3236 ;
  buffer buf_n3238( .i (n3237), .o (n3238) );
  buffer buf_n3239( .i (n3238), .o (n3239) );
  assign n3240 = n314 & ~n3238 ;
  assign n3241 = ( n3224 & n3239 ) | ( n3224 & ~n3240 ) | ( n3239 & ~n3240 ) ;
  assign n3242 = ( n177 & n2015 ) | ( n177 & ~n3241 ) | ( n2015 & ~n3241 ) ;
  assign n3243 = ( n2202 & n3223 ) | ( n2202 & ~n3242 ) | ( n3223 & ~n3242 ) ;
  assign n3244 = n237 & ~n3243 ;
  assign n3245 = ( n2715 & n3039 ) | ( n2715 & ~n3129 ) | ( n3039 & ~n3129 ) ;
  buffer buf_n3246( .i (n3245), .o (n3246) );
  buffer buf_n3247( .i (n3246), .o (n3247) );
  buffer buf_n3248( .i (n3247), .o (n3248) );
  buffer buf_n3249( .i (n3248), .o (n3249) );
  assign n3250 = n3209 & n3246 ;
  buffer buf_n3251( .i (n3250), .o (n3251) );
  buffer buf_n3252( .i (n3251), .o (n3252) );
  buffer buf_n3253( .i (n2970), .o (n3253) );
  buffer buf_n3254( .i (n3253), .o (n3254) );
  assign n3255 = ( n3136 & n3251 ) | ( n3136 & ~n3254 ) | ( n3251 & ~n3254 ) ;
  assign n3256 = ( n3249 & n3252 ) | ( n3249 & n3255 ) | ( n3252 & n3255 ) ;
  buffer buf_n3257( .i (n3256), .o (n3257) );
  buffer buf_n3258( .i (n3257), .o (n3258) );
  buffer buf_n3259( .i (n3085), .o (n3259) );
  assign n3260 = n3257 & ~n3259 ;
  buffer buf_n3261( .i (n2625), .o (n3261) );
  assign n3262 = ( n3128 & ~n3225 ) | ( n3128 & n3261 ) | ( ~n3225 & n3261 ) ;
  buffer buf_n3263( .i (n3262), .o (n3263) );
  buffer buf_n3264( .i (n3263), .o (n3264) );
  buffer buf_n3265( .i (n3264), .o (n3265) );
  buffer buf_n3267( .i (n2715), .o (n3267) );
  buffer buf_n3268( .i (n2967), .o (n3268) );
  assign n3269 = ( n2982 & ~n3267 ) | ( n2982 & n3268 ) | ( ~n3267 & n3268 ) ;
  assign n3270 = ~n3209 & n3269 ;
  assign n3271 = n3265 | n3270 ;
  buffer buf_n3272( .i (n3271), .o (n3272) );
  buffer buf_n3273( .i (n3272), .o (n3273) );
  buffer buf_n3274( .i (n3135), .o (n3274) );
  buffer buf_n3275( .i (n3274), .o (n3275) );
  assign n3276 = ( n3084 & ~n3272 ) | ( n3084 & n3275 ) | ( ~n3272 & n3275 ) ;
  assign n3277 = n1752 | n3267 ;
  buffer buf_n3278( .i (n3277), .o (n3278) );
  assign n3288 = n2594 & ~n3278 ;
  assign n3289 = n3177 & n3288 ;
  assign n3290 = ~n3275 & n3289 ;
  assign n3291 = ( n3273 & n3276 ) | ( n3273 & ~n3290 ) | ( n3276 & ~n3290 ) ;
  buffer buf_n2930( .i (n2929), .o (n2930) );
  buffer buf_n2931( .i (n2930), .o (n2931) );
  buffer buf_n2932( .i (n2931), .o (n2932) );
  assign n3292 = n2932 & ~n2976 ;
  assign n3293 = ~n2197 & n3292 ;
  assign n3294 = n3291 & ~n3293 ;
  assign n3295 = ( ~n3258 & n3260 ) | ( ~n3258 & n3294 ) | ( n3260 & n3294 ) ;
  buffer buf_n3296( .i (n2920), .o (n3296) );
  assign n3297 = ~n3295 & n3296 ;
  buffer buf_n2307( .i (n2306), .o (n2307) );
  buffer buf_n2308( .i (n2307), .o (n2308) );
  buffer buf_n2309( .i (n2308), .o (n2309) );
  buffer buf_n2310( .i (n2309), .o (n2310) );
  assign n3298 = ( n1312 & n2309 ) | ( n1312 & ~n2970 ) | ( n2309 & ~n2970 ) ;
  assign n3299 = ~n2310 & n3298 ;
  buffer buf_n3300( .i (n3299), .o (n3300) );
  buffer buf_n3301( .i (n3300), .o (n3301) );
  buffer buf_n3302( .i (n3301), .o (n3302) );
  assign n3303 = ( n2005 & n3117 ) | ( n2005 & n3300 ) | ( n3117 & n3300 ) ;
  assign n3304 = n3089 & ~n3303 ;
  assign n3305 = ( n3090 & n3302 ) | ( n3090 & ~n3304 ) | ( n3302 & ~n3304 ) ;
  assign n3306 = ( n2540 & n2959 ) | ( n2540 & n3127 ) | ( n2959 & n3127 ) ;
  buffer buf_n3307( .i (n3306), .o (n3307) );
  buffer buf_n3308( .i (n3307), .o (n3308) );
  buffer buf_n3309( .i (n3308), .o (n3309) );
  buffer buf_n3310( .i (n3268), .o (n3310) );
  assign n3311 = n3309 & n3310 ;
  buffer buf_n3312( .i (n3182), .o (n3312) );
  buffer buf_n3313( .i (n3129), .o (n3313) );
  assign n3314 = ( n3308 & n3312 ) | ( n3308 & n3313 ) | ( n3312 & n3313 ) ;
  assign n3315 = n3310 | n3314 ;
  assign n3316 = ~n3311 & n3315 ;
  assign n3317 = n3274 | n3316 ;
  buffer buf_n3318( .i (n2987), .o (n3318) );
  assign n3319 = n1046 & n3318 ;
  assign n3320 = n3274 & ~n3319 ;
  assign n3321 = n3317 & ~n3320 ;
  assign n3322 = n3089 | n3321 ;
  assign n3323 = ~n2356 & n3117 ;
  assign n3324 = n3089 & ~n3323 ;
  assign n3325 = n3322 & ~n3324 ;
  assign n3326 = n3305 | n3325 ;
  assign n3327 = ~n3296 & n3326 ;
  assign n3328 = n3297 | n3327 ;
  assign n3329 = ~n2109 & n3328 ;
  assign n3330 = n237 | n3329 ;
  assign n3331 = ~n3244 & n3330 ;
  buffer buf_n3332( .i (n2905), .o (n3332) );
  buffer buf_n3333( .i (n3332), .o (n3333) );
  assign n3334 = ( n21 & n3127 ) | ( n21 & n3333 ) | ( n3127 & n3333 ) ;
  buffer buf_n3335( .i (n3334), .o (n3335) );
  buffer buf_n3340( .i (n2978), .o (n3340) );
  assign n3341 = ( n3129 & ~n3335 ) | ( n3129 & n3340 ) | ( ~n3335 & n3340 ) ;
  buffer buf_n3342( .i (n3341), .o (n3342) );
  buffer buf_n3343( .i (n3342), .o (n3343) );
  buffer buf_n3344( .i (n3343), .o (n3344) );
  buffer buf_n3345( .i (n3344), .o (n3345) );
  assign n3346 = ( n25 & n3211 ) | ( n25 & ~n3342 ) | ( n3211 & ~n3342 ) ;
  buffer buf_n3347( .i (n3346), .o (n3347) );
  buffer buf_n3348( .i (n3347), .o (n3348) );
  buffer buf_n3336( .i (n3335), .o (n3336) );
  buffer buf_n3337( .i (n3336), .o (n3337) );
  buffer buf_n3338( .i (n3337), .o (n3338) );
  buffer buf_n3339( .i (n3338), .o (n3339) );
  assign n3349 = ~n3339 & n3347 ;
  assign n3350 = ( n3345 & n3348 ) | ( n3345 & n3349 ) | ( n3348 & n3349 ) ;
  buffer buf_n3351( .i (n3350), .o (n3351) );
  buffer buf_n3352( .i (n3351), .o (n3352) );
  assign n3353 = n2739 & n3351 ;
  assign n3354 = ( n1773 & n2507 ) | ( n1773 & n2594 ) | ( n2507 & n2594 ) ;
  buffer buf_n3355( .i (n3354), .o (n3355) );
  assign n3356 = ( ~n2976 & n3051 ) | ( ~n2976 & n3355 ) | ( n3051 & n3355 ) ;
  buffer buf_n3357( .i (n2643), .o (n3357) );
  assign n3358 = ( n2526 & ~n3355 ) | ( n2526 & n3357 ) | ( ~n3355 & n3357 ) ;
  assign n3359 = n3356 & ~n3358 ;
  buffer buf_n3360( .i (n2595), .o (n3360) );
  assign n3361 = n727 & ~n3360 ;
  assign n3362 = ~n1507 & n3361 ;
  assign n3363 = n3359 | n3362 ;
  assign n3364 = ( n3352 & ~n3353 ) | ( n3352 & n3363 ) | ( ~n3353 & n3363 ) ;
  assign n3365 = n88 | n3364 ;
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n3366( .i (n2735), .o (n3366) );
  assign n3367 = ( ~n1613 & n3052 ) | ( ~n1613 & n3366 ) | ( n3052 & n3366 ) ;
  buffer buf_n3368( .i (n2938), .o (n3368) );
  assign n3369 = ( n3139 & ~n3211 ) | ( n3139 & n3368 ) | ( ~n3211 & n3368 ) ;
  buffer buf_n3370( .i (n3369), .o (n3370) );
  buffer buf_n3371( .i (n3370), .o (n3371) );
  buffer buf_n3372( .i (n3371), .o (n3372) );
  assign n3373 = n3052 & ~n3372 ;
  assign n3374 = n3367 & ~n3373 ;
  buffer buf_n3375( .i (n1894), .o (n3375) );
  assign n3376 = n3374 & ~n3375 ;
  buffer buf_n3377( .i (n3259), .o (n3377) );
  buffer buf_n3378( .i (n3377), .o (n3378) );
  assign n3379 = ~n3376 & n3378 ;
  assign n3380 = n3365 & ~n3379 ;
  assign n3381 = n118 | n3380 ;
  assign n3382 = n2734 & n2766 ;
  buffer buf_n3383( .i (n3382), .o (n3383) );
  assign n3387 = ~n3085 & n3383 ;
  assign n3388 = ( n595 & ~n3259 ) | ( n595 & n3387 ) | ( ~n3259 & n3387 ) ;
  assign n3389 = n2920 & ~n3388 ;
  buffer buf_n3390( .i (n2734), .o (n3390) );
  assign n3391 = ( n1908 & n3084 ) | ( n1908 & n3390 ) | ( n3084 & n3390 ) ;
  buffer buf_n3392( .i (n3360), .o (n3392) );
  assign n3393 = n3391 & n3392 ;
  assign n3394 = ( n528 & n2634 ) | ( n528 & ~n3393 ) | ( n2634 & ~n3393 ) ;
  buffer buf_n3395( .i (n2739), .o (n3395) );
  assign n3396 = n3394 | n3395 ;
  assign n3397 = ( ~n3296 & n3389 ) | ( ~n3296 & n3396 ) | ( n3389 & n3396 ) ;
  buffer buf_n3398( .i (n2533), .o (n3398) );
  assign n3399 = n3397 | n3398 ;
  buffer buf_n3400( .i (n2689), .o (n3400) );
  assign n3401 = n3399 & n3400 ;
  assign n3402 = n3381 & ~n3401 ;
  assign n3403 = ( n208 & n266 ) | ( n208 & n3402 ) | ( n266 & n3402 ) ;
  assign n3404 = ( ~n3126 & n3331 ) | ( ~n3126 & n3403 ) | ( n3331 & n3403 ) ;
  buffer buf_n3405( .i (n3404), .o (n3405) );
  buffer buf_n3406( .i (n3405), .o (n3406) );
  assign n3407 = ( n3084 & ~n3357 ) | ( n3084 & n3390 ) | ( ~n3357 & n3390 ) ;
  buffer buf_n3408( .i (n3407), .o (n3408) );
  buffer buf_n3409( .i (n3408), .o (n3409) );
  buffer buf_n3410( .i (n3409), .o (n3410) );
  assign n3411 = ( n234 & n2535 ) | ( n234 & ~n3410 ) | ( n2535 & ~n3410 ) ;
  assign n3412 = ( n234 & ~n3378 ) | ( n234 & n3410 ) | ( ~n3378 & n3410 ) ;
  assign n3413 = n3411 & ~n3412 ;
  buffer buf_n3414( .i (n3413), .o (n3414) );
  buffer buf_n3415( .i (n3414), .o (n3415) );
  buffer buf_n3416( .i (n2109), .o (n3416) );
  assign n3417 = n3414 & n3416 ;
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n3418( .i (n233), .o (n3418) );
  assign n3419 = n708 & n3418 ;
  buffer buf_n3420( .i (n3378), .o (n3420) );
  buffer buf_n3421( .i (n2535), .o (n3421) );
  assign n3422 = ( n3419 & n3420 ) | ( n3419 & n3421 ) | ( n3420 & n3421 ) ;
  buffer buf_n3423( .i (n3420), .o (n3423) );
  assign n3424 = n3422 & ~n3423 ;
  buffer buf_n3384( .i (n3383), .o (n3384) );
  buffer buf_n3385( .i (n3384), .o (n3385) );
  buffer buf_n3386( .i (n3385), .o (n3386) );
  buffer buf_n3425( .i (n24), .o (n3425) );
  assign n3426 = ( n3139 & n3209 ) | ( n3139 & n3425 ) | ( n3209 & n3425 ) ;
  buffer buf_n3427( .i (n3426), .o (n3427) );
  assign n3428 = ( n2524 & n2644 ) | ( n2524 & ~n3427 ) | ( n2644 & ~n3427 ) ;
  buffer buf_n3429( .i (n3140), .o (n3429) );
  assign n3430 = ( n2644 & n3427 ) | ( n2644 & ~n3429 ) | ( n3427 & ~n3429 ) ;
  assign n3431 = ~n3428 & n3430 ;
  buffer buf_n3432( .i (n3431), .o (n3432) );
  buffer buf_n3433( .i (n3432), .o (n3433) );
  buffer buf_n3434( .i (n3433), .o (n3434) );
  buffer buf_n3435( .i (n2526), .o (n3435) );
  buffer buf_n3436( .i (n3435), .o (n3436) );
  buffer buf_n3437( .i (n3357), .o (n3437) );
  buffer buf_n3438( .i (n3437), .o (n3438) );
  assign n3439 = ( ~n3432 & n3436 ) | ( ~n3432 & n3438 ) | ( n3436 & n3438 ) ;
  assign n3440 = n3385 & n3439 ;
  assign n3441 = ( n3386 & n3434 ) | ( n3386 & ~n3440 ) | ( n3434 & ~n3440 ) ;
  assign n3442 = n3420 | n3441 ;
  buffer buf_n3443( .i (n3368), .o (n3443) );
  buffer buf_n3444( .i (n3443), .o (n3444) );
  buffer buf_n3445( .i (n3444), .o (n3445) );
  assign n3446 = ( n3357 & n3360 ) | ( n3357 & ~n3445 ) | ( n3360 & ~n3445 ) ;
  buffer buf_n3447( .i (n3446), .o (n3447) );
  assign n3448 = ( ~n2576 & n3090 ) | ( ~n2576 & n3447 ) | ( n3090 & n3447 ) ;
  assign n3449 = ( n3090 & n3438 ) | ( n3090 & ~n3447 ) | ( n3438 & ~n3447 ) ;
  assign n3450 = n3448 & ~n3449 ;
  buffer buf_n3451( .i (n3375), .o (n3451) );
  assign n3452 = n3450 & ~n3451 ;
  assign n3453 = n3420 & ~n3452 ;
  assign n3454 = n3442 & ~n3453 ;
  assign n3455 = n3424 | n3454 ;
  assign n3456 = ( n3415 & ~n3417 ) | ( n3415 & n3455 ) | ( ~n3417 & n3455 ) ;
  assign n3457 = n121 | n3456 ;
  assign n3458 = n3378 & ~n3418 ;
  buffer buf_n3459( .i (n3377), .o (n3459) );
  buffer buf_n3460( .i (n3459), .o (n3460) );
  assign n3461 = ( n598 & n3458 ) | ( n598 & ~n3460 ) | ( n3458 & ~n3460 ) ;
  assign n3462 = n2363 & n3461 ;
  buffer buf_n3463( .i (n2403), .o (n3463) );
  assign n3464 = ( n2923 & ~n3127 ) | ( n2923 & n3463 ) | ( ~n3127 & n3463 ) ;
  buffer buf_n3465( .i (n3464), .o (n3465) );
  buffer buf_n3466( .i (n3465), .o (n3466) );
  buffer buf_n3467( .i (n3466), .o (n3467) );
  buffer buf_n3468( .i (n3467), .o (n3468) );
  buffer buf_n3469( .i (n3468), .o (n3469) );
  buffer buf_n3470( .i (n3469), .o (n3470) );
  assign n3475 = ( n3390 & ~n3445 ) | ( n3390 & n3470 ) | ( ~n3445 & n3470 ) ;
  buffer buf_n3476( .i (n3475), .o (n3476) );
  buffer buf_n3477( .i (n3476), .o (n3477) );
  buffer buf_n3478( .i (n3477), .o (n3478) );
  buffer buf_n3479( .i (n3478), .o (n3479) );
  assign n3480 = ( ~n2576 & n3259 ) | ( ~n2576 & n3476 ) | ( n3259 & n3476 ) ;
  buffer buf_n3481( .i (n3480), .o (n3481) );
  buffer buf_n3482( .i (n3481), .o (n3482) );
  buffer buf_n3471( .i (n3470), .o (n3471) );
  buffer buf_n3472( .i (n3471), .o (n3472) );
  buffer buf_n3473( .i (n3472), .o (n3473) );
  buffer buf_n3474( .i (n3473), .o (n3474) );
  assign n3483 = ~n3474 & n3481 ;
  assign n3484 = ( ~n3479 & n3482 ) | ( ~n3479 & n3483 ) | ( n3482 & n3483 ) ;
  buffer buf_n3485( .i (n2830), .o (n3485) );
  assign n3486 = n3484 | n3485 ;
  assign n3487 = ( ~n63 & n3462 ) | ( ~n63 & n3486 ) | ( n3462 & n3486 ) ;
  assign n3488 = ~n3106 & n3487 ;
  buffer buf_n3489( .i (n120), .o (n3489) );
  assign n3490 = ~n3488 & n3489 ;
  assign n3491 = n3457 & ~n3490 ;
  assign n3492 = n3405 | n3491 ;
  assign n3493 = ( ~n2713 & n3406 ) | ( ~n2713 & n3492 ) | ( n3406 & n3492 ) ;
  buffer buf_n360( .i (n359), .o (n360) );
  assign n3494 = n24 & ~n2982 ;
  buffer buf_n3495( .i (n3494), .o (n3495) );
  buffer buf_n3496( .i (n3495), .o (n3496) );
  assign n3497 = ( ~n2595 & n3444 ) | ( ~n2595 & n3496 ) | ( n3444 & n3496 ) ;
  assign n3498 = ( n3253 & ~n3443 ) | ( n3253 & n3495 ) | ( ~n3443 & n3495 ) ;
  buffer buf_n3499( .i (n2594), .o (n3499) );
  assign n3500 = ( ~n2524 & n3498 ) | ( ~n2524 & n3499 ) | ( n3498 & n3499 ) ;
  assign n3501 = n3497 | n3500 ;
  assign n3502 = ~n2820 & n3501 ;
  buffer buf_n2031( .i (n2030), .o (n2031) );
  buffer buf_n2032( .i (n2031), .o (n2032) );
  buffer buf_n2033( .i (n2032), .o (n2033) );
  buffer buf_n2034( .i (n2033), .o (n2034) );
  buffer buf_n2035( .i (n2034), .o (n2035) );
  buffer buf_n3503( .i (n3313), .o (n3503) );
  buffer buf_n3504( .i (n3503), .o (n3504) );
  assign n3505 = n2035 & ~n3504 ;
  buffer buf_n3506( .i (n3505), .o (n3506) );
  buffer buf_n3510( .i (n2507), .o (n3510) );
  buffer buf_n3511( .i (n3510), .o (n3511) );
  assign n3512 = n3506 & ~n3511 ;
  assign n3513 = n2820 & ~n3512 ;
  assign n3514 = n3502 | n3513 ;
  assign n3515 = ~n3377 & n3514 ;
  buffer buf_n3516( .i (n3145), .o (n3516) );
  assign n3517 = ( n2925 & ~n3463 ) | ( n2925 & n3516 ) | ( ~n3463 & n3516 ) ;
  buffer buf_n3518( .i (n3517), .o (n3518) );
  buffer buf_n3519( .i (n3518), .o (n3519) );
  buffer buf_n3520( .i (n3519), .o (n3520) );
  buffer buf_n3521( .i (n3520), .o (n3521) );
  buffer buf_n3522( .i (n3521), .o (n3522) );
  buffer buf_n3523( .i (n3522), .o (n3523) );
  assign n3524 = ( n2557 & ~n3275 ) | ( n2557 & n3523 ) | ( ~n3275 & n3523 ) ;
  assign n3525 = ( ~n2557 & n3445 ) | ( ~n2557 & n3523 ) | ( n3445 & n3523 ) ;
  assign n3526 = n3524 & n3525 ;
  assign n3527 = ~n3436 & n3526 ;
  assign n3528 = n3377 & ~n3527 ;
  assign n3529 = n3515 | n3528 ;
  assign n3530 = ~n2830 & n3529 ;
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  assign n3531 = n862 & n3504 ;
  buffer buf_n3532( .i (n3531), .o (n3532) );
  buffer buf_n3533( .i (n3532), .o (n3533) );
  buffer buf_n3534( .i (n3533), .o (n3534) );
  buffer buf_n3536( .i (n3085), .o (n3536) );
  assign n3537 = ~n3534 & n3536 ;
  assign n3538 = n2120 & ~n3499 ;
  buffer buf_n3539( .i (n3538), .o (n3539) );
  assign n3540 = ~n2820 & n3539 ;
  assign n3541 = n3536 | n3540 ;
  assign n3542 = ~n3537 & n3541 ;
  assign n3543 = ~n3451 & n3542 ;
  assign n3544 = n2830 & ~n3543 ;
  assign n3545 = n3530 | n3544 ;
  buffer buf_n3546( .i (n3545), .o (n3546) );
  buffer buf_n3547( .i (n3546), .o (n3547) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  assign n3548 = n2320 | n3546 ;
  assign n3549 = ( ~n21 & n3333 ) | ( ~n21 & n3463 ) | ( n3333 & n3463 ) ;
  buffer buf_n3550( .i (n3549), .o (n3550) );
  assign n3555 = ( n2967 & n3340 ) | ( n2967 & ~n3550 ) | ( n3340 & ~n3550 ) ;
  buffer buf_n3556( .i (n3555), .o (n3556) );
  buffer buf_n3557( .i (n3556), .o (n3557) );
  buffer buf_n3558( .i (n3557), .o (n3558) );
  buffer buf_n3559( .i (n3558), .o (n3559) );
  assign n3560 = ( ~n3211 & n3425 ) | ( ~n3211 & n3556 ) | ( n3425 & n3556 ) ;
  buffer buf_n3561( .i (n3560), .o (n3561) );
  buffer buf_n3562( .i (n3561), .o (n3562) );
  buffer buf_n3551( .i (n3550), .o (n3551) );
  buffer buf_n3552( .i (n3551), .o (n3552) );
  buffer buf_n3553( .i (n3552), .o (n3553) );
  buffer buf_n3554( .i (n3553), .o (n3554) );
  assign n3563 = n3554 & n3561 ;
  assign n3564 = ( ~n3559 & n3562 ) | ( ~n3559 & n3563 ) | ( n3562 & n3563 ) ;
  assign n3565 = ~n3392 & n3564 ;
  assign n3566 = n3438 | n3565 ;
  assign n3567 = ~n2311 & n3444 ;
  assign n3568 = n3360 & n3567 ;
  assign n3569 = ~n3435 & n3568 ;
  assign n3570 = n3438 & ~n3569 ;
  assign n3571 = n3566 & ~n3570 ;
  assign n3572 = n2688 | n3571 ;
  assign n3573 = ~n594 & n3437 ;
  assign n3574 = ( n595 & n611 ) | ( n595 & n3573 ) | ( n611 & n3573 ) ;
  assign n3575 = ~n3375 & n3574 ;
  assign n3576 = n2688 & ~n3575 ;
  assign n3577 = n3572 & ~n3576 ;
  assign n3578 = n3423 | n3577 ;
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  assign n3579 = ( n610 & ~n2721 ) | ( n610 & n3392 ) | ( ~n2721 & n3392 ) ;
  assign n3580 = ~n2165 & n3579 ;
  assign n3581 = n3395 & n3580 ;
  buffer buf_n3582( .i (n1938), .o (n3582) );
  assign n3583 = ( ~n2967 & n3340 ) | ( ~n2967 & n3582 ) | ( n3340 & n3582 ) ;
  buffer buf_n3584( .i (n3583), .o (n3584) );
  buffer buf_n3585( .i (n3267), .o (n3585) );
  assign n3586 = ( ~n3310 & n3584 ) | ( ~n3310 & n3585 ) | ( n3584 & n3585 ) ;
  buffer buf_n3587( .i (n3586), .o (n3587) );
  assign n3590 = n2418 & n3587 ;
  buffer buf_n3591( .i (n3590), .o (n3591) );
  buffer buf_n3592( .i (n3591), .o (n3592) );
  buffer buf_n3588( .i (n3587), .o (n3588) );
  buffer buf_n3589( .i (n3588), .o (n3589) );
  assign n3593 = n3589 & ~n3591 ;
  assign n3594 = ( n2918 & ~n3592 ) | ( n2918 & n3593 ) | ( ~n3592 & n3593 ) ;
  assign n3595 = ( n2012 & ~n2685 ) | ( n2012 & n3594 ) | ( ~n2685 & n3594 ) ;
  assign n3596 = ( n568 & ~n3581 ) | ( n568 & n3595 ) | ( ~n3581 & n3595 ) ;
  assign n3597 = n3398 | n3596 ;
  assign n3598 = n3423 & n3597 ;
  assign n3599 = n3578 & ~n3598 ;
  assign n3600 = ( n453 & ~n2235 ) | ( n453 & n2607 ) | ( ~n2235 & n2607 ) ;
  buffer buf_n3601( .i (n3600), .o (n3601) );
  buffer buf_n3610( .i (n2780), .o (n3610) );
  assign n3611 = ~n1054 & n3610 ;
  buffer buf_n3612( .i (n3611), .o (n3612) );
  assign n3613 = ~n3601 & n3612 ;
  assign n3614 = n3114 & ~n3585 ;
  buffer buf_n3615( .i (n3614), .o (n3615) );
  assign n3618 = ( ~n1056 & n3612 ) | ( ~n1056 & n3615 ) | ( n3612 & n3615 ) ;
  buffer buf_n3619( .i (n3499), .o (n3619) );
  assign n3620 = ( n3613 & n3618 ) | ( n3613 & n3619 ) | ( n3618 & n3619 ) ;
  buffer buf_n3621( .i (n3177), .o (n3621) );
  buffer buf_n3622( .i (n3621), .o (n3622) );
  assign n3623 = n3620 | n3622 ;
  assign n3624 = n2607 & ~n3585 ;
  buffer buf_n3625( .i (n3624), .o (n3625) );
  buffer buf_n3626( .i (n3625), .o (n3626) );
  assign n3627 = n397 & n3626 ;
  assign n3628 = n3622 & ~n3627 ;
  assign n3629 = n3623 & ~n3628 ;
  buffer buf_n3630( .i (n3629), .o (n3630) );
  buffer buf_n3631( .i (n3630), .o (n3631) );
  assign n3632 = ( n653 & n2938 ) | ( n653 & n2982 ) | ( n2938 & n2982 ) ;
  buffer buf_n3633( .i (n3039), .o (n3633) );
  assign n3634 = ( n653 & ~n3268 ) | ( n653 & n3633 ) | ( ~n3268 & n3633 ) ;
  assign n3635 = ( n331 & ~n3632 ) | ( n331 & n3634 ) | ( ~n3632 & n3634 ) ;
  assign n3636 = n3212 & n3635 ;
  assign n3637 = n3024 & n3313 ;
  buffer buf_n3638( .i (n3637), .o (n3638) );
  assign n3642 = n3212 | n3638 ;
  assign n3643 = ~n3636 & n3642 ;
  assign n3644 = n3621 & ~n3643 ;
  assign n3645 = n371 & n2134 ;
  assign n3646 = n3621 | n3645 ;
  assign n3647 = ~n3644 & n3646 ;
  assign n3648 = ( n1114 & n2581 ) | ( n1114 & n2885 ) | ( n2581 & n2885 ) ;
  buffer buf_n3649( .i (n3648), .o (n3649) );
  assign n3654 = ( n2436 & n2922 ) | ( n2436 & ~n3649 ) | ( n2922 & ~n3649 ) ;
  buffer buf_n3655( .i (n3654), .o (n3655) );
  buffer buf_n3656( .i (n3655), .o (n3656) );
  buffer buf_n3657( .i (n3656), .o (n3657) );
  buffer buf_n3658( .i (n3657), .o (n3658) );
  buffer buf_n3659( .i (n3516), .o (n3659) );
  assign n3660 = ( n2978 & ~n3655 ) | ( n2978 & n3659 ) | ( ~n3655 & n3659 ) ;
  buffer buf_n3661( .i (n3660), .o (n3661) );
  buffer buf_n3662( .i (n3661), .o (n3662) );
  buffer buf_n3650( .i (n3649), .o (n3650) );
  buffer buf_n3651( .i (n3650), .o (n3651) );
  buffer buf_n3652( .i (n3651), .o (n3652) );
  buffer buf_n3653( .i (n3652), .o (n3653) );
  assign n3663 = ~n3653 & n3661 ;
  assign n3664 = ( n3658 & n3662 ) | ( n3658 & n3663 ) | ( n3662 & n3663 ) ;
  buffer buf_n3665( .i (n3664), .o (n3665) );
  buffer buf_n3666( .i (n3665), .o (n3666) );
  assign n3667 = n490 & n3267 ;
  buffer buf_n3668( .i (n3667), .o (n3668) );
  buffer buf_n3669( .i (n3668), .o (n3669) );
  assign n3670 = n3665 & n3669 ;
  assign n3671 = ( n3626 & n3666 ) | ( n3626 & n3670 ) | ( n3666 & n3670 ) ;
  buffer buf_n3672( .i (n3671), .o (n3672) );
  assign n3673 = ( ~n2165 & n3647 ) | ( ~n2165 & n3672 ) | ( n3647 & n3672 ) ;
  buffer buf_n3674( .i (n3633), .o (n3674) );
  assign n3675 = n2987 & ~n3674 ;
  assign n3676 = n523 & n3368 ;
  assign n3677 = ( n2119 & n3675 ) | ( n2119 & ~n3676 ) | ( n3675 & ~n3676 ) ;
  buffer buf_n3678( .i (n2226), .o (n3678) );
  assign n3679 = ( n73 & n131 ) | ( n73 & ~n3678 ) | ( n131 & ~n3678 ) ;
  buffer buf_n3680( .i (n3679), .o (n3680) );
  assign n3688 = ( ~n2285 & n2886 ) | ( ~n2285 & n3680 ) | ( n2886 & n3680 ) ;
  buffer buf_n3689( .i (n3688), .o (n3689) );
  assign n3692 = n2923 & ~n3689 ;
  buffer buf_n3693( .i (n3692), .o (n3693) );
  buffer buf_n3694( .i (n3693), .o (n3694) );
  buffer buf_n3690( .i (n3689), .o (n3690) );
  buffer buf_n3691( .i (n3690), .o (n3691) );
  assign n3695 = n3691 | n3693 ;
  assign n3696 = ( ~n3312 & n3694 ) | ( ~n3312 & n3695 ) | ( n3694 & n3695 ) ;
  buffer buf_n3697( .i (n3696), .o (n3697) );
  buffer buf_n3698( .i (n3697), .o (n3698) );
  assign n3699 = n3213 | n3697 ;
  assign n3700 = ( n3677 & n3698 ) | ( n3677 & n3699 ) | ( n3698 & n3699 ) ;
  assign n3701 = n3390 | n3700 ;
  assign n3702 = ( ~n3310 & n3368 ) | ( ~n3310 & n3674 ) | ( n3368 & n3674 ) ;
  buffer buf_n3703( .i (n3225), .o (n3703) );
  assign n3704 = ( ~n3039 & n3182 ) | ( ~n3039 & n3703 ) | ( n3182 & n3703 ) ;
  buffer buf_n3705( .i (n3704), .o (n3705) );
  buffer buf_n3715( .i (n2938), .o (n3715) );
  assign n3716 = ~n3705 & n3715 ;
  assign n3717 = n3702 & ~n3716 ;
  assign n3718 = ~n3499 & n3717 ;
  buffer buf_n3719( .i (n2734), .o (n3719) );
  assign n3720 = ~n3718 & n3719 ;
  assign n3721 = n3701 & ~n3720 ;
  buffer buf_n3722( .i (n3275), .o (n3722) );
  buffer buf_n3723( .i (n3722), .o (n3723) );
  assign n3724 = ( n3672 & n3721 ) | ( n3672 & n3723 ) | ( n3721 & n3723 ) ;
  assign n3725 = n3673 | n3724 ;
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  assign n3726 = n372 & n3511 ;
  assign n3727 = ( n588 & ~n1757 ) | ( n588 & n3726 ) | ( ~n1757 & n3726 ) ;
  assign n3728 = ~n589 & n3727 ;
  buffer buf_n3729( .i (n3728), .o (n3729) );
  assign n3730 = ( ~n3630 & n3725 ) | ( ~n3630 & n3729 ) | ( n3725 & n3729 ) ;
  assign n3731 = n3451 & ~n3729 ;
  assign n3732 = ( n3631 & n3730 ) | ( n3631 & ~n3731 ) | ( n3730 & ~n3731 ) ;
  assign n3733 = n3485 | n3732 ;
  buffer buf_n3734( .i (n2885), .o (n3734) );
  buffer buf_n3735( .i (n3734), .o (n3735) );
  assign n3736 = ( ~n3145 & n3332 ) | ( ~n3145 & n3735 ) | ( n3332 & n3735 ) ;
  assign n3737 = ( n2923 & ~n3463 ) | ( n2923 & n3736 ) | ( ~n3463 & n3736 ) ;
  buffer buf_n3738( .i (n3737), .o (n3738) );
  assign n3741 = n3182 & ~n3738 ;
  buffer buf_n3742( .i (n3741), .o (n3742) );
  buffer buf_n3743( .i (n3742), .o (n3743) );
  buffer buf_n3739( .i (n3738), .o (n3739) );
  buffer buf_n3740( .i (n3739), .o (n3740) );
  assign n3744 = n3740 | n3742 ;
  assign n3745 = ( ~n3318 & n3743 ) | ( ~n3318 & n3744 ) | ( n3743 & n3744 ) ;
  buffer buf_n3746( .i (n3213), .o (n3746) );
  assign n3747 = n3745 & n3746 ;
  assign n3748 = ( n2002 & ~n2717 ) | ( n2002 & n3715 ) | ( ~n2717 & n3715 ) ;
  assign n3749 = ( n2717 & n2987 ) | ( n2717 & ~n3715 ) | ( n2987 & ~n3715 ) ;
  assign n3750 = ( ~n3318 & n3748 ) | ( ~n3318 & n3749 ) | ( n3748 & n3749 ) ;
  assign n3751 = n3746 | n3750 ;
  assign n3752 = ( ~n2948 & n3747 ) | ( ~n2948 & n3751 ) | ( n3747 & n3751 ) ;
  assign n3753 = n3722 & ~n3752 ;
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n2519( .i (n2518), .o (n2519) );
  buffer buf_n3754( .i (n3268), .o (n3754) );
  assign n3755 = ( n3503 & ~n3585 ) | ( n3503 & n3754 ) | ( ~n3585 & n3754 ) ;
  assign n3756 = ~n3318 & n3755 ;
  assign n3757 = ( n1668 & n2519 ) | ( n1668 & ~n3756 ) | ( n2519 & ~n3756 ) ;
  assign n3758 = n3445 | n3757 ;
  assign n3759 = ~n3722 & n3758 ;
  assign n3760 = n3753 | n3759 ;
  assign n3761 = n2823 & ~n3760 ;
  assign n3762 = ( ~n1874 & n2924 ) | ( ~n1874 & n3261 ) | ( n2924 & n3261 ) ;
  buffer buf_n3763( .i (n3762), .o (n3763) );
  buffer buf_n3764( .i (n3763), .o (n3764) );
  buffer buf_n3765( .i (n3764), .o (n3765) );
  buffer buf_n3766( .i (n3261), .o (n3766) );
  buffer buf_n3767( .i (n3766), .o (n3767) );
  buffer buf_n3768( .i (n3340), .o (n3768) );
  assign n3769 = ( n3763 & ~n3767 ) | ( n3763 & n3768 ) | ( ~n3767 & n3768 ) ;
  assign n3770 = n1877 | n3769 ;
  buffer buf_n3771( .i (n3312), .o (n3771) );
  buffer buf_n3772( .i (n3771), .o (n3772) );
  assign n3773 = ( n3765 & n3770 ) | ( n3765 & ~n3772 ) | ( n3770 & ~n3772 ) ;
  assign n3774 = n3274 & n3773 ;
  assign n3775 = ( n2978 & ~n3225 ) | ( n2978 & n3261 ) | ( ~n3225 & n3261 ) ;
  buffer buf_n3776( .i (n3775), .o (n3776) );
  buffer buf_n3777( .i (n3776), .o (n3777) );
  buffer buf_n3783( .i (n3703), .o (n3783) );
  assign n3784 = n3776 & n3783 ;
  assign n3785 = ( ~n2629 & n3777 ) | ( ~n2629 & n3784 ) | ( n3777 & n3784 ) ;
  assign n3786 = ~n3772 & n3785 ;
  buffer buf_n3787( .i (n3135), .o (n3787) );
  assign n3788 = n3786 | n3787 ;
  assign n3789 = ~n3774 & n3788 ;
  assign n3790 = n3392 | n3789 ;
  buffer buf_n3791( .i (n2924), .o (n3791) );
  assign n3792 = ( ~n2627 & n3066 ) | ( ~n2627 & n3791 ) | ( n3066 & n3791 ) ;
  buffer buf_n3793( .i (n3792), .o (n3793) );
  buffer buf_n3794( .i (n3793), .o (n3794) );
  buffer buf_n3795( .i (n3794), .o (n3795) );
  buffer buf_n3796( .i (n3767), .o (n3796) );
  assign n3797 = ( ~n3771 & n3793 ) | ( ~n3771 & n3796 ) | ( n3793 & n3796 ) ;
  assign n3798 = ( ~n3135 & n3443 ) | ( ~n3135 & n3797 ) | ( n3443 & n3797 ) ;
  assign n3799 = n3795 & n3798 ;
  assign n3800 = ~n2948 & n3799 ;
  buffer buf_n3801( .i (n3619), .o (n3801) );
  assign n3802 = ~n3800 & n3801 ;
  assign n3803 = n3790 & ~n3802 ;
  assign n3804 = n2823 | n3803 ;
  buffer buf_n3805( .i (n2823), .o (n3805) );
  assign n3806 = ( n3761 & n3804 ) | ( n3761 & ~n3805 ) | ( n3804 & ~n3805 ) ;
  assign n3807 = ~n3398 & n3806 ;
  assign n3808 = n3485 & ~n3807 ;
  assign n3809 = n3733 & ~n3808 ;
  assign n3810 = n3599 | n3809 ;
  assign n3811 = ( ~n3547 & n3548 ) | ( ~n3547 & n3810 ) | ( n3548 & n3810 ) ;
  buffer buf_n3812( .i (n3811), .o (n3812) );
  buffer buf_n3813( .i (n3812), .o (n3813) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  assign n3814 = ~n24 & n3312 ;
  buffer buf_n3815( .i (n3814), .o (n3815) );
  buffer buf_n3816( .i (n3815), .o (n3816) );
  buffer buf_n3817( .i (n3816), .o (n3817) );
  buffer buf_n3818( .i (n3817), .o (n3818) );
  buffer buf_n3819( .i (n3818), .o (n3819) );
  buffer buf_n3820( .i (n3819), .o (n3820) );
  buffer buf_n3821( .i (n3820), .o (n3821) );
  assign n3823 = ~n2534 & n3375 ;
  assign n3824 = ( ~n960 & n3821 ) | ( ~n960 & n3823 ) | ( n3821 & n3823 ) ;
  assign n3825 = n2015 | n3824 ;
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  assign n3826 = ~n3425 & n3503 ;
  buffer buf_n3827( .i (n3826), .o (n3827) );
  buffer buf_n3828( .i (n3827), .o (n3828) );
  buffer buf_n3829( .i (n3828), .o (n3829) );
  buffer buf_n3830( .i (n3829), .o (n3830) );
  buffer buf_n3831( .i (n3830), .o (n3831) );
  assign n3832 = ( n1318 & n3820 ) | ( n1318 & ~n3831 ) | ( n3820 & ~n3831 ) ;
  assign n3833 = ~n2535 & n3832 ;
  assign n3834 = n2015 & ~n3833 ;
  assign n3835 = n3825 & ~n3834 ;
  buffer buf_n3836( .i (n3485), .o (n3836) );
  assign n3837 = n3835 | n3836 ;
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n2009( .i (n2008), .o (n2009) );
  assign n3838 = ~n2009 & n3805 ;
  assign n3839 = ( n518 & n803 ) | ( n518 & ~n3838 ) | ( n803 & ~n3838 ) ;
  buffer buf_n3840( .i (n3398), .o (n3840) );
  assign n3841 = n3839 & ~n3840 ;
  assign n3842 = n3836 & ~n3841 ;
  assign n3843 = n3837 & ~n3842 ;
  assign n3844 = n3489 | n3843 ;
  buffer buf_n2010( .i (n2009), .o (n2010) );
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n2722( .i (n2721), .o (n2722) );
  buffer buf_n2723( .i (n2722), .o (n2723) );
  buffer buf_n2724( .i (n2723), .o (n2724) );
  buffer buf_n2725( .i (n2724), .o (n2725) );
  buffer buf_n3845( .i (n3296), .o (n3845) );
  assign n3846 = ( ~n2725 & n2791 ) | ( ~n2725 & n3845 ) | ( n2791 & n3845 ) ;
  assign n3847 = ( ~n2725 & n3460 ) | ( ~n2725 & n3845 ) | ( n3460 & n3845 ) ;
  assign n3848 = ( n2011 & n3846 ) | ( n2011 & ~n3847 ) | ( n3846 & ~n3847 ) ;
  buffer buf_n3849( .i (n2558), .o (n3849) );
  assign n3850 = n374 & ~n3849 ;
  buffer buf_n3851( .i (n3850), .o (n3851) );
  assign n3852 = n1948 & n3851 ;
  buffer buf_n3853( .i (n3852), .o (n3853) );
  buffer buf_n3854( .i (n3853), .o (n3854) );
  buffer buf_n3855( .i (n3805), .o (n3855) );
  buffer buf_n3856( .i (n3855), .o (n3856) );
  assign n3857 = n3853 | n3856 ;
  assign n3858 = ( n3848 & n3854 ) | ( n3848 & n3857 ) | ( n3854 & n3857 ) ;
  assign n3859 = ~n3106 & n3858 ;
  assign n3860 = n3489 & ~n3859 ;
  assign n3861 = n3844 & ~n3860 ;
  assign n3862 = n3812 | n3861 ;
  assign n3863 = ( n360 & n3813 ) | ( n360 & n3862 ) | ( n3813 & n3862 ) ;
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n3864( .i (n3022), .o (n3864) );
  assign n3865 = n3791 | n3864 ;
  buffer buf_n3866( .i (n3865), .o (n3866) );
  buffer buf_n3867( .i (n3866), .o (n3867) );
  buffer buf_n3868( .i (n3867), .o (n3868) );
  buffer buf_n3869( .i (n3868), .o (n3869) );
  buffer buf_n3870( .i (n3869), .o (n3870) );
  buffer buf_n3871( .i (n3870), .o (n3871) );
  buffer buf_n3872( .i (n3871), .o (n3872) );
  buffer buf_n3873( .i (n3872), .o (n3873) );
  assign n3874 = ( ~n1086 & n1436 ) | ( ~n1086 & n3873 ) | ( n1436 & n3873 ) ;
  assign n3875 = n3845 & ~n3874 ;
  assign n3876 = ~n3840 & n3875 ;
  buffer buf_n3877( .i (n3876), .o (n3877) );
  buffer buf_n3878( .i (n3877), .o (n3878) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  assign n3879 = ( n710 & n1809 ) | ( n710 & n3423 ) | ( n1809 & n3423 ) ;
  assign n3880 = ~n2640 & n3879 ;
  buffer buf_n3507( .i (n3506), .o (n3507) );
  buffer buf_n3508( .i (n3507), .o (n3508) );
  buffer buf_n3509( .i (n3508), .o (n3509) );
  assign n3881 = ~n309 & n3504 ;
  assign n3882 = ( n3254 & n3444 ) | ( n3254 & n3881 ) | ( n3444 & n3881 ) ;
  buffer buf_n3883( .i (n3443), .o (n3883) );
  buffer buf_n3884( .i (n3883), .o (n3884) );
  assign n3885 = n3882 & ~n3884 ;
  buffer buf_n3886( .i (n3885), .o (n3886) );
  buffer buf_n3887( .i (n3886), .o (n3887) );
  buffer buf_n746( .i (n745), .o (n746) );
  assign n3888 = n746 | n3886 ;
  assign n3889 = ( n3509 & n3887 ) | ( n3509 & n3888 ) | ( n3887 & n3888 ) ;
  buffer buf_n3890( .i (n3889), .o (n3890) );
  buffer buf_n3891( .i (n3890), .o (n3891) );
  buffer buf_n3892( .i (n3451), .o (n3892) );
  assign n3893 = n3890 & n3892 ;
  buffer buf_n3894( .i (n2576), .o (n3894) );
  assign n3895 = n1402 & ~n3894 ;
  assign n3896 = ~n2099 & n3895 ;
  buffer buf_n3897( .i (n2403), .o (n3897) );
  buffer buf_n3898( .i (n3897), .o (n3898) );
  buffer buf_n3899( .i (n3898), .o (n3899) );
  assign n3900 = ( n3465 & n3864 ) | ( n3465 & ~n3899 ) | ( n3864 & ~n3899 ) ;
  assign n3901 = ( ~n3465 & n3791 ) | ( ~n3465 & n3864 ) | ( n3791 & n3864 ) ;
  assign n3902 = n3900 & ~n3901 ;
  assign n3903 = ( n3425 & n3754 ) | ( n3425 & n3902 ) | ( n3754 & n3902 ) ;
  assign n3904 = n21 & n3516 ;
  buffer buf_n3905( .i (n3904), .o (n3905) );
  assign n3910 = ( ~n2090 & n3791 ) | ( ~n2090 & n3905 ) | ( n3791 & n3905 ) ;
  buffer buf_n3911( .i (n3735), .o (n3911) );
  buffer buf_n3912( .i (n3911), .o (n3912) );
  buffer buf_n3913( .i (n3912), .o (n3913) );
  buffer buf_n3914( .i (n3913), .o (n3914) );
  assign n3915 = n3910 & ~n3914 ;
  assign n3916 = n3754 & n3915 ;
  buffer buf_n3917( .i (n20), .o (n3917) );
  buffer buf_n3918( .i (n3917), .o (n3918) );
  buffer buf_n3919( .i (n3918), .o (n3919) );
  buffer buf_n3920( .i (n3919), .o (n3920) );
  buffer buf_n3921( .i (n3920), .o (n3921) );
  buffer buf_n3922( .i (n3921), .o (n3922) );
  assign n3923 = ( n3903 & n3916 ) | ( n3903 & ~n3922 ) | ( n3916 & ~n3922 ) ;
  buffer buf_n3924( .i (n3923), .o (n3924) );
  buffer buf_n3925( .i (n3924), .o (n3925) );
  buffer buf_n3926( .i (n3925), .o (n3926) );
  buffer buf_n3927( .i (n3144), .o (n3927) );
  buffer buf_n3928( .i (n3056), .o (n3928) );
  buffer buf_n3929( .i (n1114), .o (n3929) );
  buffer buf_n3930( .i (n3929), .o (n3930) );
  assign n3931 = ( ~n3927 & n3928 ) | ( ~n3927 & n3930 ) | ( n3928 & n3930 ) ;
  buffer buf_n3932( .i (n3931), .o (n3932) );
  buffer buf_n3933( .i (n3932), .o (n3933) );
  buffer buf_n3934( .i (n3933), .o (n3934) );
  buffer buf_n3935( .i (n3934), .o (n3935) );
  buffer buf_n3936( .i (n3935), .o (n3936) );
  buffer buf_n3937( .i (n3936), .o (n3937) );
  assign n3938 = ( n3213 & n3253 ) | ( n3213 & ~n3504 ) | ( n3253 & ~n3504 ) ;
  assign n3939 = n3937 & ~n3938 ;
  assign n3940 = ( ~n3511 & n3924 ) | ( ~n3511 & n3939 ) | ( n3924 & n3939 ) ;
  assign n3941 = n3622 & ~n3940 ;
  assign n3942 = ( n3536 & n3926 ) | ( n3536 & ~n3941 ) | ( n3926 & ~n3941 ) ;
  assign n3943 = n3395 | n3942 ;
  assign n3944 = ( n1737 & n2948 ) | ( n1737 & ~n3621 ) | ( n2948 & ~n3621 ) ;
  assign n3945 = n1868 & n3944 ;
  assign n3946 = ~n3436 & n3945 ;
  assign n3947 = n3395 & ~n3946 ;
  assign n3948 = n3943 & ~n3947 ;
  assign n3949 = n3896 | n3948 ;
  assign n3950 = ( n3891 & ~n3893 ) | ( n3891 & n3949 ) | ( ~n3893 & n3949 ) ;
  buffer buf_n3951( .i (n3950), .o (n3951) );
  assign n3952 = ( ~n3877 & n3880 ) | ( ~n3877 & n3951 ) | ( n3880 & n3951 ) ;
  assign n3953 = n356 & ~n3951 ;
  assign n3954 = ( n3878 & n3952 ) | ( n3878 & ~n3953 ) | ( n3952 & ~n3953 ) ;
  buffer buf_n3955( .i (n3954), .o (n3955) );
  buffer buf_n3956( .i (n3955), .o (n3956) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  assign n3957 = n123 & n3955 ;
  buffer buf_n3958( .i (n3659), .o (n3958) );
  assign n3959 = ( n3582 & n3913 ) | ( n3582 & n3958 ) | ( n3913 & n3958 ) ;
  buffer buf_n3960( .i (n3959), .o (n3960) );
  buffer buf_n3961( .i (n3960), .o (n3961) );
  buffer buf_n3962( .i (n3961), .o (n3962) );
  buffer buf_n3963( .i (n3962), .o (n3963) );
  buffer buf_n3968( .i (n3177), .o (n3968) );
  assign n3969 = ( n2557 & ~n3963 ) | ( n2557 & n3968 ) | ( ~n3963 & n3968 ) ;
  buffer buf_n3970( .i (n3969), .o (n3970) );
  buffer buf_n3971( .i (n3970), .o (n3971) );
  buffer buf_n3972( .i (n3971), .o (n3972) );
  buffer buf_n3973( .i (n3972), .o (n3973) );
  buffer buf_n3974( .i (n3437), .o (n3974) );
  buffer buf_n3975( .i (n3801), .o (n3975) );
  assign n3976 = ( ~n3970 & n3974 ) | ( ~n3970 & n3975 ) | ( n3974 & n3975 ) ;
  buffer buf_n3977( .i (n3976), .o (n3977) );
  buffer buf_n3978( .i (n3977), .o (n3978) );
  buffer buf_n3964( .i (n3963), .o (n3964) );
  buffer buf_n3965( .i (n3964), .o (n3965) );
  buffer buf_n3966( .i (n3965), .o (n3966) );
  buffer buf_n3967( .i (n3966), .o (n3967) );
  assign n3979 = n3967 & ~n3977 ;
  assign n3980 = ( n3973 & n3978 ) | ( n3973 & ~n3979 ) | ( n3978 & ~n3979 ) ;
  assign n3981 = ( ~n236 & n264 ) | ( ~n236 & n3980 ) | ( n264 & n3980 ) ;
  assign n3982 = ~n3536 & n3849 ;
  buffer buf_n3983( .i (n3982), .o (n3983) );
  assign n3984 = ( n1548 & n3459 ) | ( n1548 & n3983 ) | ( n3459 & n3983 ) ;
  buffer buf_n3985( .i (n3974), .o (n3985) );
  buffer buf_n3986( .i (n3985), .o (n3986) );
  buffer buf_n3987( .i (n3894), .o (n3987) );
  assign n3988 = ( n3983 & n3986 ) | ( n3983 & n3987 ) | ( n3986 & n3987 ) ;
  assign n3989 = ( n1949 & n3984 ) | ( n1949 & ~n3988 ) | ( n3984 & ~n3988 ) ;
  assign n3990 = ( n236 & n264 ) | ( n236 & ~n3989 ) | ( n264 & ~n3989 ) ;
  assign n3991 = n3981 | n3990 ;
  buffer buf_n3992( .i (n3991), .o (n3992) );
  buffer buf_n3993( .i (n3992), .o (n3993) );
  buffer buf_n3088( .i (n3087), .o (n3088) );
  assign n3994 = ( n3088 & ~n3459 ) | ( n3088 & n3987 ) | ( ~n3459 & n3987 ) ;
  assign n3995 = ( ~n3088 & n3805 ) | ( ~n3088 & n3987 ) | ( n3805 & n3987 ) ;
  assign n3996 = n3994 & ~n3995 ;
  buffer buf_n3997( .i (n3996), .o (n3997) );
  buffer buf_n3998( .i (n3997), .o (n3998) );
  assign n3999 = ( n265 & n3836 ) | ( n265 & ~n3997 ) | ( n3836 & ~n3997 ) ;
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  assign n4000 = ( ~n627 & n2791 ) | ( ~n627 & n3460 ) | ( n2791 & n3460 ) ;
  buffer buf_n4001( .i (n3987), .o (n4001) );
  assign n4002 = ( n627 & ~n3845 ) | ( n627 & n4001 ) | ( ~n3845 & n4001 ) ;
  assign n4003 = n4000 & ~n4002 ;
  assign n4004 = n265 & n4003 ;
  assign n4005 = ( n3998 & n3999 ) | ( n3998 & n4004 ) | ( n3999 & n4004 ) ;
  assign n4006 = n3992 & n4005 ;
  assign n4007 = n3610 & ~n3921 ;
  buffer buf_n4008( .i (n4007), .o (n4008) );
  buffer buf_n4009( .i (n4008), .o (n4009) );
  buffer buf_n4010( .i (n4009), .o (n4010) );
  buffer buf_n4011( .i (n4010), .o (n4011) );
  buffer buf_n4012( .i (n4011), .o (n4012) );
  buffer buf_n4013( .i (n4012), .o (n4013) );
  buffer buf_n4014( .i (n4013), .o (n4014) );
  buffer buf_n4015( .i (n4014), .o (n4015) );
  buffer buf_n4016( .i (n4015), .o (n4016) );
  buffer buf_n4017( .i (n4016), .o (n4017) );
  buffer buf_n4018( .i (n4017), .o (n4018) );
  buffer buf_n4019( .i (n4018), .o (n4019) );
  assign n4020 = ( ~n3993 & n4006 ) | ( ~n3993 & n4019 ) | ( n4006 & n4019 ) ;
  buffer buf_n2236( .i (n2235), .o (n2236) );
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n4021( .i (n3429), .o (n4021) );
  assign n4022 = ( n397 & n2196 ) | ( n397 & ~n4021 ) | ( n2196 & ~n4021 ) ;
  buffer buf_n3165( .i (n3164), .o (n3165) );
  assign n4023 = n3165 & n4021 ;
  assign n4024 = ( n398 & ~n4022 ) | ( n398 & n4023 ) | ( ~n4022 & n4023 ) ;
  buffer buf_n4025( .i (n3622), .o (n4025) );
  assign n4026 = ( n3436 & n4024 ) | ( n3436 & ~n4025 ) | ( n4024 & ~n4025 ) ;
  buffer buf_n4027( .i (n825), .o (n4027) );
  assign n4028 = n2926 | n4027 ;
  buffer buf_n4029( .i (n4028), .o (n4029) );
  buffer buf_n4030( .i (n4029), .o (n4030) );
  buffer buf_n4031( .i (n4030), .o (n4031) );
  assign n4038 = n3922 & ~n4031 ;
  buffer buf_n4039( .i (n4038), .o (n4039) );
  assign n4046 = n2232 & n3659 ;
  buffer buf_n4047( .i (n4046), .o (n4047) );
  buffer buf_n4048( .i (n4047), .o (n4048) );
  buffer buf_n4049( .i (n4048), .o (n4049) );
  buffer buf_n4050( .i (n4049), .o (n4050) );
  buffer buf_n4051( .i (n4050), .o (n4051) );
  assign n4052 = n4039 & n4051 ;
  buffer buf_n4053( .i (n4052), .o (n4053) );
  assign n4060 = ~n4025 & n4053 ;
  buffer buf_n4061( .i (n3435), .o (n4061) );
  buffer buf_n4062( .i (n4061), .o (n4062) );
  assign n4063 = ( n4026 & n4060 ) | ( n4026 & ~n4062 ) | ( n4060 & ~n4062 ) ;
  buffer buf_n4064( .i (n4063), .o (n4064) );
  buffer buf_n4065( .i (n4064), .o (n4065) );
  buffer buf_n4066( .i (n4065), .o (n4066) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  assign n4067 = ( n756 & n1062 ) | ( n756 & n4064 ) | ( n1062 & n4064 ) ;
  assign n4068 = n2244 & ~n4067 ;
  assign n4069 = ( n2245 & n4066 ) | ( n2245 & ~n4068 ) | ( n4066 & ~n4068 ) ;
  buffer buf_n4070( .i (n4069), .o (n4070) );
  buffer buf_n4071( .i (n4070), .o (n4071) );
  assign n4072 = n357 & n4070 ;
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  assign n4073 = n713 & ~n1759 ;
  assign n4074 = n802 & n4073 ;
  buffer buf_n4075( .i (n4074), .o (n4075) );
  buffer buf_n4076( .i (n4075), .o (n4076) );
  buffer buf_n4077( .i (n4076), .o (n4077) );
  buffer buf_n4078( .i (n3503), .o (n4078) );
  assign n4079 = n2236 & ~n4078 ;
  buffer buf_n4080( .i (n4079), .o (n4080) );
  assign n4082 = ( n1156 & n4021 ) | ( n1156 & n4080 ) | ( n4021 & n4080 ) ;
  assign n4083 = ~n3437 & n4082 ;
  buffer buf_n4084( .i (n4083), .o (n4084) );
  buffer buf_n4085( .i (n4084), .o (n4085) );
  buffer buf_n4086( .i (n4085), .o (n4086) );
  assign n4087 = ( ~n3066 & n3582 ) | ( ~n3066 & n3958 ) | ( n3582 & n3958 ) ;
  buffer buf_n4088( .i (n4087), .o (n4088) );
  assign n4093 = ( n3139 & n3674 ) | ( n3139 & ~n4088 ) | ( n3674 & ~n4088 ) ;
  buffer buf_n4094( .i (n4093), .o (n4094) );
  buffer buf_n4095( .i (n4094), .o (n4095) );
  buffer buf_n4096( .i (n4095), .o (n4096) );
  buffer buf_n4097( .i (n4096), .o (n4097) );
  buffer buf_n4098( .i (n4078), .o (n4098) );
  assign n4099 = ( n3787 & n4094 ) | ( n3787 & ~n4098 ) | ( n4094 & ~n4098 ) ;
  buffer buf_n4100( .i (n4099), .o (n4100) );
  buffer buf_n4101( .i (n4100), .o (n4101) );
  buffer buf_n4089( .i (n4088), .o (n4089) );
  buffer buf_n4090( .i (n4089), .o (n4090) );
  buffer buf_n4091( .i (n4090), .o (n4091) );
  buffer buf_n4092( .i (n4091), .o (n4092) );
  assign n4102 = n4092 | n4100 ;
  assign n4103 = ( ~n4097 & n4101 ) | ( ~n4097 & n4102 ) | ( n4101 & n4102 ) ;
  buffer buf_n4104( .i (n4025), .o (n4104) );
  assign n4105 = ( ~n4084 & n4103 ) | ( ~n4084 & n4104 ) | ( n4103 & n4104 ) ;
  buffer buf_n4106( .i (n2534), .o (n4106) );
  assign n4107 = n4105 & ~n4106 ;
  assign n4108 = ( n3421 & ~n4086 ) | ( n3421 & n4107 ) | ( ~n4086 & n4107 ) ;
  assign n4109 = ( n3840 & ~n4075 ) | ( n3840 & n4108 ) | ( ~n4075 & n4108 ) ;
  assign n4110 = n265 & n4109 ;
  assign n4111 = ( n266 & n4077 ) | ( n266 & ~n4110 ) | ( n4077 & ~n4110 ) ;
  assign n4112 = ~n1940 & n3138 ;
  buffer buf_n4113( .i (n4112), .o (n4113) );
  assign n4114 = n1761 & n4113 ;
  assign n4115 = n3113 & ~n3313 ;
  buffer buf_n4116( .i (n4115), .o (n4116) );
  assign n4121 = ( ~n1942 & n4113 ) | ( ~n1942 & n4116 ) | ( n4113 & n4116 ) ;
  buffer buf_n4122( .i (n3772), .o (n4122) );
  assign n4123 = ( n4114 & n4121 ) | ( n4114 & ~n4122 ) | ( n4121 & ~n4122 ) ;
  buffer buf_n4124( .i (n4123), .o (n4124) );
  buffer buf_n4125( .i (n4124), .o (n4125) );
  assign n4126 = ( n1559 & n2462 ) | ( n1559 & ~n2780 ) | ( n2462 & ~n2780 ) ;
  buffer buf_n4127( .i (n4126), .o (n4127) );
  buffer buf_n4128( .i (n4127), .o (n4128) );
  buffer buf_n4129( .i (n4128), .o (n4129) );
  buffer buf_n4130( .i (n4129), .o (n4130) );
  assign n4135 = n4124 & n4130 ;
  assign n4136 = ( n71 & n99 ) | ( n71 & n159 ) | ( n99 & n159 ) ;
  buffer buf_n4137( .i (n4136), .o (n4137) );
  assign n4147 = ( n101 & ~n131 ) | ( n101 & n4137 ) | ( ~n131 & n4137 ) ;
  buffer buf_n4148( .i (n4147), .o (n4148) );
  assign n4151 = n2904 & ~n4148 ;
  buffer buf_n4152( .i (n4151), .o (n4152) );
  buffer buf_n4153( .i (n4152), .o (n4153) );
  buffer buf_n4149( .i (n4148), .o (n4149) );
  buffer buf_n4150( .i (n4149), .o (n4150) );
  assign n4154 = n4150 | n4152 ;
  assign n4155 = ( ~n2926 & n4153 ) | ( ~n2926 & n4154 ) | ( n4153 & n4154 ) ;
  assign n4156 = ( n3582 & ~n3703 ) | ( n3582 & n4155 ) | ( ~n3703 & n4155 ) ;
  buffer buf_n4157( .i (n4156), .o (n4157) );
  buffer buf_n4158( .i (n4157), .o (n4158) );
  buffer buf_n4159( .i (n4158), .o (n4159) );
  buffer buf_n4160( .i (n4159), .o (n4160) );
  assign n4161 = n3754 & n4157 ;
  buffer buf_n4162( .i (n4161), .o (n4162) );
  buffer buf_n4163( .i (n4162), .o (n4163) );
  assign n4164 = ( n3254 & n3429 ) | ( n3254 & ~n4162 ) | ( n3429 & ~n4162 ) ;
  assign n4165 = ( n4160 & n4163 ) | ( n4160 & ~n4164 ) | ( n4163 & ~n4164 ) ;
  assign n4166 = ( n71 & n99 ) | ( n71 & ~n129 ) | ( n99 & ~n129 ) ;
  buffer buf_n4167( .i (n4166), .o (n4167) );
  buffer buf_n4182( .i (n129), .o (n4182) );
  buffer buf_n4183( .i (n4182), .o (n4183) );
  assign n4184 = ( n3678 & n4167 ) | ( n3678 & n4183 ) | ( n4167 & n4183 ) ;
  buffer buf_n4185( .i (n4184), .o (n4185) );
  buffer buf_n4186( .i (n4185), .o (n4186) );
  buffer buf_n4187( .i (n4186), .o (n4187) );
  buffer buf_n4188( .i (n4187), .o (n4188) );
  assign n4189 = ( n2904 & n3734 ) | ( n2904 & n4185 ) | ( n3734 & n4185 ) ;
  buffer buf_n4190( .i (n4189), .o (n4190) );
  buffer buf_n4191( .i (n4190), .o (n4191) );
  buffer buf_n4168( .i (n4167), .o (n4168) );
  buffer buf_n4169( .i (n4168), .o (n4169) );
  buffer buf_n4170( .i (n4169), .o (n4170) );
  buffer buf_n4171( .i (n4170), .o (n4171) );
  assign n4192 = ~n4171 & n4190 ;
  assign n4193 = ( ~n4188 & n4191 ) | ( ~n4188 & n4192 ) | ( n4191 & n4192 ) ;
  assign n4194 = n3766 & ~n4193 ;
  buffer buf_n4195( .i (n2925), .o (n4195) );
  assign n4196 = n1731 & ~n4195 ;
  assign n4197 = n3766 | n4196 ;
  assign n4198 = ~n4194 & n4197 ;
  buffer buf_n4199( .i (n3138), .o (n4199) );
  assign n4200 = n4198 | n4199 ;
  assign n4201 = ~n583 & n4047 ;
  assign n4202 = n4199 & ~n4201 ;
  assign n4203 = n4200 & ~n4202 ;
  assign n4204 = ~n3746 & n4203 ;
  assign n4205 = ( n767 & n2328 ) | ( n767 & n2885 ) | ( n2328 & n2885 ) ;
  buffer buf_n4206( .i (n4205), .o (n4206) );
  buffer buf_n4207( .i (n4206), .o (n4207) );
  buffer buf_n4208( .i (n4207), .o (n4208) );
  assign n4209 = ( n3332 & n3928 ) | ( n3332 & ~n4206 ) | ( n3928 & ~n4206 ) ;
  assign n4210 = n770 | n4209 ;
  assign n4211 = ( n3912 & ~n4208 ) | ( n3912 & n4210 ) | ( ~n4208 & n4210 ) ;
  buffer buf_n4212( .i (n4211), .o (n4212) );
  buffer buf_n4213( .i (n4212), .o (n4213) );
  buffer buf_n4214( .i (n4027), .o (n4214) );
  buffer buf_n4215( .i (n4214), .o (n4215) );
  buffer buf_n4216( .i (n4195), .o (n4216) );
  buffer buf_n4217( .i (n4216), .o (n4217) );
  assign n4218 = ( n4212 & ~n4215 ) | ( n4212 & n4217 ) | ( ~n4215 & n4217 ) ;
  assign n4219 = n1685 & ~n2191 ;
  assign n4220 = ~n4215 & n4219 ;
  assign n4221 = ( ~n4213 & n4218 ) | ( ~n4213 & n4220 ) | ( n4218 & n4220 ) ;
  buffer buf_n4222( .i (n100), .o (n4222) );
  assign n4223 = n3678 & n4222 ;
  buffer buf_n4224( .i (n4223), .o (n4224) );
  buffer buf_n4225( .i (n4224), .o (n4225) );
  buffer buf_n4226( .i (n4225), .o (n4226) );
  assign n4238 = ( n3333 & ~n3911 ) | ( n3333 & n4226 ) | ( ~n3911 & n4226 ) ;
  assign n4239 = ( n3332 & n3928 ) | ( n3332 & ~n4225 ) | ( n3928 & ~n4225 ) ;
  assign n4240 = ( n2925 & ~n3911 ) | ( n2925 & n4239 ) | ( ~n3911 & n4239 ) ;
  assign n4241 = ~n4238 & n4240 ;
  buffer buf_n4242( .i (n4241), .o (n4242) );
  buffer buf_n4243( .i (n4242), .o (n4243) );
  buffer buf_n4244( .i (n3958), .o (n4244) );
  assign n4245 = ( ~n4215 & n4242 ) | ( ~n4215 & n4244 ) | ( n4242 & n4244 ) ;
  buffer buf_n2876( .i (n2875), .o (n2876) );
  buffer buf_n2877( .i (n2876), .o (n2877) );
  buffer buf_n4246( .i (n2905), .o (n4246) );
  assign n4247 = ( n2188 & n2877 ) | ( n2188 & ~n4246 ) | ( n2877 & ~n4246 ) ;
  buffer buf_n4248( .i (n4247), .o (n4248) );
  buffer buf_n4249( .i (n4248), .o (n4249) );
  assign n4267 = ( n391 & n3912 ) | ( n391 & n4248 ) | ( n3912 & n4248 ) ;
  assign n4268 = ~n4249 & n4267 ;
  assign n4269 = n4215 & n4268 ;
  assign n4270 = ( n4243 & ~n4245 ) | ( n4243 & n4269 ) | ( ~n4245 & n4269 ) ;
  assign n4271 = n4221 | n4270 ;
  assign n4272 = n3746 & n4271 ;
  assign n4273 = n4204 | n4272 ;
  assign n4274 = n4165 | n4273 ;
  assign n4275 = ( n4125 & ~n4135 ) | ( n4125 & n4274 ) | ( ~n4135 & n4274 ) ;
  assign n4276 = ( n233 & ~n4062 ) | ( n233 & n4275 ) | ( ~n4062 & n4275 ) ;
  assign n4277 = ( n44 & n100 ) | ( n44 & n2226 ) | ( n100 & n2226 ) ;
  buffer buf_n4278( .i (n4277), .o (n4278) );
  assign n4291 = ( n2228 & n3187 ) | ( n2228 & ~n4278 ) | ( n3187 & ~n4278 ) ;
  buffer buf_n4292( .i (n4291), .o (n4292) );
  buffer buf_n4293( .i (n4292), .o (n4293) );
  buffer buf_n4279( .i (n4278), .o (n4279) );
  buffer buf_n4280( .i (n4279), .o (n4280) );
  assign n4294 = ( ~n4246 & n4280 ) | ( ~n4246 & n4292 ) | ( n4280 & n4292 ) ;
  buffer buf_n4295( .i (n2436), .o (n4295) );
  assign n4296 = ( n4293 & n4294 ) | ( n4293 & ~n4295 ) | ( n4294 & ~n4295 ) ;
  buffer buf_n4297( .i (n4296), .o (n4297) );
  buffer buf_n4298( .i (n4297), .o (n4298) );
  assign n4299 = ( n3703 & ~n3913 ) | ( n3703 & n4297 ) | ( ~n3913 & n4297 ) ;
  assign n4300 = n303 | n3928 ;
  assign n4301 = ( n3333 & n4295 ) | ( n3333 & ~n4300 ) | ( n4295 & ~n4300 ) ;
  assign n4302 = ~n4195 & n4301 ;
  buffer buf_n4303( .i (n2959), .o (n4303) );
  buffer buf_n4304( .i (n4303), .o (n4304) );
  assign n4305 = n4302 & ~n4304 ;
  assign n4306 = ( n4298 & ~n4299 ) | ( n4298 & n4305 ) | ( ~n4299 & n4305 ) ;
  buffer buf_n4307( .i (n4306), .o (n4307) );
  buffer buf_n4308( .i (n4307), .o (n4308) );
  buffer buf_n4309( .i (n4308), .o (n4309) );
  buffer buf_n4310( .i (n4199), .o (n4310) );
  assign n4311 = ( n3668 & n4307 ) | ( n3668 & ~n4310 ) | ( n4307 & ~n4310 ) ;
  assign n4312 = n2931 & ~n4311 ;
  assign n4313 = ( n2932 & n4309 ) | ( n2932 & ~n4312 ) | ( n4309 & ~n4312 ) ;
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  assign n4314 = ( ~n3000 & n4195 ) | ( ~n3000 & n4303 ) | ( n4195 & n4303 ) ;
  buffer buf_n4315( .i (n4295), .o (n4315) );
  buffer buf_n4316( .i (n4246), .o (n4316) );
  buffer buf_n4317( .i (n4316), .o (n4317) );
  assign n4318 = ( ~n3000 & n4315 ) | ( ~n3000 & n4317 ) | ( n4315 & n4317 ) ;
  assign n4319 = ( n2300 & n4314 ) | ( n2300 & ~n4318 ) | ( n4314 & ~n4318 ) ;
  assign n4320 = ( n3633 & n3914 ) | ( n3633 & n4319 ) | ( n3914 & n4319 ) ;
  buffer buf_n4321( .i (n4320), .o (n4321) );
  assign n4322 = ( ~n3772 & n4310 ) | ( ~n3772 & n4321 ) | ( n4310 & n4321 ) ;
  assign n4323 = ( n3253 & n4310 ) | ( n3253 & ~n4321 ) | ( n4310 & ~n4321 ) ;
  assign n4324 = n4322 & ~n4323 ;
  buffer buf_n4325( .i (n4324), .o (n4325) );
  assign n4326 = ( ~n3801 & n4313 ) | ( ~n3801 & n4325 ) | ( n4313 & n4325 ) ;
  buffer buf_n2878( .i (n2877), .o (n2878) );
  buffer buf_n2879( .i (n2878), .o (n2879) );
  buffer buf_n2880( .i (n2879), .o (n2880) );
  buffer buf_n2881( .i (n2880), .o (n2881) );
  buffer buf_n2882( .i (n2881), .o (n2882) );
  buffer buf_n2883( .i (n2882), .o (n2883) );
  assign n4327 = ( n3610 & ~n3674 ) | ( n3610 & n3866 ) | ( ~n3674 & n3866 ) ;
  assign n4328 = ( n3610 & ~n3796 ) | ( n3610 & n3866 ) | ( ~n3796 & n3866 ) ;
  assign n4329 = ( n2883 & ~n4327 ) | ( n2883 & n4328 ) | ( ~n4327 & n4328 ) ;
  assign n4330 = n4214 & n4304 ;
  buffer buf_n4331( .i (n4330), .o (n4331) );
  buffer buf_n4337( .i (n3783), .o (n4337) );
  assign n4338 = ~n4331 & n4337 ;
  buffer buf_n4339( .i (n4338), .o (n4339) );
  assign n4340 = n4329 & n4339 ;
  buffer buf_n4332( .i (n4331), .o (n4332) );
  buffer buf_n4333( .i (n4332), .o (n4333) );
  buffer buf_n4138( .i (n4137), .o (n4138) );
  buffer buf_n4139( .i (n4138), .o (n4139) );
  buffer buf_n4140( .i (n4139), .o (n4140) );
  buffer buf_n4141( .i (n4140), .o (n4141) );
  buffer buf_n4142( .i (n4141), .o (n4142) );
  buffer buf_n4143( .i (n4142), .o (n4143) );
  buffer buf_n4144( .i (n4143), .o (n4144) );
  buffer buf_n4145( .i (n4144), .o (n4145) );
  buffer buf_n4146( .i (n4145), .o (n4146) );
  buffer buf_n4341( .i (n3633), .o (n4341) );
  assign n4342 = ( n3771 & n3796 ) | ( n3771 & n4341 ) | ( n3796 & n4341 ) ;
  buffer buf_n4343( .i (n3864), .o (n4343) );
  assign n4344 = ~n4217 & n4343 ;
  buffer buf_n4345( .i (n4344), .o (n4345) );
  assign n4355 = ( n4146 & ~n4342 ) | ( n4146 & n4345 ) | ( ~n4342 & n4345 ) ;
  assign n4356 = ( ~n4333 & n4339 ) | ( ~n4333 & n4355 ) | ( n4339 & n4355 ) ;
  assign n4357 = ( n4021 & n4340 ) | ( n4021 & n4356 ) | ( n4340 & n4356 ) ;
  assign n4358 = ( n3801 & n4325 ) | ( n3801 & n4357 ) | ( n4325 & n4357 ) ;
  assign n4359 = n4326 | n4358 ;
  buffer buf_n4360( .i (n232), .o (n4360) );
  assign n4361 = ( n4062 & ~n4359 ) | ( n4062 & n4360 ) | ( ~n4359 & n4360 ) ;
  assign n4362 = n4276 & ~n4361 ;
  buffer buf_n4363( .i (n4362), .o (n4363) );
  buffer buf_n4364( .i (n4363), .o (n4364) );
  buffer buf_n4365( .i (n4364), .o (n4365) );
  assign n4366 = ( n716 & n1246 ) | ( n716 & n4363 ) | ( n1246 & n4363 ) ;
  assign n4367 = n600 & ~n4366 ;
  assign n4368 = ( n601 & n4365 ) | ( n601 & ~n4367 ) | ( n4365 & ~n4367 ) ;
  assign n4369 = n4111 | n4368 ;
  assign n4370 = ( n4071 & ~n4072 ) | ( n4071 & n4369 ) | ( ~n4072 & n4369 ) ;
  assign n4371 = n4020 | n4370 ;
  assign n4372 = ( n3956 & ~n3957 ) | ( n3956 & n4371 ) | ( ~n3957 & n4371 ) ;
  buffer buf_n4250( .i (n4249), .o (n4250) );
  buffer buf_n4251( .i (n4250), .o (n4251) );
  buffer buf_n4252( .i (n4251), .o (n4252) );
  buffer buf_n4253( .i (n4252), .o (n4253) );
  buffer buf_n4254( .i (n4253), .o (n4254) );
  buffer buf_n4255( .i (n4254), .o (n4255) );
  buffer buf_n4256( .i (n4255), .o (n4256) );
  buffer buf_n4257( .i (n4256), .o (n4257) );
  buffer buf_n4258( .i (n4257), .o (n4258) );
  buffer buf_n4259( .i (n4258), .o (n4259) );
  buffer buf_n4260( .i (n4259), .o (n4260) );
  buffer buf_n4261( .i (n4260), .o (n4261) );
  buffer buf_n4262( .i (n4261), .o (n4262) );
  buffer buf_n4263( .i (n4262), .o (n4263) );
  buffer buf_n4264( .i (n4263), .o (n4264) );
  buffer buf_n4265( .i (n4264), .o (n4265) );
  buffer buf_n4266( .i (n4265), .o (n4266) );
  buffer buf_n4227( .i (n4226), .o (n4227) );
  buffer buf_n4228( .i (n4227), .o (n4228) );
  buffer buf_n4229( .i (n4228), .o (n4229) );
  buffer buf_n4230( .i (n4229), .o (n4230) );
  buffer buf_n4231( .i (n4230), .o (n4231) );
  buffer buf_n4232( .i (n4231), .o (n4232) );
  buffer buf_n4233( .i (n4232), .o (n4233) );
  buffer buf_n4234( .i (n4233), .o (n4234) );
  buffer buf_n4235( .i (n4234), .o (n4235) );
  buffer buf_n4373( .i (n4217), .o (n4373) );
  assign n4374 = n1478 & ~n4373 ;
  buffer buf_n4375( .i (n4374), .o (n4375) );
  buffer buf_n4376( .i (n4375), .o (n4376) );
  assign n4377 = ( n3429 & ~n4098 ) | ( n3429 & n4375 ) | ( ~n4098 & n4375 ) ;
  assign n4378 = ( n1481 & n4376 ) | ( n1481 & n4377 ) | ( n4376 & n4377 ) ;
  assign n4379 = n2558 & n4378 ;
  buffer buf_n2494( .i (n2493), .o (n2494) );
  buffer buf_n2495( .i (n2494), .o (n2495) );
  buffer buf_n2496( .i (n2495), .o (n2496) );
  buffer buf_n2497( .i (n2496), .o (n2497) );
  buffer buf_n2498( .i (n2497), .o (n2498) );
  buffer buf_n4380( .i (n4214), .o (n4380) );
  assign n4381 = n3783 | n4380 ;
  buffer buf_n4382( .i (n4381), .o (n4382) );
  buffer buf_n4383( .i (n4382), .o (n4383) );
  buffer buf_n4384( .i (n4383), .o (n4384) );
  assign n4388 = ( n2498 & ~n3097 ) | ( n2498 & n4384 ) | ( ~n3097 & n4384 ) ;
  buffer buf_n4389( .i (n3254), .o (n4389) );
  buffer buf_n4390( .i (n4389), .o (n4390) );
  assign n4391 = ( n3722 & ~n4388 ) | ( n3722 & n4390 ) | ( ~n4388 & n4390 ) ;
  assign n4392 = ( ~n4235 & n4379 ) | ( ~n4235 & n4391 ) | ( n4379 & n4391 ) ;
  buffer buf_n4393( .i (n3366), .o (n4393) );
  buffer buf_n4394( .i (n4393), .o (n4394) );
  assign n4395 = ~n4392 & n4394 ;
  assign n4396 = ( ~n3783 & n4244 ) | ( ~n3783 & n4343 ) | ( n4244 & n4343 ) ;
  buffer buf_n4397( .i (n4396), .o (n4397) );
  buffer buf_n4398( .i (n4397), .o (n4398) );
  buffer buf_n4399( .i (n4398), .o (n4399) );
  buffer buf_n4400( .i (n4399), .o (n4400) );
  assign n4401 = ~n4078 & n4397 ;
  buffer buf_n4402( .i (n4401), .o (n4402) );
  buffer buf_n4403( .i (n4402), .o (n4403) );
  buffer buf_n4404( .i (n3787), .o (n4404) );
  buffer buf_n4405( .i (n4337), .o (n4405) );
  buffer buf_n4406( .i (n4405), .o (n4406) );
  buffer buf_n4407( .i (n4406), .o (n4407) );
  assign n4408 = ( n4402 & ~n4404 ) | ( n4402 & n4407 ) | ( ~n4404 & n4407 ) ;
  assign n4409 = ( n4400 & n4403 ) | ( n4400 & n4408 ) | ( n4403 & n4408 ) ;
  assign n4410 = n3974 & n4409 ;
  assign n4411 = n4394 | n4410 ;
  assign n4412 = ~n4395 & n4411 ;
  assign n4413 = ( ~n2757 & n3460 ) | ( ~n2757 & n4412 ) | ( n3460 & n4412 ) ;
  assign n4414 = ~n455 & n3787 ;
  buffer buf_n4415( .i (n4341), .o (n4415) );
  assign n4416 = ( ~n454 & n3212 ) | ( ~n454 & n4415 ) | ( n3212 & n4415 ) ;
  buffer buf_n4417( .i (n4373), .o (n4417) );
  buffer buf_n4418( .i (n4417), .o (n4418) );
  assign n4419 = ( n2195 & ~n4416 ) | ( n2195 & n4418 ) | ( ~n4416 & n4418 ) ;
  assign n4420 = ( ~n4404 & n4414 ) | ( ~n4404 & n4419 ) | ( n4414 & n4419 ) ;
  buffer buf_n4421( .i (n4310), .o (n4421) );
  buffer buf_n4422( .i (n4421), .o (n4422) );
  buffer buf_n4423( .i (n4422), .o (n4423) );
  assign n4424 = n4420 | n4423 ;
  buffer buf_n4425( .i (n3796), .o (n4425) );
  assign n4426 = ~n1754 & n4425 ;
  buffer buf_n4427( .i (n4426), .o (n4427) );
  assign n4429 = ~n4404 & n4427 ;
  assign n4430 = n4423 & ~n4429 ;
  assign n4431 = n4424 & ~n4430 ;
  assign n4432 = n3894 & n4431 ;
  assign n4433 = ( n4199 & n4341 ) | ( n4199 & ~n4373 ) | ( n4341 & ~n4373 ) ;
  buffer buf_n4434( .i (n4433), .o (n4434) );
  buffer buf_n4435( .i (n4425), .o (n4435) );
  assign n4436 = ( n4418 & n4434 ) | ( n4418 & n4435 ) | ( n4434 & n4435 ) ;
  assign n4437 = n4418 & n4434 ;
  assign n4438 = n4434 | n4435 ;
  assign n4439 = ( ~n4436 & n4437 ) | ( ~n4436 & n4438 ) | ( n4437 & n4438 ) ;
  buffer buf_n4440( .i (n4407), .o (n4440) );
  assign n4441 = ~n4439 & n4440 ;
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n2152( .i (n2151), .o (n2152) );
  assign n4442 = ( n441 & n633 ) | ( n441 & ~n2152 ) | ( n633 & ~n2152 ) ;
  buffer buf_n4443( .i (n4442), .o (n4443) );
  assign n4446 = n4389 & n4443 ;
  assign n4447 = n4440 | n4446 ;
  assign n4448 = ~n4441 & n4447 ;
  assign n4449 = n3894 | n4448 ;
  buffer buf_n4450( .i (n3975), .o (n4450) );
  buffer buf_n4451( .i (n4450), .o (n4451) );
  assign n4452 = ( n4432 & n4449 ) | ( n4432 & ~n4451 ) | ( n4449 & ~n4451 ) ;
  buffer buf_n4453( .i (n3459), .o (n4453) );
  assign n4454 = ( n2757 & n4452 ) | ( n2757 & n4453 ) | ( n4452 & n4453 ) ;
  assign n4455 = n4413 & n4454 ;
  buffer buf_n4456( .i (n4455), .o (n4456) );
  buffer buf_n4457( .i (n4456), .o (n4457) );
  assign n4458 = n3106 & n4456 ;
  buffer buf_n4032( .i (n4031), .o (n4032) );
  buffer buf_n4033( .i (n4032), .o (n4033) );
  buffer buf_n4034( .i (n4033), .o (n4034) );
  assign n4459 = n3539 & ~n4034 ;
  buffer buf_n4460( .i (n4459), .o (n4460) );
  buffer buf_n4461( .i (n4460), .o (n4461) );
  buffer buf_n4462( .i (n4404), .o (n4462) );
  assign n4463 = ( n2096 & n3098 ) | ( n2096 & n4462 ) | ( n3098 & n4462 ) ;
  assign n4464 = ~n2097 & n4463 ;
  assign n4465 = n4460 | n4464 ;
  buffer buf_n4466( .i (n4062), .o (n4466) );
  assign n4467 = ( n4461 & n4465 ) | ( n4461 & ~n4466 ) | ( n4465 & ~n4466 ) ;
  buffer buf_n4468( .i (n4467), .o (n4468) );
  buffer buf_n4469( .i (n4468), .o (n4469) );
  buffer buf_n4470( .i (n4453), .o (n4470) );
  assign n4471 = ( n2318 & n4468 ) | ( n2318 & n4470 ) | ( n4468 & n4470 ) ;
  assign n4472 = ( n439 & ~n1361 ) | ( n439 & n2516 ) | ( ~n1361 & n2516 ) ;
  buffer buf_n4473( .i (n4472), .o (n4473) );
  buffer buf_n4474( .i (n3715), .o (n4474) );
  assign n4475 = n4473 & n4474 ;
  buffer buf_n4476( .i (n4475), .o (n4476) );
  buffer buf_n4477( .i (n4476), .o (n4477) );
  buffer buf_n4478( .i (n1115), .o (n4478) );
  assign n4479 = n2904 & n4478 ;
  buffer buf_n4480( .i (n4479), .o (n4480) );
  assign n4489 = ( n3516 & ~n4316 ) | ( n3516 & n4480 ) | ( ~n4316 & n4480 ) ;
  buffer buf_n4490( .i (n4489), .o (n4490) );
  buffer buf_n4491( .i (n4490), .o (n4491) );
  buffer buf_n4492( .i (n4491), .o (n4492) );
  assign n4493 = ( n3766 & ~n4216 ) | ( n3766 & n4490 ) | ( ~n4216 & n4490 ) ;
  buffer buf_n4494( .i (n4304), .o (n4494) );
  assign n4495 = ( n4244 & ~n4493 ) | ( n4244 & n4494 ) | ( ~n4493 & n4494 ) ;
  assign n4496 = ~n4492 & n4495 ;
  assign n4497 = n4474 | n4496 ;
  assign n4498 = n1042 & n4317 ;
  buffer buf_n4499( .i (n4498), .o (n4499) );
  assign n4509 = n3000 | n4317 ;
  buffer buf_n4510( .i (n4509), .o (n4510) );
  assign n4519 = ~n4499 & n4510 ;
  assign n4520 = n4373 & ~n4519 ;
  assign n4521 = n4474 & ~n4520 ;
  assign n4522 = n4497 & ~n4521 ;
  buffer buf_n4523( .i (n4217), .o (n4523) );
  assign n4524 = n1012 & ~n4523 ;
  assign n4525 = n3922 & n4524 ;
  buffer buf_n4526( .i (n4525), .o (n4526) );
  assign n4527 = ( ~n4476 & n4522 ) | ( ~n4476 & n4526 ) | ( n4522 & n4526 ) ;
  assign n4528 = n3511 & ~n4526 ;
  assign n4529 = ( n4477 & n4527 ) | ( n4477 & ~n4528 ) | ( n4527 & ~n4528 ) ;
  assign n4530 = n3849 & ~n4529 ;
  buffer buf_n3002( .i (n3001), .o (n3002) );
  buffer buf_n3003( .i (n3002), .o (n3003) );
  buffer buf_n3004( .i (n3003), .o (n3004) );
  buffer buf_n4531( .i (n2999), .o (n4531) );
  assign n4532 = ( ~n2761 & n4315 ) | ( ~n2761 & n4531 ) | ( n4315 & n4531 ) ;
  buffer buf_n4533( .i (n4532), .o (n4533) );
  buffer buf_n4534( .i (n4533), .o (n4534) );
  buffer buf_n4535( .i (n4534), .o (n4535) );
  buffer buf_n4536( .i (n4216), .o (n4536) );
  assign n4537 = ( n3768 & n4533 ) | ( n3768 & ~n4536 ) | ( n4533 & ~n4536 ) ;
  buffer buf_n4538( .i (n4244), .o (n4538) );
  assign n4539 = ( n3003 & n4537 ) | ( n3003 & ~n4538 ) | ( n4537 & ~n4538 ) ;
  assign n4540 = ( ~n3004 & n4535 ) | ( ~n3004 & n4539 ) | ( n4535 & n4539 ) ;
  assign n4541 = n4435 & n4540 ;
  assign n4542 = ( n3898 & n4303 ) | ( n3898 & n4315 ) | ( n4303 & n4315 ) ;
  buffer buf_n4543( .i (n4542), .o (n4543) );
  buffer buf_n4544( .i (n4543), .o (n4544) );
  assign n4548 = ~n4536 & n4543 ;
  assign n4549 = ( ~n606 & n4544 ) | ( ~n606 & n4548 ) | ( n4544 & n4548 ) ;
  assign n4550 = n4078 & n4549 ;
  assign n4551 = n4435 | n4550 ;
  assign n4552 = ~n4541 & n4551 ;
  assign n4553 = ~n3435 & n4552 ;
  assign n4554 = n3849 | n4553 ;
  assign n4555 = ~n4530 & n4554 ;
  assign n4556 = n3986 | n4555 ;
  buffer buf_n4557( .i (n4183), .o (n4557) );
  buffer buf_n4558( .i (n2273), .o (n4558) );
  assign n4559 = ( n3187 & ~n4557 ) | ( n3187 & n4558 ) | ( ~n4557 & n4558 ) ;
  buffer buf_n4560( .i (n4559), .o (n4560) );
  buffer buf_n4561( .i (n4560), .o (n4561) );
  assign n4566 = ( ~n2540 & n4295 ) | ( ~n2540 & n4561 ) | ( n4295 & n4561 ) ;
  buffer buf_n4567( .i (n4566), .o (n4567) );
  assign n4570 = n4216 & ~n4567 ;
  buffer buf_n4571( .i (n4570), .o (n4571) );
  buffer buf_n4572( .i (n4571), .o (n4572) );
  buffer buf_n4568( .i (n4567), .o (n4568) );
  buffer buf_n4569( .i (n4568), .o (n4569) );
  assign n4573 = n4569 | n4571 ;
  assign n4574 = ( ~n4417 & n4572 ) | ( ~n4417 & n4573 ) | ( n4572 & n4573 ) ;
  assign n4575 = n4406 & n4574 ;
  buffer buf_n4576( .i (n3056), .o (n4576) );
  buffer buf_n4577( .i (n4576), .o (n4577) );
  buffer buf_n4578( .i (n4577), .o (n4578) );
  buffer buf_n4579( .i (n4578), .o (n4579) );
  assign n4580 = ( ~n3899 & n3958 ) | ( ~n3899 & n4579 ) | ( n3958 & n4579 ) ;
  buffer buf_n4581( .i (n4580), .o (n4581) );
  buffer buf_n4582( .i (n4581), .o (n4582) );
  assign n4583 = n4538 & ~n4581 ;
  assign n4584 = ( n2035 & n4582 ) | ( n2035 & ~n4583 ) | ( n4582 & ~n4583 ) ;
  assign n4585 = ~n4406 & n4584 ;
  assign n4586 = ( n4407 & ~n4575 ) | ( n4407 & n4585 ) | ( ~n4575 & n4585 ) ;
  assign n4587 = n3366 & ~n4586 ;
  assign n4588 = n3898 | n4315 ;
  buffer buf_n4589( .i (n4588), .o (n4589) );
  buffer buf_n4590( .i (n4589), .o (n4590) );
  assign n4596 = n4341 & n4590 ;
  assign n4597 = ( n607 & n2608 ) | ( n607 & ~n4596 ) | ( n2608 & ~n4596 ) ;
  assign n4598 = ~n4098 & n4597 ;
  assign n4599 = ( n274 & n1753 ) | ( n274 & ~n2118 ) | ( n1753 & ~n2118 ) ;
  buffer buf_n4600( .i (n4599), .o (n4600) );
  assign n4613 = ( n4098 & n4418 ) | ( n4098 & n4600 ) | ( n4418 & n4600 ) ;
  assign n4614 = ( n688 & n4598 ) | ( n688 & ~n4613 ) | ( n4598 & ~n4613 ) ;
  assign n4615 = n3366 | n4614 ;
  assign n4616 = ( ~n4393 & n4587 ) | ( ~n4393 & n4615 ) | ( n4587 & n4615 ) ;
  buffer buf_n4617( .i (n4061), .o (n4617) );
  assign n4618 = n4616 & ~n4617 ;
  assign n4619 = n3986 & ~n4618 ;
  assign n4620 = n4556 & ~n4619 ;
  assign n4621 = ~n4470 & n4620 ;
  assign n4622 = ( n4469 & ~n4471 ) | ( n4469 & n4621 ) | ( ~n4471 & n4621 ) ;
  buffer buf_n3681( .i (n3680), .o (n3681) );
  buffer buf_n3682( .i (n3681), .o (n3682) );
  buffer buf_n3683( .i (n3682), .o (n3683) );
  buffer buf_n3684( .i (n3683), .o (n3684) );
  buffer buf_n3685( .i (n3684), .o (n3685) );
  buffer buf_n3686( .i (n3685), .o (n3686) );
  buffer buf_n3687( .i (n3686), .o (n3687) );
  assign n4623 = ~n1585 & n3687 ;
  assign n4624 = ( ~n3510 & n4421 ) | ( ~n3510 & n4623 ) | ( n4421 & n4623 ) ;
  assign n4625 = n510 & n4538 ;
  assign n4626 = n1942 & n4625 ;
  assign n4627 = ~n3510 & n4626 ;
  assign n4628 = ( ~n4422 & n4624 ) | ( ~n4422 & n4627 ) | ( n4624 & n4627 ) ;
  buffer buf_n4629( .i (n4628), .o (n4629) );
  assign n4630 = ( ~n753 & n1401 ) | ( ~n753 & n4629 ) | ( n1401 & n4629 ) ;
  assign n4631 = ( n372 & n513 ) | ( n372 & ~n1803 ) | ( n513 & ~n1803 ) ;
  buffer buf_n4632( .i (n4631), .o (n4632) );
  assign n4639 = n4629 | n4632 ;
  assign n4640 = ( n754 & n4630 ) | ( n754 & n4639 ) | ( n4630 & n4639 ) ;
  assign n4641 = n262 | n4640 ;
  assign n4642 = ( ~n3659 & n3912 ) | ( ~n3659 & n4578 ) | ( n3912 & n4578 ) ;
  buffer buf_n4643( .i (n4317), .o (n4643) );
  assign n4644 = ( n3913 & n4642 ) | ( n3913 & ~n4643 ) | ( n4642 & ~n4643 ) ;
  buffer buf_n4645( .i (n4644), .o (n4645) );
  assign n4648 = n3771 & ~n4645 ;
  buffer buf_n4649( .i (n4648), .o (n4649) );
  buffer buf_n4650( .i (n4649), .o (n4650) );
  buffer buf_n4646( .i (n4645), .o (n4646) );
  buffer buf_n4647( .i (n4646), .o (n4647) );
  assign n4651 = n4647 | n4649 ;
  assign n4652 = ( ~n3968 & n4650 ) | ( ~n3968 & n4651 ) | ( n4650 & n4651 ) ;
  assign n4653 = n4423 & n4652 ;
  buffer buf_n4654( .i (n3911), .o (n4654) );
  buffer buf_n4655( .i (n4654), .o (n4655) );
  buffer buf_n4656( .i (n3927), .o (n4656) );
  buffer buf_n4657( .i (n4656), .o (n4657) );
  buffer buf_n4658( .i (n4657), .o (n4658) );
  assign n4659 = ( n2542 & n4655 ) | ( n2542 & ~n4658 ) | ( n4655 & ~n4658 ) ;
  buffer buf_n4660( .i (n4659), .o (n4660) );
  buffer buf_n4661( .i (n4660), .o (n4661) );
  buffer buf_n4662( .i (n4661), .o (n4662) );
  buffer buf_n4663( .i (n4662), .o (n4663) );
  buffer buf_n4664( .i (n3767), .o (n4664) );
  buffer buf_n4665( .i (n4343), .o (n4665) );
  assign n4666 = ( n4660 & n4664 ) | ( n4660 & n4665 ) | ( n4664 & n4665 ) ;
  buffer buf_n4667( .i (n4666), .o (n4667) );
  buffer buf_n4668( .i (n4667), .o (n4668) );
  assign n4669 = n2546 & ~n4667 ;
  assign n4670 = ( n4663 & ~n4668 ) | ( n4663 & n4669 ) | ( ~n4668 & n4669 ) ;
  assign n4671 = n4423 | n4670 ;
  assign n4672 = ( ~n3974 & n4653 ) | ( ~n3974 & n4671 ) | ( n4653 & n4671 ) ;
  assign n4673 = ~n4617 & n4672 ;
  assign n4674 = n262 & ~n4673 ;
  assign n4675 = n4641 & ~n4674 ;
  assign n4676 = n3400 | n4675 ;
  assign n4677 = ( n3096 & n3625 ) | ( n3096 & n4122 ) | ( n3625 & n4122 ) ;
  assign n4678 = ~n3968 & n4677 ;
  buffer buf_n4679( .i (n4678), .o (n4679) );
  buffer buf_n4680( .i (n4679), .o (n4680) );
  buffer buf_n4681( .i (n4680), .o (n4681) );
  assign n4682 = ( n4027 & n4303 ) | ( n4027 & n4657 ) | ( n4303 & n4657 ) ;
  buffer buf_n4683( .i (n4682), .o (n4683) );
  buffer buf_n4684( .i (n4683), .o (n4684) );
  buffer buf_n4685( .i (n4684), .o (n4685) );
  buffer buf_n4686( .i (n4685), .o (n4686) );
  buffer buf_n4687( .i (n4686), .o (n4687) );
  buffer buf_n4688( .i (n4687), .o (n4688) );
  assign n4689 = ( n3097 & n4389 ) | ( n3097 & n4407 ) | ( n4389 & n4407 ) ;
  assign n4690 = n4688 & ~n4689 ;
  assign n4691 = ( n4025 & n4679 ) | ( n4025 & n4690 ) | ( n4679 & n4690 ) ;
  assign n4692 = n4394 & ~n4691 ;
  assign n4693 = ( n4106 & n4681 ) | ( n4106 & ~n4692 ) | ( n4681 & ~n4692 ) ;
  assign n4694 = ~n3892 & n4693 ;
  assign n4695 = n3400 & ~n4694 ;
  assign n4696 = n4676 & ~n4695 ;
  assign n4697 = n4622 | n4696 ;
  assign n4698 = ( n4457 & ~n4458 ) | ( n4457 & n4697 ) | ( ~n4458 & n4697 ) ;
  buffer buf_n4699( .i (n4698), .o (n4699) );
  buffer buf_n4700( .i (n4699), .o (n4700) );
  assign n4701 = ( n45 & n2273 ) | ( n45 & n4222 ) | ( n2273 & n4222 ) ;
  buffer buf_n4702( .i (n4701), .o (n4702) );
  buffer buf_n4703( .i (n4702), .o (n4703) );
  buffer buf_n4704( .i (n4703), .o (n4704) );
  buffer buf_n4705( .i (n4704), .o (n4705) );
  buffer buf_n4706( .i (n4705), .o (n4706) );
  buffer buf_n4707( .i (n4706), .o (n4707) );
  buffer buf_n4708( .i (n4707), .o (n4708) );
  buffer buf_n4709( .i (n4708), .o (n4709) );
  buffer buf_n4710( .i (n4709), .o (n4710) );
  buffer buf_n4711( .i (n4710), .o (n4711) );
  buffer buf_n4712( .i (n4711), .o (n4712) );
  buffer buf_n4713( .i (n4712), .o (n4713) );
  buffer buf_n4714( .i (n4713), .o (n4714) );
  buffer buf_n4715( .i (n4714), .o (n4715) );
  assign n4716 = ( n3985 & n4360 ) | ( n3985 & n4450 ) | ( n4360 & n4450 ) ;
  assign n4717 = ( n568 & ~n4715 ) | ( n568 & n4716 ) | ( ~n4715 & n4716 ) ;
  buffer buf_n4718( .i (n4717), .o (n4718) );
  buffer buf_n4719( .i (n4718), .o (n4719) );
  assign n4720 = ( n264 & n4470 ) | ( n264 & ~n4718 ) | ( n4470 & ~n4718 ) ;
  assign n4721 = n4380 & n4536 ;
  buffer buf_n4722( .i (n4721), .o (n4722) );
  buffer buf_n4723( .i (n4722), .o (n4723) );
  buffer buf_n4724( .i (n4723), .o (n4724) );
  buffer buf_n4725( .i (n4724), .o (n4725) );
  buffer buf_n4726( .i (n4725), .o (n4726) );
  buffer buf_n4727( .i (n4726), .o (n4727) );
  buffer buf_n4728( .i (n4727), .o (n4728) );
  buffer buf_n4729( .i (n4440), .o (n4729) );
  buffer buf_n4730( .i (n4729), .o (n4730) );
  buffer buf_n4731( .i (n4730), .o (n4731) );
  assign n4732 = ( n4451 & n4728 ) | ( n4451 & n4731 ) | ( n4728 & n4731 ) ;
  assign n4733 = ~n263 & n4732 ;
  assign n4734 = n4470 & n4733 ;
  assign n4735 = ( n4719 & n4720 ) | ( n4719 & n4734 ) | ( n4720 & n4734 ) ;
  buffer buf_n4736( .i (n4735), .o (n4736) );
  buffer buf_n4737( .i (n4736), .o (n4737) );
  buffer buf_n4738( .i (n3187), .o (n4738) );
  buffer buf_n4739( .i (n4738), .o (n4739) );
  buffer buf_n4740( .i (n4739), .o (n4740) );
  buffer buf_n4741( .i (n4740), .o (n4741) );
  buffer buf_n4742( .i (n4741), .o (n4742) );
  assign n4743 = ( n4304 & n4658 ) | ( n4304 & ~n4742 ) | ( n4658 & ~n4742 ) ;
  buffer buf_n4744( .i (n4743), .o (n4744) );
  buffer buf_n4745( .i (n4744), .o (n4745) );
  buffer buf_n4746( .i (n4745), .o (n4746) );
  buffer buf_n4747( .i (n4746), .o (n4747) );
  buffer buf_n4748( .i (n4747), .o (n4748) );
  buffer buf_n4753( .i (n3884), .o (n4753) );
  assign n4754 = ( n4462 & n4748 ) | ( n4462 & n4753 ) | ( n4748 & n4753 ) ;
  buffer buf_n4755( .i (n4754), .o (n4755) );
  buffer buf_n4756( .i (n4755), .o (n4756) );
  buffer buf_n4757( .i (n4756), .o (n4757) );
  buffer buf_n4758( .i (n4757), .o (n4758) );
  assign n4759 = ( n4450 & n4730 ) | ( n4450 & n4755 ) | ( n4730 & n4755 ) ;
  buffer buf_n4760( .i (n4759), .o (n4760) );
  buffer buf_n4761( .i (n4760), .o (n4761) );
  buffer buf_n4749( .i (n4748), .o (n4749) );
  buffer buf_n4750( .i (n4749), .o (n4750) );
  buffer buf_n4751( .i (n4750), .o (n4751) );
  buffer buf_n4752( .i (n4751), .o (n4752) );
  assign n4762 = n4752 & ~n4760 ;
  assign n4763 = ( n4758 & ~n4761 ) | ( n4758 & n4762 ) | ( ~n4761 & n4762 ) ;
  assign n4764 = ( ~n2640 & n3836 ) | ( ~n2640 & n4763 ) | ( n3836 & n4763 ) ;
  buffer buf_n4765( .i (n4478), .o (n4765) );
  buffer buf_n4766( .i (n4765), .o (n4766) );
  buffer buf_n4767( .i (n4766), .o (n4767) );
  assign n4768 = ( n4657 & n4741 ) | ( n4657 & n4767 ) | ( n4741 & n4767 ) ;
  buffer buf_n4769( .i (n4768), .o (n4769) );
  buffer buf_n4770( .i (n4769), .o (n4770) );
  buffer buf_n4771( .i (n4770), .o (n4771) );
  buffer buf_n4772( .i (n4771), .o (n4772) );
  buffer buf_n4773( .i (n4772), .o (n4773) );
  buffer buf_n4774( .i (n4773), .o (n4774) );
  buffer buf_n4775( .i (n3619), .o (n4775) );
  assign n4776 = ( ~n4753 & n4774 ) | ( ~n4753 & n4775 ) | ( n4774 & n4775 ) ;
  buffer buf_n4777( .i (n4776), .o (n4777) );
  assign n4780 = n4450 & ~n4777 ;
  buffer buf_n4781( .i (n4780), .o (n4781) );
  buffer buf_n4782( .i (n4781), .o (n4782) );
  buffer buf_n4778( .i (n4777), .o (n4778) );
  buffer buf_n4779( .i (n4778), .o (n4779) );
  assign n4783 = n4779 | n4781 ;
  assign n4784 = ( ~n148 & n4782 ) | ( ~n148 & n4783 ) | ( n4782 & n4783 ) ;
  buffer buf_n4785( .i (n3986), .o (n4785) );
  buffer buf_n4786( .i (n4785), .o (n4786) );
  buffer buf_n4787( .i (n4786), .o (n4787) );
  assign n4788 = ( n2640 & ~n4784 ) | ( n2640 & n4787 ) | ( ~n4784 & n4787 ) ;
  assign n4789 = n4764 & ~n4788 ;
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n4790( .i (n3723), .o (n4790) );
  assign n4791 = ( n747 & ~n4360 ) | ( n747 & n4790 ) | ( ~n4360 & n4790 ) ;
  buffer buf_n4792( .i (n4422), .o (n4792) );
  buffer buf_n4793( .i (n4792), .o (n4793) );
  assign n4794 = ( ~n746 & n3723 ) | ( ~n746 & n4793 ) | ( n3723 & n4793 ) ;
  assign n4795 = ( n4104 & ~n4360 ) | ( n4104 & n4794 ) | ( ~n4360 & n4794 ) ;
  assign n4796 = ~n4791 & n4795 ;
  buffer buf_n4797( .i (n4796), .o (n4797) );
  buffer buf_n4798( .i (n4797), .o (n4798) );
  assign n4799 = ( n3015 & n3840 ) | ( n3015 & n4797 ) | ( n3840 & n4797 ) ;
  buffer buf_n4800( .i (n4417), .o (n4800) );
  assign n4801 = n3883 & ~n4800 ;
  buffer buf_n4802( .i (n4801), .o (n4802) );
  buffer buf_n4803( .i (n4802), .o (n4803) );
  buffer buf_n4804( .i (n4803), .o (n4804) );
  buffer buf_n4805( .i (n4804), .o (n4805) );
  buffer buf_n4806( .i (n4104), .o (n4806) );
  assign n4807 = ( n708 & n4805 ) | ( n708 & n4806 ) | ( n4805 & n4806 ) ;
  assign n4808 = ~n4453 & n4807 ;
  assign n4809 = ~n3015 & n4808 ;
  assign n4810 = ( n4798 & ~n4799 ) | ( n4798 & n4809 ) | ( ~n4799 & n4809 ) ;
  buffer buf_n4811( .i (n4810), .o (n4811) );
  assign n4812 = ( ~n4736 & n4789 ) | ( ~n4736 & n4811 ) | ( n4789 & n4811 ) ;
  assign n4813 = n3020 & ~n4811 ;
  assign n4814 = ( n4737 & n4812 ) | ( n4737 & ~n4813 ) | ( n4812 & ~n4813 ) ;
  assign n4815 = n4699 | n4814 ;
  assign n4816 = ( ~n4266 & n4700 ) | ( ~n4266 & n4815 ) | ( n4700 & n4815 ) ;
  buffer buf_n1405( .i (n1404), .o (n1405) );
  assign n4817 = ( n688 & ~n798 ) | ( n688 & n2775 ) | ( ~n798 & n2775 ) ;
  assign n4818 = ( n689 & ~n4462 ) | ( n689 & n4817 ) | ( ~n4462 & n4817 ) ;
  assign n4819 = n4793 & ~n4818 ;
  assign n4820 = ~n4617 & n4819 ;
  buffer buf_n4821( .i (n4820), .o (n4821) );
  buffer buf_n4822( .i (n4821), .o (n4822) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  assign n4823 = n1568 & ~n4821 ;
  assign n4824 = ( n1405 & n4822 ) | ( n1405 & ~n4823 ) | ( n4822 & ~n4823 ) ;
  buffer buf_n4825( .i (n4824), .o (n4825) );
  buffer buf_n4826( .i (n4825), .o (n4826) );
  assign n4827 = n1404 & n2243 ;
  assign n4828 = n403 & n4827 ;
  assign n4829 = n540 | n4393 ;
  assign n4830 = ( ~n2723 & n3100 ) | ( ~n2723 & n4829 ) | ( n3100 & n4829 ) ;
  assign n4831 = ( n369 & n1429 ) | ( n369 & ~n2882 ) | ( n1429 & ~n2882 ) ;
  buffer buf_n4832( .i (n4380), .o (n4832) );
  buffer buf_n4833( .i (n4832), .o (n4833) );
  buffer buf_n4834( .i (n3914), .o (n4834) );
  buffer buf_n4835( .i (n4834), .o (n4835) );
  assign n4836 = ( n4831 & n4833 ) | ( n4831 & ~n4835 ) | ( n4833 & ~n4835 ) ;
  buffer buf_n4837( .i (n4836), .o (n4837) );
  buffer buf_n4838( .i (n4837), .o (n4838) );
  assign n4839 = ~n4422 & n4837 ;
  buffer buf_n4840( .i (n3968), .o (n4840) );
  assign n4841 = ( n4838 & n4839 ) | ( n4838 & n4840 ) | ( n4839 & n4840 ) ;
  buffer buf_n4842( .i (n4841), .o (n4842) );
  buffer buf_n4843( .i (n4842), .o (n4843) );
  buffer buf_n4844( .i (n4390), .o (n4844) );
  buffer buf_n4845( .i (n4844), .o (n4845) );
  assign n4846 = n4842 | n4845 ;
  assign n4847 = ( n4830 & n4843 ) | ( n4830 & n4846 ) | ( n4843 & n4846 ) ;
  assign n4848 = ( n2689 & ~n3892 ) | ( n2689 & n4847 ) | ( ~n3892 & n4847 ) ;
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n4849( .i (n4538), .o (n4849) );
  buffer buf_n4850( .i (n4849), .o (n4850) );
  assign n4851 = ( ~n310 & n4421 ) | ( ~n310 & n4850 ) | ( n4421 & n4850 ) ;
  buffer buf_n4852( .i (n4425), .o (n4852) );
  assign n4853 = ( ~n310 & n4850 ) | ( ~n310 & n4852 ) | ( n4850 & n4852 ) ;
  assign n4854 = ( n2154 & n4851 ) | ( n2154 & ~n4853 ) | ( n4851 & ~n4853 ) ;
  assign n4855 = ~n4390 & n4854 ;
  buffer buf_n4856( .i (n4855), .o (n4856) );
  buffer buf_n4857( .i (n4856), .o (n4857) );
  buffer buf_n4858( .i (n4421), .o (n4858) );
  buffer buf_n4859( .i (n4122), .o (n4859) );
  assign n4860 = ( n4389 & n4858 ) | ( n4389 & ~n4859 ) | ( n4858 & ~n4859 ) ;
  buffer buf_n4861( .i (n4860), .o (n4861) );
  assign n4865 = n3408 & n4861 ;
  assign n4866 = n4856 | n4865 ;
  assign n4867 = ( ~n4451 & n4857 ) | ( ~n4451 & n4866 ) | ( n4857 & n4866 ) ;
  buffer buf_n4868( .i (n2688), .o (n4868) );
  assign n4869 = ( n3892 & ~n4867 ) | ( n3892 & n4868 ) | ( ~n4867 & n4868 ) ;
  assign n4870 = n4848 & ~n4869 ;
  assign n4871 = ( ~n355 & n4828 ) | ( ~n355 & n4870 ) | ( n4828 & n4870 ) ;
  assign n4872 = ~n4825 & n4871 ;
  assign n4873 = ( ~n357 & n4826 ) | ( ~n357 & n4872 ) | ( n4826 & n4872 ) ;
  buffer buf_n4874( .i (n4873), .o (n4874) );
  buffer buf_n4875( .i (n4874), .o (n4875) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n2499( .i (n2498), .o (n2499) );
  buffer buf_n2500( .i (n2499), .o (n2500) );
  assign n4876 = ( n2500 & n3723 ) | ( n2500 & n4061 ) | ( n3723 & n4061 ) ;
  buffer buf_n4877( .i (n3510), .o (n4877) );
  buffer buf_n4878( .i (n4877), .o (n4878) );
  assign n4879 = ( ~n2499 & n4462 ) | ( ~n2499 & n4878 ) | ( n4462 & n4878 ) ;
  assign n4880 = ( n3975 & ~n4729 ) | ( n3975 & n4879 ) | ( ~n4729 & n4879 ) ;
  assign n4881 = ~n4876 & n4880 ;
  assign n4882 = n922 & ~n4800 ;
  assign n4883 = ( ~n3619 & n4877 ) | ( ~n3619 & n4882 ) | ( n4877 & n4882 ) ;
  assign n4884 = ~n4878 & n4883 ;
  buffer buf_n4885( .i (n4884), .o (n4885) );
  buffer buf_n4886( .i (n4885), .o (n4886) );
  buffer buf_n4887( .i (n232), .o (n4887) );
  assign n4888 = n4885 | n4887 ;
  assign n4889 = ( n4881 & n4886 ) | ( n4881 & n4888 ) | ( n4886 & n4888 ) ;
  assign n4890 = n4785 | n4889 ;
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  assign n4891 = n3898 & n4741 ;
  buffer buf_n4892( .i (n4891), .o (n4892) );
  buffer buf_n4893( .i (n4892), .o (n4893) );
  buffer buf_n4894( .i (n4893), .o (n4894) );
  buffer buf_n4895( .i (n4894), .o (n4895) );
  buffer buf_n4896( .i (n4895), .o (n4896) );
  buffer buf_n4897( .i (n4896), .o (n4897) );
  buffer buf_n4898( .i (n4897), .o (n4898) );
  buffer buf_n4899( .i (n4898), .o (n4899) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n4902( .i (n4800), .o (n4902) );
  buffer buf_n4903( .i (n4902), .o (n4903) );
  buffer buf_n4904( .i (n4903), .o (n4904) );
  assign n4905 = ~n671 & n4904 ;
  assign n4906 = ( n660 & n4899 ) | ( n660 & ~n4905 ) | ( n4899 & ~n4905 ) ;
  assign n4907 = ~n4466 & n4906 ;
  assign n4908 = n4785 & ~n4907 ;
  assign n4909 = n4890 & ~n4908 ;
  buffer buf_n4910( .i (n4453), .o (n4910) );
  buffer buf_n4911( .i (n4910), .o (n4911) );
  assign n4912 = n4909 | n4911 ;
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n4913( .i (n4850), .o (n4913) );
  assign n4914 = ( n609 & n4858 ) | ( n609 & ~n4913 ) | ( n4858 & ~n4913 ) ;
  assign n4915 = ( n608 & ~n3883 ) | ( n608 & n4850 ) | ( ~n3883 & n4850 ) ;
  buffer buf_n4916( .i (n4406), .o (n4916) );
  assign n4917 = ( n4858 & ~n4915 ) | ( n4858 & n4916 ) | ( ~n4915 & n4916 ) ;
  assign n4918 = ~n4914 & n4917 ;
  buffer buf_n4919( .i (n4918), .o (n4919) );
  buffer buf_n4920( .i (n4919), .o (n4920) );
  buffer buf_n4921( .i (n4920), .o (n4921) );
  buffer buf_n4922( .i (n3975), .o (n4922) );
  assign n4923 = ( n926 & n4919 ) | ( n926 & ~n4922 ) | ( n4919 & ~n4922 ) ;
  assign n4924 = n836 & ~n4923 ;
  assign n4925 = ( n837 & n4921 ) | ( n837 & ~n4924 ) | ( n4921 & ~n4924 ) ;
  buffer buf_n4926( .i (n4466), .o (n4926) );
  buffer buf_n4927( .i (n4926), .o (n4927) );
  assign n4928 = n4925 & ~n4927 ;
  assign n4929 = n4911 & ~n4928 ;
  assign n4930 = n4912 & ~n4929 ;
  assign n4931 = n181 | n4930 ;
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  assign n4932 = ( n281 & n1369 ) | ( n281 & ~n4805 ) | ( n1369 & ~n4805 ) ;
  assign n4933 = ~n745 & n4840 ;
  buffer buf_n4934( .i (n4933), .o (n4934) );
  buffer buf_n4935( .i (n4934), .o (n4935) );
  buffer buf_n4936( .i (n4935), .o (n4936) );
  assign n4937 = n4932 & n4936 ;
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  assign n4938 = n278 & ~n4903 ;
  buffer buf_n4939( .i (n4938), .o (n4939) );
  buffer buf_n4940( .i (n4939), .o (n4940) );
  buffer buf_n4941( .i (n4940), .o (n4941) );
  assign n4942 = ( ~n749 & n4936 ) | ( ~n749 & n4941 ) | ( n4936 & n4941 ) ;
  assign n4943 = ( n4786 & n4937 ) | ( n4786 & n4942 ) | ( n4937 & n4942 ) ;
  assign n4944 = n4934 & n4939 ;
  assign n4945 = n924 & n4903 ;
  buffer buf_n4946( .i (n4945), .o (n4946) );
  assign n4953 = ( ~n747 & n4934 ) | ( ~n747 & n4946 ) | ( n4934 & n4946 ) ;
  buffer buf_n4954( .i (n3985), .o (n4954) );
  assign n4955 = ( n4944 & n4953 ) | ( n4944 & n4954 ) | ( n4953 & n4954 ) ;
  buffer buf_n4956( .i (n4955), .o (n4956) );
  buffer buf_n4957( .i (n4956), .o (n4957) );
  assign n4958 = n148 & ~n4956 ;
  assign n4959 = ( n4943 & n4957 ) | ( n4943 & ~n4958 ) | ( n4957 & ~n4958 ) ;
  buffer buf_n4960( .i (n3416), .o (n4960) );
  assign n4961 = n4959 & ~n4960 ;
  assign n4962 = n181 & ~n4961 ;
  assign n4963 = n4931 & ~n4962 ;
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  assign n4964 = ~n340 & n1809 ;
  assign n4965 = ( n2583 & n3927 ) | ( n2583 & ~n3930 ) | ( n3927 & ~n3930 ) ;
  buffer buf_n4966( .i (n4965), .o (n4966) );
  assign n4969 = n4657 & ~n4966 ;
  buffer buf_n4970( .i (n4969), .o (n4970) );
  buffer buf_n4971( .i (n4970), .o (n4971) );
  buffer buf_n4967( .i (n4966), .o (n4967) );
  buffer buf_n4968( .i (n4967), .o (n4968) );
  assign n4972 = n4968 | n4970 ;
  buffer buf_n4973( .i (n4658), .o (n4973) );
  buffer buf_n4974( .i (n4973), .o (n4974) );
  assign n4975 = ( n4971 & n4972 ) | ( n4971 & ~n4974 ) | ( n4972 & ~n4974 ) ;
  assign n4976 = ~n4833 & n4975 ;
  assign n4977 = n4474 & ~n4833 ;
  buffer buf_n4978( .i (n4656), .o (n4978) );
  assign n4979 = ( ~n4654 & n4767 ) | ( ~n4654 & n4978 ) | ( n4767 & n4978 ) ;
  buffer buf_n4980( .i (n4979), .o (n4980) );
  buffer buf_n4981( .i (n4980), .o (n4981) );
  assign n4982 = n3914 & n4980 ;
  assign n4983 = ( ~n1045 & n4981 ) | ( ~n1045 & n4982 ) | ( n4981 & n4982 ) ;
  buffer buf_n4984( .i (n3768), .o (n4984) );
  buffer buf_n4985( .i (n4984), .o (n4985) );
  assign n4986 = ( ~n4833 & n4983 ) | ( ~n4833 & n4985 ) | ( n4983 & n4985 ) ;
  assign n4987 = ( n4976 & ~n4977 ) | ( n4976 & n4986 ) | ( ~n4977 & n4986 ) ;
  assign n4988 = n4902 & n4987 ;
  assign n4989 = ( n46 & ~n4557 ) | ( n46 & n4558 ) | ( ~n4557 & n4558 ) ;
  buffer buf_n4990( .i (n4989), .o (n4990) );
  assign n4995 = ( n3927 & ~n4765 ) | ( n3927 & n4990 ) | ( ~n4765 & n4990 ) ;
  buffer buf_n4996( .i (n4995), .o (n4996) );
  buffer buf_n4997( .i (n4996), .o (n4997) );
  buffer buf_n4998( .i (n4997), .o (n4998) );
  buffer buf_n4999( .i (n4998), .o (n4999) );
  buffer buf_n5000( .i (n3897), .o (n5000) );
  assign n5001 = ( n4027 & n4996 ) | ( n4027 & n5000 ) | ( n4996 & n5000 ) ;
  buffer buf_n5002( .i (n5001), .o (n5002) );
  buffer buf_n5003( .i (n5002), .o (n5003) );
  buffer buf_n4991( .i (n4990), .o (n4991) );
  buffer buf_n4992( .i (n4991), .o (n4992) );
  buffer buf_n4993( .i (n4992), .o (n4993) );
  buffer buf_n4994( .i (n4993), .o (n4994) );
  assign n5004 = n4994 & ~n5002 ;
  assign n5005 = ( n4999 & ~n5003 ) | ( n4999 & n5004 ) | ( ~n5003 & n5004 ) ;
  assign n5006 = n4835 & ~n5005 ;
  assign n5007 = n920 & n4832 ;
  assign n5008 = n4835 | n5007 ;
  assign n5009 = ~n5006 & n5008 ;
  assign n5010 = n4902 | n5009 ;
  assign n5011 = ( ~n4903 & n4988 ) | ( ~n4903 & n5010 ) | ( n4988 & n5010 ) ;
  assign n5012 = n4844 & n5011 ;
  buffer buf_n4562( .i (n4561), .o (n4562) );
  buffer buf_n4563( .i (n4562), .o (n4563) );
  buffer buf_n4564( .i (n4563), .o (n4564) );
  buffer buf_n4565( .i (n4564), .o (n4565) );
  assign n5013 = n4565 & n4834 ;
  assign n5014 = n4536 | n4564 ;
  assign n5015 = ( n4834 & ~n4974 ) | ( n4834 & n5014 ) | ( ~n4974 & n5014 ) ;
  assign n5016 = ~n5013 & n5015 ;
  buffer buf_n5017( .i (n4832), .o (n5017) );
  buffer buf_n5018( .i (n5017), .o (n5018) );
  buffer buf_n5019( .i (n4405), .o (n5019) );
  assign n5020 = ( n5016 & n5018 ) | ( n5016 & ~n5019 ) | ( n5018 & ~n5019 ) ;
  assign n5021 = n424 & ~n4984 ;
  buffer buf_n5022( .i (n4742), .o (n5022) );
  assign n5023 = ( ~n423 & n4973 ) | ( ~n423 & n5022 ) | ( n4973 & n5022 ) ;
  assign n5024 = ( n1054 & n4984 ) | ( n1054 & ~n5023 ) | ( n4984 & ~n5023 ) ;
  assign n5025 = ( n4985 & n5021 ) | ( n4985 & ~n5024 ) | ( n5021 & ~n5024 ) ;
  assign n5026 = ( n5018 & n5019 ) | ( n5018 & ~n5025 ) | ( n5019 & ~n5025 ) ;
  assign n5027 = n5020 & ~n5026 ;
  buffer buf_n2857( .i (n2856), .o (n2857) );
  buffer buf_n2858( .i (n2857), .o (n2858) );
  buffer buf_n2859( .i (n2858), .o (n2859) );
  buffer buf_n2860( .i (n2859), .o (n2860) );
  buffer buf_n2861( .i (n2860), .o (n2861) );
  buffer buf_n2862( .i (n2861), .o (n2862) );
  assign n5028 = ( ~n922 & n2862 ) | ( ~n922 & n5018 ) | ( n2862 & n5018 ) ;
  assign n5029 = n923 & n5028 ;
  assign n5030 = n5027 | n5029 ;
  assign n5031 = ~n4844 & n5030 ;
  assign n5032 = n5012 | n5031 ;
  assign n5033 = ~n4466 & n5032 ;
  buffer buf_n5034( .i (n5033), .o (n5034) );
  buffer buf_n5035( .i (n5034), .o (n5035) );
  assign n5036 = n716 | n5034 ;
  assign n5037 = ( n4964 & n5035 ) | ( n4964 & n5036 ) | ( n5035 & n5036 ) ;
  assign n5038 = n180 & ~n5037 ;
  assign n5039 = ( n4654 & n4767 ) | ( n4654 & ~n5000 ) | ( n4767 & ~n5000 ) ;
  buffer buf_n5040( .i (n5039), .o (n5040) );
  buffer buf_n5041( .i (n5040), .o (n5041) );
  buffer buf_n5042( .i (n5041), .o (n5042) );
  buffer buf_n5043( .i (n5042), .o (n5043) );
  buffer buf_n5044( .i (n5043), .o (n5044) );
  assign n5045 = ( ~n4859 & n4913 ) | ( ~n4859 & n5044 ) | ( n4913 & n5044 ) ;
  assign n5046 = ( n4913 & n4916 ) | ( n4913 & ~n5044 ) | ( n4916 & ~n5044 ) ;
  assign n5047 = n5045 & ~n5046 ;
  buffer buf_n5048( .i (n5047), .o (n5048) );
  buffer buf_n5049( .i (n5048), .o (n5049) );
  assign n5050 = ( n3985 & n4845 ) | ( n3985 & ~n5048 ) | ( n4845 & ~n5048 ) ;
  assign n5051 = n539 & n4775 ;
  assign n5052 = n611 & n5051 ;
  assign n5053 = n4845 & n5052 ;
  assign n5054 = ( n5049 & n5050 ) | ( n5049 & n5053 ) | ( n5050 & n5053 ) ;
  buffer buf_n5055( .i (n4775), .o (n5055) );
  assign n5056 = ( n4793 & n4844 ) | ( n4793 & n5055 ) | ( n4844 & n5055 ) ;
  buffer buf_n5057( .i (n4767), .o (n5057) );
  assign n5058 = ( n3899 & n4655 ) | ( n3899 & n5057 ) | ( n4655 & n5057 ) ;
  assign n5059 = ( n4494 & ~n5022 ) | ( n4494 & n5058 ) | ( ~n5022 & n5058 ) ;
  buffer buf_n5060( .i (n5059), .o (n5060) );
  assign n5063 = n4405 & ~n5060 ;
  buffer buf_n5064( .i (n5063), .o (n5064) );
  buffer buf_n5065( .i (n5064), .o (n5065) );
  buffer buf_n5061( .i (n5060), .o (n5061) );
  buffer buf_n5062( .i (n5061), .o (n5062) );
  assign n5066 = n5062 | n5064 ;
  assign n5067 = ( ~n4440 & n5065 ) | ( ~n4440 & n5066 ) | ( n5065 & n5066 ) ;
  assign n5068 = n4858 | n4913 ;
  buffer buf_n5069( .i (n5068), .o (n5069) );
  buffer buf_n5071( .i (n4390), .o (n5071) );
  assign n5072 = ( n5067 & n5069 ) | ( n5067 & n5071 ) | ( n5069 & n5071 ) ;
  assign n5073 = ~n5056 & n5072 ;
  buffer buf_n5074( .i (n5073), .o (n5074) );
  assign n5075 = ( ~n4868 & n5054 ) | ( ~n4868 & n5074 ) | ( n5054 & n5074 ) ;
  buffer buf_n5076( .i (n4655), .o (n5076) );
  assign n5077 = n3768 & ~n5076 ;
  buffer buf_n5078( .i (n5077), .o (n5078) );
  buffer buf_n5079( .i (n5078), .o (n5079) );
  buffer buf_n5086( .i (n4415), .o (n5086) );
  assign n5087 = ( n4122 & n5079 ) | ( n4122 & n5086 ) | ( n5079 & n5086 ) ;
  assign n5088 = ( n5018 & n5079 ) | ( n5018 & n5086 ) | ( n5079 & n5086 ) ;
  assign n5089 = ( n1944 & n5087 ) | ( n1944 & ~n5088 ) | ( n5087 & ~n5088 ) ;
  buffer buf_n5090( .i (n4916), .o (n5090) );
  assign n5091 = ~n5089 & n5090 ;
  assign n5092 = n4665 & ~n4832 ;
  buffer buf_n5093( .i (n5092), .o (n5093) );
  buffer buf_n2250( .i (n2249), .o (n2250) );
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  assign n5097 = n2255 & n5017 ;
  buffer buf_n5098( .i (n5017), .o (n5098) );
  assign n5099 = ( n5093 & ~n5097 ) | ( n5093 & n5098 ) | ( ~n5097 & n5098 ) ;
  assign n5100 = n4859 & ~n5099 ;
  assign n5101 = n5090 | n5100 ;
  assign n5102 = ~n5091 & n5101 ;
  assign n5103 = n4922 & ~n5102 ;
  assign n5104 = ( n663 & ~n4337 ) | ( n663 & n4665 ) | ( ~n4337 & n4665 ) ;
  buffer buf_n5105( .i (n5104), .o (n5105) );
  buffer buf_n5106( .i (n5105), .o (n5106) );
  buffer buf_n5107( .i (n5106), .o (n5107) );
  assign n5108 = ( n5019 & ~n5098 ) | ( n5019 & n5105 ) | ( ~n5098 & n5105 ) ;
  buffer buf_n5109( .i (n5086), .o (n5109) );
  assign n5110 = ( n3884 & ~n5108 ) | ( n3884 & n5109 ) | ( ~n5108 & n5109 ) ;
  assign n5111 = ~n5107 & n5110 ;
  buffer buf_n5112( .i (n4840), .o (n5112) );
  assign n5113 = n5111 & n5112 ;
  assign n5114 = n4922 | n5113 ;
  assign n5115 = ~n5103 & n5114 ;
  assign n5116 = ( n4868 & n5074 ) | ( n4868 & n5115 ) | ( n5074 & n5115 ) ;
  assign n5117 = n5075 | n5116 ;
  assign n5118 = ~n3416 & n5117 ;
  assign n5119 = n180 | n5118 ;
  assign n5120 = ~n5038 & n5119 ;
  assign n5121 = n431 & n802 ;
  assign n5122 = ( n2126 & n4785 ) | ( n2126 & n5121 ) | ( n4785 & n5121 ) ;
  assign n5123 = ~n4786 & n5122 ;
  buffer buf_n5124( .i (n5123), .o (n5124) );
  buffer buf_n5125( .i (n5124), .o (n5125) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n5126( .i (n4845), .o (n5126) );
  assign n5127 = ( n661 & n4806 ) | ( n661 & n5126 ) | ( n4806 & n5126 ) ;
  buffer buf_n5128( .i (n4806), .o (n5128) );
  assign n5129 = n5127 & ~n5128 ;
  assign n5130 = ( ~n3400 & n4786 ) | ( ~n3400 & n5129 ) | ( n4786 & n5129 ) ;
  assign n5131 = ( ~n3767 & n4380 ) | ( ~n3767 & n4973 ) | ( n4380 & n4973 ) ;
  buffer buf_n5132( .i (n4214), .o (n5132) );
  buffer buf_n5133( .i (n5132), .o (n5133) );
  assign n5134 = ( ~n4984 & n5131 ) | ( ~n4984 & n5133 ) | ( n5131 & n5133 ) ;
  buffer buf_n5135( .i (n5134), .o (n5135) );
  assign n5138 = n5098 & ~n5135 ;
  buffer buf_n5139( .i (n5138), .o (n5139) );
  buffer buf_n5140( .i (n5139), .o (n5140) );
  buffer buf_n5136( .i (n5135), .o (n5136) );
  buffer buf_n5137( .i (n5136), .o (n5137) );
  assign n5141 = n5137 | n5139 ;
  assign n5142 = ( ~n4793 & n5140 ) | ( ~n4793 & n5141 ) | ( n5140 & n5141 ) ;
  buffer buf_n5143( .i (n5142), .o (n5143) );
  buffer buf_n5144( .i (n5143), .o (n5144) );
  assign n5145 = ( ~n4806 & n5126 ) | ( ~n4806 & n5143 ) | ( n5126 & n5143 ) ;
  buffer buf_n5146( .i (n3144), .o (n5146) );
  assign n5147 = ( n3930 & n4246 ) | ( n3930 & ~n5146 ) | ( n4246 & ~n5146 ) ;
  buffer buf_n5148( .i (n5147), .o (n5148) );
  buffer buf_n5149( .i (n5148), .o (n5149) );
  buffer buf_n5150( .i (n4316), .o (n5150) );
  assign n5151 = n5148 & ~n5150 ;
  assign n5152 = ( n4658 & n5149 ) | ( n4658 & n5151 ) | ( n5149 & n5151 ) ;
  buffer buf_n5153( .i (n5152), .o (n5153) );
  buffer buf_n5154( .i (n5153), .o (n5154) );
  buffer buf_n5155( .i (n5154), .o (n5155) );
  buffer buf_n5156( .i (n5155), .o (n5156) );
  buffer buf_n5157( .i (n5156), .o (n5157) );
  buffer buf_n5158( .i (n5157), .o (n5158) );
  buffer buf_n5160( .i (n4792), .o (n5160) );
  assign n5161 = n5158 & ~n5160 ;
  assign n5162 = ~n4104 & n5161 ;
  assign n5163 = ~n5126 & n5162 ;
  assign n5164 = ( n5144 & ~n5145 ) | ( n5144 & n5163 ) | ( ~n5145 & n5163 ) ;
  buffer buf_n5165( .i (n4868), .o (n5165) );
  assign n5166 = n5164 & ~n5165 ;
  assign n5167 = ( ~n4787 & n5130 ) | ( ~n4787 & n5166 ) | ( n5130 & n5166 ) ;
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n2036( .i (n2035), .o (n2036) );
  buffer buf_n2037( .i (n2036), .o (n2037) );
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n5168( .i (n714), .o (n5168) );
  assign n5169 = n2042 & n5168 ;
  assign n5170 = n378 & n5169 ;
  buffer buf_n5171( .i (n5170), .o (n5171) );
  assign n5172 = ( ~n5124 & n5167 ) | ( ~n5124 & n5171 ) | ( n5167 & n5171 ) ;
  assign n5173 = n4960 & ~n5171 ;
  assign n5174 = ( n5125 & n5172 ) | ( n5125 & ~n5173 ) | ( n5172 & ~n5173 ) ;
  assign n5175 = n5120 | n5174 ;
  assign n5176 = ( ~n4874 & n4963 ) | ( ~n4874 & n5175 ) | ( n4963 & n5175 ) ;
  assign n5177 = n4875 | n5176 ;
  buffer buf_n5178( .i (n47), .o (n5178) );
  buffer buf_n5179( .i (n5178), .o (n5179) );
  assign n5180 = ~n4316 & n5179 ;
  buffer buf_n5181( .i (n5180), .o (n5181) );
  buffer buf_n5182( .i (n5181), .o (n5182) );
  buffer buf_n5183( .i (n5182), .o (n5183) );
  buffer buf_n5184( .i (n5183), .o (n5184) );
  buffer buf_n5185( .i (n5184), .o (n5185) );
  buffer buf_n5186( .i (n5185), .o (n5186) );
  buffer buf_n5187( .i (n5186), .o (n5187) );
  buffer buf_n5188( .i (n5187), .o (n5188) );
  buffer buf_n5189( .i (n5188), .o (n5189) );
  buffer buf_n5190( .i (n5189), .o (n5190) );
  buffer buf_n5191( .i (n5190), .o (n5191) );
  buffer buf_n5192( .i (n4790), .o (n5192) );
  buffer buf_n5193( .i (n5192), .o (n5193) );
  assign n5194 = ( ~n4926 & n5191 ) | ( ~n4926 & n5193 ) | ( n5191 & n5193 ) ;
  buffer buf_n5195( .i (n4954), .o (n5195) );
  assign n5196 = ( ~n5191 & n5193 ) | ( ~n5191 & n5195 ) | ( n5193 & n5195 ) ;
  assign n5197 = ( n178 & n5194 ) | ( n178 & ~n5196 ) | ( n5194 & ~n5196 ) ;
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n5198( .i (n5160), .o (n5198) );
  assign n5199 = ( n824 & ~n4887 ) | ( n824 & n5198 ) | ( ~n4887 & n5198 ) ;
  assign n5200 = ~n4954 & n5199 ;
  buffer buf_n5201( .i (n5200), .o (n5201) );
  buffer buf_n5202( .i (n5201), .o (n5202) );
  assign n5203 = n236 | n5201 ;
  assign n5204 = ( n5197 & n5202 ) | ( n5197 & n5203 ) | ( n5202 & n5203 ) ;
  assign n5205 = n92 | n5204 ;
  buffer buf_n4900( .i (n4899), .o (n4900) );
  buffer buf_n4901( .i (n4900), .o (n4901) );
  assign n5206 = ( n3421 & n4901 ) | ( n3421 & ~n5195 ) | ( n4901 & ~n5195 ) ;
  assign n5207 = ( n4900 & n4954 ) | ( n4900 & ~n5192 ) | ( n4954 & ~n5192 ) ;
  buffer buf_n5208( .i (n3418), .o (n5208) );
  assign n5209 = ( n3421 & ~n5207 ) | ( n3421 & n5208 ) | ( ~n5207 & n5208 ) ;
  assign n5210 = ~n5206 & n5209 ;
  assign n5211 = ~n3416 & n5210 ;
  assign n5212 = n92 & ~n5211 ;
  assign n5213 = n5205 & ~n5212 ;
  buffer buf_n5214( .i (n5213), .o (n5214) );
  buffer buf_n5215( .i (n5214), .o (n5215) );
  assign n5216 = ( n669 & ~n1803 ) | ( n669 & n2610 ) | ( ~n1803 & n2610 ) ;
  buffer buf_n5217( .i (n5216), .o (n5217) );
  buffer buf_n5218( .i (n5217), .o (n5218) );
  buffer buf_n5219( .i (n5218), .o (n5219) );
  buffer buf_n5220( .i (n5219), .o (n5220) );
  buffer buf_n5221( .i (n5220), .o (n5221) );
  buffer buf_n5222( .i (n5221), .o (n5222) );
  buffer buf_n5223( .i (n5222), .o (n5223) );
  buffer buf_n5224( .i (n5223), .o (n5224) );
  buffer buf_n5225( .i (n5224), .o (n5225) );
  buffer buf_n5226( .i (n5225), .o (n5226) );
  assign n5227 = n5214 & ~n5226 ;
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n3190( .i (n3189), .o (n3190) );
  buffer buf_n3191( .i (n3190), .o (n3191) );
  buffer buf_n3192( .i (n3191), .o (n3192) );
  buffer buf_n3193( .i (n3192), .o (n3193) );
  buffer buf_n3194( .i (n3193), .o (n3194) );
  buffer buf_n3195( .i (n3194), .o (n3195) );
  buffer buf_n3196( .i (n3195), .o (n3196) );
  buffer buf_n3197( .i (n3196), .o (n3197) );
  buffer buf_n3198( .i (n3197), .o (n3198) );
  buffer buf_n3199( .i (n3198), .o (n3199) );
  buffer buf_n3200( .i (n3199), .o (n3200) );
  assign n5228 = ( ~n3897 & n4740 ) | ( ~n3897 & n5179 ) | ( n4740 & n5179 ) ;
  buffer buf_n5229( .i (n5228), .o (n5229) );
  buffer buf_n5230( .i (n5229), .o (n5230) );
  buffer buf_n5231( .i (n5230), .o (n5231) );
  buffer buf_n5232( .i (n5231), .o (n5232) );
  buffer buf_n5233( .i (n5232), .o (n5233) );
  buffer buf_n5234( .i (n5233), .o (n5234) );
  buffer buf_n5235( .i (n5234), .o (n5235) );
  buffer buf_n5236( .i (n5235), .o (n5236) );
  buffer buf_n5237( .i (n5236), .o (n5237) );
  assign n5238 = n3200 & ~n5237 ;
  buffer buf_n5239( .i (n4617), .o (n5239) );
  assign n5240 = n5238 | n5239 ;
  buffer buf_n4591( .i (n4590), .o (n4591) );
  buffer buf_n4592( .i (n4591), .o (n4592) );
  buffer buf_n4593( .i (n4592), .o (n4593) );
  buffer buf_n4594( .i (n4593), .o (n4594) );
  buffer buf_n4595( .i (n4594), .o (n4595) );
  assign n5241 = n4595 | n5055 ;
  assign n5242 = n5198 | n5241 ;
  assign n5243 = n5239 & n5242 ;
  assign n5244 = n5240 & ~n5243 ;
  buffer buf_n5245( .i (n5244), .o (n5245) );
  buffer buf_n5246( .i (n5245), .o (n5246) );
  buffer buf_n3602( .i (n3601), .o (n3602) );
  buffer buf_n3603( .i (n3602), .o (n3603) );
  buffer buf_n3604( .i (n3603), .o (n3604) );
  buffer buf_n3605( .i (n3604), .o (n3605) );
  buffer buf_n3606( .i (n3605), .o (n3606) );
  buffer buf_n3607( .i (n3606), .o (n3607) );
  buffer buf_n3608( .i (n3607), .o (n3608) );
  buffer buf_n3609( .i (n3608), .o (n3609) );
  assign n5247 = n3609 & n5245 ;
  assign n5248 = n517 & n708 ;
  assign n5249 = ( n402 & ~n928 ) | ( n402 & n5248 ) | ( ~n928 & n5248 ) ;
  assign n5250 = n929 & n5249 ;
  buffer buf_n5251( .i (n4766), .o (n5251) );
  assign n5252 = ( ~n4741 & n5000 ) | ( ~n4741 & n5251 ) | ( n5000 & n5251 ) ;
  buffer buf_n5253( .i (n5252), .o (n5253) );
  buffer buf_n5254( .i (n5253), .o (n5254) );
  buffer buf_n5255( .i (n5254), .o (n5255) );
  buffer buf_n5256( .i (n5255), .o (n5256) );
  assign n5258 = ( n4800 & ~n5019 ) | ( n4800 & n5256 ) | ( ~n5019 & n5256 ) ;
  assign n5259 = ~n4415 & n5255 ;
  assign n5260 = ( ~n3883 & n5256 ) | ( ~n3883 & n5259 ) | ( n5256 & n5259 ) ;
  assign n5261 = n5258 | n5260 ;
  assign n5262 = n4792 & n5261 ;
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  assign n5263 = n551 | n4902 ;
  assign n5264 = ~n4792 & n5263 ;
  assign n5265 = n5262 | n5264 ;
  assign n5266 = n4922 & ~n5265 ;
  assign n5267 = ~n44 & n246 ;
  buffer buf_n5268( .i (n5267), .o (n5268) );
  buffer buf_n5269( .i (n5268), .o (n5269) );
  buffer buf_n5270( .i (n5269), .o (n5270) );
  buffer buf_n5271( .i (n5270), .o (n5271) );
  buffer buf_n5272( .i (n5271), .o (n5272) );
  buffer buf_n5273( .i (n5272), .o (n5273) );
  buffer buf_n5274( .i (n5273), .o (n5274) );
  buffer buf_n5275( .i (n5274), .o (n5275) );
  buffer buf_n5276( .i (n5275), .o (n5276) );
  buffer buf_n5277( .i (n5276), .o (n5277) );
  buffer buf_n5278( .i (n5277), .o (n5278) );
  buffer buf_n5279( .i (n5278), .o (n5279) );
  assign n5280 = ( n1362 & n4665 ) | ( n1362 & n5275 ) | ( n4665 & n5275 ) ;
  buffer buf_n5281( .i (n5280), .o (n5281) );
  buffer buf_n5282( .i (n5281), .o (n5282) );
  buffer buf_n5283( .i (n5282), .o (n5283) );
  buffer buf_n5284( .i (n4417), .o (n5284) );
  assign n5285 = ( ~n5086 & n5281 ) | ( ~n5086 & n5284 ) | ( n5281 & n5284 ) ;
  assign n5286 = ( ~n4916 & n5278 ) | ( ~n4916 & n5285 ) | ( n5278 & n5285 ) ;
  assign n5287 = ( ~n5279 & n5283 ) | ( ~n5279 & n5286 ) | ( n5283 & n5286 ) ;
  assign n5288 = ~n550 & n831 ;
  buffer buf_n5289( .i (n5288), .o (n5289) );
  buffer buf_n5290( .i (n5289), .o (n5290) );
  assign n5291 = n4753 | n5289 ;
  assign n5292 = ( n5287 & n5290 ) | ( n5287 & n5291 ) | ( n5290 & n5291 ) ;
  buffer buf_n5293( .i (n5055), .o (n5293) );
  assign n5294 = n5292 | n5293 ;
  assign n5295 = ( ~n4451 & n5266 ) | ( ~n4451 & n5294 ) | ( n5266 & n5294 ) ;
  buffer buf_n5296( .i (n4106), .o (n5296) );
  assign n5297 = ( ~n4926 & n5295 ) | ( ~n4926 & n5296 ) | ( n5295 & n5296 ) ;
  buffer buf_n5298( .i (n3899), .o (n5298) );
  buffer buf_n5299( .i (n5298), .o (n5299) );
  assign n5300 = ~n3006 & n5299 ;
  assign n5301 = ~n4415 & n5300 ;
  buffer buf_n5302( .i (n5301), .o (n5302) );
  buffer buf_n5303( .i (n5302), .o (n5303) );
  buffer buf_n5304( .i (n5284), .o (n5304) );
  assign n5305 = n5302 & ~n5304 ;
  buffer buf_n5306( .i (n4343), .o (n5306) );
  buffer buf_n5307( .i (n5306), .o (n5307) );
  assign n5308 = n395 & n5307 ;
  assign n5309 = ~n333 & n5308 ;
  assign n5310 = ( n4739 & n4765 ) | ( n4739 & ~n5146 ) | ( n4765 & ~n5146 ) ;
  buffer buf_n5311( .i (n5310), .o (n5311) );
  buffer buf_n5316( .i (n4740), .o (n5316) );
  assign n5317 = ( n5000 & n5311 ) | ( n5000 & ~n5316 ) | ( n5311 & ~n5316 ) ;
  buffer buf_n5318( .i (n5317), .o (n5318) );
  buffer buf_n5319( .i (n5318), .o (n5319) );
  buffer buf_n5320( .i (n5319), .o (n5320) );
  buffer buf_n5321( .i (n5320), .o (n5321) );
  assign n5322 = ( n4494 & ~n4973 ) | ( n4494 & n5318 ) | ( ~n4973 & n5318 ) ;
  buffer buf_n5323( .i (n5322), .o (n5323) );
  buffer buf_n5324( .i (n5323), .o (n5324) );
  buffer buf_n5312( .i (n5311), .o (n5312) );
  buffer buf_n5313( .i (n5312), .o (n5313) );
  buffer buf_n5314( .i (n5313), .o (n5314) );
  buffer buf_n5315( .i (n5314), .o (n5315) );
  assign n5325 = ~n5315 & n5323 ;
  assign n5326 = ( ~n5321 & n5324 ) | ( ~n5321 & n5325 ) | ( n5324 & n5325 ) ;
  assign n5327 = n5309 | n5326 ;
  assign n5328 = ( n5303 & ~n5305 ) | ( n5303 & n5327 ) | ( ~n5305 & n5327 ) ;
  assign n5329 = n5160 | n5328 ;
  buffer buf_n5330( .i (n4405), .o (n5330) );
  assign n5331 = n5284 & ~n5330 ;
  buffer buf_n5332( .i (n4523), .o (n5332) );
  assign n5333 = ( n1479 & ~n4985 ) | ( n1479 & n5332 ) | ( ~n4985 & n5332 ) ;
  assign n5334 = n1480 | n5333 ;
  assign n5335 = ~n5331 & n5334 ;
  buffer buf_n5336( .i (n5109), .o (n5336) );
  assign n5337 = n5335 & ~n5336 ;
  assign n5338 = n5160 & ~n5337 ;
  assign n5339 = n5329 & ~n5338 ;
  assign n5340 = ( n3584 & ~n4337 ) | ( n3584 & n5306 ) | ( ~n4337 & n5306 ) ;
  buffer buf_n5341( .i (n5340), .o (n5341) );
  assign n5344 = n5330 & n5341 ;
  buffer buf_n5345( .i (n5344), .o (n5345) );
  buffer buf_n5346( .i (n5345), .o (n5346) );
  buffer buf_n5342( .i (n5341), .o (n5342) );
  buffer buf_n5343( .i (n5342), .o (n5343) );
  assign n5347 = n5343 & ~n5345 ;
  assign n5348 = ( n4729 & ~n5346 ) | ( n4729 & n5347 ) | ( ~n5346 & n5347 ) ;
  assign n5349 = ( n4790 & ~n5293 ) | ( n4790 & n5348 ) | ( ~n5293 & n5348 ) ;
  assign n5350 = ( n401 & ~n5339 ) | ( n401 & n5349 ) | ( ~n5339 & n5349 ) ;
  assign n5351 = ( n4926 & n5296 ) | ( n4926 & n5350 ) | ( n5296 & n5350 ) ;
  assign n5352 = n5297 & ~n5351 ;
  assign n5353 = n5250 | n5352 ;
  assign n5354 = ( n5246 & ~n5247 ) | ( n5246 & n5353 ) | ( ~n5247 & n5353 ) ;
  assign n5355 = n93 | n5354 ;
  buffer buf_n4346( .i (n4345), .o (n4346) );
  buffer buf_n4347( .i (n4346), .o (n4347) );
  buffer buf_n4348( .i (n4347), .o (n4348) );
  buffer buf_n4349( .i (n4348), .o (n4349) );
  buffer buf_n4350( .i (n4349), .o (n4350) );
  buffer buf_n4351( .i (n4350), .o (n4351) );
  buffer buf_n4352( .i (n4351), .o (n4352) );
  buffer buf_n4353( .i (n4352), .o (n4353) );
  buffer buf_n4354( .i (n4353), .o (n4354) );
  assign n5356 = ( n1166 & ~n4742 ) | ( n1166 & n5057 ) | ( ~n4742 & n5057 ) ;
  buffer buf_n5357( .i (n5356), .o (n5357) );
  buffer buf_n5358( .i (n5357), .o (n5358) );
  buffer buf_n5359( .i (n5358), .o (n5359) );
  buffer buf_n5360( .i (n5359), .o (n5360) );
  assign n5361 = ( n4664 & n5299 ) | ( n4664 & n5357 ) | ( n5299 & n5357 ) ;
  buffer buf_n5362( .i (n5361), .o (n5362) );
  buffer buf_n5363( .i (n5362), .o (n5363) );
  assign n5364 = ~n1170 & n5362 ;
  assign n5365 = ( ~n5360 & n5363 ) | ( ~n5360 & n5364 ) | ( n5363 & n5364 ) ;
  buffer buf_n5366( .i (n5098), .o (n5366) );
  buffer buf_n5367( .i (n5366), .o (n5367) );
  assign n5368 = n5365 | n5367 ;
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  assign n5369 = n891 | n5304 ;
  assign n5370 = n5367 & n5369 ;
  assign n5371 = n5368 & ~n5370 ;
  assign n5372 = n5293 & n5371 ;
  buffer buf_n5373( .i (n4222), .o (n5373) );
  assign n5374 = ( n2327 & n4558 ) | ( n2327 & ~n5373 ) | ( n4558 & ~n5373 ) ;
  buffer buf_n5375( .i (n5374), .o (n5375) );
  buffer buf_n5381( .i (n2327), .o (n5381) );
  buffer buf_n5382( .i (n5381), .o (n5382) );
  assign n5383 = ( n5178 & ~n5375 ) | ( n5178 & n5382 ) | ( ~n5375 & n5382 ) ;
  buffer buf_n5384( .i (n5383), .o (n5384) );
  buffer buf_n5385( .i (n5384), .o (n5385) );
  buffer buf_n5386( .i (n5385), .o (n5386) );
  buffer buf_n5387( .i (n5386), .o (n5387) );
  buffer buf_n5388( .i (n5387), .o (n5388) );
  buffer buf_n5376( .i (n5375), .o (n5376) );
  buffer buf_n5377( .i (n5376), .o (n5377) );
  buffer buf_n5378( .i (n5377), .o (n5378) );
  buffer buf_n5389( .i (n3897), .o (n5389) );
  assign n5390 = ( ~n5150 & n5384 ) | ( ~n5150 & n5389 ) | ( n5384 & n5389 ) ;
  assign n5391 = n5378 & n5390 ;
  buffer buf_n5392( .i (n5391), .o (n5392) );
  buffer buf_n5393( .i (n5392), .o (n5393) );
  assign n5394 = n5133 & ~n5392 ;
  assign n5395 = ( n5388 & n5393 ) | ( n5388 & ~n5394 ) | ( n5393 & ~n5394 ) ;
  assign n5396 = n5330 & n5395 ;
  buffer buf_n5397( .i (n5396), .o (n5397) );
  buffer buf_n5398( .i (n5397), .o (n5398) );
  buffer buf_n5399( .i (n5179), .o (n5399) );
  assign n5400 = ( ~n5316 & n5389 ) | ( ~n5316 & n5399 ) | ( n5389 & n5399 ) ;
  assign n5401 = ( n5251 & n5316 ) | ( n5251 & ~n5399 ) | ( n5316 & ~n5399 ) ;
  assign n5402 = n5400 | n5401 ;
  buffer buf_n5403( .i (n5402), .o (n5403) );
  buffer buf_n5404( .i (n5403), .o (n5404) );
  buffer buf_n5405( .i (n5404), .o (n5405) );
  buffer buf_n5406( .i (n5405), .o (n5406) );
  buffer buf_n5407( .i (n5406), .o (n5407) );
  assign n5408 = ~n5397 & n5407 ;
  assign n5409 = ( n4393 & n5398 ) | ( n4393 & ~n5408 ) | ( n5398 & ~n5408 ) ;
  assign n5410 = n5293 | n5409 ;
  buffer buf_n5411( .i (n5055), .o (n5411) );
  buffer buf_n5412( .i (n5411), .o (n5412) );
  assign n5413 = ( n5372 & n5410 ) | ( n5372 & ~n5412 ) | ( n5410 & ~n5412 ) ;
  assign n5414 = n3855 & ~n5413 ;
  buffer buf_n5415( .i (n5399), .o (n5415) );
  assign n5416 = n4643 & n5415 ;
  buffer buf_n5417( .i (n5416), .o (n5417) );
  buffer buf_n5418( .i (n5417), .o (n5418) );
  buffer buf_n5419( .i (n5418), .o (n5419) );
  buffer buf_n5420( .i (n5419), .o (n5420) );
  buffer buf_n5421( .i (n5420), .o (n5421) );
  assign n5422 = n4852 & n5284 ;
  assign n5423 = ( ~n3884 & n5366 ) | ( ~n3884 & n5422 ) | ( n5366 & n5422 ) ;
  assign n5424 = ( n2633 & ~n5421 ) | ( n2633 & n5423 ) | ( ~n5421 & n5423 ) ;
  buffer buf_n5425( .i (n4775), .o (n5425) );
  assign n5426 = n5424 & n5425 ;
  buffer buf_n4444( .i (n4443), .o (n4444) );
  buffer buf_n4445( .i (n4444), .o (n4445) );
  buffer buf_n5427( .i (n4753), .o (n5427) );
  assign n5428 = ( n4445 & n5425 ) | ( n4445 & ~n5427 ) | ( n5425 & ~n5427 ) ;
  assign n5429 = ( ~n660 & n5426 ) | ( ~n660 & n5428 ) | ( n5426 & n5428 ) ;
  assign n5430 = n4731 & n5429 ;
  assign n5431 = n3855 | n5430 ;
  assign n5432 = ~n5414 & n5431 ;
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n5433( .i (n5367), .o (n5433) );
  assign n5434 = ( n1614 & n4729 ) | ( n1614 & ~n5433 ) | ( n4729 & ~n5433 ) ;
  buffer buf_n5435( .i (n4985), .o (n5435) );
  buffer buf_n5436( .i (n5435), .o (n5436) );
  buffer buf_n5437( .i (n5436), .o (n5437) );
  assign n5438 = ( ~n1613 & n5090 ) | ( ~n1613 & n5437 ) | ( n5090 & n5437 ) ;
  assign n5439 = ( n5425 & ~n5433 ) | ( n5425 & n5438 ) | ( ~n5433 & n5438 ) ;
  assign n5440 = ~n5434 & n5439 ;
  assign n5441 = n4106 & ~n5440 ;
  buffer buf_n5070( .i (n5069), .o (n5070) );
  assign n5442 = n280 & ~n5070 ;
  buffer buf_n5443( .i (n4394), .o (n5443) );
  assign n5444 = n5442 | n5443 ;
  assign n5445 = ~n5441 & n5444 ;
  assign n5446 = ( n3856 & ~n5165 ) | ( n3856 & n5445 ) | ( ~n5165 & n5445 ) ;
  assign n5447 = ( ~n4354 & n5432 ) | ( ~n4354 & n5446 ) | ( n5432 & n5446 ) ;
  assign n5448 = ~n4960 & n5447 ;
  assign n5449 = n93 & ~n5448 ;
  assign n5450 = n5355 & ~n5449 ;
  assign n5451 = ( n4978 & ~n5316 ) | ( n4978 & n5389 ) | ( ~n5316 & n5389 ) ;
  buffer buf_n5452( .i (n5451), .o (n5452) );
  buffer buf_n5453( .i (n5452), .o (n5453) );
  buffer buf_n5454( .i (n5453), .o (n5454) );
  assign n5461 = ( n5017 & n5332 ) | ( n5017 & n5454 ) | ( n5332 & n5454 ) ;
  buffer buf_n5462( .i (n5461), .o (n5462) );
  buffer buf_n5463( .i (n5462), .o (n5463) );
  buffer buf_n5464( .i (n5463), .o (n5464) );
  buffer buf_n5455( .i (n5454), .o (n5455) );
  buffer buf_n5456( .i (n5455), .o (n5456) );
  buffer buf_n5457( .i (n5456), .o (n5457) );
  assign n5465 = ( n5304 & n5436 ) | ( n5304 & ~n5462 ) | ( n5436 & ~n5462 ) ;
  assign n5466 = n5457 & n5465 ;
  assign n5467 = ( n5433 & ~n5464 ) | ( n5433 & n5466 ) | ( ~n5464 & n5466 ) ;
  buffer buf_n5468( .i (n5112), .o (n5468) );
  assign n5469 = ~n5467 & n5468 ;
  assign n5470 = ~n1474 & n5304 ;
  buffer buf_n5471( .i (n4849), .o (n5471) );
  buffer buf_n5472( .i (n5471), .o (n5472) );
  buffer buf_n5473( .i (n5472), .o (n5473) );
  assign n5474 = ( ~n1475 & n5470 ) | ( ~n1475 & n5473 ) | ( n5470 & n5473 ) ;
  assign n5475 = n5433 & n5474 ;
  assign n5476 = n5468 | n5475 ;
  assign n5477 = ~n5469 & n5476 ;
  assign n5478 = n3855 & ~n5477 ;
  buffer buf_n5479( .i (n5133), .o (n5479) );
  assign n5480 = ( ~n3961 & n5332 ) | ( ~n3961 & n5479 ) | ( n5332 & n5479 ) ;
  buffer buf_n5481( .i (n5480), .o (n5481) );
  buffer buf_n5482( .i (n5481), .o (n5482) );
  buffer buf_n5483( .i (n5482), .o (n5483) );
  buffer buf_n5484( .i (n5483), .o (n5484) );
  assign n5485 = ( n4859 & n5472 ) | ( n4859 & ~n5481 ) | ( n5472 & ~n5481 ) ;
  buffer buf_n5486( .i (n5485), .o (n5486) );
  buffer buf_n5487( .i (n5486), .o (n5487) );
  assign n5488 = ~n3965 & n5486 ;
  assign n5489 = ( n5484 & n5487 ) | ( n5484 & n5488 ) | ( n5487 & n5488 ) ;
  assign n5490 = ~n3418 & n5489 ;
  buffer buf_n5491( .i (n5126), .o (n5491) );
  assign n5492 = n5490 | n5491 ;
  assign n5493 = ~n5478 & n5492 ;
  buffer buf_n5494( .i (n4927), .o (n5494) );
  assign n5495 = n5493 | n5494 ;
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n2100( .i (n2099), .o (n2100) );
  buffer buf_n5496( .i (n401), .o (n5496) );
  assign n5497 = ~n2100 & n5496 ;
  assign n5498 = ~n317 & n5497 ;
  assign n5499 = n5494 & ~n5498 ;
  assign n5500 = n5495 & ~n5499 ;
  assign n5501 = n181 & n5500 ;
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n5502( .i (n4835), .o (n5502) );
  buffer buf_n5503( .i (n5502), .o (n5503) );
  buffer buf_n5504( .i (n5332), .o (n5504) );
  buffer buf_n5505( .i (n5504), .o (n5505) );
  assign n5506 = ( n5109 & n5503 ) | ( n5109 & ~n5505 ) | ( n5503 & ~n5505 ) ;
  buffer buf_n5507( .i (n5506), .o (n5507) );
  buffer buf_n5508( .i (n5507), .o (n5508) );
  buffer buf_n5509( .i (n5508), .o (n5509) );
  buffer buf_n5510( .i (n5509), .o (n5510) );
  assign n5511 = n5071 & ~n5507 ;
  buffer buf_n5512( .i (n5511), .o (n5512) );
  buffer buf_n5513( .i (n5512), .o (n5513) );
  buffer buf_n5514( .i (n5198), .o (n5514) );
  buffer buf_n5515( .i (n5468), .o (n5515) );
  assign n5516 = ( n5512 & n5514 ) | ( n5512 & n5515 ) | ( n5514 & n5515 ) ;
  assign n5517 = ( ~n5510 & n5513 ) | ( ~n5510 & n5516 ) | ( n5513 & n5516 ) ;
  assign n5518 = ( ~n1204 & n4927 ) | ( ~n1204 & n5517 ) | ( n4927 & n5517 ) ;
  buffer buf_n5519( .i (n707), .o (n5519) );
  assign n5520 = ( n4351 & n5515 ) | ( n4351 & n5519 ) | ( n5515 & n5519 ) ;
  assign n5521 = ~n5128 & n5520 ;
  assign n5522 = ~n1204 & n5521 ;
  assign n5523 = ( ~n5494 & n5518 ) | ( ~n5494 & n5522 ) | ( n5518 & n5522 ) ;
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n5524( .i (n4579), .o (n5524) );
  assign n5525 = n393 & ~n5524 ;
  buffer buf_n5526( .i (n5525), .o (n5526) );
  buffer buf_n5527( .i (n5526), .o (n5527) );
  buffer buf_n5528( .i (n5527), .o (n5528) );
  buffer buf_n5529( .i (n5528), .o (n5529) );
  buffer buf_n5530( .i (n5529), .o (n5530) );
  buffer buf_n5531( .i (n5530), .o (n5531) );
  buffer buf_n5532( .i (n5531), .o (n5532) );
  buffer buf_n5533( .i (n5532), .o (n5533) );
  buffer buf_n5534( .i (n5533), .o (n5534) );
  assign n5535 = n1405 & ~n5534 ;
  buffer buf_n4236( .i (n4235), .o (n4236) );
  buffer buf_n4237( .i (n4236), .o (n4237) );
  assign n5536 = ( n755 & n4237 ) | ( n755 & n5412 ) | ( n4237 & n5412 ) ;
  assign n5537 = ~n4001 & n5536 ;
  buffer buf_n5538( .i (n5299), .o (n5538) );
  assign n5539 = ( ~n4231 & n5479 ) | ( ~n4231 & n5538 ) | ( n5479 & n5538 ) ;
  buffer buf_n5540( .i (n5539), .o (n5540) );
  buffer buf_n5541( .i (n5540), .o (n5541) );
  buffer buf_n5542( .i (n5541), .o (n5542) );
  assign n5543 = ( ~n5366 & n5505 ) | ( ~n5366 & n5540 ) | ( n5505 & n5540 ) ;
  assign n5544 = ( n5336 & ~n5437 ) | ( n5336 & n5543 ) | ( ~n5437 & n5543 ) ;
  assign n5545 = n5542 & n5544 ;
  assign n5546 = n3532 & ~n5366 ;
  buffer buf_n5547( .i (n5546), .o (n5547) );
  buffer buf_n5548( .i (n5547), .o (n5548) );
  assign n5549 = n5425 & ~n5547 ;
  assign n5550 = ( n5545 & n5548 ) | ( n5545 & ~n5549 ) | ( n5548 & ~n5549 ) ;
  assign n5551 = ( ~n5239 & n5515 ) | ( ~n5239 & n5550 ) | ( n5515 & n5550 ) ;
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n5552( .i (n5479), .o (n5552) );
  buffer buf_n5553( .i (n5552), .o (n5553) );
  assign n5554 = ( ~n4593 & n5436 ) | ( ~n4593 & n5553 ) | ( n5436 & n5553 ) ;
  assign n5555 = ( ~n4593 & n5109 ) | ( ~n4593 & n5553 ) | ( n5109 & n5553 ) ;
  assign n5556 = ( n2258 & n5554 ) | ( n2258 & ~n5555 ) | ( n5554 & ~n5555 ) ;
  buffer buf_n5557( .i (n5473), .o (n5557) );
  assign n5558 = n5556 | n5557 ;
  assign n5559 = n833 & n2038 ;
  assign n5560 = n5557 & ~n5559 ;
  assign n5561 = n5558 & ~n5560 ;
  assign n5562 = ( n5239 & n5515 ) | ( n5239 & ~n5561 ) | ( n5515 & ~n5561 ) ;
  assign n5563 = n5551 & ~n5562 ;
  assign n5564 = n5537 | n5563 ;
  assign n5565 = ( n1406 & ~n5535 ) | ( n1406 & n5564 ) | ( ~n5535 & n5564 ) ;
  assign n5566 = n5523 | n5565 ;
  assign n5567 = ~n181 & n5566 ;
  assign n5568 = n5501 | n5567 ;
  assign n5569 = n5450 | n5568 ;
  assign n5570 = ( n5215 & ~n5227 ) | ( n5215 & n5569 ) | ( ~n5227 & n5569 ) ;
  buffer buf_n5571( .i (n5307), .o (n5571) );
  buffer buf_n5572( .i (n5571), .o (n5572) );
  assign n5573 = ( ~n3719 & n5505 ) | ( ~n3719 & n5572 ) | ( n5505 & n5572 ) ;
  buffer buf_n5574( .i (n5573), .o (n5574) );
  assign n5575 = ( ~n5071 & n5557 ) | ( ~n5071 & n5574 ) | ( n5557 & n5574 ) ;
  assign n5576 = ( n4904 & n5557 ) | ( n4904 & ~n5574 ) | ( n5557 & ~n5574 ) ;
  assign n5577 = n5575 & ~n5576 ;
  buffer buf_n5578( .i (n5577), .o (n5578) );
  buffer buf_n5579( .i (n5578), .o (n5579) );
  buffer buf_n5580( .i (n4061), .o (n5580) );
  buffer buf_n5581( .i (n5580), .o (n5581) );
  buffer buf_n5582( .i (n5581), .o (n5582) );
  assign n5583 = ( ~n5195 & n5578 ) | ( ~n5195 & n5582 ) | ( n5578 & n5582 ) ;
  buffer buf_n4035( .i (n4034), .o (n4035) );
  buffer buf_n4036( .i (n4035), .o (n4036) );
  buffer buf_n4037( .i (n4036), .o (n4037) );
  assign n5584 = n3851 & ~n4037 ;
  assign n5585 = ~n5582 & n5584 ;
  assign n5586 = ( n5579 & ~n5583 ) | ( n5579 & n5585 ) | ( ~n5583 & n5585 ) ;
  buffer buf_n5587( .i (n5586), .o (n5587) );
  buffer buf_n5588( .i (n5587), .o (n5588) );
  buffer buf_n4054( .i (n4053), .o (n4054) );
  buffer buf_n4055( .i (n4054), .o (n4055) );
  buffer buf_n4056( .i (n4055), .o (n4056) );
  buffer buf_n4057( .i (n4056), .o (n4057) );
  buffer buf_n4058( .i (n4057), .o (n4058) );
  buffer buf_n4059( .i (n4058), .o (n4059) );
  assign n5589 = ( n4523 & n4664 ) | ( n4523 & n5306 ) | ( n4664 & n5306 ) ;
  assign n5590 = ( ~n4849 & n5307 ) | ( ~n4849 & n5589 ) | ( n5307 & n5589 ) ;
  buffer buf_n5591( .i (n5590), .o (n5591) );
  assign n5594 = n5572 & ~n5591 ;
  buffer buf_n5595( .i (n5594), .o (n5595) );
  buffer buf_n5596( .i (n5595), .o (n5596) );
  buffer buf_n5592( .i (n5591), .o (n5592) );
  buffer buf_n5593( .i (n5592), .o (n5593) );
  assign n5597 = n5593 | n5595 ;
  buffer buf_n5598( .i (n5071), .o (n5598) );
  assign n5599 = ( n5596 & n5597 ) | ( n5596 & ~n5598 ) | ( n5597 & ~n5598 ) ;
  buffer buf_n5600( .i (n5599), .o (n5600) );
  buffer buf_n5601( .i (n5600), .o (n5601) );
  buffer buf_n3822( .i (n3821), .o (n3822) );
  assign n5602 = ( n3822 & n5195 ) | ( n3822 & ~n5600 ) | ( n5195 & ~n5600 ) ;
  assign n5603 = n5601 & n5602 ;
  buffer buf_n5604( .i (n5603), .o (n5604) );
  assign n5605 = ( n4059 & ~n5587 ) | ( n4059 & n5604 ) | ( ~n5587 & n5604 ) ;
  buffer buf_n5606( .i (n4911), .o (n5606) );
  assign n5607 = ~n5604 & n5606 ;
  assign n5608 = ( n5588 & n5605 ) | ( n5588 & ~n5607 ) | ( n5605 & ~n5607 ) ;
  buffer buf_n5609( .i (n5608), .o (n5609) );
  buffer buf_n5610( .i (n5609), .o (n5610) );
  buffer buf_n5611( .i (n358), .o (n5611) );
  assign n5612 = n5609 & ~n5611 ;
  buffer buf_n5613( .i (n4494), .o (n5613) );
  buffer buf_n5614( .i (n5613), .o (n5614) );
  assign n5615 = ( ~n1571 & n4425 ) | ( ~n1571 & n5614 ) | ( n4425 & n5614 ) ;
  assign n5616 = ( n1570 & ~n3921 ) | ( n1570 & n4664 ) | ( ~n3921 & n4664 ) ;
  buffer buf_n5617( .i (n4834), .o (n5617) );
  assign n5618 = ( n5614 & n5616 ) | ( n5614 & ~n5617 ) | ( n5616 & ~n5617 ) ;
  assign n5619 = n5615 & ~n5618 ;
  assign n5620 = ~n5436 & n5619 ;
  buffer buf_n5621( .i (n5620), .o (n5621) );
  buffer buf_n5622( .i (n5621), .o (n5622) );
  buffer buf_n2206( .i (n2205), .o (n2206) );
  buffer buf_n2207( .i (n2206), .o (n2207) );
  buffer buf_n2208( .i (n2207), .o (n2208) );
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n5080( .i (n5079), .o (n5080) );
  buffer buf_n5081( .i (n5080), .o (n5081) );
  buffer buf_n5623( .i (n3719), .o (n5623) );
  assign n5624 = ( n2210 & n5081 ) | ( n2210 & ~n5623 ) | ( n5081 & ~n5623 ) ;
  assign n5625 = n5621 | n5624 ;
  assign n5626 = ( n5580 & n5622 ) | ( n5580 & n5625 ) | ( n5622 & n5625 ) ;
  assign n5627 = n5412 & ~n5626 ;
  buffer buf_n3778( .i (n3777), .o (n3778) );
  buffer buf_n3779( .i (n3778), .o (n3779) );
  buffer buf_n3780( .i (n3779), .o (n3780) );
  buffer buf_n3781( .i (n3780), .o (n3781) );
  buffer buf_n3782( .i (n3781), .o (n3782) );
  assign n5628 = n3779 & ~n5435 ;
  buffer buf_n5629( .i (n5628), .o (n5629) );
  buffer buf_n5630( .i (n5629), .o (n5630) );
  assign n5631 = ( n4840 & n5623 ) | ( n4840 & ~n5629 ) | ( n5623 & ~n5629 ) ;
  assign n5632 = ( n3782 & n5630 ) | ( n3782 & ~n5631 ) | ( n5630 & ~n5631 ) ;
  assign n5633 = ~n5580 & n5632 ;
  assign n5634 = n5412 | n5633 ;
  assign n5635 = ~n5627 & n5634 ;
  buffer buf_n5636( .i (n5635), .o (n5636) );
  buffer buf_n5637( .i (n5636), .o (n5637) );
  assign n5638 = n4787 & n5636 ;
  buffer buf_n1003( .i (n1002), .o (n1003) );
  assign n5639 = ( n925 & n1003 ) | ( n925 & n2737 ) | ( n1003 & n2737 ) ;
  buffer buf_n5640( .i (n925), .o (n5640) );
  assign n5641 = ( ~n4730 & n5639 ) | ( ~n4730 & n5640 ) | ( n5639 & n5640 ) ;
  buffer buf_n5642( .i (n5641), .o (n5642) );
  buffer buf_n5643( .i (n5642), .o (n5643) );
  assign n5644 = ( ~n732 & n4001 ) | ( ~n732 & n5642 ) | ( n4001 & n5642 ) ;
  assign n5645 = n5643 & ~n5644 ;
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n2845( .i (n2844), .o (n2845) );
  buffer buf_n2846( .i (n2845), .o (n2846) );
  buffer buf_n2847( .i (n2846), .o (n2847) );
  assign n5646 = ( n2847 & n3008 ) | ( n2847 & n5552 ) | ( n3008 & n5552 ) ;
  assign n5647 = ~n3009 & n5646 ;
  buffer buf_n5648( .i (n5647), .o (n5648) );
  buffer buf_n5649( .i (n5648), .o (n5649) );
  buffer buf_n5650( .i (n5649), .o (n5650) );
  buffer buf_n2520( .i (n2519), .o (n2520) );
  buffer buf_n2521( .i (n2520), .o (n2521) );
  buffer buf_n2522( .i (n2521), .o (n2522) );
  buffer buf_n5651( .i (n5473), .o (n5651) );
  assign n5652 = ( n2522 & n5648 ) | ( n2522 & ~n5651 ) | ( n5648 & ~n5651 ) ;
  assign n5653 = n541 & ~n5652 ;
  assign n5654 = ( n542 & n5650 ) | ( n542 & ~n5653 ) | ( n5650 & ~n5653 ) ;
  assign n5655 = n5582 | n5654 ;
  buffer buf_n4511( .i (n4510), .o (n4511) );
  buffer buf_n4512( .i (n4511), .o (n4512) );
  buffer buf_n4513( .i (n4512), .o (n4513) );
  buffer buf_n4514( .i (n4513), .o (n4514) );
  buffer buf_n4515( .i (n4514), .o (n4515) );
  buffer buf_n4516( .i (n4515), .o (n4516) );
  buffer buf_n4517( .i (n4516), .o (n4517) );
  buffer buf_n4518( .i (n4517), .o (n4518) );
  assign n5656 = n315 | n4518 ;
  assign n5657 = n5582 & n5656 ;
  assign n5658 = n5655 & ~n5657 ;
  assign n5659 = n5645 | n5658 ;
  assign n5660 = ( n5637 & ~n5638 ) | ( n5637 & n5659 ) | ( ~n5638 & n5659 ) ;
  assign n5661 = n3489 | n5660 ;
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n5662( .i (n5623), .o (n5662) );
  assign n5663 = ( n958 & ~n5427 ) | ( n958 & n5662 ) | ( ~n5427 & n5662 ) ;
  buffer buf_n5664( .i (n5090), .o (n5664) );
  assign n5665 = ( ~n958 & n5427 ) | ( ~n958 & n5664 ) | ( n5427 & n5664 ) ;
  assign n5666 = ( ~n459 & n5663 ) | ( ~n459 & n5665 ) | ( n5663 & n5665 ) ;
  buffer buf_n5667( .i (n5411), .o (n5667) );
  assign n5668 = ~n5666 & n5667 ;
  buffer buf_n612( .i (n611), .o (n612) );
  assign n5669 = n612 & n5468 ;
  assign n5670 = n5667 | n5669 ;
  assign n5671 = ~n5668 & n5670 ;
  buffer buf_n5672( .i (n5514), .o (n5672) );
  buffer buf_n5673( .i (n5672), .o (n5673) );
  assign n5674 = n5671 & n5673 ;
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  assign n5675 = ( n1384 & n4852 ) | ( n1384 & ~n5079 ) | ( n4852 & ~n5079 ) ;
  buffer buf_n5676( .i (n5675), .o (n5676) );
  buffer buf_n5677( .i (n5676), .o (n5677) );
  buffer buf_n5678( .i (n5677), .o (n5678) );
  assign n5679 = ( n5437 & ~n5623 ) | ( n5437 & n5676 ) | ( ~n5623 & n5676 ) ;
  assign n5680 = ( n1387 & ~n5112 ) | ( n1387 & n5679 ) | ( ~n5112 & n5679 ) ;
  assign n5681 = ( ~n1388 & n5678 ) | ( ~n1388 & n5680 ) | ( n5678 & n5680 ) ;
  assign n5682 = ~n5667 & n5681 ;
  buffer buf_n5683( .i (n5112), .o (n5683) );
  assign n5684 = n1217 & ~n5683 ;
  assign n5685 = n5667 & ~n5684 ;
  assign n5686 = n5682 | n5685 ;
  assign n5687 = ~n5673 & n5686 ;
  assign n5688 = ( n4787 & ~n5674 ) | ( n4787 & n5687 ) | ( ~n5674 & n5687 ) ;
  assign n5689 = n4960 | n5688 ;
  buffer buf_n5690( .i (n120), .o (n5690) );
  assign n5691 = n5689 & n5690 ;
  assign n5692 = n5661 & ~n5691 ;
  assign n5693 = ( n3133 & n5502 ) | ( n3133 & ~n5504 ) | ( n5502 & ~n5504 ) ;
  buffer buf_n5694( .i (n5693), .o (n5694) );
  buffer buf_n5695( .i (n5503), .o (n5695) );
  assign n5696 = n5694 | n5695 ;
  assign n5697 = n5694 & n5695 ;
  assign n5698 = n5696 & ~n5697 ;
  buffer buf_n5699( .i (n5698), .o (n5699) );
  buffer buf_n5700( .i (n5699), .o (n5700) );
  buffer buf_n5701( .i (n4887), .o (n5701) );
  assign n5702 = ( n5581 & n5699 ) | ( n5581 & ~n5701 ) | ( n5699 & ~n5701 ) ;
  buffer buf_n3535( .i (n3534), .o (n3535) );
  assign n5703 = ~n314 & n3535 ;
  assign n5704 = ~n5581 & n5703 ;
  assign n5705 = ( n5700 & ~n5702 ) | ( n5700 & n5704 ) | ( ~n5702 & n5704 ) ;
  buffer buf_n5706( .i (n5705), .o (n5706) );
  buffer buf_n5707( .i (n5706), .o (n5707) );
  assign n5708 = ( n1404 & n2772 ) | ( n1404 & n5193 ) | ( n2772 & n5193 ) ;
  assign n5709 = ~n5165 & n5708 ;
  buffer buf_n2836( .i (n2835), .o (n2836) );
  buffer buf_n2837( .i (n2836), .o (n2837) );
  assign n5710 = n914 & ~n2837 ;
  buffer buf_n5711( .i (n5389), .o (n5711) );
  assign n5712 = ( n3518 & n4643 ) | ( n3518 & n5711 ) | ( n4643 & n5711 ) ;
  buffer buf_n5713( .i (n5712), .o (n5713) );
  buffer buf_n5714( .i (n5713), .o (n5714) );
  buffer buf_n5715( .i (n5714), .o (n5715) );
  assign n5716 = ( n4974 & n5299 ) | ( n4974 & ~n5713 ) | ( n5299 & ~n5713 ) ;
  assign n5717 = n3521 | n5716 ;
  assign n5718 = ( n4852 & ~n5715 ) | ( n4852 & n5717 ) | ( ~n5715 & n5717 ) ;
  assign n5719 = n5572 & ~n5718 ;
  assign n5720 = ~n5695 & n5719 ;
  buffer buf_n4172( .i (n4171), .o (n4172) );
  buffer buf_n4173( .i (n4172), .o (n4173) );
  assign n5721 = ( n4173 & n4655 ) | ( n4173 & ~n5711 ) | ( n4655 & ~n5711 ) ;
  buffer buf_n5722( .i (n5721), .o (n5722) );
  buffer buf_n5725( .i (n5076), .o (n5725) );
  assign n5726 = ~n5722 & n5725 ;
  buffer buf_n5727( .i (n5726), .o (n5727) );
  buffer buf_n5728( .i (n5727), .o (n5728) );
  buffer buf_n5723( .i (n5722), .o (n5723) );
  buffer buf_n5724( .i (n5723), .o (n5724) );
  assign n5729 = n5724 | n5727 ;
  assign n5730 = ( ~n5503 & n5728 ) | ( ~n5503 & n5729 ) | ( n5728 & n5729 ) ;
  assign n5731 = n5526 & ~n5617 ;
  buffer buf_n5732( .i (n5731), .o (n5732) );
  buffer buf_n5733( .i (n5732), .o (n5733) );
  assign n5734 = n5572 | n5732 ;
  assign n5735 = ( n5730 & n5733 ) | ( n5730 & n5734 ) | ( n5733 & n5734 ) ;
  assign n5736 = n5720 | n5735 ;
  assign n5737 = ( n915 & ~n5710 ) | ( n915 & n5736 ) | ( ~n5710 & n5736 ) ;
  assign n5738 = ( n5514 & ~n5581 ) | ( n5514 & n5737 ) | ( ~n5581 & n5737 ) ;
  assign n5739 = ( n4579 & ~n4742 ) | ( n4579 & n5711 ) | ( ~n4742 & n5711 ) ;
  buffer buf_n5740( .i (n5739), .o (n5740) );
  buffer buf_n5741( .i (n5740), .o (n5741) );
  buffer buf_n5742( .i (n5741), .o (n5742) );
  buffer buf_n5743( .i (n5298), .o (n5743) );
  assign n5744 = n5740 & n5743 ;
  buffer buf_n5745( .i (n4523), .o (n5745) );
  assign n5746 = ( n4849 & n5744 ) | ( n4849 & ~n5745 ) | ( n5744 & ~n5745 ) ;
  assign n5747 = ( n1431 & n5742 ) | ( n1431 & ~n5746 ) | ( n5742 & ~n5746 ) ;
  assign n5748 = n3719 | n5747 ;
  assign n5749 = n563 & ~n2094 ;
  buffer buf_n5750( .i (n4643), .o (n5750) );
  buffer buf_n5751( .i (n5750), .o (n5751) );
  buffer buf_n5752( .i (n5751), .o (n5752) );
  buffer buf_n5753( .i (n5752), .o (n5753) );
  buffer buf_n5754( .i (n5753), .o (n5754) );
  assign n5755 = ~n5749 & n5754 ;
  assign n5756 = n5748 & ~n5755 ;
  buffer buf_n5757( .i (n5695), .o (n5757) );
  assign n5758 = n5756 | n5757 ;
  buffer buf_n2056( .i (n2055), .o (n2056) );
  assign n5759 = n398 & n2056 ;
  assign n5760 = n5757 & ~n5759 ;
  assign n5761 = n5758 & ~n5760 ;
  buffer buf_n5762( .i (n5580), .o (n5762) );
  assign n5763 = ( n5514 & ~n5761 ) | ( n5514 & n5762 ) | ( ~n5761 & n5762 ) ;
  assign n5764 = n5738 & ~n5763 ;
  buffer buf_n5765( .i (n5764), .o (n5765) );
  assign n5766 = ( ~n5706 & n5709 ) | ( ~n5706 & n5765 ) | ( n5709 & n5765 ) ;
  assign n5767 = n4261 & ~n5765 ;
  assign n5768 = ( n5707 & n5766 ) | ( n5707 & ~n5767 ) | ( n5766 & ~n5767 ) ;
  assign n5769 = n267 & ~n5768 ;
  buffer buf_n2801( .i (n2800), .o (n2801) );
  buffer buf_n2802( .i (n2801), .o (n2802) );
  buffer buf_n2803( .i (n2802), .o (n2803) );
  buffer buf_n2804( .i (n2803), .o (n2804) );
  buffer buf_n2805( .i (n2804), .o (n2805) );
  buffer buf_n5770( .i (n5505), .o (n5770) );
  assign n5771 = n2805 | n5770 ;
  buffer buf_n2811( .i (n2810), .o (n2811) );
  assign n5772 = n2811 & n5770 ;
  assign n5773 = n5771 & ~n5772 ;
  assign n5774 = n5411 & ~n5773 ;
  assign n5775 = n1003 & n4904 ;
  assign n5776 = n5411 | n5775 ;
  assign n5777 = ~n5774 & n5776 ;
  buffer buf_n5778( .i (n5754), .o (n5778) );
  assign n5779 = n913 & ~n5778 ;
  assign n5780 = n2123 & n5779 ;
  buffer buf_n5781( .i (n5780), .o (n5781) );
  buffer buf_n5782( .i (n5781), .o (n5782) );
  buffer buf_n5783( .i (n5598), .o (n5783) );
  assign n5784 = ~n5781 & n5783 ;
  assign n5785 = ( n5777 & n5782 ) | ( n5777 & ~n5784 ) | ( n5782 & ~n5784 ) ;
  buffer buf_n5786( .i (n4740), .o (n5786) );
  assign n5787 = ( n4978 & ~n5150 ) | ( n4978 & n5786 ) | ( ~n5150 & n5786 ) ;
  buffer buf_n5788( .i (n5786), .o (n5788) );
  assign n5789 = ( ~n5711 & n5787 ) | ( ~n5711 & n5788 ) | ( n5787 & n5788 ) ;
  buffer buf_n5790( .i (n5789), .o (n5790) );
  buffer buf_n5793( .i (n5022), .o (n5793) );
  assign n5794 = ~n5790 & n5793 ;
  buffer buf_n5795( .i (n5794), .o (n5795) );
  buffer buf_n5796( .i (n5795), .o (n5796) );
  buffer buf_n5791( .i (n5790), .o (n5791) );
  buffer buf_n5792( .i (n5791), .o (n5792) );
  assign n5797 = n5792 | n5795 ;
  buffer buf_n5798( .i (n5504), .o (n5798) );
  assign n5799 = ( n5796 & n5797 ) | ( n5796 & ~n5798 ) | ( n5797 & ~n5798 ) ;
  buffer buf_n5800( .i (n5503), .o (n5800) );
  assign n5801 = ( n5336 & n5799 ) | ( n5336 & n5800 ) | ( n5799 & n5800 ) ;
  buffer buf_n5802( .i (n5801), .o (n5802) );
  assign n5803 = ( n5198 & ~n5598 ) | ( n5198 & n5802 ) | ( ~n5598 & n5802 ) ;
  buffer buf_n5804( .i (n5367), .o (n5804) );
  buffer buf_n5805( .i (n5804), .o (n5805) );
  assign n5806 = ( n5683 & ~n5802 ) | ( n5683 & n5805 ) | ( ~n5802 & n5805 ) ;
  assign n5807 = n5803 & ~n5806 ;
  buffer buf_n5808( .i (n5807), .o (n5808) );
  assign n5809 = ( ~n5673 & n5785 ) | ( ~n5673 & n5808 ) | ( n5785 & n5808 ) ;
  assign n5810 = ~n4578 & n5786 ;
  buffer buf_n5811( .i (n5810), .o (n5811) );
  buffer buf_n5812( .i (n5811), .o (n5812) );
  buffer buf_n5813( .i (n5812), .o (n5813) );
  buffer buf_n5814( .i (n5813), .o (n5814) );
  assign n5818 = ( n5435 & ~n5471 ) | ( n5435 & n5814 ) | ( ~n5471 & n5814 ) ;
  assign n5819 = ( n5307 & ~n5538 ) | ( n5307 & n5813 ) | ( ~n5538 & n5813 ) ;
  assign n5820 = ( n5471 & ~n5504 ) | ( n5471 & n5819 ) | ( ~n5504 & n5819 ) ;
  assign n5821 = n5818 | n5820 ;
  buffer buf_n5822( .i (n5821), .o (n5822) );
  buffer buf_n5823( .i (n5822), .o (n5823) );
  assign n5824 = n5757 | n5822 ;
  buffer buf_n1691( .i (n1690), .o (n1691) );
  assign n5825 = n1691 & n2038 ;
  assign n5826 = ( ~n4578 & n4654 ) | ( ~n4578 & n5786 ) | ( n4654 & n5786 ) ;
  buffer buf_n5827( .i (n5826), .o (n5827) );
  assign n5835 = ( n5076 & ~n5298 ) | ( n5076 & n5827 ) | ( ~n5298 & n5827 ) ;
  buffer buf_n5836( .i (n5835), .o (n5836) );
  assign n5839 = n5617 & ~n5836 ;
  buffer buf_n5840( .i (n5839), .o (n5840) );
  buffer buf_n5841( .i (n5840), .o (n5841) );
  buffer buf_n5837( .i (n5836), .o (n5837) );
  buffer buf_n5838( .i (n5837), .o (n5838) );
  assign n5842 = n5838 | n5840 ;
  assign n5843 = ( ~n5800 & n5841 ) | ( ~n5800 & n5842 ) | ( n5841 & n5842 ) ;
  assign n5844 = n5825 | n5843 ;
  assign n5845 = ( ~n5823 & n5824 ) | ( ~n5823 & n5844 ) | ( n5824 & n5844 ) ;
  assign n5846 = n5443 & ~n5845 ;
  assign n5847 = ( n525 & n5435 ) | ( n525 & ~n5455 ) | ( n5435 & ~n5455 ) ;
  buffer buf_n5848( .i (n5847), .o (n5848) );
  buffer buf_n5849( .i (n5848), .o (n5849) );
  assign n5850 = ( n5457 & ~n5800 ) | ( n5457 & n5848 ) | ( ~n5800 & n5848 ) ;
  assign n5851 = ( ~n5427 & n5849 ) | ( ~n5427 & n5850 ) | ( n5849 & n5850 ) ;
  assign n5852 = n5598 | n5851 ;
  assign n5853 = ~n5443 & n5852 ;
  assign n5854 = n5846 | n5853 ;
  assign n5855 = ( n5673 & n5808 ) | ( n5673 & ~n5854 ) | ( n5808 & ~n5854 ) ;
  assign n5856 = n5809 | n5855 ;
  buffer buf_n5857( .i (n5494), .o (n5857) );
  assign n5858 = n5856 & ~n5857 ;
  assign n5859 = n267 | n5858 ;
  assign n5860 = ~n5769 & n5859 ;
  assign n5861 = n5692 | n5860 ;
  assign n5862 = ( n5610 & ~n5612 ) | ( n5610 & n5861 ) | ( ~n5612 & n5861 ) ;
  assign n5863 = n3922 & n5745 ;
  buffer buf_n5864( .i (n5863), .o (n5864) );
  buffer buf_n5865( .i (n5864), .o (n5865) );
  assign n5866 = ( ~n5473 & n5778 ) | ( ~n5473 & n5865 ) | ( n5778 & n5865 ) ;
  assign n5867 = ( n5754 & n5798 ) | ( n5754 & ~n5864 ) | ( n5798 & ~n5864 ) ;
  buffer buf_n5868( .i (n5472), .o (n5868) );
  assign n5869 = ( n4878 & n5867 ) | ( n4878 & ~n5868 ) | ( n5867 & ~n5868 ) ;
  assign n5870 = ~n5866 & n5869 ;
  buffer buf_n5871( .i (n5870), .o (n5871) );
  buffer buf_n5872( .i (n5871), .o (n5872) );
  buffer buf_n5873( .i (n5805), .o (n5873) );
  buffer buf_n5874( .i (n5683), .o (n5874) );
  assign n5875 = ( n5871 & n5873 ) | ( n5871 & n5874 ) | ( n5873 & n5874 ) ;
  buffer buf_n2465( .i (n2464), .o (n2465) );
  buffer buf_n2466( .i (n2465), .o (n2466) );
  buffer buf_n2467( .i (n2466), .o (n2467) );
  buffer buf_n2468( .i (n2467), .o (n2468) );
  assign n5876 = ( n729 & n2468 ) | ( n729 & n5651 ) | ( n2468 & n5651 ) ;
  buffer buf_n5877( .i (n5651), .o (n5877) );
  assign n5878 = n5876 & ~n5877 ;
  assign n5879 = ~n5874 & n5878 ;
  assign n5880 = ( n5872 & ~n5875 ) | ( n5872 & n5879 ) | ( ~n5875 & n5879 ) ;
  buffer buf_n5881( .i (n5880), .o (n5881) );
  buffer buf_n5882( .i (n5881), .o (n5882) );
  buffer buf_n5883( .i (n5882), .o (n5883) );
  assign n5884 = ( ~n119 & n600 ) | ( ~n119 & n5881 ) | ( n600 & n5881 ) ;
  assign n5885 = n759 & ~n5884 ;
  assign n5886 = ( n760 & n5883 ) | ( n760 & ~n5885 ) | ( n5883 & ~n5885 ) ;
  buffer buf_n5887( .i (n5886), .o (n5887) );
  buffer buf_n5888( .i (n5887), .o (n5888) );
  assign n5889 = n2712 & n5887 ;
  buffer buf_n521( .i (n520), .o (n521) );
  assign n5890 = ( ~n2144 & n2295 ) | ( ~n2144 & n5268 ) | ( n2295 & n5268 ) ;
  assign n5891 = ( ~n3929 & n4738 ) | ( ~n3929 & n5890 ) | ( n4738 & n5890 ) ;
  buffer buf_n5892( .i (n5891), .o (n5892) );
  buffer buf_n5893( .i (n5892), .o (n5893) );
  buffer buf_n5894( .i (n4739), .o (n5894) );
  assign n5895 = n5892 & ~n5894 ;
  buffer buf_n5896( .i (n3930), .o (n5896) );
  buffer buf_n5897( .i (n5896), .o (n5897) );
  assign n5898 = ( n5893 & n5895 ) | ( n5893 & n5897 ) | ( n5895 & n5897 ) ;
  buffer buf_n5899( .i (n5898), .o (n5899) );
  buffer buf_n5900( .i (n5899), .o (n5900) );
  assign n5901 = n4029 & ~n5899 ;
  assign n5902 = ( n1304 & n5900 ) | ( n1304 & ~n5901 ) | ( n5900 & ~n5901 ) ;
  buffer buf_n5903( .i (n5306), .o (n5903) );
  assign n5904 = ~n5902 & n5903 ;
  assign n5905 = ~n5403 & n5751 ;
  assign n5906 = n5903 | n5905 ;
  assign n5907 = ~n5904 & n5906 ;
  buffer buf_n5908( .i (n5502), .o (n5908) );
  assign n5909 = n5907 & ~n5908 ;
  buffer buf_n5910( .i (n2225), .o (n5910) );
  buffer buf_n5911( .i (n5910), .o (n5911) );
  buffer buf_n5912( .i (n247), .o (n5912) );
  assign n5913 = ( ~n2328 & n5911 ) | ( ~n2328 & n5912 ) | ( n5911 & n5912 ) ;
  buffer buf_n5914( .i (n5913), .o (n5914) );
  buffer buf_n5915( .i (n5914), .o (n5915) );
  buffer buf_n5916( .i (n5915), .o (n5916) );
  buffer buf_n5917( .i (n5916), .o (n5917) );
  buffer buf_n5919( .i (n5897), .o (n5919) );
  assign n5920 = ( n5057 & ~n5917 ) | ( n5057 & n5919 ) | ( ~n5917 & n5919 ) ;
  buffer buf_n5921( .i (n5150), .o (n5921) );
  assign n5922 = ( n5917 & n5919 ) | ( n5917 & ~n5921 ) | ( n5919 & ~n5921 ) ;
  assign n5923 = n5920 & ~n5922 ;
  assign n5924 = ( ~n5133 & n5793 ) | ( ~n5133 & n5923 ) | ( n5793 & n5923 ) ;
  assign n5925 = n343 & n5921 ;
  assign n5926 = ~n5524 & n5925 ;
  buffer buf_n5927( .i (n5132), .o (n5927) );
  assign n5928 = ( n5793 & n5926 ) | ( n5793 & n5927 ) | ( n5926 & n5927 ) ;
  assign n5929 = n5924 & n5928 ;
  assign n5930 = n3025 & ~n5927 ;
  assign n5931 = n441 & n5930 ;
  assign n5932 = n5929 | n5931 ;
  assign n5933 = n5908 & n5932 ;
  assign n5934 = n5909 | n5933 ;
  buffer buf_n5935( .i (n5934), .o (n5935) );
  buffer buf_n5936( .i (n5935), .o (n5936) );
  buffer buf_n5937( .i (n3735), .o (n5937) );
  assign n5938 = ( n2907 & ~n4577 ) | ( n2907 & n5937 ) | ( ~n4577 & n5937 ) ;
  buffer buf_n5939( .i (n5938), .o (n5939) );
  buffer buf_n5942( .i (n5937), .o (n5942) );
  buffer buf_n5943( .i (n5942), .o (n5943) );
  assign n5944 = ~n5939 & n5943 ;
  buffer buf_n5945( .i (n5944), .o (n5945) );
  buffer buf_n5946( .i (n5945), .o (n5946) );
  buffer buf_n5940( .i (n5939), .o (n5940) );
  buffer buf_n5941( .i (n5940), .o (n5941) );
  assign n5947 = n5941 | n5945 ;
  assign n5948 = ( ~n5617 & n5946 ) | ( ~n5617 & n5947 ) | ( n5946 & n5947 ) ;
  buffer buf_n5949( .i (n5948), .o (n5949) );
  buffer buf_n5950( .i (n5949), .o (n5950) );
  assign n5951 = ( n348 & n5553 ) | ( n348 & n5949 ) | ( n5553 & n5949 ) ;
  assign n5952 = n742 & ~n5745 ;
  assign n5953 = n2237 & n5952 ;
  assign n5954 = ~n348 & n5953 ;
  assign n5955 = ( n5950 & ~n5951 ) | ( n5950 & n5954 ) | ( ~n5951 & n5954 ) ;
  assign n5956 = n534 & ~n5750 ;
  assign n5957 = ~n329 & n4579 ;
  buffer buf_n5958( .i (n5957), .o (n5958) );
  assign n5969 = n5956 & n5958 ;
  buffer buf_n5970( .i (n5969), .o (n5970) );
  buffer buf_n5971( .i (n5970), .o (n5971) );
  buffer buf_n5972( .i (n5971), .o (n5972) );
  assign n5973 = ( ~n5502 & n5552 ) | ( ~n5502 & n5970 ) | ( n5552 & n5970 ) ;
  assign n5974 = n3028 & ~n5973 ;
  assign n5975 = ( n3029 & n5972 ) | ( n3029 & ~n5974 ) | ( n5972 & ~n5974 ) ;
  buffer buf_n5976( .i (n4878), .o (n5976) );
  assign n5977 = ( n5955 & n5975 ) | ( n5955 & ~n5976 ) | ( n5975 & ~n5976 ) ;
  assign n5978 = ~n5935 & n5977 ;
  assign n5979 = ( ~n5762 & n5936 ) | ( ~n5762 & n5978 ) | ( n5936 & n5978 ) ;
  buffer buf_n5980( .i (n5979), .o (n5980) );
  buffer buf_n5981( .i (n5980), .o (n5981) );
  buffer buf_n5982( .i (n5981), .o (n5982) );
  assign n5983 = ( n716 & n929 ) | ( n716 & n5980 ) | ( n929 & n5980 ) ;
  assign n5984 = n520 & ~n5983 ;
  assign n5985 = ( n521 & n5982 ) | ( n521 & ~n5984 ) | ( n5982 & ~n5984 ) ;
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n2102( .i (n2101), .o (n2102) );
  assign n5986 = ( n965 & ~n3929 ) | ( n965 & n5381 ) | ( ~n3929 & n5381 ) ;
  buffer buf_n5987( .i (n5986), .o (n5987) );
  assign n5990 = n5896 & n5987 ;
  buffer buf_n5991( .i (n5990), .o (n5991) );
  buffer buf_n5992( .i (n5991), .o (n5992) );
  buffer buf_n5988( .i (n5987), .o (n5988) );
  buffer buf_n5989( .i (n5988), .o (n5989) );
  assign n5993 = n5989 & ~n5991 ;
  assign n5994 = ( n5298 & ~n5992 ) | ( n5298 & n5993 ) | ( ~n5992 & n5993 ) ;
  assign n5995 = n4974 & ~n5994 ;
  buffer buf_n5996( .i (n5725), .o (n5996) );
  assign n5997 = n5995 & n5996 ;
  buffer buf_n5998( .i (n5997), .o (n5998) );
  buffer buf_n5999( .i (n5998), .o (n5999) );
  assign n6000 = n2835 | n5998 ;
  assign n6001 = ( ~n2357 & n5999 ) | ( ~n2357 & n6000 ) | ( n5999 & n6000 ) ;
  assign n6002 = ( n5804 & ~n5976 ) | ( n5804 & n6001 ) | ( ~n5976 & n6001 ) ;
  buffer buf_n6003( .i (n5382), .o (n6003) );
  buffer buf_n6004( .i (n6003), .o (n6004) );
  assign n6005 = ( ~n3932 & n5897 ) | ( ~n3932 & n6004 ) | ( n5897 & n6004 ) ;
  buffer buf_n6006( .i (n6005), .o (n6006) );
  buffer buf_n6007( .i (n6006), .o (n6007) );
  buffer buf_n6008( .i (n6007), .o (n6008) );
  buffer buf_n6009( .i (n6008), .o (n6009) );
  buffer buf_n6010( .i (n4978), .o (n6010) );
  buffer buf_n6011( .i (n6010), .o (n6011) );
  assign n6012 = ( ~n5524 & n6006 ) | ( ~n5524 & n6011 ) | ( n6006 & n6011 ) ;
  buffer buf_n6013( .i (n6012), .o (n6013) );
  buffer buf_n6014( .i (n6013), .o (n6014) );
  assign n6015 = n3936 | n6013 ;
  assign n6016 = ( ~n6009 & n6014 ) | ( ~n6009 & n6015 ) | ( n6014 & n6015 ) ;
  assign n6017 = n5798 | n6016 ;
  assign n6018 = n5800 | n6017 ;
  assign n6019 = ( n5804 & n5976 ) | ( n5804 & n6018 ) | ( n5976 & n6018 ) ;
  assign n6020 = n6002 & ~n6019 ;
  buffer buf_n6021( .i (n6020), .o (n6021) );
  buffer buf_n6022( .i (n6021), .o (n6022) );
  buffer buf_n6023( .i (n6022), .o (n6023) );
  assign n6024 = ( n377 & n5168 ) | ( n377 & n6021 ) | ( n5168 & n6021 ) ;
  assign n6025 = n2101 | n6024 ;
  assign n6026 = ( ~n2102 & n6023 ) | ( ~n2102 & n6025 ) | ( n6023 & n6025 ) ;
  buffer buf_n6027( .i (n6026), .o (n6027) );
  assign n6028 = ( n151 & n5985 ) | ( n151 & n6027 ) | ( n5985 & n6027 ) ;
  buffer buf_n6029( .i (n5524), .o (n6029) );
  assign n6030 = ( n5254 & ~n5613 ) | ( n5254 & n6029 ) | ( ~n5613 & n6029 ) ;
  buffer buf_n6031( .i (n6030), .o (n6031) );
  buffer buf_n6032( .i (n6031), .o (n6032) );
  buffer buf_n6033( .i (n6032), .o (n6033) );
  buffer buf_n5257( .i (n5256), .o (n5257) );
  buffer buf_n6034( .i (n5538), .o (n6034) );
  assign n6035 = ( n5330 & n6031 ) | ( n5330 & ~n6034 ) | ( n6031 & ~n6034 ) ;
  assign n6036 = ~n5257 & n6035 ;
  assign n6037 = ( ~n5336 & n6033 ) | ( ~n5336 & n6036 ) | ( n6033 & n6036 ) ;
  assign n6038 = n5804 | n6037 ;
  assign n6039 = n1241 & ~n5770 ;
  buffer buf_n6040( .i (n5553), .o (n6040) );
  buffer buf_n6041( .i (n6040), .o (n6041) );
  assign n6042 = ~n6039 & n6041 ;
  assign n6043 = n6038 & ~n6042 ;
  assign n6044 = ( n839 & n5538 ) | ( n839 & n5614 ) | ( n5538 & n5614 ) ;
  buffer buf_n6045( .i (n6044), .o (n6045) );
  buffer buf_n6046( .i (n5571), .o (n6046) );
  buffer buf_n6047( .i (n6034), .o (n6047) );
  assign n6048 = ( n6045 & n6046 ) | ( n6045 & ~n6047 ) | ( n6046 & ~n6047 ) ;
  buffer buf_n6049( .i (n5614), .o (n6049) );
  buffer buf_n6050( .i (n6049), .o (n6050) );
  assign n6051 = ( ~n6045 & n6046 ) | ( ~n6045 & n6050 ) | ( n6046 & n6050 ) ;
  assign n6052 = n6048 & ~n6051 ;
  buffer buf_n6053( .i (n6052), .o (n6053) );
  buffer buf_n6054( .i (n6053), .o (n6054) );
  buffer buf_n6055( .i (n5976), .o (n6055) );
  assign n6056 = ~n6053 & n6055 ;
  assign n6057 = ( n6043 & n6054 ) | ( n6043 & ~n6056 ) | ( n6054 & ~n6056 ) ;
  assign n6058 = n5128 | n6057 ;
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  assign n6059 = ~n637 & n2180 ;
  buffer buf_n6060( .i (n5057), .o (n6060) );
  assign n6061 = n5022 | n6060 ;
  buffer buf_n6062( .i (n6061), .o (n6062) );
  buffer buf_n6063( .i (n6062), .o (n6063) );
  buffer buf_n6064( .i (n6063), .o (n6064) );
  buffer buf_n6065( .i (n5745), .o (n6065) );
  assign n6066 = ( n4346 & ~n5552 ) | ( n4346 & n6065 ) | ( ~n5552 & n6065 ) ;
  buffer buf_n6067( .i (n5479), .o (n6067) );
  assign n6068 = ( ~n4346 & n6049 ) | ( ~n4346 & n6067 ) | ( n6049 & n6067 ) ;
  assign n6069 = ( ~n6064 & n6066 ) | ( ~n6064 & n6068 ) | ( n6066 & n6068 ) ;
  assign n6070 = ~n5437 & n6069 ;
  buffer buf_n6071( .i (n4577), .o (n6071) );
  buffer buf_n6072( .i (n6071), .o (n6072) );
  buffer buf_n6073( .i (n6072), .o (n6073) );
  assign n6074 = ( n2091 & n2253 ) | ( n2091 & ~n6073 ) | ( n2253 & ~n6073 ) ;
  buffer buf_n6075( .i (n6074), .o (n6075) );
  buffer buf_n6086( .i (n5793), .o (n6086) );
  buffer buf_n6087( .i (n5613), .o (n6087) );
  assign n6088 = ( ~n6075 & n6086 ) | ( ~n6075 & n6087 ) | ( n6086 & n6087 ) ;
  buffer buf_n6089( .i (n6088), .o (n6089) );
  buffer buf_n6090( .i (n6067), .o (n6090) );
  assign n6091 = ( ~n5798 & n6089 ) | ( ~n5798 & n6090 ) | ( n6089 & n6090 ) ;
  assign n6092 = ( n6050 & ~n6089 ) | ( n6050 & n6090 ) | ( ~n6089 & n6090 ) ;
  assign n6093 = n6091 & ~n6092 ;
  assign n6094 = n6070 | n6093 ;
  assign n6095 = ( n2181 & ~n6059 ) | ( n2181 & n6094 ) | ( ~n6059 & n6094 ) ;
  assign n6096 = ~n5762 & n6095 ;
  assign n6097 = n5128 & ~n6096 ;
  assign n6098 = n6058 & ~n6097 ;
  assign n6099 = n179 | n6098 ;
  assign n6100 = ( n2034 & n4893 ) | ( n2034 & n5613 ) | ( n4893 & n5613 ) ;
  buffer buf_n6101( .i (n6100), .o (n6101) );
  buffer buf_n6102( .i (n6101), .o (n6102) );
  buffer buf_n6103( .i (n6102), .o (n6103) );
  assign n6104 = ( n6049 & n6065 ) | ( n6049 & ~n6101 ) | ( n6065 & ~n6101 ) ;
  assign n6105 = ( ~n2037 & n6047 ) | ( ~n2037 & n6104 ) | ( n6047 & n6104 ) ;
  assign n6106 = ( n2038 & ~n6103 ) | ( n2038 & n6105 ) | ( ~n6103 & n6105 ) ;
  assign n6107 = n6041 & ~n6106 ;
  assign n6108 = n942 & n6047 ;
  assign n6109 = n941 | n5571 ;
  assign n6110 = ( n6047 & n6050 ) | ( n6047 & n6109 ) | ( n6050 & n6109 ) ;
  assign n6111 = ~n6108 & n6110 ;
  assign n6112 = n6041 | n6111 ;
  assign n6113 = ( ~n5805 & n6107 ) | ( ~n5805 & n6112 ) | ( n6107 & n6112 ) ;
  assign n6114 = n5874 & ~n6113 ;
  buffer buf_n6115( .i (n6046), .o (n6115) );
  assign n6116 = ~n349 & n6115 ;
  assign n6117 = ( ~n350 & n4904 ) | ( ~n350 & n6116 ) | ( n4904 & n6116 ) ;
  assign n6118 = ~n5805 & n6117 ;
  assign n6119 = n5874 | n6118 ;
  assign n6120 = ~n6114 & n6119 ;
  assign n6121 = ~n4927 & n6120 ;
  assign n6122 = n179 & ~n6121 ;
  assign n6123 = n6099 & ~n6122 ;
  assign n6124 = ( ~n151 & n6027 ) | ( ~n151 & n6123 ) | ( n6027 & n6123 ) ;
  assign n6125 = n6028 | n6124 ;
  assign n6126 = n5076 & n6073 ;
  buffer buf_n6127( .i (n6126), .o (n6127) );
  buffer buf_n6131( .i (n6011), .o (n6131) );
  buffer buf_n6132( .i (n6131), .o (n6132) );
  assign n6133 = ( n6087 & n6127 ) | ( n6087 & n6132 ) | ( n6127 & n6132 ) ;
  buffer buf_n6134( .i (n6133), .o (n6134) );
  assign n6135 = n5472 | n6134 ;
  buffer buf_n6136( .i (n5471), .o (n6136) );
  assign n6137 = n6134 & n6136 ;
  assign n6138 = n6135 & ~n6137 ;
  assign n6139 = n5662 | n6138 ;
  assign n6140 = n1824 & n6049 ;
  assign n6141 = ( n2498 & n6050 ) | ( n2498 & ~n6140 ) | ( n6050 & ~n6140 ) ;
  buffer buf_n6142( .i (n5908), .o (n6142) );
  assign n6143 = n6141 | n6142 ;
  assign n6144 = n5662 & n6143 ;
  assign n6145 = n6139 & ~n6144 ;
  assign n6146 = n5873 & ~n6145 ;
  assign n6147 = ( ~n2239 & n5868 ) | ( ~n2239 & n6142 ) | ( n5868 & n6142 ) ;
  assign n6148 = ( n2238 & n5908 ) | ( n2238 & ~n6046 ) | ( n5908 & ~n6046 ) ;
  assign n6149 = ( ~n5778 & n5868 ) | ( ~n5778 & n6148 ) | ( n5868 & n6148 ) ;
  assign n6150 = n6147 & ~n6149 ;
  assign n6151 = ~n4730 & n6150 ;
  assign n6152 = n5873 | n6151 ;
  assign n6153 = ~n6146 & n6152 ;
  assign n6154 = n5165 & n6153 ;
  buffer buf_n6155( .i (n5251), .o (n6155) );
  assign n6156 = ( n5921 & n6010 ) | ( n5921 & n6155 ) | ( n6010 & n6155 ) ;
  assign n6157 = ( n6060 & ~n6073 ) | ( n6060 & n6156 ) | ( ~n6073 & n6156 ) ;
  buffer buf_n6158( .i (n6157), .o (n6158) );
  assign n6161 = n6087 & ~n6158 ;
  buffer buf_n6162( .i (n6161), .o (n6162) );
  buffer buf_n6163( .i (n6162), .o (n6163) );
  buffer buf_n6159( .i (n6158), .o (n6159) );
  buffer buf_n6160( .i (n6159), .o (n6160) );
  assign n6164 = n6160 | n6162 ;
  buffer buf_n6165( .i (n6087), .o (n6165) );
  buffer buf_n6166( .i (n6165), .o (n6166) );
  buffer buf_n6167( .i (n6166), .o (n6167) );
  assign n6168 = ( n6163 & n6164 ) | ( n6163 & ~n6167 ) | ( n6164 & ~n6167 ) ;
  assign n6169 = n6041 & ~n6168 ;
  assign n6170 = n2521 & ~n5868 ;
  buffer buf_n6171( .i (n6040), .o (n6171) );
  assign n6172 = n6170 | n6171 ;
  assign n6173 = ~n6169 & n6172 ;
  buffer buf_n6174( .i (n5571), .o (n6174) );
  assign n6175 = n2520 & ~n6174 ;
  assign n6176 = n2005 & n6090 ;
  assign n6177 = n6175 & n6176 ;
  buffer buf_n6178( .i (n6177), .o (n6178) );
  buffer buf_n6179( .i (n6178), .o (n6179) );
  assign n6180 = n5683 & ~n6178 ;
  assign n6181 = ( n6173 & n6179 ) | ( n6173 & ~n6180 ) | ( n6179 & ~n6180 ) ;
  buffer buf_n6182( .i (n5996), .o (n6182) );
  buffer buf_n6183( .i (n6132), .o (n6183) );
  assign n6184 = ( ~n6165 & n6182 ) | ( ~n6165 & n6183 ) | ( n6182 & n6183 ) ;
  buffer buf_n6185( .i (n6184), .o (n6185) );
  buffer buf_n6186( .i (n6136), .o (n6186) );
  assign n6187 = ( n6115 & n6185 ) | ( n6115 & ~n6186 ) | ( n6185 & ~n6186 ) ;
  assign n6188 = ( n6115 & n6142 ) | ( n6115 & ~n6185 ) | ( n6142 & ~n6185 ) ;
  assign n6189 = n6187 & ~n6188 ;
  buffer buf_n6190( .i (n6171), .o (n6190) );
  assign n6191 = n6189 | n6190 ;
  buffer buf_n4117( .i (n4116), .o (n4117) );
  buffer buf_n4118( .i (n4117), .o (n4118) );
  buffer buf_n4119( .i (n4118), .o (n4119) );
  buffer buf_n4120( .i (n4119), .o (n4120) );
  assign n6192 = n4120 & n5757 ;
  assign n6193 = n6190 & ~n6192 ;
  assign n6194 = n6191 & ~n6193 ;
  assign n6195 = n6181 | n6194 ;
  buffer buf_n6196( .i (n5193), .o (n6196) );
  assign n6197 = n6195 & ~n6196 ;
  assign n6198 = n6154 | n6197 ;
  buffer buf_n6199( .i (n6198), .o (n6199) );
  buffer buf_n6200( .i (n6199), .o (n6200) );
  assign n6201 = n3020 & n6199 ;
  buffer buf_n6202( .i (n4731), .o (n6202) );
  assign n6203 = ( n1268 & n5491 ) | ( n1268 & n6202 ) | ( n5491 & n6202 ) ;
  buffer buf_n6204( .i (n6203), .o (n6204) );
  assign n6205 = ( n179 & ~n207 ) | ( n179 & n6204 ) | ( ~n207 & n6204 ) ;
  buffer buf_n6206( .i (n5296), .o (n6206) );
  buffer buf_n6207( .i (n6206), .o (n6207) );
  buffer buf_n6208( .i (n6202), .o (n6208) );
  buffer buf_n6209( .i (n6208), .o (n6209) );
  assign n6210 = ( ~n6204 & n6207 ) | ( ~n6204 & n6209 ) | ( n6207 & n6209 ) ;
  assign n6211 = n6205 & ~n6210 ;
  buffer buf_n2246( .i (n2245), .o (n2246) );
  assign n6212 = ( n5754 & ~n6090 ) | ( n5754 & n6136 ) | ( ~n6090 & n6136 ) ;
  buffer buf_n6213( .i (n6067), .o (n6213) );
  buffer buf_n6214( .i (n5753), .o (n6214) );
  assign n6215 = ( n6174 & ~n6213 ) | ( n6174 & n6214 ) | ( ~n6213 & n6214 ) ;
  assign n6216 = n6212 & ~n6215 ;
  buffer buf_n6217( .i (n5770), .o (n6217) );
  assign n6218 = n6216 & n6217 ;
  buffer buf_n6219( .i (n6142), .o (n6219) );
  buffer buf_n6220( .i (n6219), .o (n6220) );
  assign n6221 = ( n6055 & n6218 ) | ( n6055 & n6220 ) | ( n6218 & n6220 ) ;
  assign n6222 = ~n5762 & n6221 ;
  buffer buf_n6223( .i (n6222), .o (n6223) );
  buffer buf_n6224( .i (n6223), .o (n6224) );
  buffer buf_n6225( .i (n6224), .o (n6225) );
  assign n6226 = ( ~n694 & n1405 ) | ( ~n694 & n6223 ) | ( n1405 & n6223 ) ;
  assign n6227 = n2245 & ~n6226 ;
  assign n6228 = ( n2246 & n6225 ) | ( n2246 & ~n6227 ) | ( n6225 & ~n6227 ) ;
  assign n6229 = n6211 | n6228 ;
  assign n6230 = ( n6200 & ~n6201 ) | ( n6200 & n6229 ) | ( ~n6201 & n6229 ) ;
  assign n6231 = n6125 | n6230 ;
  assign n6232 = ( n5888 & ~n5889 ) | ( n5888 & n6231 ) | ( ~n5889 & n6231 ) ;
  buffer buf_n733( .i (n732), .o (n733) );
  assign n6233 = ( n5651 & n5662 ) | ( n5651 & n6217 ) | ( n5662 & n6217 ) ;
  buffer buf_n6234( .i (n6233), .o (n6234) );
  buffer buf_n6235( .i (n6234), .o (n6235) );
  assign n6236 = ~n5443 & n6234 ;
  assign n6237 = ( ~n4001 & n6235 ) | ( ~n4001 & n6236 ) | ( n6235 & n6236 ) ;
  assign n6238 = n733 & n6237 ;
  buffer buf_n6239( .i (n6238), .o (n6239) );
  buffer buf_n6240( .i (n6239), .o (n6240) );
  assign n6241 = ( n4739 & n5178 ) | ( n4739 & ~n5382 ) | ( n5178 & ~n5382 ) ;
  buffer buf_n6242( .i (n6241), .o (n6242) );
  buffer buf_n6243( .i (n6242), .o (n6243) );
  buffer buf_n6244( .i (n6243), .o (n6244) );
  buffer buf_n6245( .i (n6244), .o (n6245) );
  buffer buf_n6246( .i (n6245), .o (n6246) );
  buffer buf_n6247( .i (n6246), .o (n6247) );
  buffer buf_n6248( .i (n6247), .o (n6248) );
  buffer buf_n6249( .i (n6248), .o (n6249) );
  buffer buf_n6250( .i (n6249), .o (n6250) );
  buffer buf_n6251( .i (n6250), .o (n6251) );
  assign n6255 = ( n6055 & ~n6190 ) | ( n6055 & n6251 ) | ( ~n6190 & n6251 ) ;
  buffer buf_n6256( .i (n6255), .o (n6256) );
  buffer buf_n6257( .i (n6256), .o (n6257) );
  buffer buf_n6258( .i (n6257), .o (n6258) );
  buffer buf_n6252( .i (n6251), .o (n6252) );
  buffer buf_n6253( .i (n6252), .o (n6253) );
  buffer buf_n6254( .i (n6253), .o (n6254) );
  buffer buf_n6259( .i (n5192), .o (n6259) );
  assign n6260 = ( n5672 & n6256 ) | ( n5672 & ~n6259 ) | ( n6256 & ~n6259 ) ;
  assign n6261 = ~n6254 & n6260 ;
  buffer buf_n6262( .i (n6055), .o (n6262) );
  buffer buf_n6263( .i (n6262), .o (n6263) );
  buffer buf_n6264( .i (n6263), .o (n6264) );
  buffer buf_n6265( .i (n6264), .o (n6265) );
  assign n6266 = ( n6258 & n6261 ) | ( n6258 & ~n6265 ) | ( n6261 & ~n6265 ) ;
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n3166( .i (n3165), .o (n3166) );
  buffer buf_n3167( .i (n3166), .o (n3167) );
  buffer buf_n3168( .i (n3167), .o (n3168) );
  buffer buf_n3169( .i (n3168), .o (n3169) );
  buffer buf_n3170( .i (n3169), .o (n3170) );
  assign n6267 = n3170 & ~n6263 ;
  assign n6268 = n544 & n6267 ;
  buffer buf_n6269( .i (n6268), .o (n6269) );
  assign n6270 = ( ~n6239 & n6266 ) | ( ~n6239 & n6269 ) | ( n6266 & n6269 ) ;
  assign n6271 = n5606 & ~n6269 ;
  assign n6272 = ( n6240 & n6270 ) | ( n6240 & ~n6271 ) | ( n6270 & ~n6271 ) ;
  buffer buf_n6273( .i (n6272), .o (n6273) );
  buffer buf_n6274( .i (n6273), .o (n6274) );
  buffer buf_n4601( .i (n4600), .o (n4601) );
  buffer buf_n4602( .i (n4601), .o (n4602) );
  buffer buf_n4603( .i (n4602), .o (n4603) );
  buffer buf_n4604( .i (n4603), .o (n4604) );
  buffer buf_n4605( .i (n4604), .o (n4605) );
  buffer buf_n4606( .i (n4605), .o (n4606) );
  buffer buf_n4607( .i (n4606), .o (n4607) );
  buffer buf_n4608( .i (n4607), .o (n4608) );
  buffer buf_n4609( .i (n4608), .o (n4609) );
  buffer buf_n4610( .i (n4609), .o (n4610) );
  buffer buf_n4611( .i (n4610), .o (n4611) );
  buffer buf_n4612( .i (n4611), .o (n4612) );
  assign n6275 = n4612 & n6273 ;
  buffer buf_n6276( .i (n5919), .o (n6276) );
  assign n6277 = n740 & ~n6276 ;
  assign n6278 = ( n6029 & n6131 ) | ( n6029 & n6277 ) | ( n6131 & n6277 ) ;
  assign n6279 = ~n6132 & n6278 ;
  buffer buf_n6280( .i (n6279), .o (n6280) );
  buffer buf_n6281( .i (n6280), .o (n6281) );
  buffer buf_n6282( .i (n6281), .o (n6282) );
  assign n6283 = ( ~n311 & n2037 ) | ( ~n311 & n6280 ) | ( n2037 & n6280 ) ;
  assign n6284 = n6186 & ~n6283 ;
  buffer buf_n6285( .i (n6186), .o (n6285) );
  assign n6286 = ( n6282 & ~n6284 ) | ( n6282 & n6285 ) | ( ~n6284 & n6285 ) ;
  assign n6287 = n4790 & ~n6286 ;
  buffer buf_n3134( .i (n3133), .o (n3134) );
  buffer buf_n6288( .i (n6034), .o (n6288) );
  assign n6289 = ( n3134 & n6136 ) | ( n3134 & ~n6288 ) | ( n6136 & ~n6288 ) ;
  buffer buf_n6290( .i (n6182), .o (n6290) );
  assign n6291 = ( n3134 & ~n6288 ) | ( n3134 & n6290 ) | ( ~n6288 & n6290 ) ;
  assign n6292 = ( n2006 & n6289 ) | ( n2006 & ~n6291 ) | ( n6289 & ~n6291 ) ;
  buffer buf_n6293( .i (n6115), .o (n6293) );
  assign n6294 = n6292 & n6293 ;
  buffer buf_n6295( .i (n6217), .o (n6295) );
  assign n6296 = n6294 | n6295 ;
  assign n6297 = ~n6287 & n6296 ;
  buffer buf_n6298( .i (n6297), .o (n6298) );
  buffer buf_n6299( .i (n6298), .o (n6299) );
  assign n6300 = n6208 & n6298 ;
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  assign n6301 = ~n590 & n612 ;
  assign n6302 = ( ~n1723 & n5873 ) | ( ~n1723 & n6301 ) | ( n5873 & n6301 ) ;
  assign n6303 = ~n5672 & n6302 ;
  buffer buf_n5379( .i (n5378), .o (n5379) );
  buffer buf_n5380( .i (n5379), .o (n5380) );
  assign n6304 = ( n439 & n6073 ) | ( n439 & n6276 ) | ( n6073 & n6276 ) ;
  assign n6305 = n5380 & ~n6304 ;
  buffer buf_n6306( .i (n5927), .o (n6306) );
  assign n6307 = n6305 & n6306 ;
  buffer buf_n6308( .i (n6072), .o (n6308) );
  assign n6309 = ( ~n5750 & n5811 ) | ( ~n5750 & n6308 ) | ( n5811 & n6308 ) ;
  assign n6310 = ( ~n5750 & n5811 ) | ( ~n5750 & n6276 ) | ( n5811 & n6276 ) ;
  assign n6311 = ( n2034 & n6309 ) | ( n2034 & ~n6310 ) | ( n6309 & ~n6310 ) ;
  assign n6312 = n6306 | n6311 ;
  assign n6313 = ( ~n6067 & n6307 ) | ( ~n6067 & n6312 ) | ( n6307 & n6312 ) ;
  assign n6314 = n6166 & ~n6313 ;
  assign n6315 = ( n2116 & n5229 ) | ( n2116 & ~n5788 ) | ( n5229 & ~n5788 ) ;
  buffer buf_n6316( .i (n6315), .o (n6316) );
  buffer buf_n6317( .i (n6316), .o (n6317) );
  assign n6318 = ( n5231 & n6029 ) | ( n5231 & ~n6316 ) | ( n6029 & ~n6316 ) ;
  assign n6319 = ( n6086 & n6317 ) | ( n6086 & ~n6318 ) | ( n6317 & ~n6318 ) ;
  assign n6320 = n5753 & n6319 ;
  assign n6321 = n6166 | n6320 ;
  assign n6322 = ~n6314 & n6321 ;
  assign n6323 = n6219 & n6322 ;
  assign n6324 = ( n2173 & n5181 ) | ( n2173 & n5788 ) | ( n5181 & n5788 ) ;
  buffer buf_n6325( .i (n5788), .o (n6325) );
  assign n6326 = n6324 & ~n6325 ;
  buffer buf_n6327( .i (n6326), .o (n6327) );
  buffer buf_n6328( .i (n6327), .o (n6328) );
  buffer buf_n6329( .i (n6328), .o (n6329) );
  assign n6330 = ( n3058 & n5179 ) | ( n3058 & n5896 ) | ( n5179 & n5896 ) ;
  buffer buf_n6331( .i (n6330), .o (n6331) );
  buffer buf_n6332( .i (n6331), .o (n6332) );
  buffer buf_n6333( .i (n6332), .o (n6333) );
  assign n6334 = ( n5919 & n6072 ) | ( n5919 & ~n6331 ) | ( n6072 & ~n6331 ) ;
  buffer buf_n6335( .i (n5921), .o (n6335) );
  assign n6336 = n6334 & n6335 ;
  assign n6337 = ( n5927 & ~n6333 ) | ( n5927 & n6336 ) | ( ~n6333 & n6336 ) ;
  assign n6338 = ( n6086 & n6327 ) | ( n6086 & n6337 ) | ( n6327 & n6337 ) ;
  assign n6339 = n6165 & ~n6338 ;
  assign n6340 = ( n6166 & n6329 ) | ( n6166 & ~n6339 ) | ( n6329 & ~n6339 ) ;
  buffer buf_n6341( .i (n5178), .o (n6341) );
  assign n6342 = ( n4766 & ~n5894 ) | ( n4766 & n6341 ) | ( ~n5894 & n6341 ) ;
  assign n6343 = ( n5399 & ~n5897 ) | ( n5399 & n6342 ) | ( ~n5897 & n6342 ) ;
  buffer buf_n6344( .i (n6343), .o (n6344) );
  assign n6347 = n5132 & ~n6344 ;
  buffer buf_n6348( .i (n6347), .o (n6348) );
  buffer buf_n6349( .i (n6348), .o (n6349) );
  buffer buf_n6345( .i (n6344), .o (n6345) );
  buffer buf_n6346( .i (n6345), .o (n6346) );
  assign n6350 = n6346 | n6348 ;
  buffer buf_n6351( .i (n6306), .o (n6351) );
  assign n6352 = ( n6349 & n6350 ) | ( n6349 & ~n6351 ) | ( n6350 & ~n6351 ) ;
  assign n6353 = ( n6174 & n6214 ) | ( n6174 & n6352 ) | ( n6214 & n6352 ) ;
  assign n6354 = ( ~n2239 & n6340 ) | ( ~n2239 & n6353 ) | ( n6340 & n6353 ) ;
  assign n6355 = n6219 | n6354 ;
  assign n6356 = ( ~n6220 & n6323 ) | ( ~n6220 & n6355 ) | ( n6323 & n6355 ) ;
  buffer buf_n6357( .i (n5877), .o (n6357) );
  assign n6358 = n6356 & n6357 ;
  assign n6359 = ( n5942 & ~n6004 ) | ( n5942 & n6242 ) | ( ~n6004 & n6242 ) ;
  buffer buf_n6360( .i (n6359), .o (n6360) );
  assign n6363 = n6335 & n6360 ;
  buffer buf_n6364( .i (n6363), .o (n6364) );
  buffer buf_n6365( .i (n6364), .o (n6365) );
  buffer buf_n6361( .i (n6360), .o (n6361) );
  buffer buf_n6362( .i (n6361), .o (n6362) );
  assign n6366 = n6362 & ~n6364 ;
  assign n6367 = ( n5753 & ~n6365 ) | ( n5753 & n6366 ) | ( ~n6365 & n6366 ) ;
  buffer buf_n6368( .i (n6367), .o (n6368) );
  buffer buf_n6369( .i (n6368), .o (n6369) );
  assign n6370 = n2179 & ~n6368 ;
  assign n6371 = ( n2137 & ~n6369 ) | ( n2137 & n6370 ) | ( ~n6369 & n6370 ) ;
  buffer buf_n6372( .i (n47), .o (n6372) );
  assign n6373 = ( n4765 & ~n5914 ) | ( n4765 & n6372 ) | ( ~n5914 & n6372 ) ;
  buffer buf_n6374( .i (n6373), .o (n6374) );
  buffer buf_n6375( .i (n6374), .o (n6375) );
  buffer buf_n6376( .i (n6375), .o (n6376) );
  buffer buf_n6377( .i (n6376), .o (n6377) );
  assign n6378 = ( ~n6004 & n6071 ) | ( ~n6004 & n6374 ) | ( n6071 & n6374 ) ;
  buffer buf_n6379( .i (n6378), .o (n6379) );
  buffer buf_n6380( .i (n6379), .o (n6380) );
  buffer buf_n5918( .i (n5917), .o (n5918) );
  assign n6381 = n5918 & n6379 ;
  assign n6382 = ( ~n6377 & n6380 ) | ( ~n6377 & n6381 ) | ( n6380 & n6381 ) ;
  buffer buf_n6383( .i (n6341), .o (n6383) );
  assign n6384 = n2172 & ~n6383 ;
  buffer buf_n6385( .i (n6004), .o (n6385) );
  assign n6386 = n6384 & ~n6385 ;
  buffer buf_n6387( .i (n6386), .o (n6387) );
  buffer buf_n6388( .i (n6387), .o (n6388) );
  assign n6389 = n5743 & ~n6387 ;
  assign n6390 = ( n6382 & n6388 ) | ( n6382 & ~n6389 ) | ( n6388 & ~n6389 ) ;
  assign n6391 = n6065 & ~n6390 ;
  assign n6392 = n2058 & n6306 ;
  assign n6393 = n6065 | n6392 ;
  assign n6394 = ~n6391 & n6393 ;
  buffer buf_n6395( .i (n6290), .o (n6395) );
  assign n6396 = n6394 & ~n6395 ;
  buffer buf_n6397( .i (n6060), .o (n6397) );
  buffer buf_n6398( .i (n6397), .o (n6398) );
  assign n6399 = ( n633 & ~n2833 ) | ( n633 & n6398 ) | ( ~n2833 & n6398 ) ;
  buffer buf_n6400( .i (n5896), .o (n6400) );
  buffer buf_n6401( .i (n6400), .o (n6401) );
  assign n6402 = ( n1103 & ~n6072 ) | ( n1103 & n6401 ) | ( ~n6072 & n6401 ) ;
  buffer buf_n6403( .i (n5894), .o (n6403) );
  buffer buf_n6404( .i (n6403), .o (n6404) );
  buffer buf_n6405( .i (n6071), .o (n6405) );
  assign n6406 = ( n1103 & ~n6404 ) | ( n1103 & n6405 ) | ( ~n6404 & n6405 ) ;
  assign n6407 = n6402 | n6406 ;
  buffer buf_n6408( .i (n5132), .o (n6408) );
  assign n6409 = ~n6407 & n6408 ;
  assign n6410 = n6398 & n6409 ;
  assign n6411 = ( n2834 & n6399 ) | ( n2834 & n6410 ) | ( n6399 & n6410 ) ;
  buffer buf_n6412( .i (n6408), .o (n6412) );
  assign n6413 = n2176 & n6412 ;
  assign n6414 = n442 & n6413 ;
  assign n6415 = n6411 | n6414 ;
  assign n6416 = n6395 & n6415 ;
  assign n6417 = n6396 | n6416 ;
  assign n6418 = n6371 | n6417 ;
  assign n6419 = ~n6357 & n6418 ;
  assign n6420 = n6358 | n6419 ;
  assign n6421 = n6303 | n6420 ;
  assign n6422 = ( n6299 & ~n6300 ) | ( n6299 & n6421 ) | ( ~n6300 & n6421 ) ;
  buffer buf_n6423( .i (n6422), .o (n6423) );
  buffer buf_n6424( .i (n6423), .o (n6424) );
  assign n6425 = n3020 & n6423 ;
  assign n6426 = n4744 & ~n5453 ;
  assign n6427 = n3815 & n6426 ;
  buffer buf_n6428( .i (n6427), .o (n6428) );
  buffer buf_n6429( .i (n6428), .o (n6429) );
  buffer buf_n6430( .i (n6429), .o (n6430) );
  buffer buf_n3906( .i (n3905), .o (n3906) );
  buffer buf_n3907( .i (n3906), .o (n3907) );
  buffer buf_n3908( .i (n3907), .o (n3908) );
  buffer buf_n3909( .i (n3908), .o (n3909) );
  assign n6431 = n585 & n6132 ;
  assign n6432 = ( n3909 & n4008 ) | ( n3909 & ~n6431 ) | ( n4008 & ~n6431 ) ;
  buffer buf_n6433( .i (n6165), .o (n6433) );
  assign n6434 = ( n6428 & n6432 ) | ( n6428 & ~n6433 ) | ( n6432 & ~n6433 ) ;
  buffer buf_n6435( .i (n6288), .o (n6435) );
  assign n6436 = ~n6434 & n6435 ;
  buffer buf_n6437( .i (n6435), .o (n6437) );
  assign n6438 = ( n6430 & ~n6436 ) | ( n6430 & n6437 ) | ( ~n6436 & n6437 ) ;
  buffer buf_n6439( .i (n5778), .o (n6439) );
  buffer buf_n6440( .i (n6439), .o (n6440) );
  assign n6441 = n6438 & n6440 ;
  buffer buf_n6442( .i (n6441), .o (n6442) );
  buffer buf_n6443( .i (n6442), .o (n6443) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  assign n6444 = ( n2469 & n5640 ) | ( n2469 & n5877 ) | ( n5640 & n5877 ) ;
  assign n6445 = ~n6357 & n6444 ;
  assign n6446 = n6442 | n6445 ;
  assign n6447 = ( ~n6264 & n6443 ) | ( ~n6264 & n6446 ) | ( n6443 & n6446 ) ;
  buffer buf_n6448( .i (n5672), .o (n6448) );
  buffer buf_n6449( .i (n6448), .o (n6449) );
  assign n6450 = n6447 | n6449 ;
  assign n6451 = ( n1367 & n6217 ) | ( n1367 & n6285 ) | ( n6217 & n6285 ) ;
  assign n6452 = ( n1367 & ~n6219 ) | ( n1367 & n6285 ) | ( ~n6219 & n6285 ) ;
  buffer buf_n6453( .i (n589), .o (n6453) );
  assign n6454 = ( ~n6451 & n6452 ) | ( ~n6451 & n6453 ) | ( n6452 & n6453 ) ;
  buffer buf_n2933( .i (n2932), .o (n2933) );
  buffer buf_n6455( .i (n6398), .o (n6455) );
  assign n6456 = n371 & ~n6455 ;
  buffer buf_n6457( .i (n6456), .o (n6457) );
  assign n6461 = n2933 & n6457 ;
  buffer buf_n6462( .i (n6461), .o (n6462) );
  buffer buf_n6463( .i (n6462), .o (n6463) );
  assign n6464 = n6440 & ~n6462 ;
  assign n6465 = ( n6454 & ~n6463 ) | ( n6454 & n6464 ) | ( ~n6463 & n6464 ) ;
  assign n6466 = n406 & n1309 ;
  buffer buf_n6467( .i (n6466), .o (n6467) );
  buffer buf_n6468( .i (n6467), .o (n6468) );
  assign n6469 = n5701 | n6467 ;
  assign n6470 = ( ~n6465 & n6468 ) | ( ~n6465 & n6469 ) | ( n6468 & n6469 ) ;
  assign n6471 = ~n6264 & n6470 ;
  assign n6472 = n6449 & ~n6471 ;
  assign n6473 = n6450 & ~n6472 ;
  assign n6474 = n3037 | n6473 ;
  assign n6475 = ( n6424 & ~n6425 ) | ( n6424 & n6474 ) | ( ~n6425 & n6474 ) ;
  buffer buf_n6458( .i (n6457), .o (n6458) );
  buffer buf_n6459( .i (n6458), .o (n6459) );
  buffer buf_n6460( .i (n6459), .o (n6460) );
  assign n6476 = ( ~n5192 & n6262 ) | ( ~n5192 & n6460 ) | ( n6262 & n6460 ) ;
  buffer buf_n2371( .i (n2370), .o (n2371) );
  buffer buf_n6477( .i (n6131), .o (n6477) );
  assign n6478 = ( n2371 & ~n6398 ) | ( n2371 & n6477 ) | ( ~n6398 & n6477 ) ;
  buffer buf_n6479( .i (n6478), .o (n6479) );
  buffer buf_n6482( .i (n6183), .o (n6482) );
  assign n6483 = ~n6479 & n6482 ;
  buffer buf_n6484( .i (n6483), .o (n6484) );
  buffer buf_n6485( .i (n6484), .o (n6485) );
  buffer buf_n6480( .i (n6479), .o (n6480) );
  buffer buf_n6481( .i (n6480), .o (n6481) );
  assign n6486 = n6481 | n6484 ;
  assign n6487 = ( ~n5877 & n6485 ) | ( ~n5877 & n6486 ) | ( n6485 & n6486 ) ;
  buffer buf_n6488( .i (n6295), .o (n6488) );
  assign n6489 = ( n6262 & ~n6487 ) | ( n6262 & n6488 ) | ( ~n6487 & n6488 ) ;
  assign n6490 = n6476 & ~n6489 ;
  buffer buf_n6491( .i (n6490), .o (n6491) );
  buffer buf_n6492( .i (n6491), .o (n6492) );
  buffer buf_n6493( .i (n6440), .o (n6493) );
  assign n6494 = n2614 & n6493 ;
  assign n6495 = ( n1062 & n6263 ) | ( n1062 & n6494 ) | ( n6263 & n6494 ) ;
  assign n6496 = ~n6264 & n6495 ;
  buffer buf_n6497( .i (n6214), .o (n6497) );
  assign n6498 = n4515 & ~n6497 ;
  assign n6499 = ( n4516 & ~n5217 ) | ( n4516 & n6498 ) | ( ~n5217 & n6498 ) ;
  buffer buf_n6500( .i (n6499), .o (n6500) );
  buffer buf_n6501( .i (n6500), .o (n6501) );
  buffer buf_n6502( .i (n6190), .o (n6502) );
  assign n6503 = ( n4013 & n6500 ) | ( n4013 & n6502 ) | ( n6500 & n6502 ) ;
  assign n6504 = ~n6501 & n6503 ;
  buffer buf_n6505( .i (n6504), .o (n6505) );
  assign n6506 = ( ~n6491 & n6496 ) | ( ~n6491 & n6505 ) | ( n6496 & n6505 ) ;
  assign n6507 = n6449 & ~n6505 ;
  assign n6508 = ( n6492 & n6506 ) | ( n6492 & ~n6507 ) | ( n6506 & ~n6507 ) ;
  assign n6509 = n93 | n6508 ;
  buffer buf_n3279( .i (n3278), .o (n3279) );
  buffer buf_n3280( .i (n3279), .o (n3280) );
  buffer buf_n3281( .i (n3280), .o (n3281) );
  buffer buf_n3282( .i (n3281), .o (n3282) );
  buffer buf_n3283( .i (n3282), .o (n3283) );
  buffer buf_n3284( .i (n3283), .o (n3284) );
  buffer buf_n3285( .i (n3284), .o (n3285) );
  buffer buf_n3286( .i (n3285), .o (n3286) );
  buffer buf_n3287( .i (n3286), .o (n3287) );
  buffer buf_n6510( .i (n6397), .o (n6510) );
  assign n6511 = ( n5752 & n6086 ) | ( n5752 & ~n6510 ) | ( n6086 & ~n6510 ) ;
  buffer buf_n6512( .i (n6511), .o (n6512) );
  buffer buf_n6517( .i (n6325), .o (n6517) );
  buffer buf_n6518( .i (n6517), .o (n6518) );
  buffer buf_n6519( .i (n6518), .o (n6519) );
  buffer buf_n6520( .i (n6519), .o (n6520) );
  assign n6521 = ( n6174 & n6512 ) | ( n6174 & ~n6520 ) | ( n6512 & ~n6520 ) ;
  buffer buf_n6522( .i (n5903), .o (n6522) );
  buffer buf_n6523( .i (n6522), .o (n6523) );
  assign n6524 = ( n6214 & ~n6512 ) | ( n6214 & n6523 ) | ( ~n6512 & n6523 ) ;
  assign n6525 = n6521 & ~n6524 ;
  assign n6526 = ( n6171 & ~n6285 ) | ( n6171 & n6525 ) | ( ~n6285 & n6525 ) ;
  assign n6527 = ( n5752 & n6510 ) | ( n5752 & n6518 ) | ( n6510 & n6518 ) ;
  buffer buf_n6528( .i (n6527), .o (n6528) );
  assign n6529 = ( n6520 & n6523 ) | ( n6520 & ~n6528 ) | ( n6523 & ~n6528 ) ;
  buffer buf_n6530( .i (n5752), .o (n6530) );
  buffer buf_n6531( .i (n6530), .o (n6531) );
  assign n6532 = ( n6523 & n6528 ) | ( n6523 & ~n6531 ) | ( n6528 & ~n6531 ) ;
  assign n6533 = ~n6529 & n6532 ;
  buffer buf_n6534( .i (n6186), .o (n6534) );
  assign n6535 = ( n6171 & ~n6533 ) | ( n6171 & n6534 ) | ( ~n6533 & n6534 ) ;
  assign n6536 = n6526 & ~n6535 ;
  buffer buf_n6537( .i (n6536), .o (n6537) );
  buffer buf_n6538( .i (n6537), .o (n6538) );
  buffer buf_n6539( .i (n6538), .o (n6539) );
  buffer buf_n6540( .i (n6502), .o (n6540) );
  assign n6541 = ( n5496 & n6537 ) | ( n5496 & ~n6540 ) | ( n6537 & ~n6540 ) ;
  assign n6542 = n3286 | n6541 ;
  assign n6543 = ( ~n3287 & n6539 ) | ( ~n3287 & n6542 ) | ( n6539 & n6542 ) ;
  assign n6544 = ~n5857 & n6543 ;
  assign n6545 = n93 & ~n6544 ;
  assign n6546 = n6509 & ~n6545 ;
  assign n6547 = n6475 | n6546 ;
  assign n6548 = ( n6274 & ~n6275 ) | ( n6274 & n6547 ) | ( ~n6275 & n6547 ) ;
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  assign n6549 = ( n4683 & ~n6060 ) | ( n4683 & n6335 ) | ( ~n6060 & n6335 ) ;
  buffer buf_n6550( .i (n6549), .o (n6550) );
  buffer buf_n6551( .i (n6550), .o (n6551) );
  buffer buf_n6552( .i (n6551), .o (n6552) );
  buffer buf_n6553( .i (n6552), .o (n6553) );
  assign n6554 = ( n6412 & n6477 ) | ( n6412 & n6550 ) | ( n6477 & n6550 ) ;
  buffer buf_n6555( .i (n6554), .o (n6555) );
  buffer buf_n6556( .i (n6555), .o (n6556) );
  assign n6557 = ~n4687 & n6555 ;
  assign n6558 = ( ~n6553 & n6556 ) | ( ~n6553 & n6557 ) | ( n6556 & n6557 ) ;
  buffer buf_n6559( .i (n6520), .o (n6559) );
  buffer buf_n6560( .i (n6559), .o (n6560) );
  assign n6561 = ~n6558 & n6560 ;
  buffer buf_n4500( .i (n4499), .o (n4500) );
  buffer buf_n4501( .i (n4500), .o (n4501) );
  buffer buf_n4502( .i (n4501), .o (n4502) );
  buffer buf_n4503( .i (n4502), .o (n4503) );
  buffer buf_n4504( .i (n4503), .o (n4504) );
  assign n6562 = n4504 & ~n6040 ;
  assign n6563 = n6560 | n6562 ;
  assign n6564 = ~n6561 & n6563 ;
  buffer buf_n6565( .i (n6220), .o (n6565) );
  assign n6566 = ( ~n6262 & n6564 ) | ( ~n6262 & n6565 ) | ( n6564 & n6565 ) ;
  assign n6567 = ~n4722 & n6518 ;
  buffer buf_n6568( .i (n6567), .o (n6568) );
  assign n6569 = ~n6531 & n6568 ;
  assign n6570 = ( ~n4724 & n6433 ) | ( ~n4724 & n6568 ) | ( n6433 & n6568 ) ;
  assign n6571 = ( n6040 & n6569 ) | ( n6040 & n6570 ) | ( n6569 & n6570 ) ;
  assign n6572 = n6534 | n6571 ;
  assign n6573 = n4127 | n6510 ;
  buffer buf_n6574( .i (n6573), .o (n6574) );
  buffer buf_n6575( .i (n6574), .o (n6575) );
  buffer buf_n6576( .i (n6213), .o (n6576) );
  assign n6577 = ~n6575 & n6576 ;
  assign n6578 = n6534 & ~n6577 ;
  assign n6579 = n6572 & ~n6578 ;
  buffer buf_n6580( .i (n4877), .o (n6580) );
  buffer buf_n6581( .i (n6580), .o (n6581) );
  buffer buf_n6582( .i (n6581), .o (n6582) );
  buffer buf_n6583( .i (n6582), .o (n6583) );
  assign n6584 = ( n6565 & ~n6579 ) | ( n6565 & n6583 ) | ( ~n6579 & n6583 ) ;
  assign n6585 = n6566 & ~n6584 ;
  assign n6586 = ( ~n1403 & n1786 ) | ( ~n1403 & n6493 ) | ( n1786 & n6493 ) ;
  buffer buf_n6587( .i (n1403), .o (n6587) );
  assign n6588 = n6586 & n6587 ;
  assign n6589 = n6585 | n6588 ;
  buffer buf_n6590( .i (n6589), .o (n6590) );
  buffer buf_n6591( .i (n6590), .o (n6591) );
  assign n6592 = ( ~n208 & n238 ) | ( ~n208 & n6590 ) | ( n238 & n6590 ) ;
  assign n6593 = ( n2046 & n6591 ) | ( n2046 & ~n6592 ) | ( n6591 & ~n6592 ) ;
  buffer buf_n6594( .i (n6593), .o (n6594) );
  buffer buf_n6595( .i (n6594), .o (n6595) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n6596( .i (n6155), .o (n6596) );
  assign n6597 = ( n1121 & ~n6308 ) | ( n1121 & n6596 ) | ( ~n6308 & n6596 ) ;
  buffer buf_n6598( .i (n6597), .o (n6598) );
  assign n6601 = n6510 & ~n6598 ;
  buffer buf_n6602( .i (n6601), .o (n6602) );
  buffer buf_n6603( .i (n6602), .o (n6603) );
  buffer buf_n6599( .i (n6598), .o (n6599) );
  buffer buf_n6600( .i (n6599), .o (n6600) );
  assign n6604 = n6600 | n6602 ;
  assign n6605 = ( ~n6167 & n6603 ) | ( ~n6167 & n6604 ) | ( n6603 & n6604 ) ;
  assign n6606 = n6534 & n6605 ;
  buffer buf_n6607( .i (n6576), .o (n6607) );
  buffer buf_n6608( .i (n6607), .o (n6608) );
  assign n6609 = ~n6606 & n6608 ;
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  assign n6610 = ~n553 & n566 ;
  assign n6611 = n6608 | n6610 ;
  assign n6612 = ~n6609 & n6611 ;
  buffer buf_n6613( .i (n6565), .o (n6613) );
  assign n6614 = ( ~n6263 & n6612 ) | ( ~n6263 & n6613 ) | ( n6612 & n6613 ) ;
  assign n6615 = ( n3307 & ~n6401 ) | ( n3307 & n6405 ) | ( ~n6401 & n6405 ) ;
  buffer buf_n6616( .i (n6615), .o (n6616) );
  assign n6619 = n6029 & ~n6616 ;
  buffer buf_n6620( .i (n6619), .o (n6620) );
  buffer buf_n6621( .i (n6620), .o (n6621) );
  buffer buf_n6617( .i (n6616), .o (n6617) );
  buffer buf_n6618( .i (n6617), .o (n6618) );
  assign n6622 = n6618 | n6620 ;
  assign n6623 = ( ~n6523 & n6621 ) | ( ~n6523 & n6622 ) | ( n6621 & n6622 ) ;
  assign n6624 = n6576 | n6623 ;
  buffer buf_n3639( .i (n3638), .o (n3639) );
  buffer buf_n3640( .i (n3639), .o (n3640) );
  buffer buf_n3641( .i (n3640), .o (n3641) );
  assign n6625 = ~n3641 & n6576 ;
  assign n6626 = n6624 & ~n6625 ;
  assign n6627 = n6295 | n6626 ;
  assign n6628 = ( n4399 & n6288 ) | ( n4399 & ~n6482 ) | ( n6288 & ~n6482 ) ;
  buffer buf_n6629( .i (n6034), .o (n6629) );
  assign n6630 = ( n4399 & n6433 ) | ( n4399 & ~n6629 ) | ( n6433 & ~n6629 ) ;
  assign n6631 = n6628 & n6630 ;
  assign n6632 = n6607 & n6631 ;
  assign n6633 = n6295 & ~n6632 ;
  assign n6634 = n6627 & ~n6633 ;
  buffer buf_n6635( .i (n6583), .o (n6635) );
  assign n6636 = ( n6613 & ~n6634 ) | ( n6613 & n6635 ) | ( ~n6634 & n6635 ) ;
  assign n6637 = n6614 & ~n6636 ;
  buffer buf_n6638( .i (n6637), .o (n6638) );
  buffer buf_n6639( .i (n6638), .o (n6639) );
  buffer buf_n6640( .i (n6639), .o (n6640) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n718( .i (n717), .o (n718) );
  assign n6641 = ( n285 & n718 ) | ( n285 & n6638 ) | ( n718 & n6638 ) ;
  assign n6642 = n1728 | n6641 ;
  assign n6643 = ( ~n1729 & n6640 ) | ( ~n1729 & n6642 ) | ( n6640 & n6642 ) ;
  buffer buf_n6644( .i (n4656), .o (n6644) );
  assign n6645 = ( n3918 & n6403 ) | ( n3918 & ~n6644 ) | ( n6403 & ~n6644 ) ;
  buffer buf_n6646( .i (n6645), .o (n6646) );
  buffer buf_n6647( .i (n6646), .o (n6647) );
  buffer buf_n6648( .i (n6647), .o (n6648) );
  buffer buf_n6649( .i (n6648), .o (n6649) );
  assign n6650 = ( n3919 & ~n6385 ) | ( n3919 & n6404 ) | ( ~n6385 & n6404 ) ;
  assign n6651 = n6646 & n6650 ;
  buffer buf_n6652( .i (n6651), .o (n6652) );
  buffer buf_n6653( .i (n6652), .o (n6653) );
  buffer buf_n6654( .i (n5751), .o (n6654) );
  assign n6655 = n6652 | n6654 ;
  assign n6656 = ( ~n6649 & n6653 ) | ( ~n6649 & n6655 ) | ( n6653 & n6655 ) ;
  buffer buf_n6657( .i (n6656), .o (n6657) );
  buffer buf_n6658( .i (n6657), .o (n6658) );
  buffer buf_n6659( .i (n6522), .o (n6659) );
  buffer buf_n6660( .i (n6659), .o (n6660) );
  assign n6661 = ( ~n6395 & n6657 ) | ( ~n6395 & n6660 ) | ( n6657 & n6660 ) ;
  assign n6662 = ( n3827 & n4128 ) | ( n3827 & n6182 ) | ( n4128 & n6182 ) ;
  assign n6663 = ~n4129 & n6662 ;
  assign n6664 = n6660 & n6663 ;
  assign n6665 = ( ~n6658 & n6661 ) | ( ~n6658 & n6664 ) | ( n6661 & n6664 ) ;
  buffer buf_n6666( .i (n6665), .o (n6666) );
  buffer buf_n6667( .i (n6666), .o (n6667) );
  buffer buf_n6668( .i (n6667), .o (n6668) );
  buffer buf_n5828( .i (n5827), .o (n5828) );
  buffer buf_n5829( .i (n5828), .o (n5829) );
  buffer buf_n5830( .i (n5829), .o (n5830) );
  buffer buf_n5831( .i (n5830), .o (n5831) );
  buffer buf_n5832( .i (n5831), .o (n5832) );
  buffer buf_n5833( .i (n5832), .o (n5833) );
  buffer buf_n5834( .i (n5833), .o (n5834) );
  assign n6669 = n5831 & ~n6520 ;
  buffer buf_n6670( .i (n6669), .o (n6670) );
  buffer buf_n6671( .i (n6670), .o (n6671) );
  buffer buf_n6672( .i (n6395), .o (n6672) );
  assign n6673 = ( n6439 & ~n6670 ) | ( n6439 & n6672 ) | ( ~n6670 & n6672 ) ;
  assign n6674 = ( n5834 & n6671 ) | ( n5834 & ~n6673 ) | ( n6671 & ~n6673 ) ;
  assign n6675 = ( ~n6583 & n6666 ) | ( ~n6583 & n6674 ) | ( n6666 & n6674 ) ;
  buffer buf_n6676( .i (n6357), .o (n6676) );
  assign n6677 = ~n6675 & n6676 ;
  assign n6678 = ( n148 & n6668 ) | ( n148 & ~n6677 ) | ( n6668 & ~n6677 ) ;
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  assign n6679 = ( n6290 & n6531 ) | ( n6290 & ~n6629 ) | ( n6531 & ~n6629 ) ;
  assign n6680 = ~n1172 & n6679 ;
  buffer buf_n6681( .i (n6482), .o (n6681) );
  buffer buf_n6682( .i (n6681), .o (n6682) );
  assign n6683 = n6680 & ~n6682 ;
  buffer buf_n6684( .i (n6293), .o (n6684) );
  assign n6685 = ( n6582 & n6683 ) | ( n6582 & ~n6684 ) | ( n6683 & ~n6684 ) ;
  assign n6686 = ~n6583 & n6685 ;
  buffer buf_n6687( .i (n6686), .o (n6687) );
  buffer buf_n6688( .i (n6687), .o (n6688) );
  buffer buf_n6689( .i (n5208), .o (n6689) );
  assign n6690 = n6687 | n6689 ;
  assign n6691 = ( n6678 & n6688 ) | ( n6678 & n6690 ) | ( n6688 & n6690 ) ;
  buffer buf_n6692( .i (n6449), .o (n6692) );
  assign n6693 = n6691 | n6692 ;
  buffer buf_n5458( .i (n5457), .o (n5458) );
  buffer buf_n5459( .i (n5458), .o (n5459) );
  buffer buf_n5460( .i (n5459), .o (n5460) );
  buffer buf_n6694( .i (n6682), .o (n6694) );
  assign n6695 = ( n4887 & n6440 ) | ( n4887 & n6694 ) | ( n6440 & n6694 ) ;
  assign n6696 = n5460 & ~n6695 ;
  assign n6697 = ( ~n5491 & n6613 ) | ( ~n5491 & n6696 ) | ( n6613 & n6696 ) ;
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  assign n6698 = n430 & n6694 ;
  assign n6699 = n875 & n6698 ;
  assign n6700 = ~n5491 & n6699 ;
  assign n6701 = ( ~n4910 & n6697 ) | ( ~n4910 & n6700 ) | ( n6697 & n6700 ) ;
  assign n6702 = ~n6265 & n6701 ;
  assign n6703 = n6692 & ~n6702 ;
  assign n6704 = n6693 & ~n6703 ;
  buffer buf_n4040( .i (n4039), .o (n4040) );
  buffer buf_n4041( .i (n4040), .o (n4041) );
  buffer buf_n4042( .i (n4041), .o (n4042) );
  buffer buf_n4043( .i (n4042), .o (n4043) );
  buffer buf_n4044( .i (n4043), .o (n4044) );
  buffer buf_n4045( .i (n4044), .o (n4045) );
  assign n6705 = ( n4706 & n6385 ) | ( n4706 & ~n6404 ) | ( n6385 & ~n6404 ) ;
  buffer buf_n6706( .i (n6705), .o (n6706) );
  buffer buf_n6707( .i (n6706), .o (n6707) );
  buffer buf_n6708( .i (n6707), .o (n6708) );
  buffer buf_n6709( .i (n6708), .o (n6709) );
  assign n6710 = ( n5743 & n6408 ) | ( n5743 & n6706 ) | ( n6408 & n6706 ) ;
  buffer buf_n6711( .i (n6710), .o (n6711) );
  buffer buf_n6712( .i (n6711), .o (n6712) );
  assign n6713 = ~n4710 & n6711 ;
  assign n6714 = ( ~n6709 & n6712 ) | ( ~n6709 & n6713 ) | ( n6712 & n6713 ) ;
  assign n6715 = n6681 & n6714 ;
  assign n6716 = ~n6581 & n6715 ;
  buffer buf_n6717( .i (n6716), .o (n6717) );
  buffer buf_n6718( .i (n6717), .o (n6718) );
  buffer buf_n6719( .i (n6718), .o (n6719) );
  buffer buf_n6720( .i (n6694), .o (n6720) );
  assign n6721 = ( n875 & n6717 ) | ( n875 & ~n6720 ) | ( n6717 & ~n6720 ) ;
  assign n6722 = n4044 & ~n6721 ;
  assign n6723 = ( n4045 & n6719 ) | ( n4045 & ~n6722 ) | ( n6719 & ~n6722 ) ;
  assign n6724 = ~n1505 & n2783 ;
  assign n6725 = ( ~n724 & n4893 ) | ( ~n724 & n5751 ) | ( n4893 & n5751 ) ;
  assign n6726 = n725 & n6725 ;
  assign n6727 = ( n4558 & n5373 ) | ( n4558 & ~n5911 ) | ( n5373 & ~n5911 ) ;
  buffer buf_n6728( .i (n6727), .o (n6728) );
  assign n6732 = ( n5382 & n6372 ) | ( n5382 & n6728 ) | ( n6372 & n6728 ) ;
  buffer buf_n6733( .i (n6732), .o (n6733) );
  buffer buf_n6734( .i (n6733), .o (n6734) );
  buffer buf_n6735( .i (n6734), .o (n6735) );
  buffer buf_n6729( .i (n6728), .o (n6729) );
  buffer buf_n6730( .i (n6729), .o (n6730) );
  buffer buf_n6731( .i (n6730), .o (n6731) );
  buffer buf_n6736( .i (n6003), .o (n6736) );
  assign n6737 = ( n6400 & ~n6733 ) | ( n6400 & n6736 ) | ( ~n6733 & n6736 ) ;
  assign n6738 = n6731 | n6737 ;
  buffer buf_n6739( .i (n5415), .o (n6739) );
  assign n6740 = ( ~n6735 & n6738 ) | ( ~n6735 & n6739 ) | ( n6738 & n6739 ) ;
  assign n6741 = ( n3921 & ~n6131 ) | ( n3921 & n6740 ) | ( ~n6131 & n6740 ) ;
  assign n6742 = ( n4702 & n4738 ) | ( n4702 & ~n5381 ) | ( n4738 & ~n5381 ) ;
  buffer buf_n6743( .i (n6742), .o (n6743) );
  assign n6746 = n5894 & ~n6743 ;
  buffer buf_n6747( .i (n6746), .o (n6747) );
  buffer buf_n6748( .i (n6747), .o (n6748) );
  buffer buf_n6744( .i (n6743), .o (n6744) );
  buffer buf_n6745( .i (n6744), .o (n6745) );
  assign n6749 = n6745 | n6747 ;
  assign n6750 = ( ~n6325 & n6748 ) | ( ~n6325 & n6749 ) | ( n6748 & n6749 ) ;
  buffer buf_n6751( .i (n3920), .o (n6751) );
  buffer buf_n6752( .i (n6011), .o (n6752) );
  assign n6753 = ( ~n6750 & n6751 ) | ( ~n6750 & n6752 ) | ( n6751 & n6752 ) ;
  assign n6754 = n6741 | n6753 ;
  assign n6755 = ~n6726 & n6754 ;
  assign n6756 = ~n6724 & n6755 ;
  assign n6757 = ~n6660 & n6756 ;
  buffer buf_n6758( .i (n3929), .o (n6758) );
  buffer buf_n6759( .i (n6758), .o (n6759) );
  assign n6760 = ( n6003 & n6341 ) | ( n6003 & ~n6759 ) | ( n6341 & ~n6759 ) ;
  buffer buf_n6761( .i (n6760), .o (n6761) );
  buffer buf_n6762( .i (n6761), .o (n6762) );
  buffer buf_n6763( .i (n6762), .o (n6763) );
  assign n6764 = ( ~n5415 & n6401 ) | ( ~n5415 & n6761 ) | ( n6401 & n6761 ) ;
  assign n6765 = ( n6276 & ~n6325 ) | ( n6276 & n6764 ) | ( ~n6325 & n6764 ) ;
  assign n6766 = ( ~n440 & n6763 ) | ( ~n440 & n6765 ) | ( n6763 & n6765 ) ;
  assign n6767 = ~n6477 & n6766 ;
  assign n6768 = n632 & n868 ;
  assign n6769 = n6477 & ~n6768 ;
  assign n6770 = n6767 | n6769 ;
  assign n6771 = n4877 | n6770 ;
  assign n6772 = n6660 & n6771 ;
  assign n6773 = n6757 | n6772 ;
  buffer buf_n6774( .i (n5664), .o (n6774) );
  assign n6775 = n6773 & n6774 ;
  buffer buf_n6776( .i (n6404), .o (n6776) );
  assign n6777 = ( n1608 & n6335 ) | ( n1608 & ~n6776 ) | ( n6335 & ~n6776 ) ;
  assign n6778 = ( ~n1607 & n6010 ) | ( ~n1607 & n6385 ) | ( n6010 & n6385 ) ;
  buffer buf_n6779( .i (n6401), .o (n6779) );
  assign n6780 = ( ~n6776 & n6778 ) | ( ~n6776 & n6779 ) | ( n6778 & n6779 ) ;
  assign n6781 = ~n6777 & n6780 ;
  assign n6782 = n6412 & n6781 ;
  buffer buf_n6783( .i (n4738), .o (n6783) );
  buffer buf_n6784( .i (n5381), .o (n6784) );
  assign n6785 = ( ~n4560 & n6783 ) | ( ~n4560 & n6784 ) | ( n6783 & n6784 ) ;
  buffer buf_n6786( .i (n6785), .o (n6786) );
  buffer buf_n6787( .i (n6786), .o (n6787) );
  buffer buf_n6788( .i (n6787), .o (n6788) );
  buffer buf_n6789( .i (n6788), .o (n6789) );
  assign n6790 = ( ~n6400 & n6644 ) | ( ~n6400 & n6786 ) | ( n6644 & n6786 ) ;
  buffer buf_n6791( .i (n6790), .o (n6791) );
  buffer buf_n6792( .i (n6791), .o (n6792) );
  assign n6793 = n4564 & n6791 ;
  assign n6794 = ( ~n6789 & n6792 ) | ( ~n6789 & n6793 ) | ( n6792 & n6793 ) ;
  assign n6795 = n6412 | n6794 ;
  assign n6796 = ( ~n6351 & n6782 ) | ( ~n6351 & n6795 ) | ( n6782 & n6795 ) ;
  assign n6797 = n6659 & ~n6796 ;
  assign n6798 = ~n394 & n5743 ;
  assign n6799 = ( ~n2630 & n2718 ) | ( ~n2630 & n6798 ) | ( n2718 & n6798 ) ;
  assign n6800 = n6351 & ~n6799 ;
  assign n6801 = n6659 | n6800 ;
  assign n6802 = ~n6797 & n6801 ;
  assign n6803 = ~n6581 & n6802 ;
  assign n6804 = n6774 | n6803 ;
  assign n6805 = ~n6775 & n6804 ;
  buffer buf_n6806( .i (n6805), .o (n6806) );
  buffer buf_n6807( .i (n6806), .o (n6807) );
  assign n6808 = n2707 & ~n6806 ;
  assign n6809 = ( n6723 & n6807 ) | ( n6723 & ~n6808 ) | ( n6807 & ~n6808 ) ;
  assign n6810 = n5606 | n6809 ;
  buffer buf_n6811( .i (n605), .o (n6811) );
  assign n6812 = n555 | n6811 ;
  assign n6813 = ( n511 & n556 ) | ( n511 & n6812 ) | ( n556 & n6812 ) ;
  assign n6814 = n6351 & ~n6813 ;
  assign n6815 = n2133 & n6654 ;
  buffer buf_n6816( .i (n6408), .o (n6816) );
  buffer buf_n6817( .i (n6816), .o (n6817) );
  assign n6818 = n6815 | n6817 ;
  assign n6819 = ~n6814 & n6818 ;
  buffer buf_n6820( .i (n6819), .o (n6820) );
  buffer buf_n6821( .i (n6820), .o (n6821) );
  buffer buf_n6822( .i (n6821), .o (n6822) );
  buffer buf_n6823( .i (n6308), .o (n6823) );
  assign n6824 = ( n6397 & n6517 ) | ( n6397 & ~n6823 ) | ( n6517 & ~n6823 ) ;
  buffer buf_n6825( .i (n6824), .o (n6825) );
  buffer buf_n6826( .i (n6825), .o (n6826) );
  buffer buf_n6827( .i (n6519), .o (n6827) );
  assign n6828 = ( n6659 & n6826 ) | ( n6659 & ~n6827 ) | ( n6826 & ~n6827 ) ;
  assign n6829 = ~n6817 & n6825 ;
  assign n6830 = ( ~n6433 & n6826 ) | ( ~n6433 & n6829 ) | ( n6826 & n6829 ) ;
  assign n6831 = n6828 | n6830 ;
  assign n6832 = ( n6439 & n6820 ) | ( n6439 & ~n6831 ) | ( n6820 & ~n6831 ) ;
  buffer buf_n6833( .i (n6437), .o (n6833) );
  assign n6834 = ~n6832 & n6833 ;
  assign n6835 = ( n5701 & n6822 ) | ( n5701 & ~n6834 ) | ( n6822 & ~n6834 ) ;
  assign n6836 = ~n6676 & n6835 ;
  buffer buf_n6837( .i (n6736), .o (n6837) );
  buffer buf_n6838( .i (n6837), .o (n6838) );
  assign n6839 = ( ~n605 & n6739 ) | ( ~n605 & n6838 ) | ( n6739 & n6838 ) ;
  buffer buf_n6840( .i (n6839), .o (n6840) );
  buffer buf_n6841( .i (n6840), .o (n6841) );
  buffer buf_n6842( .i (n6841), .o (n6842) );
  buffer buf_n6843( .i (n6779), .o (n6843) );
  buffer buf_n6844( .i (n6843), .o (n6844) );
  assign n6845 = ( ~n6816 & n6840 ) | ( ~n6816 & n6844 ) | ( n6840 & n6844 ) ;
  assign n6846 = ( n6455 & ~n6530 ) | ( n6455 & n6845 ) | ( ~n6530 & n6845 ) ;
  assign n6847 = n6842 & n6846 ;
  buffer buf_n6848( .i (n6847), .o (n6848) );
  buffer buf_n6849( .i (n6848), .o (n6849) );
  assign n6850 = ( n6293 & ~n6560 ) | ( n6293 & n6848 ) | ( ~n6560 & n6848 ) ;
  assign n6851 = ( n2310 & n6816 ) | ( n2310 & n6844 ) | ( n6816 & n6844 ) ;
  buffer buf_n6852( .i (n6851), .o (n6852) );
  assign n6853 = ( ~n6629 & n6827 ) | ( ~n6629 & n6852 ) | ( n6827 & n6852 ) ;
  assign n6854 = ( n6213 & n6827 ) | ( n6213 & ~n6852 ) | ( n6827 & ~n6852 ) ;
  assign n6855 = n6853 & ~n6854 ;
  assign n6856 = ~n6293 & n6855 ;
  assign n6857 = ( n6849 & ~n6850 ) | ( n6849 & n6856 ) | ( ~n6850 & n6856 ) ;
  assign n6858 = ( n4766 & n6341 ) | ( n4766 & n6759 ) | ( n6341 & n6759 ) ;
  buffer buf_n6859( .i (n6858), .o (n6859) );
  buffer buf_n6865( .i (n6403), .o (n6865) );
  assign n6866 = ( n6155 & n6859 ) | ( n6155 & ~n6865 ) | ( n6859 & ~n6865 ) ;
  buffer buf_n6867( .i (n6866), .o (n6867) );
  assign n6870 = n6397 & ~n6867 ;
  buffer buf_n6871( .i (n6870), .o (n6871) );
  buffer buf_n6872( .i (n6871), .o (n6872) );
  buffer buf_n6868( .i (n6867), .o (n6868) );
  buffer buf_n6869( .i (n6868), .o (n6869) );
  assign n6873 = n6869 | n6871 ;
  buffer buf_n6874( .i (n6455), .o (n6874) );
  assign n6875 = ( n6872 & n6873 ) | ( n6872 & ~n6874 ) | ( n6873 & ~n6874 ) ;
  buffer buf_n6876( .i (n6875), .o (n6876) );
  buffer buf_n6877( .i (n6876), .o (n6877) );
  buffer buf_n6878( .i (n6522), .o (n6878) );
  buffer buf_n6879( .i (n6878), .o (n6879) );
  buffer buf_n6880( .i (n6879), .o (n6880) );
  assign n6881 = ( n6439 & ~n6876 ) | ( n6439 & n6880 ) | ( ~n6876 & n6880 ) ;
  assign n6882 = ( ~n4473 & n6816 ) | ( ~n4473 & n6844 ) | ( n6816 & n6844 ) ;
  buffer buf_n6883( .i (n6882), .o (n6883) );
  buffer buf_n6884( .i (n6883), .o (n6884) );
  assign n6885 = n6213 & ~n6883 ;
  assign n6886 = ( n6435 & ~n6884 ) | ( n6435 & n6885 ) | ( ~n6884 & n6885 ) ;
  assign n6887 = n6880 & n6886 ;
  assign n6888 = ( n6877 & n6881 ) | ( n6877 & n6887 ) | ( n6881 & n6887 ) ;
  assign n6889 = n6857 | n6888 ;
  assign n6890 = n6676 & n6889 ;
  assign n6891 = n6836 | n6890 ;
  assign n6892 = ~n6265 & n6891 ;
  assign n6893 = n5606 & ~n6892 ;
  assign n6894 = n6810 & ~n6893 ;
  assign n6895 = n6704 | n6894 ;
  assign n6896 = ( ~n6594 & n6643 ) | ( ~n6594 & n6895 ) | ( n6643 & n6895 ) ;
  assign n6897 = n6595 | n6896 ;
  buffer buf_n239( .i (n238), .o (n239) );
  assign n6898 = n1745 & ~n6559 ;
  assign n6899 = n706 & ~n6898 ;
  assign n6900 = n726 & n6182 ;
  assign n6901 = ( n6827 & n6874 ) | ( n6827 & n6900 ) | ( n6874 & n6900 ) ;
  assign n6902 = ~n6167 & n6901 ;
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n6903( .i (n6596), .o (n6903) );
  buffer buf_n6904( .i (n6903), .o (n6904) );
  assign n6905 = ( ~n4382 & n5996 ) | ( ~n4382 & n6904 ) | ( n5996 & n6904 ) ;
  assign n6906 = ( ~n4382 & n5996 ) | ( ~n4382 & n6654 ) | ( n5996 & n6654 ) ;
  assign n6907 = ( n2304 & n6905 ) | ( n2304 & ~n6906 ) | ( n6905 & ~n6906 ) ;
  buffer buf_n6908( .i (n6751), .o (n6908) );
  buffer buf_n6909( .i (n6908), .o (n6909) );
  buffer buf_n6910( .i (n6909), .o (n6910) );
  buffer buf_n6911( .i (n6519), .o (n6911) );
  assign n6912 = ( n6907 & ~n6910 ) | ( n6907 & n6911 ) | ( ~n6910 & n6911 ) ;
  assign n6913 = ( n5251 & n6383 ) | ( n5251 & ~n6736 ) | ( n6383 & ~n6736 ) ;
  buffer buf_n6914( .i (n6913), .o (n6914) );
  buffer buf_n6915( .i (n6914), .o (n6915) );
  buffer buf_n6916( .i (n6915), .o (n6916) );
  buffer buf_n6917( .i (n6916), .o (n6917) );
  assign n6920 = ~n6739 & n6914 ;
  buffer buf_n6921( .i (n6920), .o (n6921) );
  buffer buf_n6922( .i (n6921), .o (n6922) );
  buffer buf_n6923( .i (n5725), .o (n6923) );
  assign n6924 = ( n6904 & ~n6921 ) | ( n6904 & n6923 ) | ( ~n6921 & n6923 ) ;
  assign n6925 = ( n6917 & n6922 ) | ( n6917 & ~n6924 ) | ( n6922 & ~n6924 ) ;
  assign n6926 = ( n6910 & n6911 ) | ( n6910 & ~n6925 ) | ( n6911 & ~n6925 ) ;
  assign n6927 = n6912 & ~n6926 ;
  assign n6928 = n6902 | n6927 ;
  assign n6929 = ( n707 & ~n6899 ) | ( n707 & n6928 ) | ( ~n6899 & n6928 ) ;
  assign n6930 = n6720 & n6929 ;
  buffer buf_n6931( .i (n4478), .o (n6931) );
  assign n6932 = ( n20 & n6784 ) | ( n20 & n6931 ) | ( n6784 & n6931 ) ;
  buffer buf_n6933( .i (n6932), .o (n6933) );
  assign n6938 = ( ~n3918 & n6403 ) | ( ~n3918 & n6933 ) | ( n6403 & n6933 ) ;
  buffer buf_n6939( .i (n6938), .o (n6939) );
  buffer buf_n6940( .i (n6939), .o (n6940) );
  buffer buf_n6941( .i (n6940), .o (n6941) );
  buffer buf_n6942( .i (n6941), .o (n6942) );
  assign n6943 = ( n6596 & n6838 ) | ( n6596 & n6939 ) | ( n6838 & n6939 ) ;
  buffer buf_n6944( .i (n6943), .o (n6944) );
  buffer buf_n6945( .i (n6944), .o (n6945) );
  buffer buf_n6934( .i (n6933), .o (n6934) );
  buffer buf_n6935( .i (n6934), .o (n6935) );
  buffer buf_n6936( .i (n6935), .o (n6936) );
  buffer buf_n6937( .i (n6936), .o (n6937) );
  assign n6946 = n6937 & ~n6944 ;
  assign n6947 = ( n6942 & ~n6945 ) | ( n6942 & n6946 ) | ( ~n6945 & n6946 ) ;
  buffer buf_n6948( .i (n6947), .o (n6948) );
  buffer buf_n6949( .i (n6948), .o (n6949) );
  buffer buf_n6950( .i (n6817), .o (n6950) );
  buffer buf_n6951( .i (n6950), .o (n6951) );
  buffer buf_n6952( .i (n6290), .o (n6952) );
  assign n6953 = ( n6948 & n6951 ) | ( n6948 & n6952 ) | ( n6951 & n6952 ) ;
  assign n6954 = n727 & ~n6574 ;
  assign n6955 = ~n6952 & n6954 ;
  assign n6956 = ( n6949 & ~n6953 ) | ( n6949 & n6955 ) | ( ~n6953 & n6955 ) ;
  buffer buf_n4481( .i (n4480), .o (n4481) );
  buffer buf_n4482( .i (n4481), .o (n4482) );
  buffer buf_n4483( .i (n4482), .o (n4483) );
  buffer buf_n4484( .i (n4483), .o (n4484) );
  buffer buf_n4485( .i (n4484), .o (n4485) );
  buffer buf_n4486( .i (n4485), .o (n4486) );
  buffer buf_n4487( .i (n4486), .o (n4487) );
  buffer buf_n4488( .i (n4487), .o (n4488) );
  assign n6957 = ( ~n752 & n4488 ) | ( ~n752 & n6497 ) | ( n4488 & n6497 ) ;
  assign n6958 = n753 & n6957 ;
  assign n6959 = n6956 | n6958 ;
  assign n6960 = ~n6720 & n6959 ;
  assign n6961 = n6930 | n6960 ;
  assign n6962 = ( n3856 & n6689 ) | ( n3856 & ~n6961 ) | ( n6689 & ~n6961 ) ;
  buffer buf_n6963( .i (n6962), .o (n6963) );
  buffer buf_n6964( .i (n6963), .o (n6964) );
  assign n6965 = n208 & ~n6963 ;
  assign n6966 = ( n239 & ~n6964 ) | ( n239 & n6965 ) | ( ~n6964 & n6965 ) ;
  buffer buf_n6967( .i (n6966), .o (n6967) );
  buffer buf_n6968( .i (n6967), .o (n6968) );
  assign n6969 = ~n6844 & n6908 ;
  assign n6970 = n6183 & ~n6969 ;
  assign n6971 = ( n609 & n2498 ) | ( n609 & ~n6970 ) | ( n2498 & ~n6970 ) ;
  assign n6972 = n6879 & ~n6971 ;
  assign n6973 = n3009 | n6910 ;
  assign n6974 = ~n6879 & n6973 ;
  assign n6975 = n6972 | n6974 ;
  buffer buf_n6976( .i (n6560), .o (n6976) );
  assign n6977 = n6975 & ~n6976 ;
  assign n6978 = n1191 & ~n6904 ;
  buffer buf_n6979( .i (n6978), .o (n6979) );
  buffer buf_n6980( .i (n6979), .o (n6980) );
  assign n6981 = ( ~n1192 & n6455 ) | ( ~n1192 & n6522 ) | ( n6455 & n6522 ) ;
  assign n6982 = n6979 | n6981 ;
  assign n6983 = ( n6167 & n6980 ) | ( n6167 & n6982 ) | ( n6980 & n6982 ) ;
  assign n6984 = n6581 | n6983 ;
  assign n6985 = n6976 & n6984 ;
  assign n6986 = n6977 | n6985 ;
  assign n6987 = ~n6613 & n6986 ;
  assign n6988 = ( n4593 & ~n6629 ) | ( n4593 & n6874 ) | ( ~n6629 & n6874 ) ;
  buffer buf_n6989( .i (n4592), .o (n6989) );
  assign n6990 = ( ~n6482 & n6874 ) | ( ~n6482 & n6989 ) | ( n6874 & n6989 ) ;
  assign n6991 = ( n658 & ~n6988 ) | ( n658 & n6990 ) | ( ~n6988 & n6990 ) ;
  assign n6992 = n6880 | n6991 ;
  assign n6993 = n349 & ~n6681 ;
  assign n6994 = n6880 & ~n6993 ;
  assign n6995 = n6992 & ~n6994 ;
  buffer buf_n6996( .i (n6582), .o (n6996) );
  assign n6997 = n6995 & ~n6996 ;
  buffer buf_n6998( .i (n6565), .o (n6998) );
  assign n6999 = ~n6997 & n6998 ;
  assign n7000 = n6987 | n6999 ;
  buffer buf_n7001( .i (n6448), .o (n7001) );
  assign n7002 = n7000 & ~n7001 ;
  buffer buf_n7003( .i (n6400), .o (n7003) );
  assign n7004 = ( n6405 & n6865 ) | ( n6405 & n7003 ) | ( n6865 & n7003 ) ;
  buffer buf_n7005( .i (n7004), .o (n7005) );
  assign n7009 = ( n6517 & n6903 ) | ( n6517 & ~n7005 ) | ( n6903 & ~n7005 ) ;
  buffer buf_n7010( .i (n7009), .o (n7010) );
  buffer buf_n7011( .i (n7010), .o (n7011) );
  buffer buf_n7012( .i (n7011), .o (n7012) );
  buffer buf_n7006( .i (n7005), .o (n7006) );
  buffer buf_n7007( .i (n7006), .o (n7007) );
  buffer buf_n7008( .i (n7007), .o (n7008) );
  buffer buf_n7013( .i (n5903), .o (n7013) );
  assign n7014 = ( ~n6519 & n7010 ) | ( ~n6519 & n7013 ) | ( n7010 & n7013 ) ;
  assign n7015 = n7008 | n7014 ;
  buffer buf_n7016( .i (n6904), .o (n7016) );
  buffer buf_n7017( .i (n7016), .o (n7017) );
  buffer buf_n7018( .i (n7017), .o (n7018) );
  assign n7019 = ( n7012 & n7015 ) | ( n7012 & ~n7018 ) | ( n7015 & ~n7018 ) ;
  assign n7020 = n6682 & ~n7019 ;
  assign n7021 = ( ~n1757 & n4802 ) | ( ~n1757 & n6559 ) | ( n4802 & n6559 ) ;
  assign n7022 = n6682 | n7021 ;
  assign n7023 = ( ~n6694 & n7020 ) | ( ~n6694 & n7022 ) | ( n7020 & n7022 ) ;
  buffer buf_n7024( .i (n6220), .o (n7024) );
  assign n7025 = n7023 & n7024 ;
  buffer buf_n7026( .i (n6903), .o (n7026) );
  assign n7027 = ~n921 & n7026 ;
  buffer buf_n7028( .i (n7027), .o (n7028) );
  assign n7029 = ~n6878 & n7028 ;
  assign n7030 = ( ~n923 & n6911 ) | ( ~n923 & n7028 ) | ( n6911 & n7028 ) ;
  assign n7031 = ( ~n6435 & n7029 ) | ( ~n6435 & n7030 ) | ( n7029 & n7030 ) ;
  buffer buf_n7032( .i (n6681), .o (n7032) );
  assign n7033 = ~n7031 & n7032 ;
  buffer buf_n7034( .i (n6843), .o (n7034) );
  assign n7035 = ( n2699 & n6518 ) | ( n2699 & n7034 ) | ( n6518 & n7034 ) ;
  buffer buf_n7036( .i (n7035), .o (n7036) );
  buffer buf_n7037( .i (n7036), .o (n7037) );
  assign n7038 = n6911 & ~n7036 ;
  buffer buf_n7039( .i (n7034), .o (n7039) );
  buffer buf_n7040( .i (n7039), .o (n7040) );
  buffer buf_n7041( .i (n7040), .o (n7041) );
  assign n7042 = ( ~n7037 & n7038 ) | ( ~n7037 & n7041 ) | ( n7038 & n7041 ) ;
  assign n7043 = ~n7032 & n7042 ;
  buffer buf_n7044( .i (n7032), .o (n7044) );
  assign n7045 = ( ~n7033 & n7043 ) | ( ~n7033 & n7044 ) | ( n7043 & n7044 ) ;
  assign n7046 = n7024 | n7045 ;
  assign n7047 = ( ~n6998 & n7025 ) | ( ~n6998 & n7046 ) | ( n7025 & n7046 ) ;
  buffer buf_n7048( .i (n6635), .o (n7048) );
  assign n7049 = n7047 & ~n7048 ;
  assign n7050 = n7001 & ~n7049 ;
  assign n7051 = n7002 | n7050 ;
  buffer buf_n7052( .i (n180), .o (n7052) );
  assign n7053 = n7051 & n7052 ;
  buffer buf_n7054( .i (n6517), .o (n7054) );
  buffer buf_n7055( .i (n7054), .o (n7055) );
  buffer buf_n7056( .i (n7055), .o (n7056) );
  assign n7057 = ( n6878 & ~n6950 ) | ( n6878 & n7056 ) | ( ~n6950 & n7056 ) ;
  buffer buf_n7058( .i (n7057), .o (n7058) );
  buffer buf_n7059( .i (n7058), .o (n7059) );
  buffer buf_n7060( .i (n7059), .o (n7060) );
  assign n7061 = n6608 & n7059 ;
  assign n7062 = ( ~n4237 & n7060 ) | ( ~n4237 & n7061 ) | ( n7060 & n7061 ) ;
  assign n7063 = n6405 | n6865 ;
  buffer buf_n7064( .i (n7063), .o (n7064) );
  buffer buf_n7067( .i (n6776), .o (n7067) );
  assign n7068 = ( n6843 & n7064 ) | ( n6843 & ~n7067 ) | ( n7064 & ~n7067 ) ;
  assign n7069 = ( n6843 & n6903 ) | ( n6843 & n7064 ) | ( n6903 & n7064 ) ;
  assign n7070 = ( n6062 & n7068 ) | ( n6062 & ~n7069 ) | ( n7068 & ~n7069 ) ;
  buffer buf_n7071( .i (n6923), .o (n7071) );
  assign n7072 = n7070 & n7071 ;
  assign n7073 = n1238 & n7054 ;
  assign n7074 = n7071 | n7073 ;
  assign n7075 = ~n7072 & n7074 ;
  assign n7076 = n6951 & ~n7075 ;
  buffer buf_n7065( .i (n7064), .o (n7065) );
  buffer buf_n7066( .i (n7065), .o (n7066) );
  assign n7077 = ~n2930 & n7034 ;
  assign n7078 = ( ~n2120 & n7066 ) | ( ~n2120 & n7077 ) | ( n7066 & n7077 ) ;
  assign n7079 = n7017 | n7078 ;
  assign n7080 = ~n6951 & n7079 ;
  assign n7081 = n7076 | n7080 ;
  buffer buf_n7082( .i (n7081), .o (n7082) );
  buffer buf_n7083( .i (n7082), .o (n7083) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n5082( .i (n5081), .o (n5082) );
  buffer buf_n5083( .i (n5082), .o (n5083) );
  assign n7084 = ( n280 & n1747 ) | ( n280 & ~n5083 ) | ( n1747 & ~n5083 ) ;
  assign n7085 = n7082 & ~n7084 ;
  assign n7086 = ( ~n7062 & n7083 ) | ( ~n7062 & n7085 ) | ( n7083 & n7085 ) ;
  buffer buf_n7087( .i (n6676), .o (n7087) );
  assign n7088 = ~n7086 & n7087 ;
  buffer buf_n7089( .i (n6596), .o (n7089) );
  assign n7090 = ( n5041 & ~n6823 ) | ( n5041 & n7089 ) | ( ~n6823 & n7089 ) ;
  buffer buf_n7091( .i (n7090), .o (n7091) );
  assign n7094 = n7016 & ~n7091 ;
  buffer buf_n7095( .i (n7094), .o (n7095) );
  buffer buf_n7096( .i (n7095), .o (n7096) );
  buffer buf_n7092( .i (n7091), .o (n7092) );
  buffer buf_n7093( .i (n7092), .o (n7093) );
  assign n7097 = n7093 | n7095 ;
  assign n7098 = ( ~n5664 & n7096 ) | ( ~n5664 & n7097 ) | ( n7096 & n7097 ) ;
  assign n7099 = ( ~n6608 & n6976 ) | ( ~n6608 & n7098 ) | ( n6976 & n7098 ) ;
  buffer buf_n6128( .i (n6127), .o (n6128) );
  buffer buf_n6129( .i (n6128), .o (n6129) );
  buffer buf_n6130( .i (n6129), .o (n6130) );
  assign n7100 = ( n924 & n2571 ) | ( n924 & ~n6130 ) | ( n2571 & ~n6130 ) ;
  buffer buf_n7101( .i (n924), .o (n7101) );
  assign n7102 = ( n6437 & n7100 ) | ( n6437 & n7101 ) | ( n7100 & n7101 ) ;
  buffer buf_n7103( .i (n6607), .o (n7103) );
  assign n7104 = ( n6976 & n7102 ) | ( n6976 & n7103 ) | ( n7102 & n7103 ) ;
  assign n7105 = n7099 & n7104 ;
  buffer buf_n7106( .i (n6559), .o (n7106) );
  assign n7107 = n1758 | n7106 ;
  buffer buf_n7108( .i (n6672), .o (n7108) );
  assign n7109 = ( n7103 & ~n7107 ) | ( n7103 & n7108 ) | ( ~n7107 & n7108 ) ;
  assign n7110 = ~n6502 & n7109 ;
  assign n7111 = n7105 | n7110 ;
  assign n7112 = ~n7087 & n7111 ;
  assign n7113 = n7088 | n7112 ;
  assign n7114 = ~n5857 & n7113 ;
  assign n7115 = n7052 | n7114 ;
  assign n7116 = ~n7053 & n7115 ;
  assign n7117 = ( n996 & n3919 ) | ( n996 & n6010 ) | ( n3919 & n6010 ) ;
  buffer buf_n7118( .i (n7117), .o (n7118) );
  buffer buf_n7119( .i (n7118), .o (n7119) );
  buffer buf_n7120( .i (n7119), .o (n7120) );
  buffer buf_n7121( .i (n6779), .o (n7121) );
  assign n7122 = ( n6752 & ~n7118 ) | ( n6752 & n7121 ) | ( ~n7118 & n7121 ) ;
  assign n7123 = ( ~n6654 & n6908 ) | ( ~n6654 & n7122 ) | ( n6908 & n7122 ) ;
  assign n7124 = ~n7120 & n7123 ;
  assign n7125 = n6950 | n7124 ;
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n1637( .i (n1636), .o (n1637) );
  assign n7126 = n1637 & ~n6909 ;
  assign n7127 = n6950 & ~n7126 ;
  assign n7128 = n7125 & ~n7127 ;
  assign n7129 = n6672 | n7128 ;
  assign n7130 = ( n3370 & n6183 ) | ( n3370 & ~n6817 ) | ( n6183 & ~n6817 ) ;
  buffer buf_n7131( .i (n6752), .o (n7131) );
  buffer buf_n7132( .i (n7131), .o (n7132) );
  assign n7133 = ( n3370 & n6530 ) | ( n3370 & ~n7132 ) | ( n6530 & ~n7132 ) ;
  assign n7134 = n7130 & n7133 ;
  assign n7135 = ~n6580 & n7134 ;
  assign n7136 = n6672 & ~n7135 ;
  assign n7137 = n7129 & ~n7136 ;
  assign n7138 = n6488 | n7137 ;
  buffer buf_n7139( .i (n6739), .o (n7139) );
  assign n7140 = ( n2670 & ~n5725 ) | ( n2670 & n7139 ) | ( ~n5725 & n7139 ) ;
  buffer buf_n7141( .i (n5943), .o (n7141) );
  buffer buf_n7142( .i (n7141), .o (n7142) );
  assign n7143 = ( n5153 & n7139 ) | ( n5153 & n7142 ) | ( n7139 & n7142 ) ;
  assign n7144 = ~n7140 & n7143 ;
  buffer buf_n7145( .i (n7144), .o (n7145) );
  buffer buf_n7146( .i (n7145), .o (n7146) );
  buffer buf_n7147( .i (n7146), .o (n7147) );
  buffer buf_n7148( .i (n7132), .o (n7148) );
  assign n7149 = ( n1001 & n7145 ) | ( n1001 & ~n7148 ) | ( n7145 & ~n7148 ) ;
  assign n7150 = n1945 & ~n7149 ;
  assign n7151 = ( n1946 & n7147 ) | ( n1946 & ~n7150 ) | ( n7147 & ~n7150 ) ;
  assign n7152 = ~n6582 & n7151 ;
  assign n7153 = n6488 & ~n7152 ;
  assign n7154 = n7138 & ~n7153 ;
  assign n7155 = ( n3856 & n6208 ) | ( n3856 & ~n7154 ) | ( n6208 & ~n7154 ) ;
  buffer buf_n7156( .i (n7155), .o (n7156) );
  buffer buf_n7157( .i (n7156), .o (n7157) );
  buffer buf_n7158( .i (n5783), .o (n7158) );
  buffer buf_n7159( .i (n7158), .o (n7159) );
  buffer buf_n7160( .i (n7159), .o (n7160) );
  buffer buf_n7161( .i (n7160), .o (n7161) );
  assign n7162 = ~n7156 & n7161 ;
  assign n7163 = ( n267 & ~n7157 ) | ( n267 & n7162 ) | ( ~n7157 & n7162 ) ;
  assign n7164 = ( n3919 & ~n5415 ) | ( n3919 & n5943 ) | ( ~n5415 & n5943 ) ;
  buffer buf_n7165( .i (n7164), .o (n7165) );
  buffer buf_n7170( .i (n6838), .o (n7170) );
  assign n7171 = ( n7139 & n7165 ) | ( n7139 & ~n7170 ) | ( n7165 & ~n7170 ) ;
  buffer buf_n7172( .i (n7171), .o (n7172) );
  buffer buf_n7173( .i (n7172), .o (n7173) );
  buffer buf_n7174( .i (n7173), .o (n7174) );
  buffer buf_n7175( .i (n7174), .o (n7175) );
  assign n7176 = ( n6909 & n7071 ) | ( n6909 & n7172 ) | ( n7071 & n7172 ) ;
  buffer buf_n7177( .i (n7176), .o (n7177) );
  buffer buf_n7178( .i (n7177), .o (n7178) );
  buffer buf_n7166( .i (n7165), .o (n7166) );
  buffer buf_n7167( .i (n7166), .o (n7167) );
  buffer buf_n7168( .i (n7167), .o (n7168) );
  buffer buf_n7169( .i (n7168), .o (n7169) );
  assign n7179 = n7169 & ~n7177 ;
  assign n7180 = ( n7175 & ~n7178 ) | ( n7175 & n7179 ) | ( ~n7178 & n7179 ) ;
  assign n7181 = ( n6833 & ~n7044 ) | ( n6833 & n7180 ) | ( ~n7044 & n7180 ) ;
  buffer buf_n7182( .i (n7181), .o (n7182) );
  assign n7183 = ( ~n5208 & n7158 ) | ( ~n5208 & n7182 ) | ( n7158 & n7182 ) ;
  buffer buf_n7184( .i (n6720), .o (n7184) );
  assign n7185 = ( ~n7158 & n7182 ) | ( ~n7158 & n7184 ) | ( n7182 & n7184 ) ;
  assign n7186 = n7183 & n7185 ;
  assign n7187 = ( ~n2631 & n7013 ) | ( ~n2631 & n7071 ) | ( n7013 & n7071 ) ;
  buffer buf_n7188( .i (n7187), .o (n7188) );
  buffer buf_n7189( .i (n7188), .o (n7189) );
  buffer buf_n7190( .i (n7189), .o (n7190) );
  assign n7191 = ( n6497 & ~n6952 ) | ( n6497 & n7188 ) | ( ~n6952 & n7188 ) ;
  buffer buf_n7192( .i (n6879), .o (n7192) );
  assign n7193 = ( n6437 & n7191 ) | ( n6437 & ~n7192 ) | ( n7191 & ~n7192 ) ;
  assign n7194 = n7190 & n7193 ;
  buffer buf_n7195( .i (n7194), .o (n7195) );
  buffer buf_n7196( .i (n7195), .o (n7196) );
  buffer buf_n7197( .i (n731), .o (n7197) );
  assign n7198 = ( n7184 & n7195 ) | ( n7184 & ~n7197 ) | ( n7195 & ~n7197 ) ;
  assign n7199 = n7196 & ~n7198 ;
  assign n7200 = n7186 | n7199 ;
  assign n7201 = n120 | n7200 ;
  assign n7202 = ~n2006 & n7041 ;
  assign n7203 = ( ~n2123 & n3871 ) | ( ~n2123 & n7202 ) | ( n3871 & n7202 ) ;
  assign n7204 = n7103 & ~n7203 ;
  buffer buf_n7205( .i (n7148), .o (n7205) );
  buffer buf_n7206( .i (n2037), .o (n7206) );
  assign n7207 = ( n6952 & ~n7205 ) | ( n6952 & n7206 ) | ( ~n7205 & n7206 ) ;
  buffer buf_n7208( .i (n2036), .o (n7208) );
  assign n7209 = ( n6878 & n7148 ) | ( n6878 & n7208 ) | ( n7148 & n7208 ) ;
  buffer buf_n7210( .i (n6923), .o (n7210) );
  buffer buf_n7211( .i (n7210), .o (n7211) );
  buffer buf_n7212( .i (n7211), .o (n7212) );
  assign n7213 = ( n7041 & ~n7209 ) | ( n7041 & n7212 ) | ( ~n7209 & n7212 ) ;
  assign n7214 = ~n7207 & n7213 ;
  assign n7215 = n7103 | n7214 ;
  assign n7216 = ( ~n6502 & n7204 ) | ( ~n6502 & n7215 ) | ( n7204 & n7215 ) ;
  assign n7217 = n5296 | n7216 ;
  assign n7218 = n6607 & n7192 ;
  buffer buf_n7219( .i (n7041), .o (n7219) );
  assign n7220 = n540 | n7219 ;
  assign n7221 = ( ~n2098 & n7218 ) | ( ~n2098 & n7220 ) | ( n7218 & n7220 ) ;
  buffer buf_n7222( .i (n7044), .o (n7222) );
  assign n7223 = n7221 & ~n7222 ;
  buffer buf_n7224( .i (n6493), .o (n7224) );
  assign n7225 = ~n7223 & n7224 ;
  assign n7226 = n7217 & ~n7225 ;
  assign n7227 = ~n6265 & n7226 ;
  buffer buf_n7228( .i (n6196), .o (n7228) );
  buffer buf_n7229( .i (n7228), .o (n7229) );
  assign n7230 = ~n7227 & n7229 ;
  assign n7231 = n7201 & ~n7230 ;
  assign n7232 = n7163 | n7231 ;
  assign n7233 = ( ~n6967 & n7116 ) | ( ~n6967 & n7232 ) | ( n7116 & n7232 ) ;
  assign n7234 = n6968 | n7233 ;
  buffer buf_n4947( .i (n4946), .o (n4947) );
  buffer buf_n4948( .i (n4947), .o (n4948) );
  buffer buf_n4949( .i (n4948), .o (n4949) );
  buffer buf_n4950( .i (n4949), .o (n4950) );
  buffer buf_n4951( .i (n4950), .o (n4951) );
  buffer buf_n4952( .i (n4951), .o (n4952) );
  buffer buf_n4633( .i (n4632), .o (n4633) );
  buffer buf_n4634( .i (n4633), .o (n4634) );
  buffer buf_n4635( .i (n4634), .o (n4635) );
  buffer buf_n4636( .i (n4635), .o (n4636) );
  buffer buf_n4637( .i (n4636), .o (n4637) );
  buffer buf_n4638( .i (n4637), .o (n4638) );
  assign n7235 = ( n759 & n4638 ) | ( n759 & ~n4951 ) | ( n4638 & ~n4951 ) ;
  buffer buf_n5084( .i (n5083), .o (n5084) );
  buffer buf_n5085( .i (n5084), .o (n5085) );
  assign n7236 = ( n5085 & ~n6259 ) | ( n5085 & n6540 ) | ( ~n6259 & n6540 ) ;
  assign n7237 = ~n6448 & n7236 ;
  buffer buf_n7238( .i (n7048), .o (n7238) );
  assign n7239 = n7237 & n7238 ;
  assign n7240 = n4638 & n7239 ;
  assign n7241 = ( n4952 & n7235 ) | ( n4952 & n7240 ) | ( n7235 & n7240 ) ;
  buffer buf_n7242( .i (n7241), .o (n7242) );
  buffer buf_n7243( .i (n7242), .o (n7243) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  assign n7244 = ~n266 & n572 ;
  assign n7245 = n7052 & n7244 ;
  buffer buf_n7246( .i (n6783), .o (n7246) );
  buffer buf_n7247( .i (n7246), .o (n7247) );
  assign n7248 = ( ~n6383 & n6736 ) | ( ~n6383 & n7247 ) | ( n6736 & n7247 ) ;
  buffer buf_n7249( .i (n7248), .o (n7249) );
  buffer buf_n7254( .i (n6155), .o (n7254) );
  assign n7255 = ( n6838 & ~n7249 ) | ( n6838 & n7254 ) | ( ~n7249 & n7254 ) ;
  buffer buf_n7256( .i (n7255), .o (n7256) );
  buffer buf_n7257( .i (n7256), .o (n7257) );
  buffer buf_n7258( .i (n7257), .o (n7258) );
  buffer buf_n7259( .i (n7258), .o (n7259) );
  buffer buf_n7260( .i (n7139), .o (n7260) );
  assign n7261 = ( ~n7054 & n7256 ) | ( ~n7054 & n7260 ) | ( n7256 & n7260 ) ;
  buffer buf_n7262( .i (n7261), .o (n7262) );
  buffer buf_n7263( .i (n7262), .o (n7263) );
  buffer buf_n7250( .i (n7249), .o (n7250) );
  buffer buf_n7251( .i (n7250), .o (n7251) );
  buffer buf_n7252( .i (n7251), .o (n7252) );
  buffer buf_n7253( .i (n7252), .o (n7253) );
  assign n7264 = n7253 & n7262 ;
  assign n7265 = ( ~n7259 & n7263 ) | ( ~n7259 & n7264 ) | ( n7263 & n7264 ) ;
  assign n7266 = ~n7032 & n7265 ;
  buffer buf_n7267( .i (n6580), .o (n7267) );
  buffer buf_n7268( .i (n7267), .o (n7268) );
  assign n7269 = n7266 & ~n7268 ;
  buffer buf_n7270( .i (n7269), .o (n7270) );
  buffer buf_n7271( .i (n7270), .o (n7271) );
  buffer buf_n4505( .i (n4504), .o (n4505) );
  buffer buf_n4506( .i (n4505), .o (n4506) );
  buffer buf_n4507( .i (n4506), .o (n4507) );
  buffer buf_n4508( .i (n4507), .o (n4508) );
  assign n7272 = n4508 | n7270 ;
  assign n7273 = ( n4045 & n7271 ) | ( n4045 & n7272 ) | ( n7271 & n7272 ) ;
  assign n7274 = ~n4911 & n7273 ;
  buffer buf_n7275( .i (n7274), .o (n7275) );
  buffer buf_n7276( .i (n7275), .o (n7276) );
  assign n7277 = n760 | n7275 ;
  assign n7278 = ( n7245 & n7276 ) | ( n7245 & n7277 ) | ( n7276 & n7277 ) ;
  buffer buf_n7279( .i (n6931), .o (n7279) );
  buffer buf_n7280( .i (n7279), .o (n7280) );
  assign n7281 = ( n3918 & n6071 ) | ( n3918 & ~n7280 ) | ( n6071 & ~n7280 ) ;
  buffer buf_n7282( .i (n7281), .o (n7282) );
  assign n7287 = ( n6011 & ~n6308 ) | ( n6011 & n7282 ) | ( ~n6308 & n7282 ) ;
  buffer buf_n7288( .i (n7287), .o (n7288) );
  buffer buf_n7289( .i (n7288), .o (n7289) );
  buffer buf_n7290( .i (n7289), .o (n7290) );
  buffer buf_n7291( .i (n7290), .o (n7291) );
  assign n7292 = ( n6908 & ~n7026 ) | ( n6908 & n7288 ) | ( ~n7026 & n7288 ) ;
  buffer buf_n7293( .i (n7292), .o (n7293) );
  buffer buf_n7294( .i (n7293), .o (n7294) );
  buffer buf_n7283( .i (n7282), .o (n7283) );
  buffer buf_n7284( .i (n7283), .o (n7284) );
  buffer buf_n7285( .i (n7284), .o (n7285) );
  buffer buf_n7286( .i (n7285), .o (n7286) );
  assign n7295 = ~n7286 & n7293 ;
  assign n7296 = ( ~n7291 & n7294 ) | ( ~n7291 & n7295 ) | ( n7294 & n7295 ) ;
  buffer buf_n7297( .i (n7212), .o (n7297) );
  assign n7298 = n7296 | n7297 ;
  assign n7299 = n3117 & n7148 ;
  assign n7300 = ~n6580 & n7299 ;
  assign n7301 = n7297 & ~n7300 ;
  assign n7302 = n7298 & ~n7301 ;
  buffer buf_n7303( .i (n6951), .o (n7303) );
  buffer buf_n7304( .i (n7303), .o (n7304) );
  buffer buf_n7305( .i (n7304), .o (n7305) );
  assign n7306 = n7302 | n7305 ;
  assign n7307 = n7089 & n7142 ;
  buffer buf_n7308( .i (n6823), .o (n7308) );
  assign n7309 = ( n7131 & n7307 ) | ( n7131 & n7308 ) | ( n7307 & n7308 ) ;
  buffer buf_n7310( .i (n7309), .o (n7310) );
  buffer buf_n7311( .i (n7310), .o (n7311) );
  buffer buf_n7312( .i (n7311), .o (n7312) );
  buffer buf_n7313( .i (n7013), .o (n7313) );
  assign n7314 = ( n7017 & ~n7310 ) | ( n7017 & n7313 ) | ( ~n7310 & n7313 ) ;
  assign n7315 = ( n7205 & n7212 ) | ( n7205 & n7314 ) | ( n7212 & n7314 ) ;
  assign n7316 = ~n7312 & n7315 ;
  assign n7317 = ~n7268 & n7316 ;
  assign n7318 = n7305 & ~n7317 ;
  assign n7319 = n7306 & ~n7318 ;
  assign n7320 = n6206 | n7319 ;
  buffer buf_n7321( .i (n4577), .o (n7321) );
  assign n7322 = ( n5942 & n6644 ) | ( n5942 & n7321 ) | ( n6644 & n7321 ) ;
  buffer buf_n7323( .i (n7322), .o (n7323) );
  buffer buf_n7324( .i (n7323), .o (n7324) );
  buffer buf_n7325( .i (n7324), .o (n7325) );
  buffer buf_n7326( .i (n7325), .o (n7326) );
  buffer buf_n7327( .i (n7326), .o (n7327) );
  buffer buf_n7328( .i (n7327), .o (n7328) );
  buffer buf_n7329( .i (n7328), .o (n7329) );
  buffer buf_n7330( .i (n7329), .o (n7330) );
  buffer buf_n7331( .i (n7313), .o (n7331) );
  assign n7332 = ( n7205 & ~n7328 ) | ( n7205 & n7331 ) | ( ~n7328 & n7331 ) ;
  buffer buf_n7333( .i (n7205), .o (n7333) );
  assign n7334 = ( n7303 & n7332 ) | ( n7303 & n7333 ) | ( n7332 & n7333 ) ;
  assign n7335 = ( n1947 & n7330 ) | ( n1947 & ~n7334 ) | ( n7330 & ~n7334 ) ;
  assign n7336 = n745 & n1764 ;
  buffer buf_n7337( .i (n7336), .o (n7337) );
  buffer buf_n7338( .i (n7337), .o (n7338) );
  assign n7339 = n6774 | n7337 ;
  assign n7340 = ( n7335 & n7338 ) | ( n7335 & n7339 ) | ( n7338 & n7339 ) ;
  assign n7341 = ~n6635 & n7340 ;
  assign n7342 = n6206 & ~n7341 ;
  assign n7343 = n7320 & ~n7342 ;
  assign n7344 = n7229 | n7343 ;
  buffer buf_n4334( .i (n4333), .o (n4334) );
  buffer buf_n4335( .i (n4334), .o (n4335) );
  buffer buf_n4336( .i (n4335), .o (n4336) );
  assign n7345 = ( n2210 & ~n7018 ) | ( n2210 & n7331 ) | ( ~n7018 & n7331 ) ;
  buffer buf_n7346( .i (n7260), .o (n7346) );
  buffer buf_n7347( .i (n7346), .o (n7347) );
  buffer buf_n7348( .i (n7347), .o (n7348) );
  assign n7349 = ( n2210 & n7331 ) | ( n2210 & n7348 ) | ( n7331 & n7348 ) ;
  assign n7350 = ( n4336 & n7345 ) | ( n4336 & ~n7349 ) | ( n7345 & ~n7349 ) ;
  assign n7351 = n7044 & n7350 ;
  buffer buf_n7352( .i (n6383), .o (n7352) );
  buffer buf_n7353( .i (n7321), .o (n7353) );
  buffer buf_n7354( .i (n7280), .o (n7354) );
  assign n7355 = ( n7352 & ~n7353 ) | ( n7352 & n7354 ) | ( ~n7353 & n7354 ) ;
  buffer buf_n7356( .i (n7355), .o (n7356) );
  assign n7361 = ( n7089 & ~n7170 ) | ( n7089 & n7356 ) | ( ~n7170 & n7356 ) ;
  buffer buf_n7362( .i (n7361), .o (n7362) );
  assign n7365 = n7016 & ~n7362 ;
  buffer buf_n7366( .i (n7365), .o (n7366) );
  buffer buf_n7367( .i (n7366), .o (n7367) );
  buffer buf_n7363( .i (n7362), .o (n7363) );
  buffer buf_n7364( .i (n7363), .o (n7364) );
  assign n7368 = n7364 | n7366 ;
  assign n7369 = ( ~n5664 & n7367 ) | ( ~n5664 & n7368 ) | ( n7367 & n7368 ) ;
  buffer buf_n7370( .i (n7333), .o (n7370) );
  assign n7371 = n7369 | n7370 ;
  assign n7372 = ( ~n7222 & n7351 ) | ( ~n7222 & n7371 ) | ( n7351 & n7371 ) ;
  assign n7373 = n6998 & n7372 ;
  buffer buf_n7374( .i (n7352), .o (n7374) );
  buffer buf_n7375( .i (n7374), .o (n7375) );
  assign n7376 = ( n6823 & ~n6915 ) | ( n6823 & n7375 ) | ( ~n6915 & n7375 ) ;
  buffer buf_n7377( .i (n7376), .o (n7377) );
  buffer buf_n7378( .i (n7377), .o (n7378) );
  buffer buf_n7379( .i (n7378), .o (n7379) );
  buffer buf_n7380( .i (n7379), .o (n7380) );
  assign n7381 = ( n6530 & ~n7016 ) | ( n6530 & n7377 ) | ( ~n7016 & n7377 ) ;
  buffer buf_n7382( .i (n7381), .o (n7382) );
  buffer buf_n7383( .i (n7382), .o (n7383) );
  buffer buf_n6918( .i (n6917), .o (n6918) );
  buffer buf_n6919( .i (n6918), .o (n6919) );
  assign n7384 = n6919 & n7382 ;
  assign n7385 = ( ~n7380 & n7383 ) | ( ~n7380 & n7384 ) | ( n7383 & n7384 ) ;
  assign n7386 = n7370 & ~n7385 ;
  buffer buf_n3616( .i (n3615), .o (n3616) );
  buffer buf_n3617( .i (n3616), .o (n3617) );
  buffer buf_n4428( .i (n4427), .o (n4428) );
  assign n7387 = n3617 | n4428 ;
  assign n7388 = ~n7303 & n7387 ;
  assign n7389 = n7370 | n7388 ;
  assign n7390 = ~n7386 & n7389 ;
  assign n7391 = n6998 | n7390 ;
  assign n7392 = ( ~n4910 & n7373 ) | ( ~n4910 & n7391 ) | ( n7373 & n7391 ) ;
  assign n7393 = ~n7238 & n7392 ;
  assign n7394 = n7229 & ~n7393 ;
  assign n7395 = n7344 & ~n7394 ;
  buffer buf_n445( .i (n444), .o (n445) );
  assign n7396 = n1400 & n2611 ;
  assign n7397 = n445 & n7396 ;
  buffer buf_n7398( .i (n7397), .o (n7398) );
  buffer buf_n7399( .i (n7398), .o (n7399) );
  buffer buf_n7400( .i (n7399), .o (n7400) );
  assign n7401 = ( n2209 & n7313 ) | ( n2209 & ~n7347 ) | ( n7313 & ~n7347 ) ;
  buffer buf_n7402( .i (n7026), .o (n7402) );
  assign n7403 = ( ~n2208 & n7013 ) | ( ~n2208 & n7402 ) | ( n7013 & n7402 ) ;
  assign n7404 = ( n6531 & ~n7347 ) | ( n6531 & n7403 ) | ( ~n7347 & n7403 ) ;
  assign n7405 = ~n7401 & n7404 ;
  assign n7406 = n7106 | n7405 ;
  assign n7407 = n3281 | n7348 ;
  assign n7408 = n7106 & n7407 ;
  assign n7409 = n7406 & ~n7408 ;
  assign n7410 = ( ~n6996 & n7398 ) | ( ~n6996 & n7409 ) | ( n7398 & n7409 ) ;
  buffer buf_n7411( .i (n7024), .o (n7411) );
  assign n7412 = ~n7410 & n7411 ;
  assign n7413 = ( n4910 & n7400 ) | ( n4910 & ~n7412 ) | ( n7400 & ~n7412 ) ;
  buffer buf_n7414( .i (n7413), .o (n7414) );
  buffer buf_n7415( .i (n7414), .o (n7415) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  assign n7416 = n1206 & n7414 ;
  buffer buf_n4545( .i (n4544), .o (n4545) );
  buffer buf_n4546( .i (n4545), .o (n4546) );
  buffer buf_n4547( .i (n4546), .o (n4547) );
  assign n7417 = n4547 & ~n6826 ;
  buffer buf_n7418( .i (n7417), .o (n7418) );
  buffer buf_n7419( .i (n7418), .o (n7419) );
  assign n7420 = n792 & n7321 ;
  assign n7421 = ( n2880 & n7353 ) | ( n2880 & ~n7420 ) | ( n7353 & ~n7420 ) ;
  assign n7422 = ( n6776 & ~n7254 ) | ( n6776 & n7421 ) | ( ~n7254 & n7421 ) ;
  buffer buf_n7423( .i (n7422), .o (n7423) );
  assign n7424 = ( n7026 & ~n7034 ) | ( n7026 & n7423 ) | ( ~n7034 & n7423 ) ;
  buffer buf_n7425( .i (n7121), .o (n7425) );
  assign n7426 = ( ~n7054 & n7423 ) | ( ~n7054 & n7425 ) | ( n7423 & n7425 ) ;
  assign n7427 = n7424 | n7426 ;
  buffer buf_n7428( .i (n7427), .o (n7428) );
  buffer buf_n7429( .i (n7428), .o (n7429) );
  buffer buf_n7430( .i (n7429), .o (n7430) );
  buffer buf_n7431( .i (n7132), .o (n7431) );
  buffer buf_n7432( .i (n7431), .o (n7432) );
  assign n7433 = ( n6497 & n7428 ) | ( n6497 & n7432 ) | ( n7428 & n7432 ) ;
  assign n7434 = n7418 & n7433 ;
  assign n7435 = ( ~n7419 & n7430 ) | ( ~n7419 & n7434 ) | ( n7430 & n7434 ) ;
  assign n7436 = n7024 & ~n7435 ;
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n7437( .i (n7170), .o (n7437) );
  assign n7438 = ( n7308 & ~n7425 ) | ( n7308 & n7437 ) | ( ~n7425 & n7437 ) ;
  assign n7439 = n7402 | n7438 ;
  assign n7440 = ~n2284 & n7439 ;
  buffer buf_n7441( .i (n7056), .o (n7441) );
  assign n7442 = ( ~n7432 & n7440 ) | ( ~n7432 & n7441 ) | ( n7440 & n7441 ) ;
  buffer buf_n7443( .i (n6837), .o (n7443) );
  assign n7444 = ( n490 & n919 ) | ( n490 & n7443 ) | ( n919 & n7443 ) ;
  buffer buf_n7445( .i (n7444), .o (n7445) );
  buffer buf_n7446( .i (n7445), .o (n7446) );
  buffer buf_n7447( .i (n7446), .o (n7447) );
  assign n7448 = ( n7425 & ~n7437 ) | ( n7425 & n7445 ) | ( ~n7437 & n7445 ) ;
  assign n7449 = ( n493 & ~n7402 ) | ( n493 & n7448 ) | ( ~n7402 & n7448 ) ;
  assign n7450 = ( ~n494 & n7447 ) | ( ~n494 & n7449 ) | ( n7447 & n7449 ) ;
  assign n7451 = ( n7432 & n7441 ) | ( n7432 & ~n7450 ) | ( n7441 & ~n7450 ) ;
  assign n7452 = n7442 & ~n7451 ;
  buffer buf_n7453( .i (n7353), .o (n7453) );
  assign n7454 = ( n1502 & n7254 ) | ( n1502 & n7453 ) | ( n7254 & n7453 ) ;
  buffer buf_n7455( .i (n7454), .o (n7455) );
  buffer buf_n7456( .i (n7455), .o (n7456) );
  buffer buf_n7457( .i (n7456), .o (n7457) );
  assign n7458 = ( n7308 & n7437 ) | ( n7308 & ~n7455 ) | ( n7437 & ~n7455 ) ;
  assign n7459 = ( n7039 & n7402 ) | ( n7039 & n7458 ) | ( n7402 & n7458 ) ;
  assign n7460 = n7457 & ~n7459 ;
  assign n7461 = ( n7432 & ~n7441 ) | ( n7432 & n7460 ) | ( ~n7441 & n7460 ) ;
  buffer buf_n7462( .i (n7089), .o (n7462) );
  buffer buf_n7463( .i (n7462), .o (n7463) );
  assign n7464 = ( n2256 & n7039 ) | ( n2256 & n7463 ) | ( n7039 & n7463 ) ;
  buffer buf_n7465( .i (n7437), .o (n7465) );
  assign n7466 = ( n2256 & n7463 ) | ( n2256 & n7465 ) | ( n7463 & n7465 ) ;
  assign n7467 = ( n871 & n7464 ) | ( n871 & ~n7466 ) | ( n7464 & ~n7466 ) ;
  buffer buf_n7468( .i (n7431), .o (n7468) );
  assign n7469 = ( n7441 & n7467 ) | ( n7441 & n7468 ) | ( n7467 & n7468 ) ;
  assign n7470 = n7461 & n7469 ;
  assign n7471 = n7452 | n7470 ;
  buffer buf_n7472( .i (n7108), .o (n7472) );
  assign n7473 = n7471 & ~n7472 ;
  assign n7474 = n7436 | n7473 ;
  assign n7475 = ( n6448 & ~n7048 ) | ( n6448 & n7474 ) | ( ~n7048 & n7474 ) ;
  assign n7476 = n394 & n2175 ;
  buffer buf_n7477( .i (n7476), .o (n7477) );
  buffer buf_n7478( .i (n7477), .o (n7478) );
  buffer buf_n7479( .i (n7453), .o (n7479) );
  assign n7480 = n4770 | n7479 ;
  buffer buf_n7481( .i (n7254), .o (n7481) );
  assign n7482 = ( n4770 & n7479 ) | ( n4770 & ~n7481 ) | ( n7479 & ~n7481 ) ;
  assign n7483 = ( n7462 & ~n7480 ) | ( n7462 & n7482 ) | ( ~n7480 & n7482 ) ;
  assign n7484 = n7477 | n7483 ;
  assign n7485 = ( ~n7040 & n7478 ) | ( ~n7040 & n7484 ) | ( n7478 & n7484 ) ;
  assign n7486 = n7212 | n7485 ;
  buffer buf_n7487( .i (n7354), .o (n7487) );
  assign n7488 = n1121 & ~n7487 ;
  buffer buf_n7489( .i (n7488), .o (n7489) );
  buffer buf_n7490( .i (n7489), .o (n7490) );
  buffer buf_n7491( .i (n7067), .o (n7491) );
  assign n7492 = ( n7131 & ~n7489 ) | ( n7131 & n7491 ) | ( ~n7489 & n7491 ) ;
  assign n7493 = ( n1124 & n7490 ) | ( n1124 & ~n7492 ) | ( n7490 & ~n7492 ) ;
  assign n7494 = n7313 & n7493 ;
  buffer buf_n7495( .i (n7211), .o (n7495) );
  assign n7496 = ~n7494 & n7495 ;
  assign n7497 = n7486 & ~n7496 ;
  buffer buf_n7498( .i (n6644), .o (n7498) );
  buffer buf_n7499( .i (n7498), .o (n7499) );
  assign n7500 = ( n4769 & ~n7453 ) | ( n4769 & n7499 ) | ( ~n7453 & n7499 ) ;
  buffer buf_n7501( .i (n7500), .o (n7501) );
  assign n7504 = n7131 & ~n7501 ;
  buffer buf_n7505( .i (n7504), .o (n7505) );
  buffer buf_n7506( .i (n7505), .o (n7506) );
  buffer buf_n7502( .i (n7501), .o (n7502) );
  buffer buf_n7503( .i (n7502), .o (n7503) );
  assign n7507 = n7503 | n7505 ;
  assign n7508 = ( ~n7468 & n7506 ) | ( ~n7468 & n7507 ) | ( n7506 & n7507 ) ;
  assign n7509 = ( n7219 & ~n7297 ) | ( n7219 & n7508 ) | ( ~n7297 & n7508 ) ;
  assign n7510 = ( ~n5083 & n7497 ) | ( ~n5083 & n7509 ) | ( n7497 & n7509 ) ;
  assign n7511 = ~n6493 & n7510 ;
  assign n7512 = ( n5255 & ~n7425 ) | ( n5255 & n7491 ) | ( ~n7425 & n7491 ) ;
  assign n7513 = ~n5254 & n7142 ;
  assign n7514 = ( ~n5255 & n7462 ) | ( ~n5255 & n7513 ) | ( n7462 & n7513 ) ;
  assign n7515 = n7512 & ~n7514 ;
  buffer buf_n7516( .i (n7308), .o (n7516) );
  buffer buf_n7517( .i (n7516), .o (n7517) );
  assign n7518 = n7515 | n7517 ;
  assign n7519 = n5041 | n7121 ;
  assign n7520 = ( n5042 & ~n6923 ) | ( n5042 & n7519 ) | ( ~n6923 & n7519 ) ;
  assign n7521 = n7055 & ~n7520 ;
  assign n7522 = n7517 & ~n7521 ;
  assign n7523 = n7518 & ~n7522 ;
  assign n7524 = n7333 & n7523 ;
  assign n7525 = n1256 & n7331 ;
  buffer buf_n7526( .i (n610), .o (n7526) );
  assign n7527 = n7525 & n7526 ;
  assign n7528 = n7524 | n7527 ;
  buffer buf_n7529( .i (n7465), .o (n7529) );
  buffer buf_n7530( .i (n7529), .o (n7530) );
  buffer buf_n7531( .i (n7530), .o (n7531) );
  buffer buf_n7532( .i (n7531), .o (n7532) );
  buffer buf_n7533( .i (n7532), .o (n7533) );
  assign n7534 = n7528 & n7533 ;
  assign n7535 = n7511 | n7534 ;
  buffer buf_n7536( .i (n6540), .o (n7536) );
  assign n7537 = ( n7048 & ~n7535 ) | ( n7048 & n7536 ) | ( ~n7535 & n7536 ) ;
  assign n7538 = n7475 & ~n7537 ;
  assign n7539 = ( n6779 & n7323 ) | ( n6779 & ~n7453 ) | ( n7323 & ~n7453 ) ;
  buffer buf_n7540( .i (n7539), .o (n7540) );
  buffer buf_n7541( .i (n7540), .o (n7541) );
  buffer buf_n7542( .i (n7541), .o (n7542) );
  buffer buf_n7543( .i (n7542), .o (n7543) );
  buffer buf_n7544( .i (n7142), .o (n7544) );
  buffer buf_n7545( .i (n6752), .o (n7545) );
  assign n7546 = ( n7540 & n7544 ) | ( n7540 & n7545 ) | ( n7544 & n7545 ) ;
  buffer buf_n7547( .i (n7546), .o (n7547) );
  buffer buf_n7548( .i (n7547), .o (n7548) );
  assign n7549 = n7327 & ~n7547 ;
  assign n7550 = ( n7543 & ~n7548 ) | ( n7543 & n7549 ) | ( ~n7548 & n7549 ) ;
  buffer buf_n7551( .i (n7550), .o (n7551) );
  buffer buf_n7552( .i (n7551), .o (n7552) );
  buffer buf_n4385( .i (n4384), .o (n4385) );
  buffer buf_n4386( .i (n4385), .o (n4386) );
  buffer buf_n4387( .i (n4386), .o (n4387) );
  buffer buf_n7553( .i (n7106), .o (n7553) );
  assign n7554 = ( n4387 & n7551 ) | ( n4387 & n7553 ) | ( n7551 & n7553 ) ;
  assign n7555 = n7552 & ~n7554 ;
  buffer buf_n7556( .i (n7555), .o (n7556) );
  buffer buf_n7557( .i (n7556), .o (n7557) );
  buffer buf_n7558( .i (n7499), .o (n7558) );
  assign n7559 = ( n7067 & n7479 ) | ( n7067 & n7558 ) | ( n7479 & n7558 ) ;
  buffer buf_n7560( .i (n7559), .o (n7560) );
  assign n7561 = ( n7055 & n7463 ) | ( n7055 & ~n7560 ) | ( n7463 & ~n7560 ) ;
  assign n7562 = ( n7463 & ~n7516 ) | ( n7463 & n7560 ) | ( ~n7516 & n7560 ) ;
  assign n7563 = ~n7561 & n7562 ;
  assign n7564 = n7495 & ~n7563 ;
  assign n7565 = n4118 & ~n7056 ;
  assign n7566 = n7495 | n7565 ;
  assign n7567 = ~n7564 & n7566 ;
  buffer buf_n7568( .i (n7567), .o (n7568) );
  buffer buf_n7569( .i (n7568), .o (n7569) );
  assign n7570 = ( n5701 & ~n7305 ) | ( n5701 & n7568 ) | ( ~n7305 & n7568 ) ;
  assign n7571 = n278 & ~n7468 ;
  buffer buf_n7572( .i (n7056), .o (n7572) );
  buffer buf_n7573( .i (n7572), .o (n7573) );
  assign n7574 = ( n7297 & n7571 ) | ( n7297 & n7573 ) | ( n7571 & n7573 ) ;
  assign n7575 = ~n7108 & n7574 ;
  assign n7576 = n7305 & n7575 ;
  assign n7577 = ( n7569 & ~n7570 ) | ( n7569 & n7576 ) | ( ~n7570 & n7576 ) ;
  assign n7578 = n279 & n712 ;
  assign n7579 = ( n6684 & n7370 ) | ( n6684 & n7578 ) | ( n7370 & n7578 ) ;
  assign n7580 = ~n5783 & n7579 ;
  buffer buf_n7581( .i (n7580), .o (n7581) );
  assign n7582 = ( ~n7556 & n7577 ) | ( ~n7556 & n7581 ) | ( n7577 & n7581 ) ;
  buffer buf_n7583( .i (n6635), .o (n7583) );
  assign n7584 = ~n7581 & n7583 ;
  assign n7585 = ( n7557 & n7582 ) | ( n7557 & ~n7584 ) | ( n7582 & ~n7584 ) ;
  assign n7586 = n7538 | n7585 ;
  assign n7587 = ( n7415 & ~n7416 ) | ( n7415 & n7586 ) | ( ~n7416 & n7586 ) ;
  assign n7588 = n7395 | n7587 ;
  assign n7589 = ( ~n7242 & n7278 ) | ( ~n7242 & n7588 ) | ( n7278 & n7588 ) ;
  assign n7590 = n7243 | n7589 ;
  buffer buf_n6076( .i (n6075), .o (n6076) );
  buffer buf_n6077( .i (n6076), .o (n6077) );
  buffer buf_n6078( .i (n6077), .o (n6078) );
  buffer buf_n6079( .i (n6078), .o (n6079) );
  buffer buf_n6080( .i (n6079), .o (n6080) );
  buffer buf_n6081( .i (n6080), .o (n6081) );
  buffer buf_n6082( .i (n6081), .o (n6082) );
  buffer buf_n6083( .i (n6082), .o (n6083) );
  buffer buf_n6084( .i (n6083), .o (n6084) );
  buffer buf_n6085( .i (n6084), .o (n6085) );
  assign n7591 = n1971 & ~n7529 ;
  buffer buf_n7592( .i (n7591), .o (n7592) );
  buffer buf_n7593( .i (n7592), .o (n7593) );
  buffer buf_n7594( .i (n7495), .o (n7594) );
  assign n7595 = ( ~n7573 & n7592 ) | ( ~n7573 & n7594 ) | ( n7592 & n7594 ) ;
  assign n7596 = ( n1974 & n7593 ) | ( n1974 & n7595 ) | ( n7593 & n7595 ) ;
  buffer buf_n7597( .i (n7304), .o (n7597) );
  assign n7598 = n7596 & n7597 ;
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n4174( .i (n4173), .o (n4174) );
  buffer buf_n4175( .i (n4174), .o (n4175) );
  buffer buf_n4176( .i (n4175), .o (n4176) );
  buffer buf_n4177( .i (n4176), .o (n4177) );
  buffer buf_n4178( .i (n4177), .o (n4178) );
  buffer buf_n4179( .i (n4178), .o (n4179) );
  buffer buf_n4180( .i (n4179), .o (n4180) );
  buffer buf_n4181( .i (n4180), .o (n4181) );
  buffer buf_n7599( .i (n7211), .o (n7599) );
  assign n7600 = ( n4179 & n7468 ) | ( n4179 & ~n7599 ) | ( n7468 & ~n7599 ) ;
  assign n7601 = ( n7531 & n7594 ) | ( n7531 & ~n7600 ) | ( n7594 & ~n7600 ) ;
  assign n7602 = ( n446 & n4181 ) | ( n446 & ~n7601 ) | ( n4181 & ~n7601 ) ;
  assign n7603 = n7597 | n7602 ;
  assign n7604 = ( ~n6540 & n7598 ) | ( ~n6540 & n7603 ) | ( n7598 & n7603 ) ;
  assign n7605 = n6208 & ~n7604 ;
  assign n7606 = n7348 | n7530 ;
  buffer buf_n7607( .i (n7606), .o (n7607) );
  assign n7608 = ( n7532 & n7553 ) | ( n7532 & ~n7607 ) | ( n7553 & ~n7607 ) ;
  assign n7609 = ( n7108 & n7553 ) | ( n7108 & ~n7607 ) | ( n7553 & ~n7607 ) ;
  assign n7610 = ( n960 & n7608 ) | ( n960 & ~n7609 ) | ( n7608 & ~n7609 ) ;
  assign n7611 = ~n7184 & n7610 ;
  buffer buf_n7612( .i (n6202), .o (n7612) );
  assign n7613 = n7611 | n7612 ;
  assign n7614 = ~n7605 & n7613 ;
  assign n7615 = ( n5857 & ~n6085 ) | ( n5857 & n7614 ) | ( ~n6085 & n7614 ) ;
  buffer buf_n6513( .i (n6512), .o (n6513) );
  buffer buf_n6514( .i (n6513), .o (n6514) );
  buffer buf_n6515( .i (n6514), .o (n6515) );
  buffer buf_n6516( .i (n6515), .o (n6516) );
  assign n7616 = n6516 & n7222 ;
  assign n7617 = ( ~n6488 & n6516 ) | ( ~n6488 & n7222 ) | ( n6516 & n7222 ) ;
  assign n7618 = ( n6259 & ~n7616 ) | ( n6259 & n7617 ) | ( ~n7616 & n7617 ) ;
  assign n7619 = n7536 | n7618 ;
  buffer buf_n7620( .i (n7411), .o (n7620) );
  buffer buf_n7621( .i (n7620), .o (n7621) );
  assign n7622 = n7619 | n7621 ;
  buffer buf_n7623( .i (n7238), .o (n7623) );
  assign n7624 = ( n6085 & n7622 ) | ( n6085 & n7623 ) | ( n7622 & n7623 ) ;
  assign n7625 = n7615 & ~n7624 ;
  buffer buf_n7626( .i (n7625), .o (n7626) );
  buffer buf_n7627( .i (n7626), .o (n7627) );
  buffer buf_n2677( .i (n2676), .o (n2677) );
  buffer buf_n2934( .i (n2933), .o (n2934) );
  buffer buf_n2935( .i (n2934), .o (n2935) );
  assign n7628 = ( n2676 & n2935 ) | ( n2676 & n7304 ) | ( n2935 & n7304 ) ;
  assign n7629 = ~n2677 & n7628 ;
  buffer buf_n7630( .i (n7629), .o (n7630) );
  buffer buf_n7631( .i (n7630), .o (n7631) );
  buffer buf_n5159( .i (n5158), .o (n5159) );
  assign n7632 = n5159 & ~n7553 ;
  assign n7633 = ( n7472 & n7597 ) | ( n7472 & n7632 ) | ( n7597 & n7632 ) ;
  buffer buf_n7634( .i (n7597), .o (n7634) );
  assign n7635 = n7633 & ~n7634 ;
  assign n7636 = n1402 & ~n1509 ;
  assign n7637 = n401 & n7636 ;
  buffer buf_n7638( .i (n7637), .o (n7638) );
  assign n7639 = ( ~n7630 & n7635 ) | ( ~n7630 & n7638 ) | ( n7635 & n7638 ) ;
  assign n7640 = n7583 & ~n7638 ;
  assign n7641 = ( n7631 & n7639 ) | ( n7631 & ~n7640 ) | ( n7639 & ~n7640 ) ;
  buffer buf_n7642( .i (n7641), .o (n7642) );
  buffer buf_n7643( .i (n7642), .o (n7643) );
  assign n7644 = n2710 & n7642 ;
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n5959( .i (n5958), .o (n5959) );
  buffer buf_n5960( .i (n5959), .o (n5960) );
  buffer buf_n5961( .i (n5960), .o (n5961) );
  buffer buf_n5962( .i (n5961), .o (n5962) );
  buffer buf_n5963( .i (n5962), .o (n5963) );
  buffer buf_n5964( .i (n5963), .o (n5964) );
  buffer buf_n5965( .i (n5964), .o (n5965) );
  buffer buf_n5966( .i (n5965), .o (n5966) );
  buffer buf_n5967( .i (n5966), .o (n5967) );
  buffer buf_n5968( .i (n5967), .o (n5968) );
  assign n7645 = ( ~n717 & n805 ) | ( ~n717 & n5968 ) | ( n805 & n5968 ) ;
  assign n7646 = n718 & n7645 ;
  buffer buf_n4131( .i (n4130), .o (n4131) );
  buffer buf_n4132( .i (n4131), .o (n4132) );
  buffer buf_n4133( .i (n4132), .o (n4133) );
  buffer buf_n4134( .i (n4133), .o (n4134) );
  assign n7647 = ( n5943 & n7003 ) | ( n5943 & n7353 ) | ( n7003 & n7353 ) ;
  buffer buf_n7648( .i (n7647), .o (n7648) );
  buffer buf_n7649( .i (n7141), .o (n7649) );
  assign n7650 = ( n7481 & ~n7648 ) | ( n7481 & n7649 ) | ( ~n7648 & n7649 ) ;
  assign n7651 = ( ~n7121 & n7481 ) | ( ~n7121 & n7648 ) | ( n7481 & n7648 ) ;
  assign n7652 = ~n7650 & n7651 ;
  assign n7653 = n7346 | n7652 ;
  assign n7654 = n2176 & n7544 ;
  assign n7655 = n7346 & ~n7654 ;
  assign n7656 = n7653 & ~n7655 ;
  buffer buf_n7657( .i (n7431), .o (n7657) );
  assign n7658 = n7656 & n7657 ;
  buffer buf_n7659( .i (n7658), .o (n7659) );
  buffer buf_n7660( .i (n7659), .o (n7660) );
  buffer buf_n7661( .i (n7517), .o (n7661) );
  assign n7662 = ( n349 & ~n2006 ) | ( n349 & n7661 ) | ( ~n2006 & n7661 ) ;
  assign n7663 = n350 & ~n7662 ;
  assign n7664 = n7659 | n7663 ;
  buffer buf_n7665( .i (n7304), .o (n7665) );
  assign n7666 = ( n7660 & n7664 ) | ( n7660 & n7665 ) | ( n7664 & n7665 ) ;
  assign n7667 = ~n4134 & n7666 ;
  buffer buf_n7668( .i (n7667), .o (n7668) );
  buffer buf_n7669( .i (n7668), .o (n7669) );
  buffer buf_n3266( .i (n3265), .o (n3266) );
  assign n7670 = ~n3263 & n7443 ;
  buffer buf_n7671( .i (n7670), .o (n7671) );
  buffer buf_n7672( .i (n7671), .o (n7672) );
  assign n7673 = ( ~n7491 & n7545 ) | ( ~n7491 & n7671 ) | ( n7545 & n7671 ) ;
  assign n7674 = ( ~n3266 & n7672 ) | ( ~n3266 & n7673 ) | ( n7672 & n7673 ) ;
  assign n7675 = n7040 & n7674 ;
  assign n7676 = ( n1045 & n7067 ) | ( n1045 & ~n7558 ) | ( n7067 & ~n7558 ) ;
  buffer buf_n7677( .i (n7170), .o (n7677) );
  assign n7678 = ( n395 & n7676 ) | ( n395 & ~n7677 ) | ( n7676 & ~n7677 ) ;
  assign n7679 = ( ~n4502 & n7465 ) | ( ~n4502 & n7678 ) | ( n7465 & n7678 ) ;
  assign n7680 = ~n7040 & n7679 ;
  buffer buf_n7681( .i (n7039), .o (n7681) );
  buffer buf_n7682( .i (n7681), .o (n7682) );
  assign n7683 = ( ~n7675 & n7680 ) | ( ~n7675 & n7682 ) | ( n7680 & n7682 ) ;
  assign n7684 = n7594 | n7683 ;
  assign n7685 = n922 & ~n7465 ;
  assign n7686 = n564 & n7685 ;
  assign n7687 = n397 & n1142 ;
  assign n7688 = n7686 | n7687 ;
  assign n7689 = n7594 & n7688 ;
  assign n7690 = n7684 & ~n7689 ;
  assign n7691 = ( ~n5783 & n7665 ) | ( ~n5783 & n7690 ) | ( n7665 & n7690 ) ;
  buffer buf_n1144( .i (n1143), .o (n1144) );
  assign n7692 = n406 & ~n1144 ;
  assign n7693 = ( n1861 & n7247 ) | ( n1861 & n7280 ) | ( n7247 & n7280 ) ;
  buffer buf_n7694( .i (n7693), .o (n7694) );
  buffer buf_n7695( .i (n7694), .o (n7695) );
  buffer buf_n7696( .i (n7695), .o (n7696) );
  buffer buf_n7697( .i (n7003), .o (n7697) );
  assign n7698 = ( n7487 & ~n7694 ) | ( n7487 & n7697 ) | ( ~n7694 & n7697 ) ;
  assign n7699 = n1864 & n7698 ;
  assign n7700 = ( n7491 & ~n7696 ) | ( n7491 & n7699 ) | ( ~n7696 & n7699 ) ;
  buffer buf_n7701( .i (n7700), .o (n7701) );
  buffer buf_n7702( .i (n7701), .o (n7702) );
  assign n7703 = ( n7431 & n7529 ) | ( n7431 & n7701 ) | ( n7529 & n7701 ) ;
  buffer buf_n7704( .i (n6865), .o (n7704) );
  buffer buf_n7705( .i (n7704), .o (n7705) );
  buffer buf_n7706( .i (n7705), .o (n7706) );
  assign n7707 = ( ~n346 & n1080 ) | ( ~n346 & n7706 ) | ( n1080 & n7706 ) ;
  assign n7708 = n347 & n7707 ;
  assign n7709 = ~n7529 & n7708 ;
  assign n7710 = ( n7702 & ~n7703 ) | ( n7702 & n7709 ) | ( ~n7703 & n7709 ) ;
  assign n7711 = ~n425 & n7544 ;
  buffer buf_n7712( .i (n7711), .o (n7712) );
  assign n7713 = n1307 & n7712 ;
  assign n7714 = ( n290 & ~n427 ) | ( n290 & n7712 ) | ( ~n427 & n7712 ) ;
  assign n7715 = ( n7572 & n7713 ) | ( n7572 & n7714 ) | ( n7713 & n7714 ) ;
  assign n7716 = n7710 | n7715 ;
  assign n7717 = ( n407 & ~n7692 ) | ( n407 & n7716 ) | ( ~n7692 & n7716 ) ;
  buffer buf_n7718( .i (n6684), .o (n7718) );
  assign n7719 = ( n7665 & n7717 ) | ( n7665 & n7718 ) | ( n7717 & n7718 ) ;
  assign n7720 = ~n7691 & n7719 ;
  assign n7721 = ~n1137 & n7347 ;
  buffer buf_n7722( .i (n7346), .o (n7722) );
  assign n7723 = n1543 | n7722 ;
  assign n7724 = ~n7721 & n7723 ;
  assign n7725 = n7333 & ~n7724 ;
  buffer buf_n7726( .i (n7443), .o (n7726) );
  assign n7727 = ( n1175 & n7705 ) | ( n1175 & n7726 ) | ( n7705 & n7726 ) ;
  buffer buf_n7728( .i (n7727), .o (n7728) );
  buffer buf_n7729( .i (n7728), .o (n7729) );
  assign n7730 = n1170 & ~n7728 ;
  assign n7731 = ( n1178 & ~n7729 ) | ( n1178 & n7730 ) | ( ~n7729 & n7730 ) ;
  assign n7732 = ~n7348 & n7731 ;
  buffer buf_n7733( .i (n7657), .o (n7733) );
  assign n7734 = n7732 | n7733 ;
  assign n7735 = ~n7725 & n7734 ;
  assign n7736 = ( n7472 & ~n7718 ) | ( n7472 & n7735 ) | ( ~n7718 & n7735 ) ;
  buffer buf_n7737( .i (n4656), .o (n7737) );
  assign n7738 = ( n2067 & ~n7280 ) | ( n2067 & n7737 ) | ( ~n7280 & n7737 ) ;
  buffer buf_n7739( .i (n7738), .o (n7739) );
  assign n7742 = n7499 & ~n7739 ;
  buffer buf_n7743( .i (n7742), .o (n7743) );
  buffer buf_n7744( .i (n7743), .o (n7744) );
  buffer buf_n7740( .i (n7739), .o (n7740) );
  buffer buf_n7741( .i (n7740), .o (n7741) );
  assign n7745 = n7741 | n7743 ;
  assign n7746 = ( ~n7132 & n7744 ) | ( ~n7132 & n7745 ) | ( n7744 & n7745 ) ;
  assign n7747 = n7722 & ~n7746 ;
  buffer buf_n7748( .i (n7545), .o (n7748) );
  assign n7749 = n1213 & ~n7748 ;
  assign n7750 = n7722 | n7749 ;
  assign n7751 = ~n7747 & n7750 ;
  assign n7752 = n7573 | n7751 ;
  buffer buf_n6860( .i (n6859), .o (n6860) );
  buffer buf_n6861( .i (n6860), .o (n6861) );
  buffer buf_n6862( .i (n6861), .o (n6862) );
  buffer buf_n6863( .i (n6862), .o (n6863) );
  buffer buf_n6864( .i (n6863), .o (n6864) );
  buffer buf_n7753( .i (n7260), .o (n7753) );
  buffer buf_n7754( .i (n7462), .o (n7754) );
  assign n7755 = ( n7748 & ~n7753 ) | ( n7748 & n7754 ) | ( ~n7753 & n7754 ) ;
  assign n7756 = n6864 & n7755 ;
  assign n7757 = ~n7530 & n7756 ;
  assign n7758 = n7573 & ~n7757 ;
  assign n7759 = n7752 & ~n7758 ;
  assign n7760 = ( n7472 & n7718 ) | ( n7472 & ~n7759 ) | ( n7718 & ~n7759 ) ;
  assign n7761 = n7736 & ~n7760 ;
  assign n7762 = ( ~n7583 & n7720 ) | ( ~n7583 & n7761 ) | ( n7720 & n7761 ) ;
  assign n7763 = ~n7668 & n7762 ;
  assign n7764 = ( ~n7623 & n7669 ) | ( ~n7623 & n7763 ) | ( n7669 & n7763 ) ;
  assign n7765 = n7646 | n7764 ;
  assign n7766 = ( n7643 & ~n7644 ) | ( n7643 & n7765 ) | ( ~n7644 & n7765 ) ;
  buffer buf_n4081( .i (n4080), .o (n4081) );
  buffer buf_n7767( .i (n7722), .o (n7767) );
  assign n7768 = ( ~n588 & n4081 ) | ( ~n588 & n7767 ) | ( n4081 & n7767 ) ;
  assign n7769 = ~n7303 & n7768 ;
  buffer buf_n7770( .i (n7769), .o (n7770) );
  buffer buf_n7771( .i (n7770), .o (n7771) );
  buffer buf_n7772( .i (n7771), .o (n7772) );
  buffer buf_n5094( .i (n5093), .o (n5094) );
  buffer buf_n5095( .i (n5094), .o (n5095) );
  buffer buf_n5096( .i (n5095), .o (n5096) );
  buffer buf_n7773( .i (n7572), .o (n7773) );
  assign n7774 = ( n5096 & n7531 ) | ( n5096 & ~n7773 ) | ( n7531 & ~n7773 ) ;
  assign n7775 = ( n5095 & ~n7530 ) | ( n5095 & n7767 ) | ( ~n7530 & n7767 ) ;
  assign n7776 = ( ~n7192 & n7773 ) | ( ~n7192 & n7775 ) | ( n7773 & n7775 ) ;
  assign n7777 = n7774 | n7776 ;
  buffer buf_n7778( .i (n7599), .o (n7778) );
  buffer buf_n7779( .i (n7778), .o (n7779) );
  buffer buf_n7780( .i (n7779), .o (n7780) );
  assign n7781 = ( n7770 & ~n7777 ) | ( n7770 & n7780 ) | ( ~n7777 & n7780 ) ;
  assign n7782 = n7184 & ~n7781 ;
  assign n7783 = ( n7087 & n7772 ) | ( n7087 & ~n7782 ) | ( n7772 & ~n7782 ) ;
  buffer buf_n7784( .i (n7783), .o (n7784) );
  buffer buf_n7785( .i (n7784), .o (n7785) );
  assign n7786 = ( n356 & n7623 ) | ( n356 & n7784 ) | ( n7623 & n7784 ) ;
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  assign n7787 = ( n1411 & n6206 ) | ( n1411 & n7159 ) | ( n6206 & n7159 ) ;
  assign n7788 = ~n7160 & n7787 ;
  assign n7789 = ~n356 & n7788 ;
  assign n7790 = ( n7785 & ~n7786 ) | ( n7785 & n7789 ) | ( ~n7786 & n7789 ) ;
  buffer buf_n7791( .i (n6759), .o (n7791) );
  buffer buf_n7792( .i (n7279), .o (n7792) );
  assign n7793 = ( ~n7737 & n7791 ) | ( ~n7737 & n7792 ) | ( n7791 & n7792 ) ;
  buffer buf_n7794( .i (n7793), .o (n7794) );
  assign n7799 = ( n3920 & n7487 ) | ( n3920 & ~n7794 ) | ( n7487 & ~n7794 ) ;
  buffer buf_n7800( .i (n7799), .o (n7800) );
  buffer buf_n7801( .i (n7800), .o (n7801) );
  buffer buf_n7802( .i (n7801), .o (n7802) );
  buffer buf_n7803( .i (n7802), .o (n7803) );
  buffer buf_n7804( .i (n7697), .o (n7804) );
  buffer buf_n7805( .i (n7804), .o (n7805) );
  assign n7806 = ( n7545 & n7800 ) | ( n7545 & ~n7805 ) | ( n7800 & ~n7805 ) ;
  buffer buf_n7807( .i (n7806), .o (n7807) );
  buffer buf_n7808( .i (n7807), .o (n7808) );
  buffer buf_n7795( .i (n7794), .o (n7795) );
  buffer buf_n7796( .i (n7795), .o (n7796) );
  buffer buf_n7797( .i (n7796), .o (n7797) );
  buffer buf_n7798( .i (n7797), .o (n7798) );
  assign n7809 = n7798 & n7807 ;
  assign n7810 = ( ~n7803 & n7808 ) | ( ~n7803 & n7809 ) | ( n7808 & n7809 ) ;
  buffer buf_n7811( .i (n7767), .o (n7811) );
  assign n7812 = n7810 | n7811 ;
  assign n7813 = ~n1330 & n7748 ;
  assign n7814 = ( ~n1331 & n7681 ) | ( ~n1331 & n7813 ) | ( n7681 & n7813 ) ;
  buffer buf_n7815( .i (n6910), .o (n7815) );
  assign n7816 = n7814 & ~n7815 ;
  assign n7817 = n7811 & ~n7816 ;
  assign n7818 = n7812 & ~n7817 ;
  assign n7819 = n7780 | n7818 ;
  assign n7820 = ( ~n7018 & n7657 ) | ( ~n7018 & n7682 ) | ( n7657 & n7682 ) ;
  assign n7821 = ( n7018 & n7682 ) | ( n7018 & ~n7767 ) | ( n7682 & ~n7767 ) ;
  assign n7822 = n7820 | n7821 ;
  assign n7823 = n7268 | n7822 ;
  assign n7824 = n7780 & n7823 ;
  assign n7825 = n7819 & ~n7824 ;
  assign n7826 = n6196 | n7825 ;
  buffer buf_n7827( .i (n7558), .o (n7827) );
  assign n7828 = ( ~n3961 & n7805 ) | ( ~n3961 & n7827 ) | ( n7805 & n7827 ) ;
  buffer buf_n7829( .i (n7828), .o (n7829) );
  buffer buf_n7830( .i (n7829), .o (n7830) );
  buffer buf_n7831( .i (n7830), .o (n7831) );
  buffer buf_n7832( .i (n7831), .o (n7832) );
  buffer buf_n7833( .i (n7753), .o (n7833) );
  assign n7834 = ( n7211 & ~n7829 ) | ( n7211 & n7833 ) | ( ~n7829 & n7833 ) ;
  buffer buf_n7835( .i (n7834), .o (n7835) );
  buffer buf_n7836( .i (n7835), .o (n7836) );
  assign n7837 = ~n3965 & n7835 ;
  assign n7838 = ( n7832 & n7836 ) | ( n7832 & n7837 ) | ( n7836 & n7837 ) ;
  buffer buf_n7839( .i (n7748), .o (n7839) );
  assign n7840 = n923 & n7839 ;
  buffer buf_n7841( .i (n311), .o (n7841) );
  assign n7842 = n7840 & ~n7841 ;
  buffer buf_n7843( .i (n7842), .o (n7843) );
  buffer buf_n7844( .i (n7843), .o (n7844) );
  assign n7845 = n6774 & ~n7843 ;
  assign n7846 = ( n7838 & n7844 ) | ( n7838 & ~n7845 ) | ( n7844 & ~n7845 ) ;
  buffer buf_n7847( .i (n6996), .o (n7847) );
  assign n7848 = n7846 & ~n7847 ;
  assign n7849 = n6196 & ~n7848 ;
  assign n7850 = n7826 & ~n7849 ;
  assign n7851 = n7161 & n7850 ;
  assign n7852 = ~n340 & n570 ;
  assign n7853 = ( n3920 & n7374 ) | ( n3920 & ~n7499 ) | ( n7374 & ~n7499 ) ;
  buffer buf_n7854( .i (n7853), .o (n7854) );
  buffer buf_n7855( .i (n7854), .o (n7855) );
  buffer buf_n7856( .i (n7855), .o (n7856) );
  buffer buf_n7857( .i (n7856), .o (n7857) );
  buffer buf_n7858( .i (n6751), .o (n7858) );
  assign n7859 = ~n7854 & n7858 ;
  buffer buf_n7860( .i (n7859), .o (n7860) );
  buffer buf_n7861( .i (n7860), .o (n7861) );
  assign n7862 = ( ~n7017 & n7833 ) | ( ~n7017 & n7860 ) | ( n7833 & n7860 ) ;
  assign n7863 = ( ~n7857 & n7861 ) | ( ~n7857 & n7862 ) | ( n7861 & n7862 ) ;
  assign n7864 = ( n7219 & n7773 ) | ( n7219 & n7863 ) | ( n7773 & n7863 ) ;
  assign n7865 = ( n727 & n4487 ) | ( n727 & n7839 ) | ( n4487 & n7839 ) ;
  assign n7866 = ~n7657 & n7865 ;
  assign n7867 = n7219 & n7866 ;
  buffer buf_n7868( .i (n7773), .o (n7868) );
  assign n7869 = ( n7864 & n7867 ) | ( n7864 & ~n7868 ) | ( n7867 & ~n7868 ) ;
  assign n7870 = ~n7780 & n7869 ;
  buffer buf_n7871( .i (n7870), .o (n7871) );
  buffer buf_n7872( .i (n7871), .o (n7872) );
  assign n7873 = n757 | n7871 ;
  assign n7874 = ( n7852 & n7872 ) | ( n7852 & n7873 ) | ( n7872 & n7873 ) ;
  assign n7875 = n7161 | n7874 ;
  assign n7876 = ( ~n209 & n7851 ) | ( ~n209 & n7875 ) | ( n7851 & n7875 ) ;
  assign n7877 = n7790 | n7876 ;
  assign n7878 = ( ~n7626 & n7766 ) | ( ~n7626 & n7877 ) | ( n7766 & n7877 ) ;
  assign n7879 = n7627 | n7878 ;
  assign n7880 = n7267 & ~n7778 ;
  assign n7881 = ( n4861 & ~n7267 ) | ( n4861 & n7778 ) | ( ~n7267 & n7778 ) ;
  assign n7882 = n4861 & n7811 ;
  assign n7883 = ( n7880 & n7881 ) | ( n7880 & ~n7882 ) | ( n7881 & ~n7882 ) ;
  assign n7884 = ~n4731 & n7883 ;
  buffer buf_n7885( .i (n7884), .o (n7885) );
  buffer buf_n7886( .i (n7885), .o (n7886) );
  buffer buf_n3706( .i (n3705), .o (n3706) );
  buffer buf_n3707( .i (n3706), .o (n3707) );
  buffer buf_n3708( .i (n3707), .o (n3708) );
  buffer buf_n3709( .i (n3708), .o (n3709) );
  buffer buf_n3710( .i (n3709), .o (n3710) );
  buffer buf_n3711( .i (n3710), .o (n3711) );
  buffer buf_n3712( .i (n3711), .o (n3712) );
  buffer buf_n3713( .i (n3712), .o (n3713) );
  buffer buf_n4862( .i (n4861), .o (n4862) );
  buffer buf_n4863( .i (n4862), .o (n4863) );
  buffer buf_n4864( .i (n4863), .o (n4864) );
  assign n7887 = n3713 & n4864 ;
  assign n7888 = n7885 | n7887 ;
  assign n7889 = ( ~n7238 & n7886 ) | ( ~n7238 & n7888 ) | ( n7886 & n7888 ) ;
  assign n7890 = n7229 | n7889 ;
  buffer buf_n3714( .i (n3713), .o (n3714) );
  buffer buf_n7891( .i (n7754), .o (n7891) );
  buffer buf_n7892( .i (n7891), .o (n7892) );
  buffer buf_n7893( .i (n7892), .o (n7893) );
  buffer buf_n7894( .i (n7893), .o (n7894) );
  assign n7895 = n3711 & ~n7894 ;
  buffer buf_n7896( .i (n7895), .o (n7896) );
  buffer buf_n7897( .i (n7896), .o (n7897) );
  assign n7898 = ( ~n7411 & n7634 ) | ( ~n7411 & n7896 ) | ( n7634 & n7896 ) ;
  assign n7899 = ( n3714 & n7897 ) | ( n3714 & n7898 ) | ( n7897 & n7898 ) ;
  buffer buf_n7900( .i (n7583), .o (n7900) );
  assign n7901 = n7899 & ~n7900 ;
  buffer buf_n7902( .i (n7228), .o (n7902) );
  assign n7903 = ~n7901 & n7902 ;
  assign n7904 = n7890 & ~n7903 ;
  buffer buf_n7905( .i (n7904), .o (n7905) );
  buffer buf_n7906( .i (n7905), .o (n7906) );
  buffer buf_n2678( .i (n2677), .o (n2678) );
  buffer buf_n2679( .i (n2678), .o (n2679) );
  buffer buf_n2680( .i (n2679), .o (n2680) );
  buffer buf_n2681( .i (n2680), .o (n2681) );
  buffer buf_n2682( .i (n2681), .o (n2682) );
  buffer buf_n2683( .i (n2682), .o (n2683) );
  buffer buf_n2684( .i (n2683), .o (n2684) );
  assign n7907 = n2684 & n7905 ;
  buffer buf_n4281( .i (n4280), .o (n4281) );
  buffer buf_n4282( .i (n4281), .o (n4282) );
  buffer buf_n4283( .i (n4282), .o (n4283) );
  buffer buf_n4284( .i (n4283), .o (n4284) );
  buffer buf_n4285( .i (n4284), .o (n4285) );
  buffer buf_n4286( .i (n4285), .o (n4286) );
  buffer buf_n4287( .i (n4286), .o (n4287) );
  buffer buf_n4288( .i (n4287), .o (n4288) );
  buffer buf_n4289( .i (n4288), .o (n4289) );
  buffer buf_n4290( .i (n4289), .o (n4290) );
  buffer buf_n5815( .i (n5814), .o (n5815) );
  buffer buf_n5816( .i (n5815), .o (n5816) );
  buffer buf_n5817( .i (n5816), .o (n5817) );
  assign n7908 = ( n4290 & ~n5817 ) | ( n4290 & n7893 ) | ( ~n5817 & n7893 ) ;
  assign n7909 = n7779 & ~n7908 ;
  buffer buf_n7357( .i (n7356), .o (n7357) );
  buffer buf_n7358( .i (n7357), .o (n7358) );
  buffer buf_n7359( .i (n7358), .o (n7359) );
  buffer buf_n7360( .i (n7359), .o (n7360) );
  assign n7910 = ~n7360 & n7572 ;
  assign n7911 = n7058 & ~n7910 ;
  assign n7912 = n7779 | n7911 ;
  buffer buf_n7913( .i (n7779), .o (n7913) );
  assign n7914 = ( n7909 & n7912 ) | ( n7909 & ~n7913 ) | ( n7912 & ~n7913 ) ;
  assign n7915 = n7847 | n7914 ;
  assign n7916 = n591 | n7665 ;
  assign n7917 = n7847 & n7916 ;
  assign n7918 = n7915 & ~n7917 ;
  assign n7919 = ( n237 & n6207 ) | ( n237 & n7918 ) | ( n6207 & n7918 ) ;
  buffer buf_n7920( .i (n7919), .o (n7920) );
  assign n7921 = ( n151 & ~n7052 ) | ( n151 & n7920 ) | ( ~n7052 & n7920 ) ;
  buffer buf_n7922( .i (n150), .o (n7922) );
  assign n7923 = ( n239 & ~n7920 ) | ( n239 & n7922 ) | ( ~n7920 & n7922 ) ;
  assign n7924 = n7921 & ~n7923 ;
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  assign n7925 = n930 & ~n7160 ;
  assign n7926 = n601 & n7925 ;
  assign n7927 = n719 & ~n7926 ;
  buffer buf_n7928( .i (n7321), .o (n7928) );
  assign n7929 = ( n996 & n7352 ) | ( n996 & n7928 ) | ( n7352 & n7928 ) ;
  buffer buf_n7930( .i (n7929), .o (n7930) );
  buffer buf_n7931( .i (n7930), .o (n7931) );
  buffer buf_n7932( .i (n7931), .o (n7932) );
  assign n7933 = ( n7479 & n7804 ) | ( n7479 & ~n7930 ) | ( n7804 & ~n7930 ) ;
  assign n7934 = ( n7260 & ~n7677 ) | ( n7260 & n7933 ) | ( ~n7677 & n7933 ) ;
  assign n7935 = ~n7932 & n7934 ;
  buffer buf_n7936( .i (n7055), .o (n7936) );
  assign n7937 = n7935 | n7936 ;
  assign n7938 = n2054 & n7753 ;
  assign n7939 = n7936 & ~n7938 ;
  assign n7940 = n7937 & ~n7939 ;
  assign n7941 = n7778 & n7940 ;
  buffer buf_n7942( .i (n7928), .o (n7942) );
  buffer buf_n7943( .i (n7942), .o (n7943) );
  assign n7944 = ( n998 & n7705 ) | ( n998 & n7943 ) | ( n7705 & n7943 ) ;
  assign n7945 = ( n997 & n7443 ) | ( n997 & ~n7942 ) | ( n7443 & ~n7942 ) ;
  assign n7946 = ( n7705 & n7804 ) | ( n7705 & ~n7945 ) | ( n7804 & ~n7945 ) ;
  assign n7947 = ~n7944 & n7946 ;
  assign n7948 = n7753 | n7947 ;
  assign n7949 = n2833 & ~n7706 ;
  buffer buf_n7950( .i (n7375), .o (n7950) );
  buffer buf_n7951( .i (n7950), .o (n7951) );
  assign n7952 = ~n7949 & n7951 ;
  assign n7953 = n7948 & ~n7952 ;
  buffer buf_n7954( .i (n7706), .o (n7954) );
  buffer buf_n7955( .i (n2119), .o (n7955) );
  assign n7956 = ( n7951 & ~n7954 ) | ( n7951 & n7955 ) | ( ~n7954 & n7955 ) ;
  buffer buf_n7957( .i (n7943), .o (n7957) );
  assign n7958 = ( n2119 & n7706 ) | ( n2119 & ~n7957 ) | ( n7706 & ~n7957 ) ;
  buffer buf_n7959( .i (n7805), .o (n7959) );
  assign n7960 = ( n7951 & ~n7958 ) | ( n7951 & n7959 ) | ( ~n7958 & n7959 ) ;
  assign n7961 = ~n7956 & n7960 ;
  assign n7962 = n7953 | n7961 ;
  buffer buf_n7963( .i (n7599), .o (n7963) );
  assign n7964 = n7962 & ~n7963 ;
  assign n7965 = n7941 | n7964 ;
  buffer buf_n7966( .i (n7733), .o (n7966) );
  buffer buf_n7967( .i (n7966), .o (n7967) );
  assign n7968 = n7965 & ~n7967 ;
  assign n7969 = n5418 & ~n7805 ;
  assign n7970 = ( ~n5417 & n7375 ) | ( ~n5417 & n7649 ) | ( n7375 & n7649 ) ;
  buffer buf_n7971( .i (n7804), .o (n7971) );
  assign n7972 = ( n742 & ~n7970 ) | ( n742 & n7971 ) | ( ~n7970 & n7971 ) ;
  assign n7973 = ( n7959 & n7969 ) | ( n7959 & ~n7972 ) | ( n7969 & ~n7972 ) ;
  buffer buf_n7974( .i (n7973), .o (n7974) );
  buffer buf_n7975( .i (n7974), .o (n7975) );
  buffer buf_n7976( .i (n7936), .o (n7976) );
  assign n7977 = ( n7661 & n7974 ) | ( n7661 & n7976 ) | ( n7974 & n7976 ) ;
  buffer buf_n7978( .i (n7677), .o (n7978) );
  assign n7979 = ( ~n743 & n4895 ) | ( ~n743 & n7978 ) | ( n4895 & n7978 ) ;
  assign n7980 = n744 & n7979 ;
  assign n7981 = ~n7661 & n7980 ;
  assign n7982 = ( n7975 & ~n7977 ) | ( n7975 & n7981 ) | ( ~n7977 & n7981 ) ;
  assign n7983 = ( ~n3735 & n6372 ) | ( ~n3735 & n6758 ) | ( n6372 & n6758 ) ;
  buffer buf_n7984( .i (n7983), .o (n7984) );
  assign n7989 = ( n7247 & ~n7791 ) | ( n7247 & n7984 ) | ( ~n7791 & n7984 ) ;
  buffer buf_n7990( .i (n7989), .o (n7990) );
  buffer buf_n7991( .i (n7990), .o (n7991) );
  buffer buf_n7992( .i (n7991), .o (n7992) );
  buffer buf_n7993( .i (n7992), .o (n7993) );
  assign n7994 = ( ~n7141 & n7374 ) | ( ~n7141 & n7990 ) | ( n7374 & n7990 ) ;
  buffer buf_n7995( .i (n7994), .o (n7995) );
  buffer buf_n7996( .i (n7995), .o (n7996) );
  buffer buf_n7985( .i (n7984), .o (n7985) );
  buffer buf_n7986( .i (n7985), .o (n7986) );
  buffer buf_n7987( .i (n7986), .o (n7987) );
  buffer buf_n7988( .i (n7987), .o (n7988) );
  assign n7997 = ~n7988 & n7995 ;
  assign n7998 = ( ~n7993 & n7996 ) | ( ~n7993 & n7997 ) | ( n7996 & n7997 ) ;
  buffer buf_n7999( .i (n7998), .o (n7999) );
  buffer buf_n8000( .i (n7999), .o (n8000) );
  buffer buf_n8001( .i (n7978), .o (n8001) );
  buffer buf_n8002( .i (n8001), .o (n8002) );
  assign n8003 = ( n7661 & ~n7999 ) | ( n7661 & n8002 ) | ( ~n7999 & n8002 ) ;
  assign n8004 = ( n5937 & n6003 ) | ( n5937 & ~n7246 ) | ( n6003 & ~n7246 ) ;
  buffer buf_n8005( .i (n8004), .o (n8005) );
  assign n8010 = ( ~n6837 & n7003 ) | ( ~n6837 & n8005 ) | ( n7003 & n8005 ) ;
  buffer buf_n8011( .i (n8010), .o (n8011) );
  buffer buf_n8012( .i (n8011), .o (n8012) );
  buffer buf_n8013( .i (n8012), .o (n8013) );
  buffer buf_n8014( .i (n8013), .o (n8014) );
  buffer buf_n8015( .i (n7704), .o (n8015) );
  assign n8016 = ( n7649 & n8011 ) | ( n7649 & ~n8015 ) | ( n8011 & ~n8015 ) ;
  buffer buf_n8017( .i (n8016), .o (n8017) );
  buffer buf_n8018( .i (n8017), .o (n8018) );
  buffer buf_n8006( .i (n8005), .o (n8006) );
  buffer buf_n8007( .i (n8006), .o (n8007) );
  buffer buf_n8008( .i (n8007), .o (n8008) );
  buffer buf_n8009( .i (n8008), .o (n8009) );
  assign n8019 = ~n8009 & n8017 ;
  assign n8020 = ( ~n8014 & n8018 ) | ( ~n8014 & n8019 ) | ( n8018 & n8019 ) ;
  buffer buf_n8021( .i (n7517), .o (n8021) );
  assign n8022 = n8020 & n8021 ;
  assign n8023 = ( n8000 & n8003 ) | ( n8000 & n8022 ) | ( n8003 & n8022 ) ;
  assign n8024 = n7982 | n8023 ;
  assign n8025 = n7967 & n8024 ;
  assign n8026 = n7968 | n8025 ;
  buffer buf_n8027( .i (n8026), .o (n8027) );
  buffer buf_n8028( .i (n8027), .o (n8028) );
  assign n8029 = ( ~n6209 & n7900 ) | ( ~n6209 & n8027 ) | ( n7900 & n8027 ) ;
  assign n8030 = n315 | n2200 ;
  assign n8031 = ( n282 & n693 ) | ( n282 & n8030 ) | ( n693 & n8030 ) ;
  assign n8032 = n283 & ~n8031 ;
  assign n8033 = ~n7900 & n8032 ;
  assign n8034 = ( n8028 & ~n8029 ) | ( n8028 & n8033 ) | ( ~n8029 & n8033 ) ;
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n8035( .i (n7827), .o (n8035) );
  assign n8036 = ( ~n743 & n4232 ) | ( ~n743 & n8035 ) | ( n4232 & n8035 ) ;
  assign n8037 = n744 & n8036 ;
  assign n8038 = ~n7892 & n8037 ;
  buffer buf_n8039( .i (n8038), .o (n8039) );
  buffer buf_n8040( .i (n8039), .o (n8040) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  assign n8041 = ( n7375 & n7649 ) | ( n7375 & ~n7943 ) | ( n7649 & ~n7943 ) ;
  buffer buf_n8042( .i (n8041), .o (n8042) );
  buffer buf_n8043( .i (n8042), .o (n8043) );
  buffer buf_n8044( .i (n8043), .o (n8044) );
  assign n8045 = ( ~n7210 & n7516 ) | ( ~n7210 & n8042 ) | ( n7516 & n8042 ) ;
  buffer buf_n8046( .i (n7210), .o (n8046) );
  assign n8047 = ( n7839 & ~n8045 ) | ( n7839 & n8046 ) | ( ~n8045 & n8046 ) ;
  assign n8048 = ( n1497 & n8044 ) | ( n1497 & ~n8047 ) | ( n8044 & ~n8047 ) ;
  buffer buf_n8049( .i (n8048), .o (n8049) );
  buffer buf_n8050( .i (n8049), .o (n8050) );
  assign n8051 = ( n7868 & n7894 ) | ( n7868 & n8049 ) | ( n7894 & n8049 ) ;
  assign n8052 = ( n8040 & n8050 ) | ( n8040 & ~n8051 ) | ( n8050 & ~n8051 ) ;
  assign n8053 = ~n7224 & n8052 ;
  assign n8054 = n4287 & n8035 ;
  assign n8055 = ( n4232 & ~n7951 ) | ( n4232 & n8035 ) | ( ~n7951 & n8035 ) ;
  buffer buf_n8056( .i (n7950), .o (n8056) );
  assign n8057 = ~n4232 & n8056 ;
  assign n8058 = ( ~n8054 & n8055 ) | ( ~n8054 & n8057 ) | ( n8055 & n8057 ) ;
  buffer buf_n8059( .i (n8058), .o (n8059) );
  buffer buf_n8060( .i (n8059), .o (n8060) );
  assign n8061 = ( n7893 & n7963 ) | ( n7893 & ~n8059 ) | ( n7963 & ~n8059 ) ;
  assign n8062 = ( ~n8039 & n8060 ) | ( ~n8039 & n8061 ) | ( n8060 & n8061 ) ;
  assign n8063 = ( n1384 & n2609 ) | ( n1384 & ~n6128 ) | ( n2609 & ~n6128 ) ;
  assign n8064 = ( n7833 & n7839 ) | ( n7833 & ~n8063 ) | ( n7839 & ~n8063 ) ;
  buffer buf_n8065( .i (n8064), .o (n8065) );
  buffer buf_n8066( .i (n7976), .o (n8066) );
  assign n8067 = ( ~n7733 & n8065 ) | ( ~n7733 & n8066 ) | ( n8065 & n8066 ) ;
  assign n8068 = ( n7811 & ~n8065 ) | ( n7811 & n8066 ) | ( ~n8065 & n8066 ) ;
  assign n8069 = n8067 & ~n8068 ;
  assign n8070 = n8062 & ~n8069 ;
  assign n8071 = n7224 & ~n8070 ;
  assign n8072 = n8053 | n8071 ;
  buffer buf_n2155( .i (n2154), .o (n2155) );
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n8073( .i (n7833), .o (n8073) );
  buffer buf_n8074( .i (n8073), .o (n8074) );
  assign n8075 = n7192 | n8074 ;
  assign n8076 = ( n596 & n2157 ) | ( n596 & n8075 ) | ( n2157 & n8075 ) ;
  assign n8077 = ( n597 & ~n7967 ) | ( n597 & n8076 ) | ( ~n7967 & n8076 ) ;
  buffer buf_n8078( .i (n8035), .o (n8078) );
  buffer buf_n8079( .i (n8078), .o (n8079) );
  assign n8080 = n4428 & ~n8079 ;
  assign n8081 = n8074 & n8080 ;
  buffer buf_n8082( .i (n8081), .o (n8082) );
  buffer buf_n8083( .i (n8082), .o (n8083) );
  buffer buf_n8084( .i (n7894), .o (n8084) );
  assign n8085 = n8082 | n8084 ;
  assign n8086 = ( n8077 & n8083 ) | ( n8077 & n8085 ) | ( n8083 & n8085 ) ;
  buffer buf_n8087( .i (n6259), .o (n8087) );
  assign n8088 = ( n7620 & n8086 ) | ( n7620 & n8087 ) | ( n8086 & n8087 ) ;
  assign n8089 = ( ~n434 & n8072 ) | ( ~n434 & n8088 ) | ( n8072 & n8088 ) ;
  assign n8090 = ( n7141 & n7374 ) | ( n7141 & n7942 ) | ( n7374 & n7942 ) ;
  buffer buf_n8091( .i (n8090), .o (n8091) );
  buffer buf_n8092( .i (n8015), .o (n8092) );
  assign n8093 = ( n7950 & ~n8091 ) | ( n7950 & n8092 ) | ( ~n8091 & n8092 ) ;
  assign n8094 = ( ~n7544 & n8091 ) | ( ~n7544 & n8092 ) | ( n8091 & n8092 ) ;
  assign n8095 = ~n8093 & n8094 ;
  buffer buf_n8096( .i (n6909), .o (n8096) );
  assign n8097 = n8095 | n8096 ;
  assign n8098 = n3867 | n8092 ;
  assign n8099 = n8056 | n8098 ;
  assign n8100 = n8096 & n8099 ;
  assign n8101 = n8097 & ~n8100 ;
  assign n8102 = ( n7733 & n7893 ) | ( n7733 & n8101 ) | ( n7893 & n8101 ) ;
  buffer buf_n8103( .i (n8102), .o (n8103) );
  assign n8104 = ( n7533 & ~n8084 ) | ( n7533 & n8103 ) | ( ~n8084 & n8103 ) ;
  assign n8105 = ( n7533 & n7967 ) | ( n7533 & ~n8103 ) | ( n7967 & ~n8103 ) ;
  assign n8106 = n8104 & ~n8105 ;
  buffer buf_n8107( .i (n8106), .o (n8107) );
  buffer buf_n8108( .i (n8107), .o (n8108) );
  assign n8109 = n7900 & ~n8107 ;
  assign n8110 = ( n8089 & n8108 ) | ( n8089 & ~n8109 ) | ( n8108 & ~n8109 ) ;
  assign n8111 = n8034 | n8110 ;
  assign n8112 = ( n720 & ~n7927 ) | ( n720 & n8111 ) | ( ~n7927 & n8111 ) ;
  assign n8113 = n7924 | n8112 ;
  assign n8114 = ( n7906 & ~n7907 ) | ( n7906 & n8113 ) | ( ~n7907 & n8113 ) ;
  assign y0 = n420 ;
  assign y1 = n765 ;
  assign y2 = n1098 ;
  assign y3 = n1422 ;
  assign y4 = n1957 ;
  assign y5 = n2624 ;
  assign y6 = n3111 ;
  assign y7 = n3493 ;
  assign y8 = n3863 ;
  assign y9 = n4372 ;
  assign y10 = n4816 ;
  assign y11 = n5177 ;
  assign y12 = n5570 ;
  assign y13 = n5862 ;
  assign y14 = n6232 ;
  assign y15 = n6548 ;
  assign y16 = n6897 ;
  assign y17 = n7234 ;
  assign y18 = n7590 ;
  assign y19 = n7879 ;
  assign y20 = n8114 ;
endmodule
