module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 ;
  wire n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 ;
  buffer buf_n833( .i (x28), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n776( .i (x26), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n608( .i (x21), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n508( .i (x18), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n541( .i (x19), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  assign n1320 = ~n521 & n554 ;
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  assign n1338 = n628 & n1326 ;
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  assign n1343 = n799 & n1340 ;
  buffer buf_n865( .i (x29), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n900( .i (x30), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  assign n1344 = ~n884 & n919 ;
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  assign n1355 = ( n857 & n1343 ) | ( n857 & n1348 ) | ( n1343 & n1348 ) ;
  assign n1356 = ~n858 & n1355 ;
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n46( .i (x0), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  assign n1369 = ~n72 & n534 ;
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n573( .i (x20), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  assign n1372 = ~n588 & n623 ;
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  assign n1385 = ( n569 & n1370 ) | ( n569 & n1384 ) | ( n1370 & n1384 ) ;
  assign n1386 = ~n570 & n1385 ;
  assign n1387 = ( n863 & n1354 ) | ( n863 & n1386 ) | ( n1354 & n1386 ) ;
  assign n1388 = ~n864 & n1387 ;
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  assign n1394 = n559 & n626 ;
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  assign n1404 = ( n601 & ~n1370 ) | ( n601 & n1403 ) | ( ~n1370 & n1403 ) ;
  assign n1405 = n1371 & n1404 ;
  buffer buf_n710( .i (x24), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  assign n1406 = n732 & n922 ;
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  assign n1414 = ( n895 & n1405 ) | ( n895 & n1413 ) | ( n1405 & n1413 ) ;
  assign n1415 = ~n896 & n1414 ;
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n320( .i (x10), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  assign n1420 = n340 & n628 ;
  assign n1421 = ( n529 & n562 ) | ( n529 & n1420 ) | ( n562 & n1420 ) ;
  assign n1422 = ~n530 & n1421 ;
  buffer buf_n741( .i (x25), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  assign n1423 = n763 & ~n887 ;
  assign n1424 = ( n856 & n1422 ) | ( n856 & n1423 ) | ( n1422 & n1423 ) ;
  assign n1425 = ~n857 & n1424 ;
  assign n1426 = n925 & n1425 ;
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  assign n1436 = n735 & n1342 ;
  assign n1437 = ( n859 & n1350 ) | ( n859 & n1436 ) | ( n1350 & n1436 ) ;
  assign n1438 = ~n860 & n1437 ;
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  assign n1445 = ~n522 & n587 ;
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  buffer buf_n1455( .i (n1454), .o (n1455) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  assign n1458 = ( n73 & ~n568 ) | ( n73 & n1457 ) | ( ~n568 & n1457 ) ;
  assign n1459 = ~n74 & n1458 ;
  assign n1460 = n637 & n1459 ;
  assign n1461 = ( n740 & n895 ) | ( n740 & n1460 ) | ( n895 & n1460 ) ;
  assign n1462 = ~n896 & n1461 ;
  assign n1463 = n932 & n1462 ;
  buffer buf_n1464( .i (n1463), .o (n1464) );
  assign n1465 = n1444 | n1464 ;
  assign n1466 = n1435 | n1465 ;
  assign n1467 = n1419 | n1466 ;
  assign n1468 = ( ~n1367 & n1393 ) | ( ~n1367 & n1467 ) | ( n1393 & n1467 ) ;
  assign n1469 = n1368 | n1468 ;
  assign n1470 = n1417 | n1464 ;
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  assign n1475 = n1357 | n1427 ;
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  assign n1487 = n1363 | n1416 ;
  assign n1488 = n1444 | n1487 ;
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  assign n1493 = ~n554 & n586 ;
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  assign n1510 = ( n65 & n527 ) | ( n65 & n1498 ) | ( n527 & n1498 ) ;
  assign n1511 = ~n528 & n1510 ;
  buffer buf_n1512( .i (n1511), .o (n1512) );
  assign n1513 = n630 & n1512 ;
  buffer buf_n1514( .i (n1513), .o (n1514) );
  assign n1516 = ( n889 & n1407 ) | ( n889 & n1514 ) | ( n1407 & n1514 ) ;
  assign n1517 = ~n890 & n1516 ;
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n1522( .i (n1521), .o (n1522) );
  assign n1523 = n63 & n558 ;
  buffer buf_n1524( .i (n1523), .o (n1524) );
  assign n1527 = n527 & n1524 ;
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  assign n1534 = n599 & n1533 ;
  assign n1535 = n627 & n919 ;
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  assign n1544 = ( n892 & n1534 ) | ( n892 & n1542 ) | ( n1534 & n1542 ) ;
  assign n1545 = ~n893 & n1544 ;
  buffer buf_n1546( .i (n1545), .o (n1546) );
  assign n1549 = n61 & ~n556 ;
  buffer buf_n1550( .i (n1549), .o (n1550) );
  assign n1556 = n525 & n1550 ;
  assign n1557 = ~n851 & n1556 ;
  assign n1558 = ( n592 & n627 ) | ( n592 & n1557 ) | ( n627 & n1557 ) ;
  assign n1559 = ~n593 & n1558 ;
  assign n1560 = n1345 & n1559 ;
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  assign n1569 = n68 & n630 ;
  assign n1570 = ( n531 & n564 ) | ( n531 & n1569 ) | ( n564 & n1569 ) ;
  assign n1571 = ~n532 & n1570 ;
  assign n1572 = n852 & n919 ;
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  assign n1579 = ( n890 & n1571 ) | ( n890 & n1577 ) | ( n1571 & n1577 ) ;
  assign n1580 = ~n891 & n1579 ;
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  assign n1586 = n1567 | n1582 ;
  assign n1587 = ( ~n1521 & n1546 ) | ( ~n1521 & n1586 ) | ( n1546 & n1586 ) ;
  assign n1588 = n1522 | n1587 ;
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n346( .i (x11), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  assign n1596 = n336 & n524 ;
  buffer buf_n1597( .i (n1596), .o (n1597) );
  assign n1600 = ( n64 & n364 ) | ( n64 & n1597 ) | ( n364 & n1597 ) ;
  assign n1601 = ~n365 & n1600 ;
  assign n1602 = n554 & ~n621 ;
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  assign n1611 = ( n593 & n1601 ) | ( n593 & n1608 ) | ( n1601 & n1608 ) ;
  assign n1612 = ~n594 & n1611 ;
  assign n1613 = n763 & n1612 ;
  assign n1614 = ( n888 & n923 ) | ( n888 & n1613 ) | ( n923 & n1613 ) ;
  assign n1615 = ~n924 & n1614 ;
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n146( .i (x3), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  assign n1627 = n165 & n560 ;
  assign n1628 = ( ~n66 & n528 ) | ( ~n66 & n1627 ) | ( n528 & n1627 ) ;
  assign n1629 = n67 & n1628 ;
  buffer buf_n804( .i (x27), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  assign n1630 = n594 & n825 ;
  assign n1631 = ( n630 & n1629 ) | ( n630 & n1630 ) | ( n1629 & n1630 ) ;
  assign n1632 = ~n631 & n1631 ;
  assign n1633 = ~n889 & n1632 ;
  assign n1634 = ~n925 & n1633 ;
  buffer buf_n1635( .i (n1634), .o (n1635) );
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n1637( .i (n1636), .o (n1637) );
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n203( .i (x5), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n1643 = n57 & ~n214 ;
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  assign n1652 = n560 & n1650 ;
  assign n1653 = n528 & n1652 ;
  assign n1654 = n592 & ~n823 ;
  buffer buf_n1655( .i (n1654), .o (n1655) );
  assign n1657 = ( n629 & n1653 ) | ( n629 & n1655 ) | ( n1653 & n1655 ) ;
  buffer buf_n1658( .i (n629), .o (n1658) );
  assign n1659 = n1657 & ~n1658 ;
  assign n1660 = n923 & n1659 ;
  assign n1661 = ( n857 & n889 ) | ( n857 & n1660 ) | ( n889 & n1660 ) ;
  assign n1662 = ~n858 & n1661 ;
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n177( .i (x4), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  assign n1670 = ~n196 & n560 ;
  buffer buf_n1671( .i (n527), .o (n1671) );
  assign n1672 = ( n66 & n1670 ) | ( n66 & n1671 ) | ( n1670 & n1671 ) ;
  assign n1673 = ~n67 & n1672 ;
  assign n1674 = ( n1656 & n1658 ) | ( n1656 & n1673 ) | ( n1658 & n1673 ) ;
  assign n1675 = ~n631 & n1674 ;
  buffer buf_n1676( .i (n856), .o (n1676) );
  assign n1677 = n1675 & n1676 ;
  assign n1678 = ( n890 & n925 ) | ( n890 & n1677 ) | ( n925 & n1677 ) ;
  assign n1679 = ~n926 & n1678 ;
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  assign n1687 = n1669 | n1685 ;
  assign n1688 = n1642 | n1687 ;
  assign n1689 = ~n627 & n795 ;
  buffer buf_n1690( .i (n1689), .o (n1690) );
  assign n1694 = ( n594 & n1528 ) | ( n594 & n1690 ) | ( n1528 & n1690 ) ;
  assign n1695 = ~n595 & n1694 ;
  assign n1696 = ~n923 & n1695 ;
  buffer buf_n1697( .i (n888), .o (n1697) );
  assign n1698 = ( n1676 & n1696 ) | ( n1676 & n1697 ) | ( n1696 & n1697 ) ;
  assign n1699 = ~n858 & n1698 ;
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  assign n1709 = n367 & n562 ;
  assign n1710 = ( ~n68 & n530 ) | ( ~n68 & n1709 ) | ( n530 & n1709 ) ;
  assign n1711 = n69 & n1710 ;
  assign n1712 = ( n597 & n1693 ) | ( n597 & n1711 ) | ( n1693 & n1711 ) ;
  assign n1713 = ~n598 & n1712 ;
  assign n1714 = ( n891 & n1578 ) | ( n891 & n1713 ) | ( n1578 & n1713 ) ;
  assign n1715 = ~n892 & n1714 ;
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  assign n1722 = ( n367 & n529 ) | ( n367 & n1526 ) | ( n529 & n1526 ) ;
  assign n1723 = ~n368 & n1722 ;
  assign n1724 = ( n596 & n1692 ) | ( n596 & n1723 ) | ( n1692 & n1723 ) ;
  assign n1725 = ~n597 & n1724 ;
  buffer buf_n1726( .i (n1697), .o (n1726) );
  assign n1727 = ( n1577 & n1725 ) | ( n1577 & n1726 ) | ( n1725 & n1726 ) ;
  assign n1728 = ~n891 & n1727 ;
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  assign n1734 = n1718 | n1732 ;
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  assign n1737 = n1707 | n1736 ;
  assign n1738 = ( ~n1625 & n1688 ) | ( ~n1625 & n1737 ) | ( n1688 & n1737 ) ;
  assign n1739 = n1626 | n1738 ;
  buffer buf_n117( .i (x2), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  assign n1740 = n62 & ~n162 ;
  assign n1741 = ( n134 & ~n525 ) | ( n134 & n1740 ) | ( ~n525 & n1740 ) ;
  assign n1742 = ~n135 & n1741 ;
  buffer buf_n1743( .i (n626), .o (n1743) );
  assign n1744 = n1742 & ~n1743 ;
  assign n1745 = ( n561 & n593 ) | ( n561 & n1744 ) | ( n593 & n1744 ) ;
  assign n1746 = ~n562 & n1745 ;
  assign n1747 = ( n887 & n1574 ) | ( n887 & n1746 ) | ( n1574 & n1746 ) ;
  assign n1748 = ~n888 & n1747 ;
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n680( .i (x23), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  assign n1758 = ~n855 & n1512 ;
  assign n1759 = ( n631 & n703 ) | ( n631 & n1758 ) | ( n703 & n1758 ) ;
  assign n1760 = ~n632 & n1759 ;
  buffer buf_n1761( .i (n924), .o (n1761) );
  assign n1762 = n1760 & ~n1761 ;
  buffer buf_n1763( .i (n1726), .o (n1763) );
  assign n1764 = n1762 & n1763 ;
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  assign n1773 = n134 & ~n525 ;
  assign n1774 = ( n64 & n164 ) | ( n64 & n1773 ) | ( n164 & n1773 ) ;
  assign n1775 = ~n165 & n1774 ;
  buffer buf_n1776( .i (n592), .o (n1776) );
  assign n1777 = n1775 & ~n1776 ;
  buffer buf_n1778( .i (n561), .o (n1778) );
  assign n1779 = ( ~n629 & n1777 ) | ( ~n629 & n1778 ) | ( n1777 & n1778 ) ;
  assign n1780 = ~n563 & n1779 ;
  buffer buf_n1781( .i (n887), .o (n1781) );
  assign n1782 = ( n1575 & n1780 ) | ( n1575 & n1781 ) | ( n1780 & n1781 ) ;
  assign n1783 = ~n1697 & n1782 ;
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n438( .i (x15), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  assign n1793 = ~n457 & n1650 ;
  assign n1794 = n366 & n1793 ;
  assign n1795 = n522 & n587 ;
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  assign n1811 = ( n1778 & n1794 ) | ( n1778 & n1801 ) | ( n1794 & n1801 ) ;
  assign n1812 = ~n563 & n1811 ;
  buffer buf_n1813( .i (n1658), .o (n1813) );
  assign n1814 = n1812 & n1813 ;
  assign n1815 = ( n800 & n1676 ) | ( n800 & n1814 ) | ( n1676 & n1814 ) ;
  buffer buf_n1816( .i (n1676), .o (n1816) );
  assign n1817 = n1815 & ~n1816 ;
  assign n1818 = n1350 & n1817 ;
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  assign n1825 = ~n359 & n1644 ;
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  assign n1828 = ~n454 & n1827 ;
  assign n1829 = ( n558 & n1797 ) | ( n558 & n1828 ) | ( n1797 & n1828 ) ;
  assign n1830 = ~n559 & n1829 ;
  assign n1831 = n1743 & n1830 ;
  assign n1832 = ( n796 & n853 ) | ( n796 & n1831 ) | ( n853 & n1831 ) ;
  assign n1833 = ~n854 & n1832 ;
  assign n1834 = n1346 & n1833 ;
  buffer buf_n1835( .i (n1834), .o (n1835) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n458( .i (n457), .o (n458) );
  assign n1847 = n362 & n1647 ;
  assign n1848 = n337 & n1847 ;
  assign n1849 = ~n559 & n1848 ;
  buffer buf_n1850( .i (n526), .o (n1850) );
  assign n1851 = ( n457 & n1849 ) | ( n457 & n1850 ) | ( n1849 & n1850 ) ;
  assign n1852 = ~n458 & n1851 ;
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  assign n1855 = n591 & n759 ;
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  assign n1859 = ( n1658 & ~n1853 ) | ( n1658 & n1858 ) | ( ~n1853 & n1858 ) ;
  assign n1860 = n1854 & n1859 ;
  buffer buf_n1861( .i (n856), .o (n1861) );
  assign n1862 = ( n1348 & n1860 ) | ( n1348 & n1861 ) | ( n1860 & n1861 ) ;
  assign n1863 = ~n1816 & n1862 ;
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1871( .i (n524), .o (n1871) );
  assign n1872 = ( n163 & n1648 ) | ( n163 & ~n1871 ) | ( n1648 & ~n1871 ) ;
  assign n1873 = ~n164 & n1872 ;
  buffer buf_n1874( .i (n591), .o (n1874) );
  assign n1875 = n1873 & ~n1874 ;
  assign n1876 = ( n561 & ~n628 ) | ( n561 & n1875 ) | ( ~n628 & n1875 ) ;
  assign n1877 = ~n1778 & n1876 ;
  assign n1878 = ~n922 & n1877 ;
  buffer buf_n1879( .i (n855), .o (n1879) );
  assign n1880 = ( n1781 & n1878 ) | ( n1781 & n1879 ) | ( n1878 & n1879 ) ;
  assign n1881 = ~n1861 & n1880 ;
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  assign n1890 = n1864 | n1883 ;
  assign n1891 = ( ~n1819 & n1839 ) | ( ~n1819 & n1890 ) | ( n1839 & n1890 ) ;
  assign n1892 = n1820 | n1891 ;
  assign n1893 = n1788 | n1892 ;
  assign n1894 = ( ~n1755 & n1768 ) | ( ~n1755 & n1893 ) | ( n1768 & n1893 ) ;
  assign n1895 = n1756 | n1894 ;
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n644( .i (x22), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  assign n1898 = n665 & n921 ;
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  assign n1902 = ( n1515 & n1726 ) | ( n1515 & n1901 ) | ( n1726 & n1901 ) ;
  assign n1903 = ~n1763 & n1902 ;
  buffer buf_n1904( .i (n1903), .o (n1904) );
  assign n1905 = n339 & ~n1850 ;
  assign n1906 = ( n66 & n366 ) | ( n66 & n1905 ) | ( n366 & n1905 ) ;
  assign n1907 = ~n367 & n1906 ;
  buffer buf_n1908( .i (n1743), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  assign n1911 = n1907 & n1910 ;
  assign n1912 = ( n564 & n596 ) | ( n564 & n1911 ) | ( n596 & n1911 ) ;
  assign n1913 = ~n565 & n1912 ;
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n1914( .i (n922), .o (n1914) );
  assign n1915 = n764 & n1914 ;
  buffer buf_n1916( .i (n1915), .o (n1916) );
  assign n1918 = ( n1726 & n1913 ) | ( n1726 & n1916 ) | ( n1913 & n1916 ) ;
  assign n1919 = ~n1763 & n1918 ;
  buffer buf_n1920( .i (n1919), .o (n1920) );
  assign n1926 = n1904 | n1920 ;
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  buffer buf_n1930( .i (n1929), .o (n1930) );
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1932( .i (n558), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  assign n1934 = n365 & ~n1933 ;
  buffer buf_n1935( .i (n65), .o (n1935) );
  assign n1936 = ( n1671 & n1934 ) | ( n1671 & n1935 ) | ( n1934 & n1935 ) ;
  assign n1937 = ~n529 & n1936 ;
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  assign n1940 = n590 & n793 ;
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  assign n1952 = ( n1813 & ~n1938 ) | ( n1813 & n1945 ) | ( ~n1938 & n1945 ) ;
  assign n1953 = n1939 & n1952 ;
  assign n1954 = n1349 & n1953 ;
  buffer buf_n1955( .i (n1954), .o (n1955) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  buffer buf_n1960( .i (n1959), .o (n1960) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  assign n1961 = ( n458 & n1326 ) | ( n458 & n1651 ) | ( n1326 & n1651 ) ;
  assign n1962 = ~n459 & n1961 ;
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  assign n1965 = n590 & n661 ;
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n1967( .i (n1966), .o (n1967) );
  buffer buf_n1968( .i (n1967), .o (n1968) );
  buffer buf_n1969( .i (n1968), .o (n1969) );
  buffer buf_n1970( .i (n1969), .o (n1970) );
  assign n1971 = ( n1813 & ~n1963 ) | ( n1813 & n1970 ) | ( ~n1963 & n1970 ) ;
  assign n1972 = n1964 & n1971 ;
  assign n1973 = ( n1349 & n1816 ) | ( n1349 & n1972 ) | ( n1816 & n1972 ) ;
  assign n1974 = ~n859 & n1973 ;
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  assign n1987 = n335 & n1826 ;
  assign n1988 = ~n557 & n1987 ;
  assign n1989 = ( n455 & n1871 ) | ( n455 & n1988 ) | ( n1871 & n1988 ) ;
  assign n1990 = ~n456 & n1989 ;
  buffer buf_n1991( .i (n1990), .o (n1991) );
  buffer buf_n1992( .i (n1991), .o (n1992) );
  assign n1993 = ( n1856 & n1908 ) | ( n1856 & ~n1991 ) | ( n1908 & ~n1991 ) ;
  assign n1994 = n1992 & n1993 ;
  assign n1995 = ( n855 & n1346 ) | ( n855 & n1994 ) | ( n1346 & n1994 ) ;
  assign n1996 = ~n1879 & n1995 ;
  buffer buf_n1997( .i (n1996), .o (n1997) );
  buffer buf_n1998( .i (n1997), .o (n1998) );
  buffer buf_n1999( .i (n1998), .o (n1999) );
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n2001( .i (n2000), .o (n2001) );
  assign n2005 = n1650 & ~n1933 ;
  assign n2006 = ( n458 & n1671 ) | ( n458 & n2005 ) | ( n1671 & n2005 ) ;
  assign n2007 = ~n459 & n2006 ;
  buffer buf_n2008( .i (n2007), .o (n2008) );
  buffer buf_n2009( .i (n2008), .o (n2009) );
  assign n2010 = ( n1813 & n1970 ) | ( n1813 & ~n2008 ) | ( n1970 & ~n2008 ) ;
  assign n2011 = n2009 & n2010 ;
  assign n2012 = ( n1349 & n1816 ) | ( n1349 & n2011 ) | ( n1816 & n2011 ) ;
  assign n2013 = ~n859 & n2012 ;
  buffer buf_n2014( .i (n2013), .o (n2014) );
  buffer buf_n2015( .i (n2014), .o (n2015) );
  assign n2016 = n2001 | n2015 ;
  buffer buf_n2017( .i (n2016), .o (n2017) );
  assign n2019 = n1978 | n2017 ;
  assign n2020 = n1960 | n2019 ;
  buffer buf_n1917( .i (n1916), .o (n1917) );
  assign n2021 = n340 & n1935 ;
  buffer buf_n2022( .i (n366), .o (n2022) );
  buffer buf_n2023( .i (n1671), .o (n2023) );
  assign n2024 = ( n2021 & n2022 ) | ( n2021 & n2023 ) | ( n2022 & n2023 ) ;
  assign n2025 = ~n530 & n2024 ;
  buffer buf_n2026( .i (n1910), .o (n2026) );
  assign n2027 = n2025 & n2026 ;
  assign n2028 = ( n565 & n597 ) | ( n565 & n2027 ) | ( n597 & n2027 ) ;
  assign n2029 = ~n566 & n2028 ;
  assign n2030 = ( n1763 & n1917 ) | ( n1763 & n2029 ) | ( n1917 & n2029 ) ;
  assign n2031 = ~n892 & n2030 ;
  buffer buf_n2032( .i (n2031), .o (n2032) );
  assign n2034 = n65 & ~n1850 ;
  buffer buf_n2035( .i (n365), .o (n2035) );
  buffer buf_n2036( .i (n1933), .o (n2036) );
  assign n2037 = ( n2034 & n2035 ) | ( n2034 & ~n2036 ) | ( n2035 & ~n2036 ) ;
  assign n2038 = ~n2022 & n2037 ;
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  assign n2041 = ( n1945 & n2026 ) | ( n1945 & ~n2039 ) | ( n2026 & ~n2039 ) ;
  assign n2042 = n2040 & n2041 ;
  buffer buf_n2043( .i (n1348), .o (n2043) );
  assign n2044 = n2042 & n2043 ;
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  assign n2051 = n2032 | n2047 ;
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  assign n2055 = n2020 | n2054 ;
  assign n2056 = ( ~n1896 & n1931 ) | ( ~n1896 & n2055 ) | ( n1931 & n2055 ) ;
  assign n2057 = n1897 | n2056 ;
  assign n2058 = ~n626 & n662 ;
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  assign n2062 = ( n595 & n1529 ) | ( n595 & n2061 ) | ( n1529 & n2061 ) ;
  assign n2063 = ~n596 & n2062 ;
  assign n2064 = ~n924 & n2063 ;
  buffer buf_n2065( .i (n1697), .o (n2065) );
  assign n2066 = n2064 & n2065 ;
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n2073( .i (n2072), .o (n2073) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n2075( .i (n2074), .o (n2075) );
  assign n2076 = n63 & n590 ;
  assign n2077 = ( n526 & n1932 ) | ( n526 & n2076 ) | ( n1932 & n2076 ) ;
  assign n2078 = ~n1850 & n2077 ;
  assign n2079 = n2059 & n2078 ;
  assign n2080 = n854 & n2079 ;
  buffer buf_n2081( .i (n886), .o (n2081) );
  buffer buf_n2082( .i (n921), .o (n2082) );
  assign n2083 = ( n2080 & n2081 ) | ( n2080 & n2082 ) | ( n2081 & n2082 ) ;
  assign n2084 = ~n1914 & n2083 ;
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2089( .i (n2088), .o (n2089) );
  buffer buf_n2090( .i (n2089), .o (n2090) );
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  assign n2094 = n1324 & n1649 ;
  assign n2095 = ( n1743 & n1966 ) | ( n1743 & n2094 ) | ( n1966 & n2094 ) ;
  assign n2096 = ~n1908 & n2095 ;
  assign n2097 = ~n921 & n2096 ;
  buffer buf_n2098( .i (n854), .o (n2098) );
  assign n2099 = ( n2081 & n2097 ) | ( n2081 & n2098 ) | ( n2097 & n2098 ) ;
  assign n2100 = ~n1879 & n2099 ;
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n2102( .i (n2101), .o (n2102) );
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n488( .i (x17), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  assign n2111 = n62 & n504 ;
  buffer buf_n2112( .i (n557), .o (n2112) );
  assign n2113 = ( n1871 & n2111 ) | ( n1871 & n2112 ) | ( n2111 & n2112 ) ;
  assign n2114 = ~n1932 & n2113 ;
  buffer buf_n2115( .i (n625), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  assign n2117 = ( n1941 & n2114 ) | ( n1941 & n2116 ) | ( n2114 & n2116 ) ;
  assign n2118 = ~n1908 & n2117 ;
  buffer buf_n2119( .i (n920), .o (n2119) );
  assign n2120 = n2118 & ~n2119 ;
  assign n2121 = ( n2081 & n2098 ) | ( n2081 & n2120 ) | ( n2098 & n2120 ) ;
  assign n2122 = ~n1879 & n2121 ;
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  assign n2131 = ( n505 & n1550 ) | ( n505 & n1871 ) | ( n1550 & n1871 ) ;
  assign n2132 = ~n506 & n2131 ;
  assign n2133 = ( n1941 & n2116 ) | ( n1941 & n2132 ) | ( n2116 & n2132 ) ;
  buffer buf_n2134( .i (n2116), .o (n2134) );
  assign n2135 = n2133 & ~n2134 ;
  assign n2136 = ~n2119 & n2135 ;
  assign n2137 = ( n2081 & n2098 ) | ( n2081 & n2136 ) | ( n2098 & n2136 ) ;
  buffer buf_n2138( .i (n2098), .o (n2138) );
  assign n2139 = n2137 & ~n2138 ;
  buffer buf_n2140( .i (n2139), .o (n2140) );
  assign n2149 = n2123 | n2140 ;
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  buffer buf_n2152( .i (n2151), .o (n2152) );
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n2155( .i (n2154), .o (n2155) );
  assign n2156 = n2108 | n2155 ;
  assign n2157 = n2093 | n2156 ;
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  assign n2158 = ( n1599 & ~n1935 ) | ( n1599 & n2035 ) | ( ~n1935 & n2035 ) ;
  assign n2159 = n67 & n2158 ;
  assign n2160 = ( n595 & n1610 ) | ( n595 & n2159 ) | ( n1610 & n2159 ) ;
  buffer buf_n2161( .i (n1776), .o (n2161) );
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n2163( .i (n2162), .o (n2163) );
  assign n2164 = n2160 & ~n2163 ;
  assign n2165 = n765 & n2164 ;
  assign n2166 = ( n1761 & n2065 ) | ( n1761 & n2165 ) | ( n2065 & n2165 ) ;
  assign n2167 = ~n926 & n2166 ;
  buffer buf_n2168( .i (n2167), .o (n2168) );
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  buffer buf_n2171( .i (n2170), .o (n2171) );
  buffer buf_n2172( .i (n2171), .o (n2172) );
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n2174( .i (n2023), .o (n2174) );
  assign n2175 = ( n368 & n1555 ) | ( n368 & n2174 ) | ( n1555 & n2174 ) ;
  assign n2176 = ~n369 & n2175 ;
  assign n2177 = ( n632 & n1946 ) | ( n632 & n2176 ) | ( n1946 & n2176 ) ;
  assign n2178 = ~n633 & n2177 ;
  buffer buf_n2179( .i (n2065), .o (n2179) );
  assign n2180 = ( n1578 & n2178 ) | ( n1578 & n2179 ) | ( n2178 & n2179 ) ;
  buffer buf_n2181( .i (n2179), .o (n2181) );
  assign n2182 = n2180 & ~n2181 ;
  buffer buf_n2183( .i (n2182), .o (n2183) );
  buffer buf_n2187( .i (n1935), .o (n2187) );
  assign n2188 = n2022 & n2187 ;
  assign n2189 = ( n563 & n2174 ) | ( n563 & n2188 ) | ( n2174 & n2188 ) ;
  assign n2190 = ~n564 & n2189 ;
  assign n2191 = ( n632 & n1946 ) | ( n632 & n2190 ) | ( n1946 & n2190 ) ;
  assign n2192 = ~n633 & n2191 ;
  assign n2193 = ( n1578 & n2179 ) | ( n1578 & n2192 ) | ( n2179 & n2192 ) ;
  assign n2194 = ~n2181 & n2193 ;
  buffer buf_n2195( .i (n2194), .o (n2195) );
  assign n2200 = n2183 | n2195 ;
  buffer buf_n2201( .i (n2200), .o (n2201) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  buffer buf_n2203( .i (n2202), .o (n2203) );
  assign n2204 = n2173 | n2203 ;
  assign n2205 = ( ~n2074 & n2157 ) | ( ~n2074 & n2204 ) | ( n2157 & n2204 ) ;
  assign n2206 = n2075 | n2205 ;
  assign n2207 = n2057 | n2206 ;
  assign n2208 = n1739 | n2207 ;
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  assign n2210 = n2001 | n2032 ;
  assign n2211 = n1922 | n2210 ;
  assign n2212 = n1621 | n2211 ;
  assign n2213 = ( ~n1869 & n2172 ) | ( ~n1869 & n2212 ) | ( n2172 & n2212 ) ;
  assign n2214 = n1870 | n2213 ;
  buffer buf_n2215( .i (n2214), .o (n2215) );
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  assign n2220 = n1928 | n1978 ;
  assign n2221 = n2050 | n2220 ;
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n1888( .i (n1887), .o (n1888) );
  buffer buf_n2018( .i (n2017), .o (n2018) );
  assign n2222 = n1888 | n2018 ;
  assign n2223 = ( ~n1844 & n2221 ) | ( ~n1844 & n2222 ) | ( n2221 & n2222 ) ;
  assign n2224 = n1845 | n2223 ;
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  assign n2225 = n1753 | n2195 ;
  assign n2226 = ( ~n2070 & n2090 ) | ( ~n2070 & n2225 ) | ( n2090 & n2225 ) ;
  assign n2227 = n2071 | n2226 ;
  assign n2228 = n1733 | n2227 ;
  assign n2229 = ( n1623 & ~n1685 ) | ( n1623 & n2228 ) | ( ~n1685 & n2228 ) ;
  assign n2230 = n1686 | n2229 ;
  assign n2231 = n2224 | n2230 ;
  buffer buf_n2232( .i (n2231), .o (n2232) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  assign n2235 = n1637 | n1766 ;
  assign n2236 = n1788 | n2235 ;
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  assign n2245 = ~n552 & n619 ;
  buffer buf_n2246( .i (n2245), .o (n2246) );
  assign n2249 = ( n521 & ~n586 ) | ( n521 & n2246 ) | ( ~n586 & n2246 ) ;
  assign n2250 = ~n522 & n2249 ;
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  assign n2260 = n662 & n883 ;
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  assign n2265 = ( n2138 & n2258 ) | ( n2138 & n2264 ) | ( n2258 & n2264 ) ;
  assign n2266 = ~n1861 & n2265 ;
  assign n2267 = n1761 & n2266 ;
  buffer buf_n2268( .i (n2267), .o (n2268) );
  buffer buf_n2269( .i (n2268), .o (n2269) );
  buffer buf_n2270( .i (n2269), .o (n2270) );
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2273( .i (n2272), .o (n2273) );
  buffer buf_n1199( .i (x40), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1247( .i (x42), .o (n1247) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1220( .i (x41), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1173( .i (x39), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1158( .i (x38), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n302( .i (x9), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  assign n2274 = n512 | n577 ;
  assign n2275 = ( ~n307 & n546 ) | ( ~n307 & n2274 ) | ( n546 & n2274 ) ;
  assign n2276 = n308 | n2275 ;
  assign n2277 = n615 & ~n2276 ;
  assign n2278 = ( n652 & n841 ) | ( n652 & n2277 ) | ( n841 & n2277 ) ;
  assign n2279 = ~n842 & n2278 ;
  buffer buf_n2280( .i (n2279), .o (n2280) );
  assign n2295 = ~n911 & n2280 ;
  assign n2296 = n877 & n2295 ;
  buffer buf_n2297( .i (n2296), .o (n2297) );
  assign n2298 = ~n1172 & n2297 ;
  buffer buf_n2299( .i (n2298), .o (n2299) );
  assign n2309 = ~n1189 & n2299 ;
  buffer buf_n2310( .i (n2309), .o (n2310) );
  assign n2317 = ~n1238 & n2310 ;
  assign n2318 = ( n1218 & ~n1266 ) | ( n1218 & n2317 ) | ( ~n1266 & n2317 ) ;
  assign n2319 = ~n1219 & n2318 ;
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n1272( .i (x43), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1296( .i (x44), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  assign n2321 = ~n1293 & n1317 ;
  assign n2322 = n2320 & n2321 ;
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2325( .i (n2324), .o (n2325) );
  buffer buf_n2326( .i (n2325), .o (n2326) );
  buffer buf_n2327( .i (n2326), .o (n2327) );
  buffer buf_n2328( .i (n2327), .o (n2328) );
  buffer buf_n2329( .i (n2328), .o (n2329) );
  buffer buf_n2330( .i (n2329), .o (n2330) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  buffer buf_n2307( .i (n2306), .o (n2307) );
  buffer buf_n2308( .i (n2307), .o (n2308) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  assign n2335 = n1197 & n1271 ;
  assign n2336 = ( n1245 & n2308 ) | ( n1245 & n2335 ) | ( n2308 & n2335 ) ;
  assign n2337 = ~n1246 & n2336 ;
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  assign n2343 = ~n1243 & n1270 ;
  assign n2344 = n2316 & n2343 ;
  buffer buf_n2345( .i (n2344), .o (n2345) );
  buffer buf_n2346( .i (n2345), .o (n2346) );
  buffer buf_n2347( .i (n2346), .o (n2347) );
  assign n2352 = n1196 & ~n1270 ;
  assign n2353 = ( n1244 & n2307 ) | ( n1244 & n2352 ) | ( n2307 & n2352 ) ;
  assign n2354 = ~n1245 & n2353 ;
  buffer buf_n2355( .i (n2354), .o (n2355) );
  buffer buf_n2356( .i (n2355), .o (n2356) );
  assign n2358 = n2347 | n2356 ;
  assign n2359 = n2339 | n2358 ;
  buffer buf_n2360( .i (n2359), .o (n2360) );
  assign n2363 = n2330 | n2360 ;
  assign n2364 = n2273 | n2363 ;
  buffer buf_n2365( .i (n2364), .o (n2365) );
  buffer buf_n2366( .i (n2365), .o (n2366) );
  buffer buf_n507( .i (n506), .o (n507) );
  assign n2370 = ( n507 & n1799 ) | ( n507 & n1933 ) | ( n1799 & n1933 ) ;
  assign n2371 = ~n2036 & n2370 ;
  assign n2372 = n1690 & n2371 ;
  buffer buf_n2373( .i (n2372), .o (n2373) );
  assign n2375 = ~n2138 & n2373 ;
  buffer buf_n2376( .i (n2375), .o (n2376) );
  assign n2377 = ~n1761 & n2376 ;
  assign n2378 = n2179 & n2377 ;
  buffer buf_n2379( .i (n2378), .o (n2379) );
  buffer buf_n2380( .i (n2379), .o (n2380) );
  buffer buf_n2381( .i (n2380), .o (n2381) );
  buffer buf_n2382( .i (n2381), .o (n2382) );
  buffer buf_n2383( .i (n2382), .o (n2383) );
  buffer buf_n2384( .i (n2383), .o (n2384) );
  assign n2388 = ( n503 & n523 ) | ( n503 & n1494 ) | ( n523 & n1494 ) ;
  assign n2389 = ~n504 & n2388 ;
  assign n2390 = ~n850 & n2389 ;
  assign n2391 = ( n794 & n2115 ) | ( n794 & n2390 ) | ( n2115 & n2390 ) ;
  assign n2392 = ~n2116 & n2391 ;
  buffer buf_n2393( .i (n2392), .o (n2393) );
  assign n2397 = n2119 & n2393 ;
  buffer buf_n2398( .i (n886), .o (n2398) );
  assign n2399 = n2397 & n2398 ;
  buffer buf_n2400( .i (n2399), .o (n2400) );
  buffer buf_n2401( .i (n2400), .o (n2401) );
  buffer buf_n2402( .i (n2401), .o (n2402) );
  buffer buf_n2403( .i (n2402), .o (n2403) );
  buffer buf_n2404( .i (n2403), .o (n2404) );
  buffer buf_n2405( .i (n2404), .o (n2405) );
  buffer buf_n2406( .i (n2405), .o (n2406) );
  buffer buf_n2407( .i (n2406), .o (n2407) );
  buffer buf_n2408( .i (n2407), .o (n2408) );
  assign n2416 = n524 & ~n624 ;
  buffer buf_n2417( .i (n589), .o (n2417) );
  assign n2418 = ( n2112 & n2416 ) | ( n2112 & n2417 ) | ( n2416 & n2417 ) ;
  assign n2419 = ~n1932 & n2418 ;
  buffer buf_n2420( .i (n2419), .o (n2420) );
  buffer buf_n2421( .i (n2420), .o (n2421) );
  assign n2423 = n794 & n883 ;
  buffer buf_n2424( .i (n2423), .o (n2424) );
  assign n2425 = ( n853 & ~n2420 ) | ( n853 & n2424 ) | ( ~n2420 & n2424 ) ;
  assign n2426 = n2421 & n2425 ;
  assign n2427 = ~n2082 & n2426 ;
  buffer buf_n2428( .i (n2427), .o (n2428) );
  buffer buf_n2429( .i (n2428), .o (n2429) );
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  buffer buf_n2432( .i (n2431), .o (n2432) );
  buffer buf_n2433( .i (n2432), .o (n2433) );
  buffer buf_n2434( .i (n2433), .o (n2434) );
  buffer buf_n2435( .i (n2434), .o (n2435) );
  buffer buf_n666( .i (n665), .o (n666) );
  assign n2444 = ~n623 & n1321 ;
  assign n2445 = n589 & n2444 ;
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n2448( .i (n2447), .o (n2448) );
  buffer buf_n2449( .i (n2448), .o (n2449) );
  buffer buf_n2450( .i (n853), .o (n2450) );
  assign n2451 = n2449 & ~n2450 ;
  assign n2452 = n666 & n2451 ;
  buffer buf_n2453( .i (n2452), .o (n2453) );
  buffer buf_n2455( .i (n1914), .o (n2455) );
  assign n2456 = n2453 & n2455 ;
  assign n2457 = n2065 & n2456 ;
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n2460( .i (n2459), .o (n2460) );
  assign n2465 = n851 & n2446 ;
  assign n2466 = n663 & n2465 ;
  buffer buf_n2467( .i (n2466), .o (n2467) );
  assign n2472 = n2119 & n2467 ;
  assign n2473 = n2398 & n2472 ;
  buffer buf_n2474( .i (n2473), .o (n2474) );
  buffer buf_n2475( .i (n2474), .o (n2475) );
  buffer buf_n2476( .i (n2475), .o (n2476) );
  buffer buf_n2477( .i (n2476), .o (n2477) );
  buffer buf_n2478( .i (n2477), .o (n2478) );
  buffer buf_n84( .i (x1), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  assign n2485 = n99 & ~n588 ;
  buffer buf_n2486( .i (n523), .o (n2486) );
  assign n2487 = ( n557 & n2485 ) | ( n557 & n2486 ) | ( n2485 & n2486 ) ;
  buffer buf_n2488( .i (n2486), .o (n2488) );
  assign n2489 = n2487 & ~n2488 ;
  buffer buf_n2490( .i (n2489), .o (n2490) );
  buffer buf_n2491( .i (n2490), .o (n2491) );
  buffer buf_n2492( .i (n2491), .o (n2492) );
  assign n2493 = ~n1909 & n2492 ;
  buffer buf_n2494( .i (n2493), .o (n2494) );
  assign n2495 = n703 & n2494 ;
  buffer buf_n2496( .i (n1781), .o (n2496) );
  assign n2497 = ( n2455 & n2495 ) | ( n2455 & n2496 ) | ( n2495 & n2496 ) ;
  buffer buf_n2498( .i (n2455), .o (n2498) );
  assign n2499 = n2497 & ~n2498 ;
  buffer buf_n2500( .i (n2499), .o (n2500) );
  buffer buf_n2501( .i (n2500), .o (n2501) );
  assign n2508 = n2478 | n2501 ;
  assign n2509 = n2460 | n2508 ;
  buffer buf_n2510( .i (n2509), .o (n2510) );
  assign n2514 = n2435 | n2510 ;
  assign n2515 = ( ~n2383 & n2408 ) | ( ~n2383 & n2514 ) | ( n2408 & n2514 ) ;
  assign n2516 = n2384 | n2515 ;
  assign n2517 = n1244 & n2307 ;
  buffer buf_n2518( .i (n2517), .o (n2518) );
  buffer buf_n2519( .i (n2518), .o (n2519) );
  buffer buf_n2520( .i (n2519), .o (n2520) );
  buffer buf_n2521( .i (n2520), .o (n2521) );
  buffer buf_n2522( .i (n2521), .o (n2522) );
  buffer buf_n2523( .i (n2522), .o (n2523) );
  buffer buf_n2524( .i (n2523), .o (n2524) );
  assign n2529 = n1172 & n2297 ;
  buffer buf_n2530( .i (n2529), .o (n2530) );
  buffer buf_n2531( .i (n2530), .o (n2531) );
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n2532), .o (n2533) );
  buffer buf_n2534( .i (n2533), .o (n2534) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  buffer buf_n2536( .i (n2535), .o (n2536) );
  buffer buf_n2537( .i (n2536), .o (n2537) );
  buffer buf_n2538( .i (n2537), .o (n2538) );
  buffer buf_n2539( .i (n2538), .o (n2539) );
  buffer buf_n2540( .i (n2539), .o (n2540) );
  buffer buf_n2541( .i (n2540), .o (n2541) );
  buffer buf_n2542( .i (n2541), .o (n2542) );
  buffer buf_n2543( .i (n2542), .o (n2543) );
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n933( .i (x31), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  assign n2547 = n319 & ~n2112 ;
  assign n2548 = ( n526 & ~n591 ) | ( n526 & n2547 ) | ( ~n591 & n2547 ) ;
  buffer buf_n2549( .i (n2488), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  assign n2551 = n2548 & ~n2550 ;
  assign n2552 = n2134 & n2551 ;
  assign n2553 = ( n665 & n2450 ) | ( n665 & n2552 ) | ( n2450 & n2552 ) ;
  buffer buf_n2554( .i (n2450), .o (n2554) );
  assign n2555 = n2553 & ~n2554 ;
  assign n2556 = n1347 & n2555 ;
  buffer buf_n2557( .i (n2556), .o (n2557) );
  buffer buf_n2558( .i (n2557), .o (n2558) );
  buffer buf_n993( .i (x33), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  assign n2565 = ~n1018 & n1198 ;
  assign n2566 = ( n959 & n2558 ) | ( n959 & n2565 ) | ( n2558 & n2565 ) ;
  assign n2567 = ~n960 & n2566 ;
  buffer buf_n2568( .i (n2567), .o (n2568) );
  buffer buf_n2569( .i (n2568), .o (n2569) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n2574( .i (n521), .o (n2574) );
  assign n2575 = n555 & n2574 ;
  assign n2576 = ( n588 & n623 ) | ( n588 & n2575 ) | ( n623 & n2575 ) ;
  assign n2577 = ~n624 & n2576 ;
  buffer buf_n2578( .i (n2577), .o (n2578) );
  buffer buf_n2579( .i (n2578), .o (n2579) );
  buffer buf_n2580( .i (n2579), .o (n2580) );
  buffer buf_n2581( .i (n2580), .o (n2581) );
  assign n2584 = n886 & n2581 ;
  assign n2585 = ( n826 & n2554 ) | ( n826 & n2584 ) | ( n2554 & n2584 ) ;
  assign n2586 = ~n827 & n2585 ;
  assign n2587 = n2455 & n2586 ;
  buffer buf_n2588( .i (n2587), .o (n2588) );
  buffer buf_n2589( .i (n2588), .o (n2589) );
  buffer buf_n2590( .i (n2589), .o (n2590) );
  buffer buf_n2591( .i (n2590), .o (n2591) );
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n2289( .i (n2288), .o (n2289) );
  buffer buf_n2290( .i (n2289), .o (n2290) );
  buffer buf_n2291( .i (n2290), .o (n2291) );
  buffer buf_n2292( .i (n2291), .o (n2292) );
  buffer buf_n2293( .i (n2292), .o (n2293) );
  buffer buf_n2294( .i (n2293), .o (n2294) );
  assign n2599 = n2043 & n2294 ;
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  buffer buf_n2582( .i (n2581), .o (n2582) );
  buffer buf_n2583( .i (n2582), .o (n2583) );
  assign n2606 = n826 & n2082 ;
  assign n2607 = ( n1781 & n2583 ) | ( n1781 & n2606 ) | ( n2583 & n2606 ) ;
  assign n2608 = ~n2496 & n2607 ;
  buffer buf_n2609( .i (n2608), .o (n2609) );
  buffer buf_n2610( .i (n2609), .o (n2610) );
  buffer buf_n2611( .i (n2610), .o (n2611) );
  assign n2619 = n2601 | n2611 ;
  assign n2620 = n2591 | n2619 ;
  assign n2621 = n2569 | n2620 ;
  assign n2622 = ( ~n2523 & n2545 ) | ( ~n2523 & n2621 ) | ( n2545 & n2621 ) ;
  assign n2623 = n2524 | n2622 ;
  buffer buf_n2624( .i (n885), .o (n2624) );
  assign n2625 = n2581 & ~n2624 ;
  assign n2626 = ( n826 & n2554 ) | ( n826 & n2625 ) | ( n2554 & n2625 ) ;
  assign n2627 = ~n827 & n2626 ;
  buffer buf_n2628( .i (n2627), .o (n2628) );
  assign n2631 = ~n2498 & n2628 ;
  buffer buf_n2632( .i (n2631), .o (n2632) );
  buffer buf_n2633( .i (n2632), .o (n2633) );
  buffer buf_n2634( .i (n2633), .o (n2634) );
  buffer buf_n2635( .i (n2634), .o (n2635) );
  buffer buf_n2636( .i (n2635), .o (n2636) );
  buffer buf_n2637( .i (n2636), .o (n2637) );
  buffer buf_n2638( .i (n587), .o (n2638) );
  assign n2639 = ( n523 & n1603 ) | ( n523 & n2638 ) | ( n1603 & n2638 ) ;
  assign n2640 = ~n589 & n2639 ;
  buffer buf_n2641( .i (n2640), .o (n2641) );
  assign n2650 = n851 & n2641 ;
  assign n2651 = n795 & n2650 ;
  buffer buf_n2652( .i (n2651), .o (n2652) );
  buffer buf_n2653( .i (n920), .o (n2653) );
  assign n2654 = n2652 & ~n2653 ;
  assign n2655 = n2398 & n2654 ;
  buffer buf_n2656( .i (n2655), .o (n2656) );
  buffer buf_n2657( .i (n2656), .o (n2657) );
  buffer buf_n2658( .i (n2657), .o (n2658) );
  buffer buf_n2659( .i (n2658), .o (n2659) );
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2660), .o (n2661) );
  buffer buf_n2662( .i (n2661), .o (n2662) );
  buffer buf_n2663( .i (n2662), .o (n2663) );
  buffer buf_n2642( .i (n2641), .o (n2642) );
  buffer buf_n2643( .i (n2642), .o (n2643) );
  buffer buf_n2644( .i (n2643), .o (n2644) );
  buffer buf_n2645( .i (n2644), .o (n2645) );
  buffer buf_n2646( .i (n2645), .o (n2646) );
  buffer buf_n2647( .i (n2646), .o (n2647) );
  buffer buf_n2666( .i (n2398), .o (n2666) );
  assign n2667 = ( n1899 & ~n2646 ) | ( n1899 & n2666 ) | ( ~n2646 & n2666 ) ;
  assign n2668 = n2647 & n2667 ;
  buffer buf_n2669( .i (n2668), .o (n2669) );
  buffer buf_n2670( .i (n2669), .o (n2670) );
  buffer buf_n2671( .i (n2670), .o (n2671) );
  buffer buf_n2672( .i (n2671), .o (n2672) );
  buffer buf_n2673( .i (n2672), .o (n2673) );
  buffer buf_n2676( .i (n852), .o (n2676) );
  assign n2677 = n2643 & ~n2676 ;
  assign n2678 = n797 & n2677 ;
  buffer buf_n2679( .i (n2678), .o (n2679) );
  assign n2681 = n1914 & n2679 ;
  assign n2682 = n2496 & n2681 ;
  buffer buf_n2683( .i (n2682), .o (n2683) );
  buffer buf_n2684( .i (n2683), .o (n2684) );
  buffer buf_n2685( .i (n2684), .o (n2685) );
  buffer buf_n2686( .i (n2685), .o (n2686) );
  buffer buf_n2648( .i (n2647), .o (n2648) );
  buffer buf_n2649( .i (n2648), .o (n2649) );
  buffer buf_n2692( .i (n2496), .o (n2692) );
  assign n2693 = ( n1916 & ~n2648 ) | ( n1916 & n2692 ) | ( ~n2648 & n2692 ) ;
  assign n2694 = n2649 & n2693 ;
  buffer buf_n2695( .i (n2694), .o (n2695) );
  buffer buf_n2696( .i (n2695), .o (n2696) );
  assign n2703 = n2686 | n2696 ;
  assign n2704 = n2673 | n2703 ;
  assign n2705 = n2663 | n2704 ;
  assign n2706 = n2637 | n2705 ;
  assign n2707 = n2623 | n2706 ;
  assign n2708 = ( ~n2365 & n2516 ) | ( ~n2365 & n2707 ) | ( n2516 & n2707 ) ;
  assign n2709 = n2366 | n2708 ;
  buffer buf_n2710( .i (n2709), .o (n2710) );
  buffer buf_n2711( .i (n2710), .o (n2711) );
  buffer buf_n2712( .i (n2550), .o (n2712) );
  assign n2713 = ( n1395 & n1776 ) | ( n1395 & ~n2712 ) | ( n1776 & ~n2712 ) ;
  assign n2714 = n2023 & n2713 ;
  buffer buf_n2715( .i (n2714), .o (n2715) );
  buffer buf_n2716( .i (n2082), .o (n2716) );
  assign n2717 = n2715 & ~n2716 ;
  buffer buf_n2718( .i (n2666), .o (n2718) );
  assign n2719 = n2717 & n2718 ;
  buffer buf_n2720( .i (n2719), .o (n2720) );
  buffer buf_n2721( .i (n2720), .o (n2721) );
  buffer buf_n2722( .i (n2721), .o (n2722) );
  buffer buf_n2723( .i (n2722), .o (n2723) );
  buffer buf_n2724( .i (n2723), .o (n2724) );
  buffer buf_n2725( .i (n2724), .o (n2725) );
  buffer buf_n2726( .i (n2725), .o (n2726) );
  buffer buf_n2727( .i (n2726), .o (n2727) );
  buffer buf_n2728( .i (n2727), .o (n2728) );
  buffer buf_n2729( .i (n2728), .o (n2729) );
  buffer buf_n2730( .i (n2729), .o (n2730) );
  assign n2731 = n759 & n883 ;
  buffer buf_n2732( .i (n2731), .o (n2732) );
  buffer buf_n2733( .i (n556), .o (n2733) );
  assign n2734 = ( n362 & n1796 ) | ( n362 & n2733 ) | ( n1796 & n2733 ) ;
  assign n2735 = ~n2112 & n2734 ;
  assign n2736 = n2115 & n2735 ;
  buffer buf_n2737( .i (n2736), .o (n2737) );
  assign n2738 = ( n2676 & n2732 ) | ( n2676 & n2737 ) | ( n2732 & n2737 ) ;
  assign n2739 = ~n2450 & n2738 ;
  buffer buf_n2740( .i (n2739), .o (n2740) );
  buffer buf_n2741( .i (n2740), .o (n2741) );
  buffer buf_n2742( .i (n2741), .o (n2742) );
  buffer buf_n2743( .i (n2742), .o (n2743) );
  buffer buf_n2744( .i (n2743), .o (n2744) );
  buffer buf_n2745( .i (n2744), .o (n2745) );
  buffer buf_n2746( .i (n2745), .o (n2746) );
  buffer buf_n2747( .i (n2746), .o (n2747) );
  buffer buf_n2748( .i (n2747), .o (n2748) );
  buffer buf_n2749( .i (n2748), .o (n2749) );
  buffer buf_n2750( .i (n2749), .o (n2750) );
  buffer buf_n2751( .i (n2750), .o (n2751) );
  assign n2753 = ( n362 & n1495 ) | ( n362 & n2486 ) | ( n1495 & n2486 ) ;
  assign n2754 = ~n363 & n2753 ;
  assign n2755 = n2115 & n2754 ;
  buffer buf_n2756( .i (n2755), .o (n2756) );
  assign n2757 = ( n2424 & n2676 ) | ( n2424 & n2756 ) | ( n2676 & n2756 ) ;
  buffer buf_n2758( .i (n2676), .o (n2758) );
  assign n2759 = n2757 & ~n2758 ;
  buffer buf_n2760( .i (n2759), .o (n2760) );
  buffer buf_n2761( .i (n2760), .o (n2761) );
  buffer buf_n2762( .i (n2761), .o (n2762) );
  buffer buf_n2763( .i (n2762), .o (n2763) );
  buffer buf_n2764( .i (n2763), .o (n2764) );
  buffer buf_n2765( .i (n2764), .o (n2765) );
  buffer buf_n2766( .i (n2765), .o (n2766) );
  buffer buf_n2767( .i (n2766), .o (n2767) );
  buffer buf_n2768( .i (n2767), .o (n2768) );
  buffer buf_n2769( .i (n2768), .o (n2769) );
  buffer buf_n2770( .i (n2769), .o (n2770) );
  buffer buf_n2771( .i (n2770), .o (n2771) );
  assign n2772 = n927 & ~n2764 ;
  buffer buf_n2773( .i (n2772), .o (n2773) );
  buffer buf_n2774( .i (n2773), .o (n2774) );
  buffer buf_n2775( .i (n2774), .o (n2775) );
  buffer buf_n2776( .i (n2775), .o (n2776) );
  buffer buf_n2777( .i (n2776), .o (n2777) );
  buffer buf_n2778( .i (n2777), .o (n2778) );
  assign n2779 = ( n2751 & n2771 ) | ( n2751 & ~n2778 ) | ( n2771 & ~n2778 ) ;
  buffer buf_n2780( .i (n852), .o (n2780) );
  assign n2781 = ( n2424 & n2737 ) | ( n2424 & n2780 ) | ( n2737 & n2780 ) ;
  assign n2782 = ~n2758 & n2781 ;
  buffer buf_n2783( .i (n2782), .o (n2783) );
  buffer buf_n2784( .i (n2783), .o (n2784) );
  buffer buf_n2785( .i (n2784), .o (n2785) );
  buffer buf_n2786( .i (n2785), .o (n2786) );
  buffer buf_n2787( .i (n2786), .o (n2787) );
  buffer buf_n2788( .i (n2787), .o (n2788) );
  buffer buf_n2789( .i (n2788), .o (n2789) );
  buffer buf_n2790( .i (n2789), .o (n2790) );
  buffer buf_n2791( .i (n2790), .o (n2791) );
  buffer buf_n2792( .i (n2791), .o (n2792) );
  buffer buf_n2793( .i (n2792), .o (n2793) );
  buffer buf_n2794( .i (n2793), .o (n2794) );
  buffer buf_n667( .i (n666), .o (n667) );
  assign n2795 = n667 & n2494 ;
  buffer buf_n2796( .i (n2716), .o (n2796) );
  assign n2797 = ( n2718 & n2795 ) | ( n2718 & n2796 ) | ( n2795 & n2796 ) ;
  assign n2798 = ~n2498 & n2797 ;
  buffer buf_n2799( .i (n2798), .o (n2799) );
  buffer buf_n2800( .i (n2799), .o (n2800) );
  buffer buf_n2801( .i (n2800), .o (n2801) );
  buffer buf_n2802( .i (n2801), .o (n2802) );
  buffer buf_n2803( .i (n2802), .o (n2803) );
  buffer buf_n2804( .i (n2803), .o (n2804) );
  buffer buf_n2805( .i (n2804), .o (n2805) );
  buffer buf_n2808( .i (n625), .o (n2808) );
  assign n2809 = ( n1497 & n2549 ) | ( n1497 & ~n2808 ) | ( n2549 & ~n2808 ) ;
  assign n2810 = ~n2550 & n2809 ;
  buffer buf_n2811( .i (n2810), .o (n2811) );
  buffer buf_n2812( .i (n2811), .o (n2812) );
  buffer buf_n2813( .i (n2812), .o (n2813) );
  buffer buf_n2814( .i (n2813), .o (n2814) );
  assign n2819 = n2796 & n2814 ;
  buffer buf_n2820( .i (n1861), .o (n2820) );
  assign n2821 = ( n2692 & n2819 ) | ( n2692 & n2820 ) | ( n2819 & n2820 ) ;
  buffer buf_n2822( .i (n2820), .o (n2822) );
  assign n2823 = n2821 & ~n2822 ;
  buffer buf_n2824( .i (n2823), .o (n2824) );
  buffer buf_n2825( .i (n2824), .o (n2825) );
  buffer buf_n2826( .i (n2825), .o (n2826) );
  buffer buf_n2827( .i (n2826), .o (n2827) );
  buffer buf_n2828( .i (n2827), .o (n2828) );
  assign n2833 = n2138 & n2813 ;
  assign n2834 = ( n2718 & n2796 ) | ( n2718 & n2833 ) | ( n2796 & n2833 ) ;
  assign n2835 = ~n2498 & n2834 ;
  buffer buf_n2836( .i (n2835), .o (n2836) );
  buffer buf_n2837( .i (n2836), .o (n2837) );
  buffer buf_n2838( .i (n2837), .o (n2838) );
  buffer buf_n2839( .i (n2838), .o (n2839) );
  buffer buf_n2840( .i (n2839), .o (n2840) );
  buffer buf_n2845( .i (n2733), .o (n2845) );
  buffer buf_n2846( .i (n2845), .o (n2846) );
  buffer buf_n2847( .i (n2846), .o (n2847) );
  buffer buf_n2848( .i (n2808), .o (n2848) );
  assign n2849 = n2847 | n2848 ;
  assign n2850 = ( n1776 & ~n2712 ) | ( n1776 & n2849 ) | ( ~n2712 & n2849 ) ;
  assign n2851 = n2023 | n2850 ;
  buffer buf_n2852( .i (n2851), .o (n2852) );
  assign n2854 = n2716 & ~n2852 ;
  buffer buf_n2855( .i (n2554), .o (n2855) );
  buffer buf_n2856( .i (n2855), .o (n2856) );
  assign n2857 = ( n2718 & n2854 ) | ( n2718 & n2856 ) | ( n2854 & n2856 ) ;
  assign n2858 = ~n2820 & n2857 ;
  buffer buf_n2859( .i (n2858), .o (n2859) );
  buffer buf_n2860( .i (n2859), .o (n2860) );
  assign n2866 = ~n2852 & n2855 ;
  buffer buf_n2867( .i (n2666), .o (n2867) );
  assign n2868 = ( n2796 & n2866 ) | ( n2796 & n2867 ) | ( n2866 & n2867 ) ;
  buffer buf_n2869( .i (n2716), .o (n2869) );
  buffer buf_n2870( .i (n2869), .o (n2870) );
  assign n2871 = n2868 & ~n2870 ;
  buffer buf_n2872( .i (n2871), .o (n2872) );
  buffer buf_n2873( .i (n2872), .o (n2873) );
  assign n2880 = n2860 | n2873 ;
  buffer buf_n2881( .i (n2880), .o (n2881) );
  buffer buf_n2882( .i (n2881), .o (n2882) );
  assign n2883 = n2840 | n2882 ;
  assign n2884 = ( ~n2804 & n2828 ) | ( ~n2804 & n2883 ) | ( n2828 & n2883 ) ;
  assign n2885 = n2805 | n2884 ;
  assign n2886 = n2794 | n2885 ;
  assign n2887 = ( ~n2729 & n2779 ) | ( ~n2729 & n2886 ) | ( n2779 & n2886 ) ;
  assign n2888 = n2730 | n2887 ;
  assign n2889 = n1339 & n2162 ;
  assign n2890 = ( n2264 & n2855 ) | ( n2264 & n2889 ) | ( n2855 & n2889 ) ;
  assign n2891 = ~n2856 & n2890 ;
  buffer buf_n2892( .i (n2891), .o (n2892) );
  assign n2895 = ~n926 & n2892 ;
  buffer buf_n2896( .i (n2895), .o (n2896) );
  buffer buf_n2897( .i (n2896), .o (n2897) );
  buffer buf_n2898( .i (n2897), .o (n2898) );
  buffer buf_n2899( .i (n2898), .o (n2899) );
  buffer buf_n2900( .i (n2899), .o (n2900) );
  buffer buf_n2901( .i (n2900), .o (n2901) );
  buffer buf_n2902( .i (n2901), .o (n2902) );
  buffer buf_n2903( .i (n2902), .o (n2903) );
  assign n2904 = ( n1373 & n2488 ) | ( n1373 & n2845 ) | ( n2488 & n2845 ) ;
  assign n2905 = ~n2846 & n2904 ;
  buffer buf_n2906( .i (n2905), .o (n2906) );
  assign n2911 = ~n920 & n2906 ;
  assign n2912 = ( n2624 & n2758 ) | ( n2624 & n2911 ) | ( n2758 & n2911 ) ;
  buffer buf_n2913( .i (n2758), .o (n2913) );
  assign n2914 = n2912 & ~n2913 ;
  buffer buf_n2915( .i (n2914), .o (n2915) );
  buffer buf_n2916( .i (n2915), .o (n2916) );
  buffer buf_n2917( .i (n2916), .o (n2917) );
  buffer buf_n2918( .i (n2917), .o (n2918) );
  buffer buf_n2919( .i (n2918), .o (n2919) );
  buffer buf_n2920( .i (n2919), .o (n2920) );
  buffer buf_n2921( .i (n2920), .o (n2921) );
  buffer buf_n2922( .i (n2921), .o (n2922) );
  buffer buf_n2923( .i (n2922), .o (n2923) );
  buffer buf_n2924( .i (n2923), .o (n2924) );
  buffer buf_n2925( .i (n2924), .o (n2925) );
  assign n2926 = n1339 & n2913 ;
  buffer buf_n2927( .i (n2653), .o (n2927) );
  buffer buf_n2928( .i (n2927), .o (n2928) );
  assign n2929 = ( n2666 & n2926 ) | ( n2666 & n2928 ) | ( n2926 & n2928 ) ;
  assign n2930 = ~n2869 & n2929 ;
  buffer buf_n2931( .i (n2930), .o (n2931) );
  buffer buf_n2932( .i (n2931), .o (n2932) );
  buffer buf_n2933( .i (n2932), .o (n2933) );
  buffer buf_n2934( .i (n2933), .o (n2934) );
  buffer buf_n2935( .i (n2934), .o (n2935) );
  buffer buf_n2936( .i (n2935), .o (n2936) );
  buffer buf_n2937( .i (n2936), .o (n2937) );
  buffer buf_n2938( .i (n2937), .o (n2938) );
  assign n2939 = ( n2732 & n2756 ) | ( n2732 & n2780 ) | ( n2756 & n2780 ) ;
  buffer buf_n2940( .i (n2780), .o (n2940) );
  assign n2941 = n2939 & ~n2940 ;
  buffer buf_n2942( .i (n2941), .o (n2942) );
  assign n2948 = ~n2928 & n2942 ;
  buffer buf_n2949( .i (n2948), .o (n2949) );
  buffer buf_n2950( .i (n2949), .o (n2950) );
  buffer buf_n2951( .i (n2950), .o (n2951) );
  buffer buf_n2952( .i (n2951), .o (n2952) );
  buffer buf_n2953( .i (n2952), .o (n2953) );
  assign n2956 = n625 & n2488 ;
  buffer buf_n2957( .i (n2417), .o (n2957) );
  assign n2958 = ( n2846 & n2956 ) | ( n2846 & n2957 ) | ( n2956 & n2957 ) ;
  assign n2959 = ~n2847 & n2958 ;
  assign n2960 = ( n2261 & n2780 ) | ( n2261 & n2959 ) | ( n2780 & n2959 ) ;
  assign n2961 = ~n2940 & n2960 ;
  buffer buf_n2962( .i (n2961), .o (n2962) );
  buffer buf_n2963( .i (n2962), .o (n2963) );
  buffer buf_n2964( .i (n2963), .o (n2964) );
  assign n2968 = ~n2870 & n2964 ;
  buffer buf_n2969( .i (n2968), .o (n2969) );
  buffer buf_n2970( .i (n2969), .o (n2970) );
  buffer buf_n2971( .i (n2970), .o (n2971) );
  assign n2976 = n2953 | n2971 ;
  buffer buf_n2977( .i (n2976), .o (n2977) );
  buffer buf_n2978( .i (n2977), .o (n2978) );
  buffer buf_n2979( .i (n2978), .o (n2979) );
  assign n2980 = n2938 | n2979 ;
  assign n2981 = ( ~n2902 & n2925 ) | ( ~n2902 & n2980 ) | ( n2925 & n2980 ) ;
  assign n2982 = n2903 | n2981 ;
  assign n2983 = n2490 & n2848 ;
  buffer buf_n2984( .i (n2983), .o (n2984) );
  assign n2985 = ( n701 & n2940 ) | ( n701 & n2984 ) | ( n2940 & n2984 ) ;
  assign n2986 = ~n2913 & n2985 ;
  assign n2987 = n1347 & n2986 ;
  buffer buf_n2988( .i (n2987), .o (n2988) );
  buffer buf_n2989( .i (n2988), .o (n2989) );
  buffer buf_n2990( .i (n2989), .o (n2990) );
  buffer buf_n2991( .i (n2990), .o (n2991) );
  buffer buf_n2992( .i (n2991), .o (n2992) );
  buffer buf_n2993( .i (n2992), .o (n2993) );
  buffer buf_n2994( .i (n2993), .o (n2994) );
  buffer buf_n2995( .i (n2994), .o (n2995) );
  buffer buf_n2996( .i (n2995), .o (n2996) );
  buffer buf_n2997( .i (n2996), .o (n2997) );
  buffer buf_n2998( .i (n2997), .o (n2998) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2999( .i (n2574), .o (n2999) );
  assign n3000 = ( n2248 & n2638 ) | ( n2248 & n2999 ) | ( n2638 & n2999 ) ;
  assign n3001 = ~n2486 & n3000 ;
  buffer buf_n3002( .i (n3001), .o (n3002) );
  buffer buf_n3003( .i (n3002), .o (n3003) );
  buffer buf_n3004( .i (n3003), .o (n3004) );
  buffer buf_n3005( .i (n3004), .o (n3005) );
  assign n3014 = ~n2653 & n3005 ;
  buffer buf_n3015( .i (n2624), .o (n3015) );
  assign n3016 = ( n798 & n3014 ) | ( n798 & n3015 ) | ( n3014 & n3015 ) ;
  assign n3017 = ~n799 & n3016 ;
  buffer buf_n3018( .i (n3017), .o (n3018) );
  assign n3027 = n797 & n3005 ;
  assign n3028 = ( n2927 & n3015 ) | ( n2927 & n3027 ) | ( n3015 & n3027 ) ;
  assign n3029 = ~n2928 & n3028 ;
  buffer buf_n3030( .i (n3029), .o (n3030) );
  assign n3038 = n3018 | n3030 ;
  buffer buf_n3039( .i (n3038), .o (n3039) );
  buffer buf_n3040( .i (n3039), .o (n3040) );
  buffer buf_n3041( .i (n3040), .o (n3041) );
  buffer buf_n3042( .i (n3041), .o (n3042) );
  buffer buf_n3043( .i (n3042), .o (n3043) );
  buffer buf_n3044( .i (n3043), .o (n3044) );
  buffer buf_n3045( .i (n3044), .o (n3045) );
  buffer buf_n3046( .i (n3045), .o (n3046) );
  buffer buf_n3006( .i (n3005), .o (n3006) );
  buffer buf_n3007( .i (n3006), .o (n3007) );
  buffer buf_n3008( .i (n3007), .o (n3008) );
  buffer buf_n3048( .i (n918), .o (n3048) );
  buffer buf_n3049( .i (n3048), .o (n3049) );
  assign n3050 = n796 & n3049 ;
  buffer buf_n3051( .i (n3050), .o (n3051) );
  buffer buf_n3052( .i (n3051), .o (n3052) );
  buffer buf_n3053( .i (n3015), .o (n3053) );
  assign n3054 = ( ~n3007 & n3052 ) | ( ~n3007 & n3053 ) | ( n3052 & n3053 ) ;
  assign n3055 = n3008 & n3054 ;
  buffer buf_n3056( .i (n3055), .o (n3056) );
  buffer buf_n3057( .i (n3056), .o (n3057) );
  buffer buf_n3058( .i (n3057), .o (n3058) );
  buffer buf_n3059( .i (n3058), .o (n3059) );
  buffer buf_n3060( .i (n3059), .o (n3060) );
  buffer buf_n3061( .i (n3060), .o (n3061) );
  buffer buf_n3062( .i (n3061), .o (n3062) );
  buffer buf_n3063( .i (n3062), .o (n3063) );
  assign n3068 = ( n665 & n2940 ) | ( n665 & n2984 ) | ( n2940 & n2984 ) ;
  assign n3069 = ~n2913 & n3068 ;
  assign n3070 = n1347 & n3069 ;
  buffer buf_n3071( .i (n3070), .o (n3071) );
  assign n3080 = n731 & n3005 ;
  assign n3081 = ( n2927 & n3015 ) | ( n2927 & n3080 ) | ( n3015 & n3080 ) ;
  assign n3082 = ~n2928 & n3081 ;
  buffer buf_n3083( .i (n3082), .o (n3083) );
  assign n3095 = n3071 | n3083 ;
  buffer buf_n3096( .i (n3095), .o (n3096) );
  buffer buf_n3097( .i (n3096), .o (n3097) );
  buffer buf_n3098( .i (n3097), .o (n3098) );
  buffer buf_n3099( .i (n3098), .o (n3099) );
  buffer buf_n3100( .i (n3099), .o (n3100) );
  buffer buf_n3101( .i (n3100), .o (n3101) );
  buffer buf_n3102( .i (n3101), .o (n3102) );
  assign n3103 = n3063 | n3102 ;
  assign n3104 = ( ~n2997 & n3046 ) | ( ~n2997 & n3103 ) | ( n3046 & n3103 ) ;
  assign n3105 = n2998 | n3104 ;
  assign n3106 = n2982 | n3105 ;
  assign n3107 = ( ~n2710 & n2888 ) | ( ~n2710 & n3106 ) | ( n2888 & n3106 ) ;
  assign n3108 = n2711 | n3107 ;
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  assign n3109 = ~n1318 & n2320 ;
  assign n3110 = n1295 & n3109 ;
  buffer buf_n3111( .i (n3110), .o (n3111) );
  buffer buf_n3112( .i (n3111), .o (n3112) );
  buffer buf_n3113( .i (n3112), .o (n3113) );
  buffer buf_n3114( .i (n3113), .o (n3114) );
  buffer buf_n3115( .i (n3114), .o (n3115) );
  buffer buf_n3116( .i (n3115), .o (n3116) );
  buffer buf_n3117( .i (n3116), .o (n3117) );
  buffer buf_n3118( .i (n3117), .o (n3118) );
  buffer buf_n3119( .i (n3118), .o (n3119) );
  buffer buf_n3120( .i (n3119), .o (n3120) );
  buffer buf_n3121( .i (n3120), .o (n3121) );
  buffer buf_n166( .i (n165), .o (n166) );
  assign n3122 = ( n165 & n1799 ) | ( n165 & n2847 ) | ( n1799 & n2847 ) ;
  assign n3123 = ~n166 & n3122 ;
  assign n3124 = ~n2624 & n3123 ;
  buffer buf_n3125( .i (n825), .o (n3125) );
  assign n3126 = ( n1910 & n3124 ) | ( n1910 & n3125 ) | ( n3124 & n3125 ) ;
  assign n3127 = ~n2026 & n3126 ;
  assign n3128 = ~n2869 & n3127 ;
  buffer buf_n3129( .i (n3128), .o (n3129) );
  buffer buf_n3130( .i (n3129), .o (n3130) );
  buffer buf_n3131( .i (n3130), .o (n3131) );
  buffer buf_n3132( .i (n3131), .o (n3132) );
  buffer buf_n3133( .i (n3132), .o (n3133) );
  assign n3139 = n2635 | n3133 ;
  buffer buf_n3140( .i (n3139), .o (n3140) );
  buffer buf_n3141( .i (n3140), .o (n3141) );
  buffer buf_n3142( .i (n3141), .o (n3142) );
  buffer buf_n2612( .i (n2611), .o (n2612) );
  buffer buf_n2613( .i (n2612), .o (n2613) );
  buffer buf_n2614( .i (n2613), .o (n2614) );
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  buffer buf_n2374( .i (n2373), .o (n2374) );
  buffer buf_n3143( .i (n850), .o (n3143) );
  buffer buf_n3144( .i (n3143), .o (n3144) );
  buffer buf_n3145( .i (n3144), .o (n3145) );
  assign n3146 = ~n3049 & n3145 ;
  buffer buf_n3147( .i (n3146), .o (n3147) );
  buffer buf_n3148( .i (n3147), .o (n3148) );
  buffer buf_n3149( .i (n3148), .o (n3149) );
  assign n3154 = ( n2374 & n2867 ) | ( n2374 & n3149 ) | ( n2867 & n3149 ) ;
  assign n3155 = ~n2692 & n3154 ;
  buffer buf_n3156( .i (n3155), .o (n3156) );
  buffer buf_n3157( .i (n3156), .o (n3157) );
  buffer buf_n3158( .i (n3157), .o (n3158) );
  buffer buf_n3159( .i (n3158), .o (n3159) );
  buffer buf_n3160( .i (n3159), .o (n3160) );
  buffer buf_n2461( .i (n2460), .o (n2461) );
  buffer buf_n3165( .i (n885), .o (n3165) );
  assign n3166 = n2652 & ~n3165 ;
  assign n3167 = ~n2927 & n3166 ;
  buffer buf_n3168( .i (n3167), .o (n3168) );
  buffer buf_n3169( .i (n3168), .o (n3169) );
  buffer buf_n3170( .i (n3169), .o (n3170) );
  buffer buf_n3171( .i (n3170), .o (n3171) );
  buffer buf_n3172( .i (n3171), .o (n3172) );
  assign n3178 = n2685 | n3172 ;
  buffer buf_n3179( .i (n3178), .o (n3179) );
  assign n3182 = n2461 | n3179 ;
  assign n3183 = ( ~n2382 & n3160 ) | ( ~n2382 & n3182 ) | ( n3160 & n3182 ) ;
  assign n3184 = n2383 | n3183 ;
  assign n3185 = n2616 | n3184 ;
  assign n3186 = ( ~n3120 & n3142 ) | ( ~n3120 & n3185 ) | ( n3142 & n3185 ) ;
  assign n3187 = n3121 | n3186 ;
  buffer buf_n3188( .i (n3187), .o (n3188) );
  buffer buf_n3189( .i (n3188), .o (n3189) );
  buffer buf_n2829( .i (n2828), .o (n2829) );
  buffer buf_n2830( .i (n2829), .o (n2830) );
  buffer buf_n2831( .i (n2830), .o (n2831) );
  buffer buf_n2832( .i (n2831), .o (n2832) );
  buffer buf_n2841( .i (n2840), .o (n2841) );
  buffer buf_n2842( .i (n2841), .o (n2842) );
  buffer buf_n2843( .i (n2842), .o (n2843) );
  buffer buf_n2844( .i (n2843), .o (n2844) );
  buffer buf_n2874( .i (n2873), .o (n2874) );
  buffer buf_n2875( .i (n2874), .o (n2875) );
  buffer buf_n2876( .i (n2875), .o (n2876) );
  buffer buf_n2877( .i (n2876), .o (n2877) );
  buffer buf_n2878( .i (n2877), .o (n2878) );
  buffer buf_n2879( .i (n2878), .o (n2879) );
  buffer buf_n2861( .i (n2860), .o (n2861) );
  buffer buf_n2862( .i (n2861), .o (n2862) );
  buffer buf_n2863( .i (n2862), .o (n2863) );
  buffer buf_n2864( .i (n2863), .o (n2864) );
  buffer buf_n2865( .i (n2864), .o (n2865) );
  assign n3190 = n2727 | n2865 ;
  assign n3191 = n2879 | n3190 ;
  assign n3192 = n2844 | n3191 ;
  assign n3193 = n2832 | n3192 ;
  buffer buf_n3194( .i (n2870), .o (n3194) );
  assign n3195 = n2892 & n3194 ;
  buffer buf_n3196( .i (n3195), .o (n3196) );
  buffer buf_n3197( .i (n3196), .o (n3197) );
  buffer buf_n3198( .i (n3197), .o (n3198) );
  buffer buf_n3199( .i (n3198), .o (n3199) );
  buffer buf_n3200( .i (n3199), .o (n3200) );
  assign n3202 = ( ~n1341 & n1576 ) | ( ~n1341 & n2867 ) | ( n1576 & n2867 ) ;
  assign n3203 = n1342 & n3202 ;
  buffer buf_n3204( .i (n3203), .o (n3204) );
  buffer buf_n3205( .i (n3204), .o (n3205) );
  buffer buf_n3206( .i (n3205), .o (n3206) );
  assign n3209 = n2897 | n3206 ;
  assign n3210 = n2935 | n3209 ;
  buffer buf_n2907( .i (n2906), .o (n2907) );
  assign n3211 = n2653 & n2907 ;
  buffer buf_n3212( .i (n3145), .o (n3212) );
  buffer buf_n3213( .i (n3212), .o (n3213) );
  buffer buf_n3214( .i (n3165), .o (n3214) );
  assign n3215 = ( n3211 & n3213 ) | ( n3211 & n3214 ) | ( n3213 & n3214 ) ;
  assign n3216 = ~n2855 & n3215 ;
  buffer buf_n3217( .i (n3216), .o (n3217) );
  buffer buf_n3218( .i (n3217), .o (n3218) );
  buffer buf_n3219( .i (n3218), .o (n3219) );
  buffer buf_n3220( .i (n3219), .o (n3220) );
  buffer buf_n3221( .i (n3220), .o (n3221) );
  buffer buf_n2943( .i (n2942), .o (n2943) );
  buffer buf_n2944( .i (n2943), .o (n2944) );
  buffer buf_n2945( .i (n2944), .o (n2945) );
  buffer buf_n2946( .i (n2945), .o (n2946) );
  buffer buf_n2947( .i (n2946), .o (n2947) );
  buffer buf_n2965( .i (n2964), .o (n2965) );
  buffer buf_n2966( .i (n2965), .o (n2966) );
  buffer buf_n2967( .i (n2966), .o (n2967) );
  assign n3222 = n2947 | n2967 ;
  assign n3223 = n3221 | n3222 ;
  assign n3224 = n2921 | n3223 ;
  assign n3225 = ( ~n3199 & n3210 ) | ( ~n3199 & n3224 ) | ( n3210 & n3224 ) ;
  assign n3226 = n3200 | n3225 ;
  buffer buf_n3227( .i (n3226), .o (n3227) );
  buffer buf_n3228( .i (n3227), .o (n3228) );
  buffer buf_n3084( .i (n3083), .o (n3084) );
  buffer buf_n3085( .i (n3084), .o (n3085) );
  assign n3229 = n3057 | n3085 ;
  buffer buf_n3230( .i (n3229), .o (n3230) );
  buffer buf_n3231( .i (n3230), .o (n3231) );
  buffer buf_n3232( .i (n3231), .o (n3232) );
  buffer buf_n3233( .i (n3232), .o (n3233) );
  buffer buf_n3234( .i (n3233), .o (n3234) );
  buffer buf_n3235( .i (n3234), .o (n3235) );
  assign n3236 = n700 & n1326 ;
  assign n3237 = ( n1909 & n2161 ) | ( n1909 & n3236 ) | ( n2161 & n3236 ) ;
  assign n3238 = ~n2162 & n3237 ;
  buffer buf_n3239( .i (n3049), .o (n3239) );
  buffer buf_n3240( .i (n3239), .o (n3240) );
  buffer buf_n3241( .i (n3240), .o (n3241) );
  assign n3242 = n3238 & ~n3241 ;
  assign n3243 = ( n2856 & n2867 ) | ( n2856 & n3242 ) | ( n2867 & n3242 ) ;
  assign n3244 = ~n2820 & n3243 ;
  buffer buf_n3245( .i (n3244), .o (n3245) );
  buffer buf_n3246( .i (n3245), .o (n3246) );
  buffer buf_n3247( .i (n3246), .o (n3247) );
  buffer buf_n3248( .i (n3247), .o (n3248) );
  buffer buf_n3249( .i (n3248), .o (n3249) );
  assign n3251 = n663 & n1325 ;
  buffer buf_n3252( .i (n1874), .o (n3252) );
  assign n3253 = ( n2134 & n3251 ) | ( n2134 & n3252 ) | ( n3251 & n3252 ) ;
  assign n3254 = ~n2161 & n3253 ;
  assign n3255 = ~n3240 & n3254 ;
  buffer buf_n3256( .i (n3213), .o (n3256) );
  assign n3257 = ( n3053 & n3255 ) | ( n3053 & n3256 ) | ( n3255 & n3256 ) ;
  assign n3258 = ~n2856 & n3257 ;
  buffer buf_n3259( .i (n3258), .o (n3259) );
  buffer buf_n3260( .i (n3259), .o (n3260) );
  buffer buf_n3261( .i (n3260), .o (n3261) );
  buffer buf_n3262( .i (n3261), .o (n3262) );
  buffer buf_n3263( .i (n3262), .o (n3263) );
  buffer buf_n3072( .i (n3071), .o (n3072) );
  buffer buf_n3073( .i (n3072), .o (n3073) );
  buffer buf_n3009( .i (n3008), .o (n3009) );
  buffer buf_n3267( .i (n3053), .o (n3267) );
  assign n3268 = ( n1407 & ~n3008 ) | ( n1407 & n3267 ) | ( ~n3008 & n3267 ) ;
  assign n3269 = n3009 & n3268 ;
  buffer buf_n3270( .i (n3269), .o (n3270) );
  assign n3277 = n3073 | n3270 ;
  buffer buf_n3278( .i (n3277), .o (n3278) );
  buffer buf_n3279( .i (n3278), .o (n3279) );
  assign n3280 = n3263 | n3279 ;
  assign n3281 = ( ~n2994 & n3249 ) | ( ~n2994 & n3280 ) | ( n3249 & n3280 ) ;
  assign n3282 = n2995 | n3281 ;
  buffer buf_n3031( .i (n3030), .o (n3031) );
  buffer buf_n3032( .i (n3031), .o (n3032) );
  buffer buf_n3033( .i (n3032), .o (n3033) );
  buffer buf_n3034( .i (n3033), .o (n3034) );
  buffer buf_n3035( .i (n3034), .o (n3035) );
  buffer buf_n3036( .i (n3035), .o (n3036) );
  buffer buf_n3037( .i (n3036), .o (n3037) );
  buffer buf_n3019( .i (n3018), .o (n3019) );
  buffer buf_n3020( .i (n3019), .o (n3020) );
  buffer buf_n3021( .i (n3020), .o (n3021) );
  buffer buf_n3022( .i (n3021), .o (n3022) );
  buffer buf_n3023( .i (n3022), .o (n3023) );
  buffer buf_n3024( .i (n3023), .o (n3024) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  assign n3283 = n2869 & n3008 ;
  assign n3284 = ( n801 & n2692 ) | ( n801 & n3283 ) | ( n2692 & n3283 ) ;
  assign n3285 = ~n802 & n3284 ;
  buffer buf_n3286( .i (n3285), .o (n3286) );
  buffer buf_n3287( .i (n3286), .o (n3287) );
  buffer buf_n3288( .i (n3287), .o (n3288) );
  buffer buf_n3289( .i (n3288), .o (n3289) );
  assign n3291 = n3024 | n3289 ;
  assign n3292 = n3037 | n3291 ;
  assign n3293 = n3282 | n3292 ;
  assign n3294 = ( ~n3227 & n3235 ) | ( ~n3227 & n3293 ) | ( n3235 & n3293 ) ;
  assign n3295 = n3228 | n3294 ;
  buffer buf_n2752( .i (n2751), .o (n2752) );
  assign n3296 = n2742 & ~n2870 ;
  buffer buf_n3297( .i (n3296), .o (n3297) );
  buffer buf_n3298( .i (n3297), .o (n3298) );
  buffer buf_n3299( .i (n3298), .o (n3299) );
  buffer buf_n3300( .i (n3299), .o (n3300) );
  buffer buf_n3301( .i (n3300), .o (n3301) );
  buffer buf_n3302( .i (n3301), .o (n3302) );
  buffer buf_n3303( .i (n3302), .o (n3303) );
  buffer buf_n3304( .i (n3303), .o (n3304) );
  buffer buf_n3305( .i (n3304), .o (n3305) );
  assign n3306 = n2771 | n2794 ;
  assign n3307 = ( n2752 & ~n3305 ) | ( n2752 & n3306 ) | ( ~n3305 & n3306 ) ;
  assign n3308 = n3295 | n3307 ;
  assign n3309 = ( ~n3188 & n3193 ) | ( ~n3188 & n3308 ) | ( n3193 & n3308 ) ;
  assign n3310 = n3189 | n3309 ;
  buffer buf_n2617( .i (n2616), .o (n2617) );
  buffer buf_n2618( .i (n2617), .o (n2618) );
  assign n3311 = n2588 | n3129 ;
  buffer buf_n3312( .i (n3311), .o (n3312) );
  buffer buf_n3313( .i (n3312), .o (n3313) );
  buffer buf_n3314( .i (n3313), .o (n3314) );
  buffer buf_n3315( .i (n3314), .o (n3315) );
  buffer buf_n3316( .i (n3315), .o (n3316) );
  buffer buf_n3317( .i (n3316), .o (n3317) );
  buffer buf_n3318( .i (n3317), .o (n3318) );
  buffer buf_n2687( .i (n2686), .o (n2687) );
  buffer buf_n2688( .i (n2687), .o (n2688) );
  assign n3319 = n2433 | n2696 ;
  assign n3320 = ( n2673 & ~n2687 ) | ( n2673 & n3319 ) | ( ~n2687 & n3319 ) ;
  assign n3321 = n2688 | n3320 ;
  assign n3322 = n2656 | n3168 ;
  buffer buf_n3323( .i (n3322), .o (n3323) );
  buffer buf_n3324( .i (n3323), .o (n3324) );
  buffer buf_n3325( .i (n3324), .o (n3325) );
  buffer buf_n3326( .i (n3325), .o (n3326) );
  buffer buf_n3327( .i (n3326), .o (n3327) );
  buffer buf_n3328( .i (n3327), .o (n3328) );
  assign n3333 = n2636 | n3328 ;
  assign n3334 = n3321 | n3333 ;
  buffer buf_n1319( .i (n1318), .o (n1319) );
  assign n3335 = ~n1294 & n2320 ;
  assign n3336 = ~n1319 & n3335 ;
  buffer buf_n3337( .i (n3336), .o (n3337) );
  buffer buf_n3338( .i (n3337), .o (n3338) );
  buffer buf_n3339( .i (n3338), .o (n3339) );
  buffer buf_n3340( .i (n3339), .o (n3340) );
  buffer buf_n3341( .i (n3340), .o (n3341) );
  buffer buf_n3342( .i (n3341), .o (n3342) );
  buffer buf_n3343( .i (n3342), .o (n3343) );
  buffer buf_n3344( .i (n3343), .o (n3344) );
  buffer buf_n2602( .i (n2601), .o (n2602) );
  buffer buf_n2603( .i (n2602), .o (n2603) );
  buffer buf_n2604( .i (n2603), .o (n2604) );
  assign n3345 = n2330 | n2604 ;
  assign n3346 = n3344 | n3345 ;
  assign n3347 = n3334 | n3346 ;
  assign n3348 = ( ~n2617 & n3318 ) | ( ~n2617 & n3347 ) | ( n3318 & n3347 ) ;
  assign n3349 = n2618 | n3348 ;
  buffer buf_n3350( .i (n3349), .o (n3350) );
  buffer buf_n3351( .i (n3350), .o (n3351) );
  buffer buf_n2385( .i (n2384), .o (n2385) );
  buffer buf_n2386( .i (n2385), .o (n2386) );
  buffer buf_n2387( .i (n2386), .o (n2387) );
  buffer buf_n3161( .i (n3160), .o (n3161) );
  buffer buf_n3162( .i (n3161), .o (n3162) );
  buffer buf_n3163( .i (n3162), .o (n3163) );
  buffer buf_n3164( .i (n3163), .o (n3164) );
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  buffer buf_n2511( .i (n2510), .o (n2511) );
  buffer buf_n2512( .i (n2511), .o (n2512) );
  buffer buf_n2513( .i (n2512), .o (n2513) );
  assign n3352 = n2410 | n2513 ;
  assign n3353 = ( ~n2386 & n3164 ) | ( ~n2386 & n3352 ) | ( n3164 & n3352 ) ;
  assign n3354 = n2387 | n3353 ;
  assign n3355 = n2740 & n3241 ;
  buffer buf_n3356( .i (n3355), .o (n3356) );
  buffer buf_n3357( .i (n3356), .o (n3357) );
  buffer buf_n3358( .i (n3357), .o (n3358) );
  buffer buf_n3359( .i (n3358), .o (n3359) );
  buffer buf_n3360( .i (n3359), .o (n3360) );
  buffer buf_n3361( .i (n3360), .o (n3361) );
  buffer buf_n3362( .i (n3361), .o (n3362) );
  buffer buf_n3363( .i (n3362), .o (n3363) );
  assign n3365 = n2945 & n3194 ;
  buffer buf_n3366( .i (n3365), .o (n3366) );
  assign n3371 = n3298 | n3366 ;
  buffer buf_n3372( .i (n3371), .o (n3372) );
  buffer buf_n3373( .i (n3372), .o (n3373) );
  assign n3376 = n2962 & n3241 ;
  buffer buf_n3377( .i (n3376), .o (n3377) );
  buffer buf_n3378( .i (n3377), .o (n3378) );
  assign n3388 = n2950 | n3378 ;
  buffer buf_n3389( .i (n3388), .o (n3389) );
  buffer buf_n3390( .i (n3389), .o (n3390) );
  buffer buf_n3391( .i (n3390), .o (n3391) );
  assign n3392 = n2971 | n3221 ;
  assign n3393 = n3391 | n3392 ;
  assign n3394 = ( ~n3362 & n3373 ) | ( ~n3362 & n3393 ) | ( n3373 & n3393 ) ;
  assign n3395 = n3363 | n3394 ;
  buffer buf_n3396( .i (n3395), .o (n3396) );
  buffer buf_n3397( .i (n3396), .o (n3397) );
  assign n3398 = n2932 | n3245 ;
  buffer buf_n3399( .i (n3398), .o (n3399) );
  assign n3400 = n3206 | n3399 ;
  buffer buf_n3401( .i (n3400), .o (n3401) );
  assign n3405 = n3199 | n3401 ;
  assign n3406 = ( ~n2900 & n2923 ) | ( ~n2900 & n3405 ) | ( n2923 & n3405 ) ;
  assign n3407 = n2901 | n3406 ;
  assign n3408 = n2783 & n3241 ;
  buffer buf_n3409( .i (n3408), .o (n3409) );
  buffer buf_n3410( .i (n3409), .o (n3410) );
  buffer buf_n3411( .i (n3410), .o (n3411) );
  buffer buf_n3412( .i (n3411), .o (n3412) );
  buffer buf_n3413( .i (n3412), .o (n3413) );
  buffer buf_n3414( .i (n3413), .o (n3414) );
  buffer buf_n3415( .i (n3414), .o (n3415) );
  buffer buf_n3416( .i (n3415), .o (n3416) );
  assign n3417 = ( n1597 & n2846 ) | ( n1597 & n2957 ) | ( n2846 & n2957 ) ;
  assign n3418 = ~n1874 & n3417 ;
  buffer buf_n3419( .i (n3418), .o (n3419) );
  buffer buf_n3420( .i (n3419), .o (n3420) );
  assign n3423 = ( n762 & n1536 ) | ( n762 & ~n3419 ) | ( n1536 & ~n3419 ) ;
  assign n3424 = n3420 & n3423 ;
  buffer buf_n3425( .i (n3424), .o (n3425) );
  buffer buf_n3426( .i (n3425), .o (n3426) );
  buffer buf_n3427( .i (n3426), .o (n3427) );
  buffer buf_n3428( .i (n3427), .o (n3428) );
  buffer buf_n3429( .i (n3428), .o (n3429) );
  buffer buf_n3430( .i (n3429), .o (n3430) );
  buffer buf_n3431( .i (n3430), .o (n3431) );
  buffer buf_n3432( .i (n3431), .o (n3432) );
  assign n3435 = ( n1395 & n2712 ) | ( n1395 & n3252 ) | ( n2712 & n3252 ) ;
  assign n3436 = ~n2161 & n3435 ;
  buffer buf_n3437( .i (n3436), .o (n3437) );
  buffer buf_n3441( .i (n3240), .o (n3441) );
  assign n3442 = n3437 & n3441 ;
  assign n3443 = n800 & n3442 ;
  buffer buf_n3444( .i (n3443), .o (n3444) );
  buffer buf_n3445( .i (n3444), .o (n3445) );
  buffer buf_n3446( .i (n3445), .o (n3446) );
  buffer buf_n3447( .i (n3446), .o (n3447) );
  buffer buf_n3448( .i (n3447), .o (n3448) );
  assign n3451 = ( n2766 & ~n2773 ) | ( n2766 & n2789 ) | ( ~n2773 & n2789 ) ;
  assign n3452 = n3448 | n3451 ;
  assign n3453 = ( ~n3415 & n3432 ) | ( ~n3415 & n3452 ) | ( n3432 & n3452 ) ;
  assign n3454 = n3416 | n3453 ;
  buffer buf_n3264( .i (n3263), .o (n3264) );
  buffer buf_n3265( .i (n3264), .o (n3265) );
  buffer buf_n3271( .i (n3270), .o (n3271) );
  buffer buf_n3272( .i (n3271), .o (n3272) );
  buffer buf_n3273( .i (n3272), .o (n3273) );
  buffer buf_n3274( .i (n3273), .o (n3274) );
  buffer buf_n3086( .i (n3085), .o (n3086) );
  buffer buf_n3087( .i (n3086), .o (n3087) );
  buffer buf_n3088( .i (n3087), .o (n3088) );
  buffer buf_n3010( .i (n3009), .o (n3010) );
  buffer buf_n3011( .i (n3010), .o (n3011) );
  buffer buf_n3012( .i (n3011), .o (n3012) );
  buffer buf_n3013( .i (n3012), .o (n3013) );
  assign n3455 = n894 & n3013 ;
  assign n3456 = n3088 | n3455 ;
  assign n3457 = ( ~n3264 & n3274 ) | ( ~n3264 & n3456 ) | ( n3274 & n3456 ) ;
  assign n3458 = n3265 | n3457 ;
  assign n3459 = n3454 | n3458 ;
  assign n3460 = ( ~n3396 & n3407 ) | ( ~n3396 & n3459 ) | ( n3407 & n3459 ) ;
  assign n3461 = n3397 | n3460 ;
  buffer buf_n2806( .i (n2805), .o (n2806) );
  buffer buf_n2807( .i (n2806), .o (n2807) );
  assign n3462 = n2715 & n3441 ;
  buffer buf_n3463( .i (n3462), .o (n3463) );
  buffer buf_n3468( .i (n3267), .o (n3468) );
  assign n3469 = n3463 & n3468 ;
  buffer buf_n3470( .i (n3469), .o (n3470) );
  buffer buf_n3471( .i (n3470), .o (n3471) );
  buffer buf_n3472( .i (n3471), .o (n3472) );
  buffer buf_n3473( .i (n3472), .o (n3473) );
  buffer buf_n3474( .i (n3473), .o (n3474) );
  assign n3475 = n2724 | n2881 ;
  assign n3476 = n3474 | n3475 ;
  buffer buf_n3477( .i (n3476), .o (n3477) );
  assign n3478 = n2842 | n3477 ;
  assign n3479 = ( ~n2806 & n2830 ) | ( ~n2806 & n3478 ) | ( n2830 & n3478 ) ;
  assign n3480 = n2807 | n3479 ;
  assign n3481 = n3461 | n3480 ;
  assign n3482 = ( ~n3350 & n3354 ) | ( ~n3350 & n3481 ) | ( n3354 & n3481 ) ;
  assign n3483 = n3351 | n3482 ;
  buffer buf_n2367( .i (n2366), .o (n2367) );
  buffer buf_n2368( .i (n2367), .o (n2368) );
  buffer buf_n2369( .i (n2368), .o (n2369) );
  assign n3484 = ( n1901 & n2648 ) | ( n1901 & n3468 ) | ( n2648 & n3468 ) ;
  buffer buf_n3485( .i (n3468), .o (n3485) );
  assign n3486 = n3484 & ~n3485 ;
  buffer buf_n3487( .i (n3486), .o (n3487) );
  buffer buf_n3488( .i (n3487), .o (n3488) );
  buffer buf_n3489( .i (n3488), .o (n3489) );
  buffer buf_n3490( .i (n3489), .o (n3490) );
  buffer buf_n3491( .i (n3490), .o (n3491) );
  buffer buf_n3492( .i (n3491), .o (n3492) );
  buffer buf_n3493( .i (n3492), .o (n3493) );
  buffer buf_n3494( .i (n3493), .o (n3494) );
  buffer buf_n3495( .i (n3494), .o (n3495) );
  assign n3496 = n2400 | n2428 ;
  buffer buf_n3497( .i (n3496), .o (n3497) );
  buffer buf_n3498( .i (n3497), .o (n3498) );
  buffer buf_n3499( .i (n3498), .o (n3499) );
  buffer buf_n3500( .i (n3499), .o (n3500) );
  buffer buf_n3501( .i (n3500), .o (n3501) );
  buffer buf_n3502( .i (n3501), .o (n3502) );
  buffer buf_n3503( .i (n3502), .o (n3503) );
  buffer buf_n3504( .i (n3503), .o (n3504) );
  buffer buf_n3505( .i (n3504), .o (n3505) );
  buffer buf_n3506( .i (n3505), .o (n3506) );
  assign n3507 = n2043 & n2376 ;
  buffer buf_n3508( .i (n3507), .o (n3508) );
  buffer buf_n2394( .i (n2393), .o (n2394) );
  buffer buf_n2395( .i (n2394), .o (n2395) );
  buffer buf_n2396( .i (n2395), .o (n2396) );
  buffer buf_n3515( .i (n1346), .o (n3515) );
  buffer buf_n3516( .i (n3515), .o (n3516) );
  assign n3517 = n2396 & n3516 ;
  buffer buf_n3518( .i (n3517), .o (n3518) );
  buffer buf_n3519( .i (n3518), .o (n3519) );
  assign n3529 = n3508 | n3519 ;
  assign n3530 = n3157 | n3529 ;
  buffer buf_n3531( .i (n3530), .o (n3531) );
  buffer buf_n3532( .i (n3531), .o (n3532) );
  buffer buf_n3533( .i (n3532), .o (n3533) );
  buffer buf_n3534( .i (n3533), .o (n3534) );
  buffer buf_n3535( .i (n3534), .o (n3535) );
  buffer buf_n2680( .i (n2679), .o (n2680) );
  assign n3536 = n2680 & n3516 ;
  buffer buf_n3537( .i (n3536), .o (n3537) );
  buffer buf_n3538( .i (n3537), .o (n3538) );
  buffer buf_n3539( .i (n3538), .o (n3539) );
  buffer buf_n3540( .i (n3539), .o (n3540) );
  buffer buf_n3541( .i (n3540), .o (n3541) );
  buffer buf_n3542( .i (n3541), .o (n3542) );
  buffer buf_n3543( .i (n3542), .o (n3543) );
  buffer buf_n3544( .i (n3543), .o (n3544) );
  buffer buf_n3173( .i (n3172), .o (n3173) );
  buffer buf_n3174( .i (n3173), .o (n3174) );
  buffer buf_n3175( .i (n3174), .o (n3175) );
  buffer buf_n3176( .i (n3175), .o (n3176) );
  buffer buf_n2674( .i (n2673), .o (n2674) );
  buffer buf_n2697( .i (n2696), .o (n2697) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n3421( .i (n3420), .o (n3421) );
  buffer buf_n3422( .i (n3421), .o (n3422) );
  assign n3548 = ~n3267 & n3422 ;
  assign n3549 = ( n633 & n766 ) | ( n633 & n3548 ) | ( n766 & n3548 ) ;
  assign n3550 = ~n634 & n3549 ;
  buffer buf_n3551( .i (n3550), .o (n3551) );
  assign n3553 = n928 & n3551 ;
  buffer buf_n3554( .i (n3553), .o (n3554) );
  assign n3559 = n2697 | n3554 ;
  assign n3560 = n2674 | n3559 ;
  assign n3561 = n3176 | n3560 ;
  assign n3562 = n3544 | n3561 ;
  assign n3563 = n3535 | n3562 ;
  assign n3564 = ( ~n3494 & n3506 ) | ( ~n3494 & n3563 ) | ( n3506 & n3563 ) ;
  assign n3565 = n3495 | n3564 ;
  buffer buf_n2479( .i (n2478), .o (n2479) );
  buffer buf_n2480( .i (n2479), .o (n2480) );
  buffer buf_n2481( .i (n2480), .o (n2481) );
  buffer buf_n2482( .i (n2481), .o (n2482) );
  buffer buf_n2483( .i (n2482), .o (n2483) );
  buffer buf_n2484( .i (n2483), .o (n2484) );
  assign n3566 = n161 & n2638 ;
  buffer buf_n3567( .i (n2999), .o (n3567) );
  assign n3568 = ( n2733 & n3566 ) | ( n2733 & n3567 ) | ( n3566 & n3567 ) ;
  buffer buf_n3569( .i (n3567), .o (n3569) );
  assign n3570 = n3568 & ~n3569 ;
  assign n3571 = n3143 & n3570 ;
  assign n3572 = ( n663 & n2848 ) | ( n663 & n3571 ) | ( n2848 & n3571 ) ;
  assign n3573 = ~n2134 & n3572 ;
  assign n3574 = n1345 & n3573 ;
  buffer buf_n3575( .i (n3574), .o (n3575) );
  buffer buf_n3576( .i (n3575), .o (n3576) );
  buffer buf_n3577( .i (n3576), .o (n3577) );
  buffer buf_n3578( .i (n3577), .o (n3578) );
  buffer buf_n3579( .i (n3578), .o (n3579) );
  buffer buf_n3580( .i (n3579), .o (n3580) );
  buffer buf_n3581( .i (n3580), .o (n3581) );
  buffer buf_n3582( .i (n3581), .o (n3582) );
  buffer buf_n3583( .i (n3582), .o (n3583) );
  buffer buf_n3584( .i (n3583), .o (n3584) );
  buffer buf_n3585( .i (n3584), .o (n3585) );
  assign n3586 = ~n162 & n2733 ;
  assign n3587 = ( n134 & ~n3569 ) | ( n134 & n3586 ) | ( ~n3569 & n3586 ) ;
  assign n3588 = ~n135 & n3587 ;
  assign n3589 = ( n1966 & n2848 ) | ( n1966 & n3588 ) | ( n2848 & n3588 ) ;
  buffer buf_n3590( .i (n2808), .o (n3590) );
  buffer buf_n3591( .i (n3590), .o (n3591) );
  assign n3592 = n3589 & ~n3591 ;
  assign n3593 = ( n1573 & n3165 ) | ( n1573 & n3592 ) | ( n3165 & n3592 ) ;
  assign n3594 = ~n3214 & n3593 ;
  buffer buf_n3595( .i (n3594), .o (n3595) );
  buffer buf_n3596( .i (n3595), .o (n3596) );
  buffer buf_n3597( .i (n3596), .o (n3597) );
  buffer buf_n3598( .i (n3597), .o (n3598) );
  buffer buf_n3599( .i (n3598), .o (n3599) );
  buffer buf_n3600( .i (n3599), .o (n3600) );
  buffer buf_n3601( .i (n3600), .o (n3601) );
  buffer buf_n3602( .i (n3601), .o (n3602) );
  buffer buf_n3603( .i (n3602), .o (n3603) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n2422( .i (n2421), .o (n2422) );
  assign n3604 = n2422 & n3240 ;
  buffer buf_n3605( .i (n3604), .o (n3605) );
  assign n3606 = n668 & n3605 ;
  buffer buf_n3607( .i (n3606), .o (n3607) );
  buffer buf_n704( .i (n703), .o (n704) );
  assign n3616 = n704 & n3605 ;
  buffer buf_n3617( .i (n3616), .o (n3617) );
  assign n3623 = n3607 | n3617 ;
  buffer buf_n3624( .i (n3623), .o (n3624) );
  buffer buf_n3625( .i (n3624), .o (n3625) );
  buffer buf_n3626( .i (n3625), .o (n3626) );
  buffer buf_n3627( .i (n3626), .o (n3627) );
  buffer buf_n3628( .i (n3627), .o (n3628) );
  assign n3629 = n3603 | n3628 ;
  assign n3630 = ( ~n2483 & n3585 ) | ( ~n2483 & n3629 ) | ( n3585 & n3629 ) ;
  assign n3631 = n2484 | n3630 ;
  buffer buf_n3074( .i (n3073), .o (n3074) );
  buffer buf_n3075( .i (n3074), .o (n3075) );
  buffer buf_n3076( .i (n3075), .o (n3076) );
  buffer buf_n3077( .i (n3076), .o (n3077) );
  buffer buf_n3078( .i (n3077), .o (n3078) );
  buffer buf_n3079( .i (n3078), .o (n3079) );
  assign n3632 = n3300 | n3431 ;
  assign n3633 = n2994 | n3632 ;
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n3634( .i (n3252), .o (n3634) );
  assign n3635 = n1327 & ~n3634 ;
  assign n3636 = ~n1910 & n3635 ;
  buffer buf_n3637( .i (n3636), .o (n3637) );
  assign n3638 = ( n1900 & n3267 ) | ( n1900 & n3637 ) | ( n3267 & n3637 ) ;
  assign n3639 = ~n3468 & n3638 ;
  buffer buf_n3640( .i (n3639), .o (n3640) );
  buffer buf_n3641( .i (n3640), .o (n3641) );
  buffer buf_n3642( .i (n3641), .o (n3642) );
  buffer buf_n3643( .i (n3642), .o (n3643) );
  assign n3649 = n699 & ~n884 ;
  buffer buf_n3650( .i (n3649), .o (n3650) );
  buffer buf_n3651( .i (n3650), .o (n3651) );
  assign n3652 = ( n2812 & n3213 ) | ( n2812 & n3651 ) | ( n3213 & n3651 ) ;
  assign n3653 = ~n3256 & n3652 ;
  buffer buf_n3654( .i (n3441), .o (n3654) );
  assign n3655 = n3653 & n3654 ;
  buffer buf_n3656( .i (n3655), .o (n3656) );
  buffer buf_n3657( .i (n3656), .o (n3657) );
  buffer buf_n3658( .i (n3657), .o (n3658) );
  buffer buf_n3659( .i (n3658), .o (n3659) );
  assign n3663 = ( ~n2852 & n3256 ) | ( ~n2852 & n3515 ) | ( n3256 & n3515 ) ;
  buffer buf_n3664( .i (n3256), .o (n3664) );
  assign n3665 = n3663 & ~n3664 ;
  buffer buf_n3666( .i (n3665), .o (n3666) );
  buffer buf_n3667( .i (n3666), .o (n3667) );
  assign n3674 = n3470 | n3667 ;
  assign n3675 = n3446 | n3674 ;
  assign n3676 = n3659 | n3675 ;
  assign n3677 = n3643 | n3676 ;
  buffer buf_n414( .i (x14), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  assign n3678 = n434 & ~n3145 ;
  assign n3679 = ( n825 & ~n3165 ) | ( n825 & n3678 ) | ( ~n3165 & n3678 ) ;
  assign n3680 = ~n3125 & n3679 ;
  assign n3681 = ~n3441 & n3680 ;
  buffer buf_n3682( .i (n3681), .o (n3682) );
  buffer buf_n392( .i (x13), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  assign n3689 = n410 & ~n822 ;
  assign n3690 = ( n433 & n3590 ) | ( n433 & n3689 ) | ( n3590 & n3689 ) ;
  assign n3691 = ~n434 & n3690 ;
  buffer buf_n3692( .i (n885), .o (n3692) );
  assign n3693 = n3691 & ~n3692 ;
  buffer buf_n3694( .i (n3239), .o (n3694) );
  assign n3695 = ( n3213 & n3693 ) | ( n3213 & ~n3694 ) | ( n3693 & ~n3694 ) ;
  buffer buf_n3696( .i (n3212), .o (n3696) );
  buffer buf_n3697( .i (n3696), .o (n3697) );
  assign n3698 = n3695 & ~n3697 ;
  buffer buf_n3699( .i (n3698), .o (n3699) );
  assign n3709 = n3682 | n3699 ;
  buffer buf_n3710( .i (n3709), .o (n3710) );
  buffer buf_n3711( .i (n3710), .o (n3711) );
  buffer buf_n3712( .i (n3711), .o (n3712) );
  buffer buf_n3713( .i (n3712), .o (n3713) );
  buffer buf_n3714( .i (n3713), .o (n3714) );
  assign n3715 = n3677 | n3714 ;
  assign n3716 = ( ~n3078 & n3633 ) | ( ~n3078 & n3715 ) | ( n3633 & n3715 ) ;
  assign n3717 = n3079 | n3716 ;
  buffer buf_n3718( .i (n884), .o (n3718) );
  assign n3719 = n796 & ~n3718 ;
  assign n3720 = ( n2449 & n3212 ) | ( n2449 & n3719 ) | ( n3212 & n3719 ) ;
  assign n3721 = ~n3696 & n3720 ;
  buffer buf_n3722( .i (n3694), .o (n3722) );
  assign n3723 = n3721 & n3722 ;
  buffer buf_n3724( .i (n3723), .o (n3724) );
  buffer buf_n3725( .i (n3724), .o (n3725) );
  buffer buf_n3726( .i (n3725), .o (n3726) );
  buffer buf_n3727( .i (n3726), .o (n3727) );
  buffer buf_n3728( .i (n3727), .o (n3728) );
  buffer buf_n3729( .i (n3728), .o (n3729) );
  buffer buf_n3730( .i (n3729), .o (n3730) );
  buffer buf_n3731( .i (n3730), .o (n3731) );
  assign n3732 = ( n2449 & n3212 ) | ( n2449 & n3650 ) | ( n3212 & n3650 ) ;
  assign n3733 = ~n3696 & n3732 ;
  assign n3734 = n3722 & n3733 ;
  buffer buf_n3735( .i (n3734), .o (n3735) );
  buffer buf_n3736( .i (n3735), .o (n3736) );
  buffer buf_n3737( .i (n3736), .o (n3737) );
  buffer buf_n3738( .i (n3737), .o (n3738) );
  buffer buf_n3739( .i (n3738), .o (n3739) );
  buffer buf_n3740( .i (n3739), .o (n3740) );
  buffer buf_n3741( .i (n3740), .o (n3741) );
  buffer buf_n2454( .i (n2453), .o (n2454) );
  assign n3744 = n2043 & n2454 ;
  buffer buf_n3745( .i (n3744), .o (n3745) );
  buffer buf_n3746( .i (n3745), .o (n3746) );
  buffer buf_n3747( .i (n3746), .o (n3747) );
  buffer buf_n3748( .i (n3747), .o (n3748) );
  assign n3755 = n700 & n3049 ;
  buffer buf_n3756( .i (n3755), .o (n3756) );
  buffer buf_n3757( .i (n3756), .o (n3757) );
  buffer buf_n3758( .i (n3757), .o (n3758) );
  buffer buf_n3759( .i (n3053), .o (n3759) );
  assign n3760 = ( n3637 & n3758 ) | ( n3637 & n3759 ) | ( n3758 & n3759 ) ;
  buffer buf_n3761( .i (n3759), .o (n3761) );
  assign n3762 = n3760 & ~n3761 ;
  buffer buf_n3763( .i (n3762), .o (n3763) );
  buffer buf_n3764( .i (n3763), .o (n3764) );
  assign n3771 = n2501 | n3764 ;
  assign n3772 = n2801 | n3771 ;
  assign n3773 = n3748 | n3772 ;
  assign n3774 = ( ~n3730 & n3741 ) | ( ~n3730 & n3773 ) | ( n3741 & n3773 ) ;
  assign n3775 = n3731 | n3774 ;
  buffer buf_n3776( .i (n3775), .o (n3776) );
  assign n3779 = n3717 | n3776 ;
  assign n3780 = n3631 | n3779 ;
  buffer buf_n3134( .i (n3133), .o (n3134) );
  buffer buf_n3135( .i (n3134), .o (n3135) );
  buffer buf_n3136( .i (n3135), .o (n3136) );
  buffer buf_n3137( .i (n3136), .o (n3137) );
  buffer buf_n3138( .i (n3137), .o (n3138) );
  buffer buf_n2570( .i (n2569), .o (n2570) );
  buffer buf_n2571( .i (n2570), .o (n2571) );
  buffer buf_n2572( .i (n2571), .o (n2572) );
  buffer buf_n2573( .i (n2572), .o (n2573) );
  buffer buf_n2664( .i (n2663), .o (n2664) );
  buffer buf_n2665( .i (n2664), .o (n2665) );
  buffer buf_n2592( .i (n2591), .o (n2592) );
  buffer buf_n2593( .i (n2592), .o (n2593) );
  buffer buf_n2594( .i (n2593), .o (n2594) );
  assign n3781 = ~n823 & n2579 ;
  assign n3782 = ~n3145 & n3781 ;
  buffer buf_n3783( .i (n3782), .o (n3783) );
  buffer buf_n3784( .i (n3783), .o (n3784) );
  assign n3785 = n3515 & n3784 ;
  buffer buf_n3786( .i (n3785), .o (n3786) );
  buffer buf_n3787( .i (n3786), .o (n3787) );
  buffer buf_n3788( .i (n3787), .o (n3788) );
  buffer buf_n3789( .i (n3788), .o (n3789) );
  buffer buf_n3790( .i (n3789), .o (n3790) );
  buffer buf_n3791( .i (n3790), .o (n3791) );
  buffer buf_n3792( .i (n3791), .o (n3792) );
  buffer buf_n3793( .i (n3792), .o (n3793) );
  assign n3795 = n2594 | n3793 ;
  assign n3796 = n2665 | n3795 ;
  assign n3797 = n2573 | n3796 ;
  assign n3798 = n3138 | n3797 ;
  assign n3799 = n3780 | n3798 ;
  assign n3800 = ( ~n2368 & n3565 ) | ( ~n2368 & n3799 ) | ( n3565 & n3799 ) ;
  assign n3801 = n2369 | n3800 ;
  buffer buf_n2357( .i (n2356), .o (n2357) );
  assign n3802 = n1219 & ~n1267 ;
  assign n3803 = ( n1241 & n2313 ) | ( n1241 & n3802 ) | ( n2313 & n3802 ) ;
  assign n3804 = ~n1242 & n3803 ;
  buffer buf_n3805( .i (n3804), .o (n3805) );
  buffer buf_n3806( .i (n3805), .o (n3806) );
  buffer buf_n3807( .i (n3806), .o (n3807) );
  buffer buf_n3808( .i (n3807), .o (n3808) );
  buffer buf_n3809( .i (n3808), .o (n3809) );
  assign n3814 = n2269 | n3809 ;
  assign n3815 = n2357 | n3814 ;
  buffer buf_n3816( .i (n3815), .o (n3816) );
  buffer buf_n3817( .i (n3816), .o (n3817) );
  buffer buf_n3818( .i (n3817), .o (n3818) );
  buffer buf_n3819( .i (n3818), .o (n3819) );
  buffer buf_n3820( .i (n3819), .o (n3820) );
  buffer buf_n3821( .i (n3820), .o (n3821) );
  buffer buf_n3822( .i (n3821), .o (n3822) );
  buffer buf_n3823( .i (n3822), .o (n3823) );
  buffer buf_n2525( .i (n2524), .o (n2525) );
  buffer buf_n2526( .i (n2525), .o (n2526) );
  buffer buf_n2527( .i (n2526), .o (n2527) );
  buffer buf_n2528( .i (n2527), .o (n2528) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n2559( .i (n2558), .o (n2559) );
  buffer buf_n2560( .i (n2559), .o (n2560) );
  assign n3824 = n1021 & n2560 ;
  buffer buf_n3825( .i (n3824), .o (n3825) );
  buffer buf_n3826( .i (n3825), .o (n3826) );
  buffer buf_n3827( .i (n3826), .o (n3827) );
  buffer buf_n3828( .i (n3827), .o (n3828) );
  buffer buf_n3829( .i (n3828), .o (n3829) );
  buffer buf_n3830( .i (n3829), .o (n3830) );
  assign n3831 = n2573 | n3137 ;
  assign n3832 = ( ~n2527 & n3830 ) | ( ~n2527 & n3831 ) | ( n3830 & n3831 ) ;
  assign n3833 = n2528 | n3832 ;
  buffer buf_n2502( .i (n2501), .o (n2502) );
  buffer buf_n2503( .i (n2502), .o (n2503) );
  buffer buf_n2504( .i (n2503), .o (n2504) );
  buffer buf_n2505( .i (n2504), .o (n2505) );
  buffer buf_n2506( .i (n2505), .o (n2506) );
  buffer buf_n3449( .i (n3448), .o (n3449) );
  assign n3834 = n2803 | n3449 ;
  assign n3835 = ( ~n2505 & n3584 ) | ( ~n2505 & n3834 ) | ( n3584 & n3834 ) ;
  assign n3836 = n2506 | n3835 ;
  assign n3837 = n2478 | n3599 ;
  buffer buf_n3838( .i (n3837), .o (n3838) );
  buffer buf_n3839( .i (n3838), .o (n3839) );
  buffer buf_n3840( .i (n3839), .o (n3840) );
  buffer buf_n3841( .i (n3840), .o (n3841) );
  assign n3844 = n927 & n2764 ;
  buffer buf_n3845( .i (n3844), .o (n3845) );
  buffer buf_n3846( .i (n3845), .o (n3846) );
  assign n3849 = n2990 | n3057 ;
  assign n3850 = ( ~n3196 & n3205 ) | ( ~n3196 & n3849 ) | ( n3205 & n3849 ) ;
  assign n3851 = n3197 | n3850 ;
  assign n3852 = n3846 | n3851 ;
  assign n3853 = ( n3301 & ~n3415 ) | ( n3301 & n3852 ) | ( ~n3415 & n3852 ) ;
  assign n3854 = n3416 | n3853 ;
  assign n3855 = n3841 | n3854 ;
  assign n3856 = ( ~n3163 & n3836 ) | ( ~n3163 & n3855 ) | ( n3836 & n3855 ) ;
  assign n3857 = n3164 | n3856 ;
  buffer buf_n3329( .i (n3328), .o (n3329) );
  buffer buf_n3330( .i (n3329), .o (n3330) );
  buffer buf_n3331( .i (n3330), .o (n3331) );
  buffer buf_n3332( .i (n3331), .o (n3332) );
  buffer buf_n2595( .i (n2594), .o (n2595) );
  buffer buf_n2596( .i (n2595), .o (n2596) );
  assign n3858 = n2669 | n3497 ;
  buffer buf_n3859( .i (n3858), .o (n3859) );
  buffer buf_n3860( .i (n3859), .o (n3860) );
  assign n3861 = n2696 | n3860 ;
  buffer buf_n3862( .i (n3861), .o (n3862) );
  buffer buf_n3863( .i (n3862), .o (n3863) );
  buffer buf_n3864( .i (n3863), .o (n3864) );
  buffer buf_n3865( .i (n3864), .o (n3865) );
  assign n3866 = n2596 | n3865 ;
  assign n3867 = n3332 | n3866 ;
  assign n3868 = n3857 | n3867 ;
  assign n3869 = ( ~n3822 & n3833 ) | ( ~n3822 & n3868 ) | ( n3833 & n3868 ) ;
  assign n3870 = n3823 | n3869 ;
  buffer buf_n962( .i (x32), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  assign n3871 = n696 & n2251 ;
  assign n3872 = ( n882 & n917 ) | ( n882 & n3871 ) | ( n917 & n3871 ) ;
  assign n3873 = ~n918 & n3872 ;
  buffer buf_n3874( .i (n3873), .o (n3874) );
  buffer buf_n3875( .i (n3874), .o (n3875) );
  buffer buf_n3876( .i (n3875), .o (n3876) );
  buffer buf_n3877( .i (n3876), .o (n3877) );
  buffer buf_n3878( .i (n3877), .o (n3878) );
  buffer buf_n3879( .i (n3878), .o (n3879) );
  buffer buf_n3880( .i (n3879), .o (n3880) );
  buffer buf_n3881( .i (n3880), .o (n3881) );
  buffer buf_n3882( .i (n3881), .o (n3882) );
  assign n3888 = n960 & n3881 ;
  assign n3889 = ( n990 & n3882 ) | ( n990 & n3888 ) | ( n3882 & n3888 ) ;
  buffer buf_n3890( .i (n3889), .o (n3890) );
  buffer buf_n3891( .i (n3890), .o (n3891) );
  assign n3892 = ( n2257 & n3214 ) | ( n2257 & n3756 ) | ( n3214 & n3756 ) ;
  buffer buf_n3893( .i (n3214), .o (n3893) );
  assign n3894 = n3892 & ~n3893 ;
  buffer buf_n3895( .i (n3894), .o (n3895) );
  buffer buf_n3896( .i (n3895), .o (n3896) );
  buffer buf_n3897( .i (n3896), .o (n3897) );
  buffer buf_n3898( .i (n3897), .o (n3898) );
  buffer buf_n3899( .i (n3898), .o (n3899) );
  buffer buf_n3900( .i (n3899), .o (n3900) );
  buffer buf_n1125( .i (x37), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1060( .i (x35), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  assign n3904 = ~n982 & n3874 ;
  assign n3905 = ( n954 & ~n1014 ) | ( n954 & n3904 ) | ( ~n1014 & n3904 ) ;
  assign n3906 = ~n955 & n3905 ;
  buffer buf_n3907( .i (n3906), .o (n3907) );
  buffer buf_n3908( .i (n3907), .o (n3908) );
  buffer buf_n1026( .i (x34), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  assign n3916 = n1050 & n3907 ;
  assign n3917 = ( n1085 & n3908 ) | ( n1085 & n3916 ) | ( n3908 & n3916 ) ;
  buffer buf_n3918( .i (n3917), .o (n3918) );
  buffer buf_n3919( .i (n3918), .o (n3919) );
  buffer buf_n3920( .i (n3919), .o (n3920) );
  buffer buf_n1093( .i (x36), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  assign n3921 = ~n1050 & n3907 ;
  assign n3922 = ~n1085 & n3921 ;
  buffer buf_n3923( .i (n3922), .o (n3923) );
  assign n3929 = ( ~n1120 & n3918 ) | ( ~n1120 & n3923 ) | ( n3918 & n3923 ) ;
  assign n3930 = n1153 & ~n3929 ;
  assign n3931 = ( n1154 & n3920 ) | ( n1154 & ~n3930 ) | ( n3920 & ~n3930 ) ;
  assign n3932 = n3900 | n3931 ;
  assign n3933 = ( ~n3117 & n3891 ) | ( ~n3117 & n3932 ) | ( n3891 & n3932 ) ;
  assign n3934 = n3118 | n3933 ;
  buffer buf_n3935( .i (n3934), .o (n3935) );
  buffer buf_n3936( .i (n3935), .o (n3936) );
  buffer buf_n3937( .i (n3692), .o (n3937) );
  assign n3938 = n3125 & n3937 ;
  assign n3939 = ( n2583 & n3697 ) | ( n2583 & n3938 ) | ( n3697 & n3938 ) ;
  assign n3940 = ~n3664 & n3939 ;
  buffer buf_n3941( .i (n3654), .o (n3941) );
  assign n3942 = n3940 & ~n3941 ;
  buffer buf_n3943( .i (n3942), .o (n3943) );
  buffer buf_n3944( .i (n3943), .o (n3944) );
  buffer buf_n3945( .i (n3944), .o (n3945) );
  buffer buf_n3946( .i (n3945), .o (n3946) );
  buffer buf_n3947( .i (n3946), .o (n3947) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  assign n3949 = ( n1899 & ~n2258 ) | ( n1899 & n3697 ) | ( ~n2258 & n3697 ) ;
  assign n3950 = n2259 & n3949 ;
  buffer buf_n3951( .i (n3950), .o (n3951) );
  buffer buf_n3952( .i (n3951), .o (n3952) );
  buffer buf_n3953( .i (n3952), .o (n3953) );
  buffer buf_n3954( .i (n3953), .o (n3954) );
  buffer buf_n3955( .i (n3954), .o (n3955) );
  buffer buf_n3956( .i (n3955), .o (n3956) );
  assign n3958 = n3947 | n3956 ;
  buffer buf_n3959( .i (n3958), .o (n3959) );
  buffer buf_n3960( .i (n3959), .o (n3960) );
  assign n3961 = n1636 | n2611 ;
  buffer buf_n3962( .i (n3961), .o (n3962) );
  buffer buf_n3963( .i (n3962), .o (n3963) );
  buffer buf_n3964( .i (n3963), .o (n3964) );
  buffer buf_n3965( .i (n3964), .o (n3965) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n3966( .i (n1778), .o (n3966) );
  assign n3967 = ( ~n199 & n1802 ) | ( ~n199 & n3966 ) | ( n1802 & n3966 ) ;
  assign n3968 = n200 & n3967 ;
  assign n3969 = ~n827 & n3697 ;
  buffer buf_n3970( .i (n2026), .o (n3970) );
  assign n3971 = ( n3968 & n3969 ) | ( n3968 & n3970 ) | ( n3969 & n3970 ) ;
  buffer buf_n3972( .i (n3970), .o (n3972) );
  assign n3973 = n3971 & ~n3972 ;
  assign n3974 = ~n3194 & n3973 ;
  assign n3975 = n2181 & n3974 ;
  buffer buf_n3976( .i (n3975), .o (n3976) );
  buffer buf_n3977( .i (n3976), .o (n3977) );
  buffer buf_n3978( .i (n3977), .o (n3978) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  assign n3982 = ( ~n222 & n1799 ) | ( ~n222 & n2847 ) | ( n1799 & n2847 ) ;
  assign n3983 = n223 & n3982 ;
  buffer buf_n3984( .i (n824), .o (n3984) );
  assign n3985 = n3983 & ~n3984 ;
  buffer buf_n3986( .i (n1909), .o (n3986) );
  assign n3987 = ( ~n3696 & n3985 ) | ( ~n3696 & n3986 ) | ( n3985 & n3986 ) ;
  buffer buf_n3988( .i (n3986), .o (n3988) );
  assign n3989 = n3987 & ~n3988 ;
  assign n3990 = n3654 & n3989 ;
  assign n3991 = n3761 & n3990 ;
  buffer buf_n3992( .i (n3991), .o (n3992) );
  buffer buf_n3993( .i (n3992), .o (n3993) );
  buffer buf_n3994( .i (n3993), .o (n3994) );
  assign n3998 = n2634 | n3994 ;
  buffer buf_n3999( .i (n3998), .o (n3999) );
  assign n4003 = ( ~n2593 & n3978 ) | ( ~n2593 & n3999 ) | ( n3978 & n3999 ) ;
  assign n4004 = n2594 | n4003 ;
  assign n4005 = n3965 | n4004 ;
  assign n4006 = ( ~n3935 & n3960 ) | ( ~n3935 & n4005 ) | ( n3960 & n4005 ) ;
  assign n4007 = n3936 | n4006 ;
  buffer buf_n4008( .i (n4007), .o (n4008) );
  buffer buf_n4009( .i (n4008), .o (n4009) );
  assign n4010 = n2786 & ~n3194 ;
  buffer buf_n4011( .i (n4010), .o (n4011) );
  buffer buf_n4012( .i (n4011), .o (n4012) );
  buffer buf_n4013( .i (n4012), .o (n4013) );
  buffer buf_n4014( .i (n4013), .o (n4014) );
  buffer buf_n4015( .i (n4014), .o (n4015) );
  buffer buf_n4016( .i (n4015), .o (n4016) );
  buffer buf_n4017( .i (n4016), .o (n4017) );
  buffer buf_n4018( .i (n4017), .o (n4018) );
  buffer buf_n4019( .i (n164), .o (n4019) );
  assign n4020 = ~n2550 & n4019 ;
  buffer buf_n4021( .i (n4020), .o (n4021) );
  buffer buf_n4025( .i (n2036), .o (n4025) );
  assign n4026 = n4021 & ~n4025 ;
  assign n4027 = ~n3986 & n4026 ;
  buffer buf_n4028( .i (n3144), .o (n4028) );
  buffer buf_n4029( .i (n4028), .o (n4029) );
  buffer buf_n4030( .i (n4029), .o (n4030) );
  buffer buf_n4031( .i (n4030), .o (n4031) );
  assign n4032 = ( n2163 & n4027 ) | ( n2163 & ~n4031 ) | ( n4027 & ~n4031 ) ;
  buffer buf_n4033( .i (n2163), .o (n4033) );
  assign n4034 = n4032 & ~n4033 ;
  assign n4035 = ~n3941 & n4034 ;
  assign n4036 = n3485 & n4035 ;
  buffer buf_n4037( .i (n4036), .o (n4037) );
  buffer buf_n4038( .i (n4037), .o (n4038) );
  buffer buf_n4039( .i (n4038), .o (n4039) );
  buffer buf_n4040( .i (n4039), .o (n4040) );
  buffer buf_n4041( .i (n4040), .o (n4041) );
  buffer buf_n4042( .i (n4041), .o (n4042) );
  buffer buf_n4043( .i (n4042), .o (n4043) );
  assign n4044 = n2760 & ~n3722 ;
  buffer buf_n4045( .i (n4044), .o (n4045) );
  buffer buf_n4046( .i (n4045), .o (n4046) );
  buffer buf_n4047( .i (n4046), .o (n4047) );
  buffer buf_n4048( .i (n4047), .o (n4048) );
  buffer buf_n4049( .i (n4048), .o (n4049) );
  buffer buf_n4050( .i (n4049), .o (n4050) );
  buffer buf_n4051( .i (n4050), .o (n4051) );
  buffer buf_n4052( .i (n4051), .o (n4052) );
  buffer buf_n4053( .i (n4052), .o (n4053) );
  assign n4056 = n2727 | n4053 ;
  assign n4057 = ( ~n4017 & n4043 ) | ( ~n4017 & n4056 ) | ( n4043 & n4056 ) ;
  assign n4058 = n4018 | n4057 ;
  buffer buf_n3644( .i (n3643), .o (n3644) );
  buffer buf_n3645( .i (n3644), .o (n3645) );
  assign n4059 = n1755 | n2840 ;
  assign n4060 = n3645 | n4059 ;
  assign n4061 = ( n1407 & n2814 ) | ( n1407 & n3759 ) | ( n2814 & n3759 ) ;
  assign n4062 = ~n3761 & n4061 ;
  buffer buf_n4063( .i (n4062), .o (n4063) );
  buffer buf_n4064( .i (n4063), .o (n4064) );
  buffer buf_n4065( .i (n4064), .o (n4065) );
  buffer buf_n4066( .i (n4065), .o (n4066) );
  buffer buf_n4067( .i (n4066), .o (n4067) );
  buffer buf_n4068( .i (n4067), .o (n4068) );
  buffer buf_n233( .i (x6), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n4069( .i (n2845), .o (n4069) );
  buffer buf_n4070( .i (n4069), .o (n4070) );
  assign n4071 = n252 & ~n4070 ;
  assign n4072 = ( n166 & n2712 ) | ( n166 & n4071 ) | ( n2712 & n4071 ) ;
  buffer buf_n4073( .i (n2549), .o (n4073) );
  buffer buf_n4074( .i (n4073), .o (n4074) );
  buffer buf_n4075( .i (n4074), .o (n4075) );
  assign n4076 = n4072 & ~n4075 ;
  assign n4077 = n3252 & n4028 ;
  buffer buf_n4078( .i (n4077), .o (n4078) );
  assign n4083 = ( n3986 & n4076 ) | ( n3986 & n4078 ) | ( n4076 & n4078 ) ;
  assign n4084 = ~n3988 & n4083 ;
  assign n4085 = n3516 & n4084 ;
  buffer buf_n4086( .i (n4085), .o (n4086) );
  buffer buf_n136( .i (n135), .o (n136) );
  assign n4093 = ~n163 & n250 ;
  assign n4094 = ( n135 & ~n2549 ) | ( n135 & n4093 ) | ( ~n2549 & n4093 ) ;
  assign n4095 = ~n136 & n4094 ;
  assign n4096 = ~n3591 & n4095 ;
  assign n4097 = ( n3634 & n4025 ) | ( n3634 & n4096 ) | ( n4025 & n4096 ) ;
  assign n4098 = ~n3966 & n4097 ;
  assign n4099 = ( n1575 & n3893 ) | ( n1575 & n4098 ) | ( n3893 & n4098 ) ;
  assign n4100 = ~n3759 & n4099 ;
  buffer buf_n4101( .i (n4100), .o (n4101) );
  assign n4106 = n4086 | n4101 ;
  buffer buf_n4107( .i (n4106), .o (n4107) );
  buffer buf_n4108( .i (n4107), .o (n4108) );
  buffer buf_n4109( .i (n4108), .o (n4109) );
  buffer buf_n4110( .i (n4109), .o (n4110) );
  buffer buf_n4111( .i (n4110), .o (n4111) );
  assign n4112 = n4068 | n4111 ;
  assign n4113 = ( ~n2829 & n4060 ) | ( ~n2829 & n4112 ) | ( n4060 & n4112 ) ;
  assign n4114 = n2830 | n4113 ;
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n224( .i (n223), .o (n224) );
  assign n4115 = n224 & ~n4075 ;
  assign n4116 = ( n168 & ~n3966 ) | ( n168 & n4115 ) | ( ~n3966 & n4115 ) ;
  assign n4117 = ~n169 & n4116 ;
  assign n4118 = ~n3970 & n4117 ;
  buffer buf_n4119( .i (n3664), .o (n4119) );
  assign n4120 = ( n598 & n4118 ) | ( n598 & ~n4119 ) | ( n4118 & ~n4119 ) ;
  assign n4121 = ~n599 & n4120 ;
  assign n4122 = ~n927 & n4121 ;
  assign n4123 = n893 & n4122 ;
  buffer buf_n4124( .i (n4123), .o (n4124) );
  buffer buf_n4125( .i (n4124), .o (n4125) );
  buffer buf_n4126( .i (n4125), .o (n4126) );
  assign n4129 = n2877 | n4126 ;
  assign n4130 = ( ~n1791 & n2865 ) | ( ~n1791 & n4129 ) | ( n2865 & n4129 ) ;
  assign n4131 = n1792 | n4130 ;
  assign n4132 = n4114 | n4131 ;
  assign n4133 = n4058 | n4132 ;
  buffer buf_n3509( .i (n3508), .o (n3509) );
  buffer buf_n3510( .i (n3509), .o (n3510) );
  buffer buf_n3511( .i (n3510), .o (n3511) );
  buffer buf_n3512( .i (n3511), .o (n3512) );
  buffer buf_n3513( .i (n3512), .o (n3513) );
  buffer buf_n3514( .i (n3513), .o (n3514) );
  buffer buf_n4134( .i (n133), .o (n4134) );
  assign n4135 = ( n163 & n1323 ) | ( n163 & n4134 ) | ( n1323 & n4134 ) ;
  buffer buf_n4136( .i (n162), .o (n4136) );
  buffer buf_n4137( .i (n4136), .o (n4137) );
  assign n4138 = n4135 & ~n4137 ;
  assign n4139 = ( n1966 & n3590 ) | ( n1966 & n4138 ) | ( n3590 & n4138 ) ;
  assign n4140 = ~n3591 & n4139 ;
  assign n4141 = ( n1573 & n3692 ) | ( n1573 & n4140 ) | ( n3692 & n4140 ) ;
  assign n4142 = ~n3937 & n4141 ;
  buffer buf_n4143( .i (n4142), .o (n4143) );
  buffer buf_n4144( .i (n4143), .o (n4144) );
  buffer buf_n4145( .i (n4144), .o (n4145) );
  buffer buf_n4146( .i (n4145), .o (n4146) );
  buffer buf_n4147( .i (n4146), .o (n4147) );
  buffer buf_n4148( .i (n4147), .o (n4148) );
  buffer buf_n4149( .i (n4148), .o (n4149) );
  buffer buf_n4150( .i (n4149), .o (n4150) );
  buffer buf_n4151( .i (n4150), .o (n4151) );
  assign n4152 = n2482 | n4151 ;
  assign n4153 = ( ~n2384 & n3514 ) | ( ~n2384 & n4152 ) | ( n3514 & n4152 ) ;
  assign n4154 = n2385 | n4153 ;
  assign n4155 = n2688 | n3862 ;
  assign n4156 = ( ~n2664 & n3543 ) | ( ~n2664 & n4155 ) | ( n3543 & n4155 ) ;
  assign n4157 = n2665 | n4156 ;
  buffer buf_n2462( .i (n2461), .o (n2462) );
  buffer buf_n2463( .i (n2462), .o (n2463) );
  buffer buf_n2464( .i (n2463), .o (n2464) );
  buffer buf_n4158( .i (n2638), .o (n4158) );
  assign n4159 = n219 & n4158 ;
  assign n4160 = ( n2845 & n3569 ) | ( n2845 & n4159 ) | ( n3569 & n4159 ) ;
  buffer buf_n4161( .i (n3569), .o (n4161) );
  assign n4162 = n4160 & ~n4161 ;
  buffer buf_n4163( .i (n4162), .o (n4163) );
  assign n4168 = ~n4028 & n4163 ;
  buffer buf_n4169( .i (n3591), .o (n4169) );
  buffer buf_n4170( .i (n664), .o (n4170) );
  assign n4171 = ( n4168 & n4169 ) | ( n4168 & n4170 ) | ( n4169 & n4170 ) ;
  buffer buf_n4172( .i (n4169), .o (n4172) );
  assign n4173 = n4171 & ~n4172 ;
  assign n4174 = ~n3722 & n4173 ;
  buffer buf_n4175( .i (n3893), .o (n4175) );
  assign n4176 = n4174 & n4175 ;
  buffer buf_n4177( .i (n4176), .o (n4177) );
  buffer buf_n4178( .i (n4177), .o (n4178) );
  buffer buf_n4179( .i (n4178), .o (n4179) );
  buffer buf_n4180( .i (n4179), .o (n4180) );
  buffer buf_n4181( .i (n4180), .o (n4181) );
  buffer buf_n4182( .i (n4181), .o (n4182) );
  assign n4185 = n2504 | n4182 ;
  assign n4186 = ( ~n2463 & n2804 ) | ( ~n2463 & n4185 ) | ( n2804 & n4185 ) ;
  assign n4187 = n2464 | n4186 ;
  assign n4188 = n4157 | n4187 ;
  assign n4189 = n4154 | n4188 ;
  assign n4190 = n2931 | n2989 ;
  buffer buf_n4191( .i (n4190), .o (n4191) );
  buffer buf_n4192( .i (n4191), .o (n4192) );
  buffer buf_n4193( .i (n4192), .o (n4193) );
  buffer buf_n4194( .i (n4193), .o (n4194) );
  assign n4195 = n3714 | n4194 ;
  assign n4196 = ( n3044 & ~n3101 ) | ( n3044 & n4195 ) | ( ~n3101 & n4195 ) ;
  assign n4197 = n3102 | n4196 ;
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n2908( .i (n2907), .o (n2908) );
  assign n4198 = ( n2908 & n3147 ) | ( n2908 & n3937 ) | ( n3147 & n3937 ) ;
  assign n4199 = ~n3893 & n4198 ;
  buffer buf_n4200( .i (n4199), .o (n4200) );
  buffer buf_n4201( .i (n4200), .o (n4201) );
  buffer buf_n4202( .i (n4201), .o (n4202) );
  buffer buf_n4203( .i (n4202), .o (n4203) );
  buffer buf_n4204( .i (n4203), .o (n4204) );
  buffer buf_n4205( .i (n4204), .o (n4205) );
  assign n4208 = n1568 | n4205 ;
  assign n4209 = ( ~n2899 & n2922 ) | ( ~n2899 & n4208 ) | ( n2922 & n4208 ) ;
  assign n4210 = n2900 | n4209 ;
  assign n4211 = n2979 | n4210 ;
  assign n4212 = ( ~n3304 & n4197 ) | ( ~n3304 & n4211 ) | ( n4197 & n4211 ) ;
  assign n4213 = n3305 | n4212 ;
  assign n4214 = n4189 | n4213 ;
  assign n4215 = ( ~n4008 & n4133 ) | ( ~n4008 & n4214 ) | ( n4133 & n4214 ) ;
  assign n4216 = n4009 | n4215 ;
  buffer buf_n2331( .i (n2330), .o (n2331) );
  buffer buf_n2332( .i (n2331), .o (n2332) );
  buffer buf_n2333( .i (n2332), .o (n2333) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  assign n4217 = n2270 | n2339 ;
  buffer buf_n4218( .i (n4217), .o (n4218) );
  buffer buf_n4219( .i (n4218), .o (n4219) );
  buffer buf_n4220( .i (n4219), .o (n4220) );
  buffer buf_n4221( .i (n4220), .o (n4221) );
  assign n4222 = n2345 | n2518 ;
  assign n4223 = n2355 | n4222 ;
  buffer buf_n4224( .i (n4223), .o (n4224) );
  buffer buf_n4225( .i (n4224), .o (n4225) );
  buffer buf_n4226( .i (n4225), .o (n4226) );
  buffer buf_n4227( .i (n4226), .o (n4227) );
  buffer buf_n4228( .i (n4227), .o (n4228) );
  assign n4229 = n1636 | n3312 ;
  assign n4230 = n3945 | n4229 ;
  assign n4231 = n2544 | n4230 ;
  assign n4232 = ( ~n2570 & n2604 ) | ( ~n2570 & n4231 ) | ( n2604 & n4231 ) ;
  assign n4233 = n2571 | n4232 ;
  assign n4234 = n4228 | n4233 ;
  assign n4235 = ( ~n2333 & n4221 ) | ( ~n2333 & n4234 ) | ( n4221 & n4234 ) ;
  assign n4236 = n2334 | n4235 ;
  buffer buf_n4237( .i (n4236), .o (n4237) );
  buffer buf_n4238( .i (n4237), .o (n4238) );
  buffer buf_n3545( .i (n3544), .o (n3545) );
  buffer buf_n3546( .i (n3545), .o (n3546) );
  buffer buf_n3547( .i (n3546), .o (n3547) );
  buffer buf_n2698( .i (n2697), .o (n2698) );
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n2700( .i (n2699), .o (n2700) );
  buffer buf_n2701( .i (n2700), .o (n2701) );
  buffer buf_n2702( .i (n2701), .o (n2702) );
  buffer buf_n3555( .i (n3554), .o (n3555) );
  buffer buf_n3556( .i (n3555), .o (n3556) );
  buffer buf_n3557( .i (n3556), .o (n3557) );
  buffer buf_n3558( .i (n3557), .o (n3558) );
  assign n4239 = n3487 | n3859 ;
  buffer buf_n4240( .i (n4239), .o (n4240) );
  buffer buf_n4241( .i (n4240), .o (n4241) );
  buffer buf_n4242( .i (n4241), .o (n4242) );
  buffer buf_n4243( .i (n4242), .o (n4243) );
  buffer buf_n4244( .i (n4243), .o (n4244) );
  assign n4245 = n3558 | n4244 ;
  assign n4246 = ( n2702 & ~n3546 ) | ( n2702 & n4245 ) | ( ~n3546 & n4245 ) ;
  assign n4247 = n3547 | n4246 ;
  buffer buf_n3608( .i (n3607), .o (n3608) );
  buffer buf_n3609( .i (n3608), .o (n3609) );
  buffer buf_n3610( .i (n3609), .o (n3610) );
  buffer buf_n3611( .i (n3610), .o (n3611) );
  buffer buf_n3612( .i (n3611), .o (n3612) );
  buffer buf_n3613( .i (n3612), .o (n3613) );
  assign n4248 = n3595 | n4143 ;
  buffer buf_n4249( .i (n4248), .o (n4249) );
  buffer buf_n4250( .i (n4249), .o (n4250) );
  buffer buf_n4251( .i (n4250), .o (n4251) );
  buffer buf_n4252( .i (n4251), .o (n4252) );
  buffer buf_n4253( .i (n4252), .o (n4253) );
  buffer buf_n4254( .i (n4253), .o (n4254) );
  assign n4255 = n2476 | n4177 ;
  assign n4256 = n3579 | n4255 ;
  assign n4257 = n3724 | n3735 ;
  buffer buf_n4258( .i (n4257), .o (n4258) );
  assign n4267 = n2799 | n4258 ;
  assign n4268 = ( ~n2501 & n4256 ) | ( ~n2501 & n4267 ) | ( n4256 & n4267 ) ;
  assign n4269 = n2502 | n4268 ;
  assign n4270 = n3531 | n4269 ;
  assign n4271 = ( ~n3612 & n4254 ) | ( ~n3612 & n4270 ) | ( n4254 & n4270 ) ;
  assign n4272 = n3613 | n4271 ;
  buffer buf_n4273( .i (n4272), .o (n4273) );
  buffer buf_n4274( .i (n4273), .o (n4274) );
  assign n4275 = n1752 | n4107 ;
  buffer buf_n4276( .i (n4275), .o (n4276) );
  buffer buf_n4277( .i (n4276), .o (n4277) );
  buffer buf_n4278( .i (n4277), .o (n4278) );
  buffer buf_n4279( .i (n4278), .o (n4279) );
  buffer buf_n4280( .i (n4279), .o (n4280) );
  assign n4281 = n4011 | n4037 ;
  assign n4282 = n4049 | n4281 ;
  assign n4283 = n3035 | n4282 ;
  assign n4284 = ( ~n3301 & n3714 ) | ( ~n3301 & n4283 ) | ( n3714 & n4283 ) ;
  assign n4285 = n3302 | n4284 ;
  assign n4286 = ( n1900 & n2814 ) | ( n1900 & n4175 ) | ( n2814 & n4175 ) ;
  assign n4287 = ~n3761 & n4286 ;
  buffer buf_n4288( .i (n4287), .o (n4288) );
  buffer buf_n4289( .i (n4288), .o (n4289) );
  buffer buf_n4290( .i (n4289), .o (n4290) );
  buffer buf_n4291( .i (n4290), .o (n4291) );
  buffer buf_n4292( .i (n4291), .o (n4292) );
  assign n4301 = n731 & n2811 ;
  assign n4302 = ( n3694 & n3937 ) | ( n3694 & n4301 ) | ( n3937 & n4301 ) ;
  buffer buf_n4303( .i (n3694), .o (n4303) );
  assign n4304 = n4302 & ~n4303 ;
  buffer buf_n4305( .i (n4304), .o (n4305) );
  buffer buf_n4306( .i (n4305), .o (n4306) );
  buffer buf_n4307( .i (n4306), .o (n4307) );
  buffer buf_n4308( .i (n4307), .o (n4308) );
  buffer buf_n4309( .i (n4308), .o (n4309) );
  buffer buf_n4310( .i (n4309), .o (n4310) );
  assign n4312 = n4124 | n4310 ;
  assign n4313 = ( ~n1789 & n4292 ) | ( ~n1789 & n4312 ) | ( n4292 & n4312 ) ;
  assign n4314 = n1790 | n4313 ;
  assign n4315 = n4285 | n4314 ;
  assign n4316 = ( ~n4273 & n4280 ) | ( ~n4273 & n4315 ) | ( n4280 & n4315 ) ;
  assign n4317 = n4274 | n4316 ;
  buffer buf_n3979( .i (n3978), .o (n3979) );
  buffer buf_n3980( .i (n3979), .o (n3980) );
  buffer buf_n3981( .i (n3980), .o (n3981) );
  buffer buf_n4000( .i (n3999), .o (n4000) );
  buffer buf_n4001( .i (n4000), .o (n4001) );
  buffer buf_n4002( .i (n4001), .o (n4002) );
  assign n4318 = n3981 | n4002 ;
  buffer buf_n4319( .i (n3239), .o (n4319) );
  assign n4320 = n3783 & ~n4319 ;
  buffer buf_n4321( .i (n3692), .o (n4321) );
  buffer buf_n4322( .i (n4321), .o (n4322) );
  assign n4323 = n4320 & n4322 ;
  buffer buf_n4324( .i (n4323), .o (n4324) );
  buffer buf_n4325( .i (n4324), .o (n4325) );
  buffer buf_n4326( .i (n4325), .o (n4326) );
  assign n4334 = n3788 | n4326 ;
  buffer buf_n4335( .i (n4334), .o (n4335) );
  buffer buf_n4336( .i (n4335), .o (n4336) );
  buffer buf_n4337( .i (n4336), .o (n4337) );
  buffer buf_n4338( .i (n4337), .o (n4338) );
  buffer buf_n4339( .i (n4338), .o (n4339) );
  buffer buf_n4340( .i (n4339), .o (n4340) );
  assign n4341 = n3331 | n4340 ;
  assign n4342 = n4318 | n4341 ;
  assign n4343 = n4317 | n4342 ;
  assign n4344 = ( ~n4237 & n4247 ) | ( ~n4237 & n4343 ) | ( n4247 & n4343 ) ;
  assign n4345 = n4238 | n4344 ;
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n3924( .i (n3923), .o (n3924) );
  buffer buf_n3925( .i (n3924), .o (n3925) );
  buffer buf_n3926( .i (n3925), .o (n3926) );
  buffer buf_n3927( .i (n3926), .o (n3927) );
  buffer buf_n3928( .i (n3927), .o (n3928) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  assign n4346 = n1124 & n3927 ;
  assign n4347 = ( n1157 & n3928 ) | ( n1157 & n4346 ) | ( n3928 & n4346 ) ;
  buffer buf_n4348( .i (n4347), .o (n4348) );
  buffer buf_n3901( .i (n3900), .o (n3901) );
  buffer buf_n3902( .i (n3901), .o (n3902) );
  buffer buf_n3903( .i (n3902), .o (n3903) );
  buffer buf_n3810( .i (n3809), .o (n3810) );
  buffer buf_n3811( .i (n3810), .o (n3811) );
  assign n4349 = n3811 | n3955 ;
  assign n4350 = ( ~n3343 & n3826 ) | ( ~n3343 & n4349 ) | ( n3826 & n4349 ) ;
  assign n4351 = n3344 | n4350 ;
  assign n4352 = n3903 | n4351 ;
  assign n4353 = ( ~n3120 & n4348 ) | ( ~n3120 & n4352 ) | ( n4348 & n4352 ) ;
  assign n4354 = n3121 | n4353 ;
  buffer buf_n4355( .i (n4354), .o (n4355) );
  buffer buf_n4356( .i (n4355), .o (n4356) );
  buffer buf_n2597( .i (n2596), .o (n2597) );
  buffer buf_n2598( .i (n2597), .o (n2598) );
  buffer buf_n2689( .i (n2688), .o (n2689) );
  buffer buf_n2690( .i (n2689), .o (n2690) );
  buffer buf_n2691( .i (n2690), .o (n2691) );
  assign n4357 = n3329 | n3543 ;
  assign n4358 = ( ~n2690 & n2700 ) | ( ~n2690 & n4357 ) | ( n2700 & n4357 ) ;
  assign n4359 = n2691 | n4358 ;
  buffer buf_n4327( .i (n4326), .o (n4327) );
  buffer buf_n4328( .i (n4327), .o (n4328) );
  buffer buf_n4329( .i (n4328), .o (n4329) );
  buffer buf_n4330( .i (n4329), .o (n4330) );
  buffer buf_n4331( .i (n4330), .o (n4331) );
  buffer buf_n4332( .i (n4331), .o (n4332) );
  buffer buf_n4333( .i (n4332), .o (n4333) );
  assign n4360 = n2610 | n3943 ;
  buffer buf_n4361( .i (n4360), .o (n4361) );
  buffer buf_n4362( .i (n4361), .o (n4362) );
  buffer buf_n4363( .i (n4362), .o (n4363) );
  buffer buf_n4364( .i (n4363), .o (n4364) );
  buffer buf_n4365( .i (n4364), .o (n4365) );
  buffer buf_n4366( .i (n4365), .o (n4366) );
  assign n4367 = n4333 | n4366 ;
  assign n4368 = ( ~n2597 & n4359 ) | ( ~n2597 & n4367 ) | ( n4359 & n4367 ) ;
  assign n4369 = n2598 | n4368 ;
  buffer buf_n3847( .i (n3846), .o (n3847) );
  buffer buf_n3848( .i (n3847), .o (n3848) );
  buffer buf_n2972( .i (n2971), .o (n2972) );
  buffer buf_n2909( .i (n2908), .o (n2909) );
  buffer buf_n2910( .i (n2909), .o (n2910) );
  assign n4370 = ( n1576 & n2910 ) | ( n1576 & n4175 ) | ( n2910 & n4175 ) ;
  buffer buf_n4371( .i (n4175), .o (n4371) );
  assign n4372 = n4370 & ~n4371 ;
  buffer buf_n4373( .i (n4372), .o (n4373) );
  buffer buf_n4374( .i (n4373), .o (n4374) );
  buffer buf_n4375( .i (n4374), .o (n4375) );
  assign n4380 = n3220 | n3389 ;
  assign n4381 = ( ~n2971 & n4375 ) | ( ~n2971 & n4380 ) | ( n4375 & n4380 ) ;
  assign n4382 = n2972 | n4381 ;
  assign n4383 = n3361 | n3372 ;
  assign n4384 = ( ~n3847 & n4382 ) | ( ~n3847 & n4383 ) | ( n4382 & n4383 ) ;
  assign n4385 = n3848 | n4384 ;
  buffer buf_n4386( .i (n4385), .o (n4386) );
  buffer buf_n4387( .i (n4386), .o (n4387) );
  buffer buf_n3433( .i (n3432), .o (n3433) );
  buffer buf_n3434( .i (n3433), .o (n3434) );
  buffer buf_n3450( .i (n3449), .o (n3450) );
  buffer buf_n3438( .i (n3437), .o (n3438) );
  buffer buf_n3439( .i (n3438), .o (n3439) );
  buffer buf_n3440( .i (n3439), .o (n3440) );
  buffer buf_n669( .i (n668), .o (n669) );
  assign n4388 = ( n669 & ~n3439 ) | ( n669 & n3941 ) | ( ~n3439 & n3941 ) ;
  assign n4389 = ( n3410 & n3440 ) | ( n3410 & n4388 ) | ( n3440 & n4388 ) ;
  buffer buf_n4390( .i (n4389), .o (n4390) );
  buffer buf_n4391( .i (n4390), .o (n4391) );
  buffer buf_n4392( .i (n4391), .o (n4392) );
  buffer buf_n4393( .i (n4392), .o (n4393) );
  buffer buf_n4394( .i (n4393), .o (n4394) );
  assign n4395 = n3450 | n4394 ;
  assign n4396 = n3434 | n4395 ;
  assign n4397 = n3230 | n3278 ;
  buffer buf_n4398( .i (n4397), .o (n4398) );
  buffer buf_n4399( .i (n4398), .o (n4399) );
  assign n4400 = ( ~n2992 & n3262 ) | ( ~n2992 & n3399 ) | ( n3262 & n3399 ) ;
  assign n4401 = n2993 | n4400 ;
  buffer buf_n2893( .i (n2892), .o (n2893) );
  buffer buf_n2894( .i (n2893), .o (n2894) );
  assign n4402 = n2894 | n3205 ;
  assign n4403 = n2920 | n4402 ;
  assign n4404 = n3032 | n3710 ;
  assign n4405 = ( ~n3021 & n3286 ) | ( ~n3021 & n4404 ) | ( n3286 & n4404 ) ;
  assign n4406 = n3022 | n4405 ;
  assign n4407 = n4403 | n4406 ;
  assign n4408 = ( ~n4398 & n4401 ) | ( ~n4398 & n4407 ) | ( n4401 & n4407 ) ;
  assign n4409 = n4399 | n4408 ;
  assign n4410 = n3477 | n4409 ;
  assign n4411 = ( ~n4386 & n4396 ) | ( ~n4386 & n4410 ) | ( n4396 & n4410 ) ;
  assign n4412 = n4387 | n4411 ;
  buffer buf_n3842( .i (n3841), .o (n3842) );
  buffer buf_n3843( .i (n3842), .o (n3843) );
  assign n4413 = n2458 | n3579 ;
  buffer buf_n4414( .i (n4413), .o (n4414) );
  buffer buf_n4415( .i (n4414), .o (n4415) );
  buffer buf_n4416( .i (n4415), .o (n4416) );
  buffer buf_n4417( .i (n4416), .o (n4417) );
  buffer buf_n4418( .i (n4417), .o (n4418) );
  buffer buf_n4419( .i (n4418), .o (n4419) );
  assign n4420 = n2404 | n2671 ;
  assign n4421 = ( ~n2433 & n3158 ) | ( ~n2433 & n4420 ) | ( n3158 & n4420 ) ;
  assign n4422 = n2434 | n4421 ;
  assign n4423 = n3511 | n3626 ;
  assign n4424 = ( ~n2382 & n4422 ) | ( ~n2382 & n4423 ) | ( n4422 & n4423 ) ;
  assign n4425 = n2383 | n4424 ;
  assign n4426 = n2838 | n4065 ;
  assign n4427 = n2826 | n4426 ;
  assign n4428 = n3741 | n4427 ;
  assign n4429 = n3645 | n4428 ;
  assign n4430 = n4425 | n4429 ;
  assign n4431 = ( ~n3842 & n4419 ) | ( ~n3842 & n4430 ) | ( n4419 & n4430 ) ;
  assign n4432 = n3843 | n4431 ;
  assign n4433 = n4412 | n4432 ;
  assign n4434 = ( ~n4355 & n4369 ) | ( ~n4355 & n4433 ) | ( n4369 & n4433 ) ;
  assign n4435 = n4356 | n4434 ;
  buffer buf_n3668( .i (n3667), .o (n3668) );
  buffer buf_n3669( .i (n3668), .o (n3669) );
  buffer buf_n3670( .i (n3669), .o (n3670) );
  assign n4436 = n2862 | n3670 ;
  assign n4437 = n2876 | n4436 ;
  assign n4438 = n2725 | n2977 ;
  assign n4439 = n4437 | n4438 ;
  buffer buf_n4440( .i (n4439), .o (n4440) );
  buffer buf_n4441( .i (n4440), .o (n4441) );
  buffer buf_n3646( .i (n3645), .o (n3646) );
  assign n4442 = n3659 | n4065 ;
  buffer buf_n4443( .i (n4442), .o (n4443) );
  assign n4447 = n2840 | n4443 ;
  assign n4448 = ( n2828 & ~n3645 ) | ( n2828 & n4447 ) | ( ~n3645 & n4447 ) ;
  assign n4449 = n3646 | n4448 ;
  buffer buf_n4376( .i (n4375), .o (n4376) );
  buffer buf_n4377( .i (n4376), .o (n4377) );
  buffer buf_n4378( .i (n4377), .o (n4378) );
  assign n4450 = n2897 | n2934 ;
  assign n4451 = n1568 | n4450 ;
  assign n4452 = n2922 | n4451 ;
  assign n4453 = n4378 | n4452 ;
  assign n4454 = n3023 | n3099 ;
  assign n4455 = ( ~n2994 & n3714 ) | ( ~n2994 & n4454 ) | ( n3714 & n4454 ) ;
  assign n4456 = n2995 | n4455 ;
  assign n4457 = n4453 | n4456 ;
  assign n4458 = ( ~n4440 & n4449 ) | ( ~n4440 & n4457 ) | ( n4449 & n4457 ) ;
  assign n4459 = n4441 | n4458 ;
  buffer buf_n4460( .i (n4459), .o (n4460) );
  buffer buf_n4461( .i (n4460), .o (n4461) );
  buffer buf_n3520( .i (n3519), .o (n3520) );
  buffer buf_n3521( .i (n3520), .o (n3521) );
  buffer buf_n3522( .i (n3521), .o (n3522) );
  buffer buf_n3523( .i (n3522), .o (n3523) );
  buffer buf_n3524( .i (n3523), .o (n3524) );
  buffer buf_n3525( .i (n3524), .o (n3525) );
  buffer buf_n3526( .i (n3525), .o (n3526) );
  buffer buf_n3527( .i (n3526), .o (n3527) );
  buffer buf_n3528( .i (n3527), .o (n3528) );
  buffer buf_n3614( .i (n3613), .o (n3614) );
  buffer buf_n3615( .i (n3614), .o (n3615) );
  assign n4462 = ~n2957 & n4161 ;
  buffer buf_n4463( .i (n4462), .o (n4463) );
  assign n4466 = ( n340 & n2036 ) | ( n340 & n4463 ) | ( n2036 & n4463 ) ;
  buffer buf_n4467( .i (n4466), .o (n4467) );
  assign n4468 = ~n3966 & n4467 ;
  assign n4469 = n4303 & n4468 ;
  assign n4470 = ( n765 & n3970 ) | ( n765 & n4469 ) | ( n3970 & n4469 ) ;
  assign n4471 = ~n3972 & n4470 ;
  buffer buf_n4472( .i (n4471), .o (n4472) );
  buffer buf_n4473( .i (n4472), .o (n4473) );
  buffer buf_n4474( .i (n4473), .o (n4474) );
  buffer buf_n4475( .i (n4474), .o (n4475) );
  buffer buf_n4476( .i (n4475), .o (n4476) );
  buffer buf_n4477( .i (n4476), .o (n4477) );
  buffer buf_n4478( .i (n4477), .o (n4478) );
  assign n4479 = n2464 | n4478 ;
  assign n4480 = n3615 | n4479 ;
  assign n4481 = n2386 | n4480 ;
  assign n4482 = n3528 | n4481 ;
  buffer buf_n3777( .i (n3776), .o (n3777) );
  buffer buf_n3778( .i (n3777), .o (n3778) );
  assign n4483 = n2687 | n3489 ;
  assign n4484 = n3555 | n4483 ;
  assign n4485 = n3793 | n4484 ;
  assign n4486 = ( n2616 & ~n3136 ) | ( n2616 & n4485 ) | ( ~n3136 & n4485 ) ;
  assign n4487 = n3137 | n4486 ;
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n3948( .i (n3947), .o (n3948) );
  assign n4488 = ( ~n1058 & n1092 ) | ( ~n1058 & n3948 ) | ( n1092 & n3948 ) ;
  buffer buf_n3909( .i (n3908), .o (n3909) );
  buffer buf_n3910( .i (n3909), .o (n3910) );
  buffer buf_n3911( .i (n3910), .o (n3911) );
  buffer buf_n3912( .i (n3911), .o (n3912) );
  buffer buf_n3913( .i (n3912), .o (n3913) );
  buffer buf_n3914( .i (n3913), .o (n3914) );
  buffer buf_n3915( .i (n3914), .o (n3915) );
  assign n4489 = n3915 | n3948 ;
  assign n4490 = ( n1059 & n4488 ) | ( n1059 & n4489 ) | ( n4488 & n4489 ) ;
  assign n4491 = n4348 | n4490 ;
  assign n4492 = n4487 | n4491 ;
  assign n4493 = n3778 | n4492 ;
  assign n4494 = ( ~n4460 & n4482 ) | ( ~n4460 & n4493 ) | ( n4482 & n4493 ) ;
  assign n4495 = n4461 | n4494 ;
  buffer buf_n3794( .i (n3793), .o (n3794) );
  buffer buf_n3180( .i (n3179), .o (n3180) );
  assign n4496 = n2614 | n3180 ;
  assign n4497 = ( n3140 & ~n3793 ) | ( n3140 & n4496 ) | ( ~n3793 & n4496 ) ;
  assign n4498 = n3794 | n4497 ;
  assign n4499 = ~n1051 & n1085 ;
  assign n4500 = n3909 & n4499 ;
  buffer buf_n4501( .i (n4500), .o (n4501) );
  buffer buf_n4502( .i (n4501), .o (n4502) );
  buffer buf_n4503( .i (n4502), .o (n4503) );
  buffer buf_n4504( .i (n4503), .o (n4504) );
  buffer buf_n4505( .i (n4504), .o (n4505) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  assign n4506 = ~n986 & n1017 ;
  buffer buf_n4507( .i (n4506), .o (n4507) );
  buffer buf_n4508( .i (n4507), .o (n4508) );
  buffer buf_n4509( .i (n4508), .o (n4509) );
  buffer buf_n4510( .i (n4509), .o (n4510) );
  buffer buf_n4511( .i (n4510), .o (n4511) );
  buffer buf_n961( .i (n960), .o (n961) );
  assign n4512 = ~n961 & n3882 ;
  buffer buf_n4513( .i (n4512), .o (n4513) );
  assign n4517 = ( n992 & n4511 ) | ( n992 & n4513 ) | ( n4511 & n4513 ) ;
  buffer buf_n4518( .i (n4517), .o (n4518) );
  assign n4521 = n4505 | n4518 ;
  assign n4522 = n3959 | n4521 ;
  assign n4523 = ( ~n3120 & n4498 ) | ( ~n3120 & n4522 ) | ( n4498 & n4522 ) ;
  assign n4524 = n3121 | n4523 ;
  buffer buf_n4525( .i (n4524), .o (n4525) );
  buffer buf_n4526( .i (n4525), .o (n4526) );
  assign n4527 = n2379 | n3520 ;
  buffer buf_n4528( .i (n4527), .o (n4528) );
  buffer buf_n4529( .i (n4528), .o (n4529) );
  buffer buf_n4530( .i (n4529), .o (n4530) );
  assign n4531 = n3161 | n4530 ;
  buffer buf_n4532( .i (n4531), .o (n4532) );
  assign n4533 = n3558 | n4532 ;
  assign n4534 = ( n3494 & ~n3546 ) | ( n3494 & n4533 ) | ( ~n3546 & n4533 ) ;
  assign n4535 = n3547 | n4534 ;
  buffer buf_n2507( .i (n2506), .o (n2507) );
  buffer buf_n3765( .i (n3764), .o (n3765) );
  buffer buf_n3766( .i (n3765), .o (n3766) );
  buffer buf_n3767( .i (n3766), .o (n3767) );
  buffer buf_n3768( .i (n3767), .o (n3768) );
  buffer buf_n3660( .i (n3659), .o (n3660) );
  assign n4536 = n2826 | n3660 ;
  buffer buf_n4537( .i (n2839), .o (n4537) );
  assign n4538 = n4536 | n4537 ;
  assign n4539 = n3768 | n4538 ;
  assign n4540 = ( ~n2506 & n3646 ) | ( ~n2506 & n4539 ) | ( n3646 & n4539 ) ;
  assign n4541 = n2507 | n4540 ;
  buffer buf_n2973( .i (n2972), .o (n2973) );
  buffer buf_n2974( .i (n2973), .o (n2974) );
  buffer buf_n2975( .i (n2974), .o (n2975) );
  assign n4542 = n1562 | n2915 ;
  buffer buf_n4543( .i (n4542), .o (n4543) );
  buffer buf_n4544( .i (n4543), .o (n4544) );
  buffer buf_n4545( .i (n4544), .o (n4545) );
  buffer buf_n4546( .i (n4545), .o (n4546) );
  buffer buf_n4547( .i (n4546), .o (n4547) );
  buffer buf_n4548( .i (n4547), .o (n4548) );
  buffer buf_n4549( .i (n4548), .o (n4549) );
  assign n4552 = n3039 | n3096 ;
  assign n4553 = ( ~n2896 & n4191 ) | ( ~n2896 & n4552 ) | ( n4191 & n4552 ) ;
  assign n4554 = n2897 | n4553 ;
  buffer buf_n4555( .i (n4554), .o (n4555) );
  assign n4560 = n2953 | n4012 ;
  assign n4561 = n4050 | n4560 ;
  assign n4562 = n4555 | n4561 ;
  assign n4563 = ( ~n2974 & n4549 ) | ( ~n2974 & n4562 ) | ( n4549 & n4562 ) ;
  assign n4564 = n2975 | n4563 ;
  assign n4565 = n2874 | n4290 ;
  buffer buf_n4566( .i (n4565), .o (n4566) );
  buffer buf_n4567( .i (n4566), .o (n4567) );
  buffer buf_n4311( .i (n4310), .o (n4311) );
  assign n4568 = n2720 | n3666 ;
  buffer buf_n4569( .i (n4568), .o (n4569) );
  buffer buf_n4570( .i (n4569), .o (n4570) );
  buffer buf_n4571( .i (n4570), .o (n4571) );
  buffer buf_n4572( .i (n4571), .o (n4572) );
  assign n4573 = n4311 | n4572 ;
  assign n4574 = ( ~n2864 & n4567 ) | ( ~n2864 & n4573 ) | ( n4567 & n4573 ) ;
  assign n4575 = n2865 | n4574 ;
  assign n4576 = n4564 | n4575 ;
  assign n4577 = n4541 | n4576 ;
  buffer buf_n3749( .i (n3748), .o (n3749) );
  buffer buf_n3750( .i (n3749), .o (n3750) );
  buffer buf_n3751( .i (n3750), .o (n3751) );
  buffer buf_n3752( .i (n3751), .o (n3752) );
  buffer buf_n3753( .i (n3752), .o (n3753) );
  buffer buf_n3742( .i (n3741), .o (n3742) );
  buffer buf_n3743( .i (n3742), .o (n3743) );
  buffer buf_n3618( .i (n3617), .o (n3618) );
  buffer buf_n3619( .i (n3618), .o (n3619) );
  buffer buf_n3620( .i (n3619), .o (n3620) );
  buffer buf_n3621( .i (n3620), .o (n3621) );
  buffer buf_n3622( .i (n3621), .o (n3622) );
  assign n4578 = n3512 | n3622 ;
  assign n4579 = n3603 | n4578 ;
  assign n4580 = n3743 | n4579 ;
  assign n4581 = ( ~n3752 & n4419 ) | ( ~n3752 & n4580 ) | ( n4419 & n4580 ) ;
  assign n4582 = n3753 | n4581 ;
  assign n4583 = n4577 | n4582 ;
  assign n4584 = ( ~n4525 & n4535 ) | ( ~n4525 & n4583 ) | ( n4535 & n4583 ) ;
  assign n4585 = n4526 | n4584 ;
  buffer buf_n2411( .i (n2410), .o (n2411) );
  buffer buf_n2412( .i (n2411), .o (n2412) );
  buffer buf_n2413( .i (n2412), .o (n2413) );
  buffer buf_n2414( .i (n2413), .o (n2414) );
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n2436( .i (n2435), .o (n2436) );
  buffer buf_n2437( .i (n2436), .o (n2437) );
  buffer buf_n2438( .i (n2437), .o (n2438) );
  buffer buf_n2439( .i (n2438), .o (n2439) );
  buffer buf_n2440( .i (n2439), .o (n2440) );
  buffer buf_n2441( .i (n2440), .o (n2441) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  buffer buf_n2443( .i (n2442), .o (n2443) );
  assign n4586 = n3111 | n3895 ;
  assign n4587 = n3338 | n4586 ;
  buffer buf_n4588( .i (n4587), .o (n4588) );
  assign n4591 = n2324 | n3806 ;
  buffer buf_n4592( .i (n4591), .o (n4592) );
  assign n4596 = n3952 | n4592 ;
  assign n4597 = ( ~n2269 & n4588 ) | ( ~n2269 & n4596 ) | ( n4588 & n4596 ) ;
  assign n4598 = n2270 | n4597 ;
  buffer buf_n4599( .i (n4598), .o (n4599) );
  buffer buf_n4600( .i (n4599), .o (n4600) );
  assign n4601 = ( n959 & n3880 ) | ( n959 & n4507 ) | ( n3880 & n4507 ) ;
  assign n4602 = ~n960 & n4601 ;
  buffer buf_n4603( .i (n4602), .o (n4603) );
  buffer buf_n4604( .i (n4603), .o (n4604) );
  assign n4607 = n1055 | n4603 ;
  assign n4608 = ( n3913 & n4604 ) | ( n3913 & n4607 ) | ( n4604 & n4607 ) ;
  assign n4609 = ( ~n1121 & n1153 ) | ( ~n1121 & n4501 ) | ( n1153 & n4501 ) ;
  assign n4610 = n3924 | n4501 ;
  assign n4611 = ( n1122 & n4609 ) | ( n1122 & n4610 ) | ( n4609 & n4610 ) ;
  assign n4612 = n3890 | n4611 ;
  assign n4613 = ( ~n4599 & n4608 ) | ( ~n4599 & n4612 ) | ( n4608 & n4612 ) ;
  assign n4614 = n4600 | n4613 ;
  buffer buf_n4615( .i (n4614), .o (n4615) );
  buffer buf_n4616( .i (n4615), .o (n4616) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  assign n4617 = n2570 | n3826 ;
  assign n4618 = ( ~n2524 & n2546 ) | ( ~n2524 & n4617 ) | ( n2546 & n4617 ) ;
  assign n4619 = n2525 | n4618 ;
  buffer buf_n2361( .i (n2360), .o (n2361) );
  buffer buf_n2362( .i (n2361), .o (n2362) );
  buffer buf_n2605( .i (n2604), .o (n2605) );
  assign n4620 = n2634 | n3313 ;
  assign n4621 = n3977 | n4620 ;
  assign n4622 = n3946 | n3962 ;
  assign n4623 = ( ~n2604 & n4621 ) | ( ~n2604 & n4622 ) | ( n4621 & n4622 ) ;
  assign n4624 = n2605 | n4623 ;
  assign n4625 = n2362 | n4624 ;
  assign n4626 = ( ~n4615 & n4619 ) | ( ~n4615 & n4625 ) | ( n4619 & n4625 ) ;
  assign n4627 = n4616 | n4626 ;
  buffer buf_n4628( .i (n4627), .o (n4628) );
  buffer buf_n4629( .i (n4628), .o (n4629) );
  buffer buf_n3364( .i (n3363), .o (n3364) );
  assign n4630 = n3217 | n4200 ;
  buffer buf_n4631( .i (n4630), .o (n4631) );
  assign n4638 = n2969 | n4631 ;
  assign n4639 = n4374 | n4638 ;
  assign n4640 = n3197 | n4639 ;
  assign n4641 = ( ~n2898 & n4547 ) | ( ~n2898 & n4640 ) | ( n4547 & n4640 ) ;
  assign n4642 = n2899 | n4641 ;
  assign n4643 = ~n338 & n1649 ;
  assign n4644 = ~n457 & n4643 ;
  buffer buf_n4645( .i (n4070), .o (n4645) );
  assign n4646 = ( n1800 & n4644 ) | ( n1800 & n4645 ) | ( n4644 & n4645 ) ;
  assign n4647 = ~n4025 & n4646 ;
  assign n4648 = n4172 & n4647 ;
  assign n4649 = ( n764 & n4031 ) | ( n764 & n4648 ) | ( n4031 & n4648 ) ;
  assign n4650 = ~n3664 & n4649 ;
  buffer buf_n4651( .i (n3516), .o (n4651) );
  assign n4652 = n4650 & n4651 ;
  buffer buf_n4653( .i (n4652), .o (n4653) );
  buffer buf_n4654( .i (n4653), .o (n4654) );
  buffer buf_n4655( .i (n4654), .o (n4655) );
  buffer buf_n4656( .i (n4655), .o (n4656) );
  buffer buf_n3379( .i (n3378), .o (n3379) );
  buffer buf_n3380( .i (n3379), .o (n3380) );
  buffer buf_n3381( .i (n3380), .o (n3381) );
  assign n4663 = n221 & ~n4069 ;
  assign n4664 = ( n339 & n4073 ) | ( n339 & n4663 ) | ( n4073 & n4663 ) ;
  buffer buf_n4665( .i (n339), .o (n4665) );
  assign n4666 = n4664 & ~n4665 ;
  buffer buf_n4667( .i (n4666), .o (n4667) );
  buffer buf_n4668( .i (n4667), .o (n4668) );
  assign n4669 = ( n1858 & n4172 ) | ( n1858 & ~n4667 ) | ( n4172 & ~n4667 ) ;
  assign n4670 = n4668 & n4669 ;
  buffer buf_n4671( .i (n4031), .o (n4671) );
  buffer buf_n4672( .i (n3515), .o (n4672) );
  assign n4673 = ( n4670 & n4671 ) | ( n4670 & n4672 ) | ( n4671 & n4672 ) ;
  assign n4674 = ~n4119 & n4673 ;
  buffer buf_n4675( .i (n4674), .o (n4675) );
  buffer buf_n4676( .i (n4675), .o (n4676) );
  assign n4684 = n2952 | n4676 ;
  assign n4685 = ( n3381 & ~n4655 ) | ( n3381 & n4684 ) | ( ~n4655 & n4684 ) ;
  assign n4686 = n4656 | n4685 ;
  assign n4687 = n3373 | n4686 ;
  assign n4688 = ( ~n3363 & n4642 ) | ( ~n3363 & n4687 ) | ( n4642 & n4687 ) ;
  assign n4689 = n3364 | n4688 ;
  buffer buf_n4690( .i (n4689), .o (n4690) );
  buffer buf_n4691( .i (n4690), .o (n4691) );
  buffer buf_n3266( .i (n3265), .o (n3266) );
  assign n4692 = ~n338 & n4069 ;
  assign n4693 = ~n4073 & n4692 ;
  buffer buf_n4694( .i (n3590), .o (n4694) );
  assign n4695 = n4693 & n4694 ;
  assign n4696 = ( n762 & n4029 ) | ( n762 & n4695 ) | ( n4029 & n4695 ) ;
  assign n4697 = ~n4030 & n4696 ;
  buffer buf_n4698( .i (n1345), .o (n4698) );
  buffer buf_n4699( .i (n4698), .o (n4699) );
  assign n4700 = n4697 & n4699 ;
  buffer buf_n4701( .i (n4700), .o (n4701) );
  buffer buf_n4702( .i (n4701), .o (n4702) );
  buffer buf_n4703( .i (n4702), .o (n4703) );
  buffer buf_n4704( .i (n4703), .o (n4704) );
  buffer buf_n4705( .i (n4704), .o (n4705) );
  buffer buf_n4706( .i (n4705), .o (n4706) );
  buffer buf_n4707( .i (n4706), .o (n4707) );
  buffer buf_n4708( .i (n4707), .o (n4708) );
  assign n4711 = n3078 | n4708 ;
  assign n4712 = ( ~n2996 & n3266 ) | ( ~n2996 & n4711 ) | ( n3266 & n4711 ) ;
  assign n4713 = n2997 | n4712 ;
  buffer buf_n3402( .i (n3401), .o (n3402) );
  buffer buf_n3403( .i (n3402), .o (n3403) );
  buffer buf_n3404( .i (n3403), .o (n3404) );
  buffer buf_n3025( .i (n3024), .o (n3025) );
  buffer buf_n3026( .i (n3025), .o (n3026) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  assign n4714 = ( n344 & ~n565 ) | ( n344 & n1454 ) | ( ~n565 & n1454 ) ;
  assign n4715 = ~n345 & n4714 ;
  assign n4716 = n767 & n4715 ;
  assign n4717 = n635 & n4716 ;
  buffer buf_n4718( .i (n4717), .o (n4718) );
  buffer buf_n4719( .i (n4718), .o (n4719) );
  assign n4723 = n3288 | n4719 ;
  buffer buf_n4724( .i (n4723), .o (n4724) );
  buffer buf_n3683( .i (n3682), .o (n3683) );
  buffer buf_n3684( .i (n3683), .o (n3684) );
  buffer buf_n3685( .i (n3684), .o (n3685) );
  buffer buf_n3686( .i (n3685), .o (n3686) );
  buffer buf_n3687( .i (n3686), .o (n3687) );
  buffer buf_n3688( .i (n3687), .o (n3688) );
  assign n4729 = n3058 | n3271 ;
  assign n4730 = ( n3034 & ~n3087 ) | ( n3034 & n4729 ) | ( ~n3087 & n4729 ) ;
  assign n4731 = n3088 | n4730 ;
  assign n4732 = n3688 | n4731 ;
  assign n4733 = ( ~n3025 & n4724 ) | ( ~n3025 & n4732 ) | ( n4724 & n4732 ) ;
  assign n4734 = n3026 | n4733 ;
  assign n4735 = n3404 | n4734 ;
  assign n4736 = ( ~n4690 & n4713 ) | ( ~n4690 & n4735 ) | ( n4713 & n4735 ) ;
  assign n4737 = n4691 | n4736 ;
  buffer buf_n3552( .i (n3551), .o (n3552) );
  assign n4738 = ~n342 & n4467 ;
  buffer buf_n4739( .i (n4738), .o (n4739) );
  buffer buf_n4740( .i (n4739), .o (n4740) );
  assign n4741 = ~n4371 & n4740 ;
  assign n4742 = ( n634 & n767 ) | ( n634 & n4741 ) | ( n767 & n4741 ) ;
  assign n4743 = ~n635 & n4742 ;
  assign n4744 = n928 & n4743 ;
  assign n4745 = ( n929 & n3552 ) | ( n929 & n4744 ) | ( n3552 & n4744 ) ;
  buffer buf_n4746( .i (n4745), .o (n4746) );
  assign n4748 = n2683 | n3323 ;
  assign n4749 = n3538 | n4748 ;
  assign n4750 = n3993 | n4749 ;
  assign n4751 = n4335 | n4750 ;
  assign n4752 = n4240 | n4751 ;
  assign n4753 = ( ~n2698 & n4746 ) | ( ~n2698 & n4752 ) | ( n4746 & n4752 ) ;
  assign n4754 = n2699 | n4753 ;
  buffer buf_n4755( .i (n4754), .o (n4755) );
  buffer buf_n4756( .i (n4755), .o (n4756) );
  assign n4757 = n3728 | n4414 ;
  assign n4758 = n4181 | n4757 ;
  assign n4759 = n3838 | n4475 ;
  assign n4760 = ( ~n4150 & n4758 ) | ( ~n4150 & n4759 ) | ( n4758 & n4759 ) ;
  assign n4761 = n4151 | n4760 ;
  buffer buf_n4762( .i (n3567), .o (n4762) );
  buffer buf_n4763( .i (n556), .o (n4763) );
  buffer buf_n4764( .i (n4763), .o (n4764) );
  assign n4765 = n4762 & ~n4764 ;
  buffer buf_n4766( .i (n4765), .o (n4766) );
  buffer buf_n4767( .i (n4766), .o (n4767) );
  buffer buf_n4768( .i (n4767), .o (n4768) );
  buffer buf_n4769( .i (n4768), .o (n4769) );
  assign n4770 = ( n342 & ~n2162 ) | ( n342 & n4769 ) | ( ~n2162 & n4769 ) ;
  assign n4771 = ~n343 & n4770 ;
  assign n4772 = n3654 & n4771 ;
  assign n4773 = ( n766 & n3972 ) | ( n766 & n4772 ) | ( n3972 & n4772 ) ;
  assign n4774 = ~n634 & n4773 ;
  buffer buf_n4775( .i (n4774), .o (n4775) );
  buffer buf_n4776( .i (n4775), .o (n4776) );
  assign n4777 = n3610 | n4776 ;
  assign n4778 = ( ~n3511 & n3621 ) | ( ~n3511 & n4777 ) | ( n3621 & n4777 ) ;
  assign n4779 = n3512 | n4778 ;
  buffer buf_n4780( .i (n4779), .o (n4780) );
  assign n4781 = n4761 | n4780 ;
  assign n4782 = ( n4532 & ~n4755 ) | ( n4532 & n4781 ) | ( ~n4755 & n4781 ) ;
  assign n4783 = n4756 | n4782 ;
  assign n4784 = ( n3471 & ~n4037 ) | ( n3471 & n4569 ) | ( ~n4037 & n4569 ) ;
  assign n4785 = n4038 | n4784 ;
  assign n4786 = n4124 | n4785 ;
  assign n4787 = ( ~n1789 & n2863 ) | ( ~n1789 & n4786 ) | ( n2863 & n4786 ) ;
  assign n4788 = n1790 | n4787 ;
  buffer buf_n4789( .i (n4788), .o (n4789) );
  buffer buf_n4790( .i (n4789), .o (n4790) );
  assign n4791 = n2800 | n3641 ;
  assign n4792 = ( ~n1753 & n3765 ) | ( ~n1753 & n4791 ) | ( n3765 & n4791 ) ;
  assign n4793 = n1754 | n4792 ;
  assign n4794 = n3741 | n4793 ;
  assign n4795 = ( n2505 & ~n3750 ) | ( n2505 & n4794 ) | ( ~n3750 & n4794 ) ;
  assign n4796 = n3751 | n4795 ;
  assign n4797 = ( n765 & n1539 ) | ( n765 & ~n4739 ) | ( n1539 & ~n4739 ) ;
  assign n4798 = n4740 & n4797 ;
  buffer buf_n4799( .i (n4798), .o (n4799) );
  buffer buf_n4800( .i (n4799), .o (n4800) );
  buffer buf_n4801( .i (n4800), .o (n4801) );
  assign n4807 = ( n669 & n3426 ) | ( n669 & n3439 ) | ( n3426 & n3439 ) ;
  buffer buf_n4808( .i (n3941), .o (n4808) );
  assign n4809 = ~n4807 & n4808 ;
  buffer buf_n4810( .i (n4808), .o (n4810) );
  assign n4811 = ( n3428 & ~n4809 ) | ( n3428 & n4810 ) | ( ~n4809 & n4810 ) ;
  assign n4812 = n3446 | n4811 ;
  assign n4813 = n4801 | n4812 ;
  assign n4814 = n4050 | n4813 ;
  assign n4815 = ( n2791 & ~n3847 ) | ( n2791 & n4814 ) | ( ~n3847 & n4814 ) ;
  assign n4816 = n3848 | n4815 ;
  buffer buf_n4087( .i (n4086), .o (n4087) );
  buffer buf_n4088( .i (n4087), .o (n4088) );
  buffer buf_n4089( .i (n4088), .o (n4089) );
  buffer buf_n4090( .i (n4089), .o (n4090) );
  buffer buf_n4091( .i (n4090), .o (n4091) );
  buffer buf_n4092( .i (n4091), .o (n4092) );
  buffer buf_n4102( .i (n4101), .o (n4102) );
  buffer buf_n4103( .i (n4102), .o (n4103) );
  buffer buf_n4104( .i (n4103), .o (n4104) );
  buffer buf_n4105( .i (n4104), .o (n4105) );
  assign n4817 = n4063 | n4288 ;
  buffer buf_n4818( .i (n4817), .o (n4818) );
  assign n4829 = n3658 | n4308 ;
  assign n4830 = n4818 | n4829 ;
  assign n4831 = n4105 | n4830 ;
  assign n4832 = ( n2827 & ~n4091 ) | ( n2827 & n4831 ) | ( ~n4091 & n4831 ) ;
  assign n4833 = n4092 | n4832 ;
  assign n4834 = n4816 | n4833 ;
  assign n4835 = ( ~n4789 & n4796 ) | ( ~n4789 & n4834 ) | ( n4796 & n4834 ) ;
  assign n4836 = n4790 | n4835 ;
  assign n4837 = n4783 | n4836 ;
  assign n4838 = ( ~n4628 & n4737 ) | ( ~n4628 & n4837 ) | ( n4737 & n4837 ) ;
  assign n4839 = n4629 | n4838 ;
  assign n4840 = n3034 | n4012 ;
  assign n4841 = n4050 | n4840 ;
  buffer buf_n4842( .i (n4841), .o (n4842) );
  buffer buf_n4843( .i (n4842), .o (n4843) );
  buffer buf_n4844( .i (n4843), .o (n4844) );
  buffer buf_n4845( .i (n4844), .o (n4845) );
  buffer buf_n4846( .i (n4845), .o (n4846) );
  buffer buf_n4847( .i (n4846), .o (n4847) );
  buffer buf_n4848( .i (n4847), .o (n4848) );
  buffer buf_n4849( .i (n4848), .o (n4849) );
  buffer buf_n4293( .i (n4292), .o (n4293) );
  buffer buf_n4294( .i (n4293), .o (n4294) );
  buffer buf_n4295( .i (n4294), .o (n4295) );
  buffer buf_n4296( .i (n4295), .o (n4296) );
  buffer buf_n4297( .i (n4296), .o (n4297) );
  buffer buf_n4298( .i (n4297), .o (n4298) );
  buffer buf_n4299( .i (n4298), .o (n4299) );
  buffer buf_n4300( .i (n4299), .o (n4300) );
  buffer buf_n4259( .i (n4258), .o (n4259) );
  buffer buf_n4260( .i (n4259), .o (n4260) );
  buffer buf_n4261( .i (n4260), .o (n4261) );
  buffer buf_n4262( .i (n4261), .o (n4262) );
  buffer buf_n4263( .i (n4262), .o (n4263) );
  buffer buf_n4264( .i (n4263), .o (n4264) );
  buffer buf_n4265( .i (n4264), .o (n4265) );
  buffer buf_n4266( .i (n4265), .o (n4266) );
  buffer buf_n4747( .i (n4746), .o (n4747) );
  assign n4850 = n3540 | n3899 ;
  assign n4851 = n3791 | n4850 ;
  assign n4852 = n3490 | n4851 ;
  assign n4853 = ( ~n3524 & n4747 ) | ( ~n3524 & n4852 ) | ( n4747 & n4852 ) ;
  assign n4854 = n3525 | n4853 ;
  buffer buf_n4464( .i (n4463), .o (n4464) );
  buffer buf_n4465( .i (n4464), .o (n4465) );
  buffer buf_n4855( .i (n4025), .o (n4855) );
  assign n4856 = ( ~n4172 & n4465 ) | ( ~n4172 & n4855 ) | ( n4465 & n4855 ) ;
  buffer buf_n4857( .i (n4855), .o (n4857) );
  assign n4858 = n4856 & ~n4857 ;
  buffer buf_n4859( .i (n4303), .o (n4859) );
  assign n4860 = n4858 & n4859 ;
  assign n4861 = n669 & n4860 ;
  buffer buf_n4862( .i (n4861), .o (n4862) );
  assign n4866 = n4472 | n4862 ;
  buffer buf_n4867( .i (n4866), .o (n4867) );
  buffer buf_n4868( .i (n4867), .o (n4868) );
  buffer buf_n4869( .i (n4868), .o (n4869) );
  buffer buf_n4870( .i (n4869), .o (n4870) );
  buffer buf_n4871( .i (n4870), .o (n4871) );
  assign n4872 = n4780 | n4871 ;
  assign n4873 = ( ~n4265 & n4854 ) | ( ~n4265 & n4872 ) | ( n4854 & n4872 ) ;
  assign n4874 = n4266 | n4873 ;
  buffer buf_n4875( .i (n4874), .o (n4875) );
  buffer buf_n4876( .i (n4875), .o (n4876) );
  buffer buf_n3754( .i (n3753), .o (n3754) );
  buffer buf_n3647( .i (n3646), .o (n3647) );
  buffer buf_n3648( .i (n3647), .o (n3648) );
  buffer buf_n3769( .i (n3768), .o (n3769) );
  buffer buf_n3770( .i (n3769), .o (n3770) );
  buffer buf_n4819( .i (n4818), .o (n4819) );
  buffer buf_n4820( .i (n4819), .o (n4820) );
  buffer buf_n4821( .i (n4820), .o (n4821) );
  buffer buf_n4822( .i (n4821), .o (n4822) );
  buffer buf_n3661( .i (n3660), .o (n3661) );
  buffer buf_n3662( .i (n3661), .o (n3662) );
  assign n4877 = ( n2812 & n3051 ) | ( n2812 & n4321 ) | ( n3051 & n4321 ) ;
  assign n4878 = ~n4322 & n4877 ;
  buffer buf_n4879( .i (n4878), .o (n4879) );
  buffer buf_n4880( .i (n4879), .o (n4880) );
  buffer buf_n4881( .i (n4880), .o (n4881) );
  buffer buf_n4882( .i (n4881), .o (n4882) );
  buffer buf_n4883( .i (n4882), .o (n4883) );
  buffer buf_n4884( .i (n4883), .o (n4884) );
  buffer buf_n4885( .i (n4884), .o (n4885) );
  buffer buf_n4886( .i (n4885), .o (n4886) );
  assign n4887 = n3662 | n4886 ;
  assign n4888 = n4822 | n4887 ;
  assign n4889 = n3770 | n4888 ;
  assign n4890 = ( n3648 & ~n3753 ) | ( n3648 & n4889 ) | ( ~n3753 & n4889 ) ;
  assign n4891 = n3754 | n4890 ;
  buffer buf_n4657( .i (n4656), .o (n4657) );
  buffer buf_n4658( .i (n4657), .o (n4658) );
  buffer buf_n4659( .i (n4658), .o (n4659) );
  buffer buf_n4660( .i (n4659), .o (n4660) );
  buffer buf_n4661( .i (n4660), .o (n4661) );
  buffer buf_n4802( .i (n4801), .o (n4802) );
  buffer buf_n4803( .i (n4802), .o (n4803) );
  buffer buf_n4804( .i (n4803), .o (n4804) );
  buffer buf_n4805( .i (n4804), .o (n4805) );
  buffer buf_n4806( .i (n4805), .o (n4806) );
  buffer buf_n3671( .i (n3670), .o (n3671) );
  buffer buf_n3672( .i (n3671), .o (n3672) );
  buffer buf_n3673( .i (n3672), .o (n3673) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n3464( .i (n3463), .o (n3464) );
  buffer buf_n3465( .i (n3464), .o (n3465) );
  buffer buf_n3466( .i (n3465), .o (n3466) );
  buffer buf_n3467( .i (n3466), .o (n3467) );
  assign n4892 = n673 & n3467 ;
  buffer buf_n4893( .i (n4892), .o (n4893) );
  buffer buf_n4894( .i (n4893), .o (n4894) );
  buffer buf_n4895( .i (n4894), .o (n4895) );
  assign n4896 = n3673 | n4895 ;
  assign n4897 = ( ~n4660 & n4806 ) | ( ~n4660 & n4896 ) | ( n4806 & n4896 ) ;
  assign n4898 = n4661 | n4897 ;
  buffer buf_n4677( .i (n4676), .o (n4677) );
  buffer buf_n4678( .i (n4677), .o (n4678) );
  buffer buf_n4679( .i (n4678), .o (n4679) );
  buffer buf_n4680( .i (n4679), .o (n4680) );
  buffer buf_n4681( .i (n4680), .o (n4681) );
  buffer buf_n4682( .i (n4681), .o (n4682) );
  buffer buf_n4683( .i (n4682), .o (n4683) );
  buffer buf_n3700( .i (n3699), .o (n3700) );
  buffer buf_n3701( .i (n3700), .o (n3701) );
  buffer buf_n3702( .i (n3701), .o (n3702) );
  buffer buf_n3703( .i (n3702), .o (n3703) );
  buffer buf_n3704( .i (n3703), .o (n3704) );
  buffer buf_n3705( .i (n3704), .o (n3705) );
  buffer buf_n3706( .i (n3705), .o (n3706) );
  buffer buf_n3707( .i (n3706), .o (n3707) );
  buffer buf_n3708( .i (n3707), .o (n3708) );
  buffer buf_n4709( .i (n4708), .o (n4709) );
  buffer buf_n4720( .i (n4719), .o (n4720) );
  buffer buf_n4721( .i (n4720), .o (n4721) );
  buffer buf_n4722( .i (n4721), .o (n4722) );
  assign n4899 = n4709 | n4722 ;
  assign n4900 = ( n3708 & ~n4682 ) | ( n3708 & n4899 ) | ( ~n4682 & n4899 ) ;
  assign n4901 = n4683 | n4900 ;
  assign n4902 = n4898 | n4901 ;
  assign n4903 = ( ~n4875 & n4891 ) | ( ~n4875 & n4902 ) | ( n4891 & n4902 ) ;
  assign n4904 = n4876 | n4903 ;
  assign n4905 = n3656 | n3666 ;
  assign n4906 = ( ~n3745 & n3788 ) | ( ~n3745 & n4905 ) | ( n3788 & n4905 ) ;
  assign n4907 = n3746 | n4906 ;
  buffer buf_n4908( .i (n4907), .o (n4908) );
  buffer buf_n4909( .i (n4908), .o (n4909) );
  buffer buf_n4910( .i (n4909), .o (n4910) );
  buffer buf_n4911( .i (n4910), .o (n4911) );
  buffer buf_n4912( .i (n4911), .o (n4912) );
  buffer buf_n4913( .i (n4912), .o (n4913) );
  buffer buf_n4914( .i (n4913), .o (n4914) );
  buffer buf_n4915( .i (n4914), .o (n4915) );
  buffer buf_n4916( .i (n4915), .o (n4916) );
  buffer buf_n4917( .i (n4916), .o (n4917) );
  assign n4918 = n4124 | n4276 ;
  assign n4919 = ( ~n1789 & n4040 ) | ( ~n1789 & n4918 ) | ( n4040 & n4918 ) ;
  assign n4920 = n1790 | n4919 ;
  buffer buf_n3995( .i (n3994), .o (n3995) );
  assign n4921 = n3995 | n4181 ;
  assign n4922 = n4150 | n4921 ;
  assign n4923 = n3979 | n4922 ;
  assign n4924 = ( ~n1641 & n4920 ) | ( ~n1641 & n4923 ) | ( n4920 & n4923 ) ;
  assign n4925 = n1642 | n4924 ;
  buffer buf_n4926( .i (n4925), .o (n4926) );
  buffer buf_n4927( .i (n4926), .o (n4927) );
  buffer buf_n4928( .i (n4927), .o (n4928) );
  buffer buf_n4929( .i (n4928), .o (n4929) );
  buffer buf_n3064( .i (n3063), .o (n3064) );
  buffer buf_n3065( .i (n3064), .o (n3065) );
  buffer buf_n3066( .i (n3065), .o (n3066) );
  buffer buf_n3067( .i (n3066), .o (n3067) );
  buffer buf_n4725( .i (n4724), .o (n4725) );
  buffer buf_n4726( .i (n4725), .o (n4726) );
  buffer buf_n4727( .i (n4726), .o (n4727) );
  buffer buf_n4728( .i (n4727), .o (n4728) );
  buffer buf_n4710( .i (n4709), .o (n4710) );
  buffer buf_n3275( .i (n3274), .o (n3275) );
  buffer buf_n3276( .i (n3275), .o (n3276) );
  assign n4930 = n3266 | n3276 ;
  assign n4931 = n4710 | n4930 ;
  buffer buf_n464( .i (x16), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n259( .i (x7), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  assign n4932 = ( n277 & n482 ) | ( n277 & n1324 ) | ( n482 & n1324 ) ;
  assign n4933 = ~n483 & n4932 ;
  buffer buf_n4934( .i (n4933), .o (n4934) );
  buffer buf_n4935( .i (n4934), .o (n4935) );
  assign n4936 = ( n1968 & n4169 ) | ( n1968 & ~n4934 ) | ( n4169 & ~n4934 ) ;
  assign n4937 = n4935 & n4936 ;
  assign n4938 = ( n3148 & n4322 ) | ( n3148 & n4937 ) | ( n4322 & n4937 ) ;
  buffer buf_n4939( .i (n4322), .o (n4939) );
  assign n4940 = n4938 & ~n4939 ;
  buffer buf_n4941( .i (n4940), .o (n4941) );
  buffer buf_n4942( .i (n4941), .o (n4942) );
  buffer buf_n4943( .i (n4942), .o (n4943) );
  buffer buf_n4944( .i (n4943), .o (n4944) );
  buffer buf_n4945( .i (n4944), .o (n4945) );
  buffer buf_n4946( .i (n4945), .o (n4946) );
  buffer buf_n4947( .i (n4946), .o (n4947) );
  buffer buf_n4948( .i (n4947), .o (n4948) );
  buffer buf_n4949( .i (n4948), .o (n4949) );
  buffer buf_n3150( .i (n3149), .o (n3150) );
  buffer buf_n281( .i (x8), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  assign n4950 = n483 & n4070 ;
  assign n4951 = ( n301 & n4074 ) | ( n301 & n4950 ) | ( n4074 & n4950 ) ;
  assign n4952 = ~n4075 & n4951 ;
  buffer buf_n4953( .i (n4952), .o (n4953) );
  buffer buf_n4954( .i (n4953), .o (n4954) );
  assign n4955 = ( n1970 & n3988 ) | ( n1970 & ~n4953 ) | ( n3988 & ~n4953 ) ;
  assign n4956 = n4954 & n4955 ;
  assign n4957 = ( n3150 & n4371 ) | ( n3150 & n4956 ) | ( n4371 & n4956 ) ;
  assign n4958 = ~n3485 & n4957 ;
  buffer buf_n4959( .i (n4958), .o (n4959) );
  buffer buf_n4960( .i (n4959), .o (n4960) );
  buffer buf_n4961( .i (n4960), .o (n4961) );
  buffer buf_n4962( .i (n4961), .o (n4962) );
  buffer buf_n4963( .i (n4962), .o (n4963) );
  buffer buf_n4964( .i (n4963), .o (n4964) );
  buffer buf_n3250( .i (n3249), .o (n3250) );
  buffer buf_n3207( .i (n3206), .o (n3207) );
  buffer buf_n3208( .i (n3207), .o (n3208) );
  buffer buf_n4164( .i (n4163), .o (n4164) );
  buffer buf_n4165( .i (n4164), .o (n4165) );
  buffer buf_n4166( .i (n4165), .o (n4166) );
  buffer buf_n4167( .i (n4166), .o (n4167) );
  buffer buf_n4965( .i (n3988), .o (n4965) );
  assign n4966 = n4167 & n4965 ;
  buffer buf_n4967( .i (n668), .o (n4967) );
  assign n4968 = ( n4119 & n4966 ) | ( n4119 & n4967 ) | ( n4966 & n4967 ) ;
  assign n4969 = ~n2822 & n4968 ;
  assign n4970 = n1351 & n4969 ;
  buffer buf_n4971( .i (n4970), .o (n4971) );
  buffer buf_n4972( .i (n4971), .o (n4972) );
  buffer buf_n4973( .i (n4972), .o (n4973) );
  assign n4974 = n3208 | n4973 ;
  assign n4975 = n3250 | n4974 ;
  assign n4976 = n4964 | n4975 ;
  assign n4977 = n4949 | n4976 ;
  assign n4978 = n4931 | n4977 ;
  assign n4979 = ( ~n3066 & n4728 ) | ( ~n3066 & n4978 ) | ( n4728 & n4978 ) ;
  assign n4980 = n3067 | n4979 ;
  buffer buf_n3883( .i (n3882), .o (n3883) );
  buffer buf_n3884( .i (n3883), .o (n3884) );
  buffer buf_n3885( .i (n3884), .o (n3885) );
  buffer buf_n3886( .i (n3885), .o (n3886) );
  buffer buf_n3887( .i (n3886), .o (n3887) );
  buffer buf_n4514( .i (n4513), .o (n4514) );
  buffer buf_n4515( .i (n4514), .o (n4515) );
  buffer buf_n4516( .i (n4515), .o (n4516) );
  buffer buf_n3957( .i (n3956), .o (n3957) );
  assign n4981 = n3344 | n3957 ;
  assign n4982 = ( n3887 & ~n4516 ) | ( n3887 & n4981 ) | ( ~n4516 & n4981 ) ;
  buffer buf_n4983( .i (n4982), .o (n4983) );
  buffer buf_n4984( .i (n4983), .o (n4984) );
  assign n4985 = n3445 | n4799 ;
  assign n4986 = n3429 | n4985 ;
  buffer buf_n4987( .i (n4986), .o (n4987) );
  buffer buf_n4988( .i (n4987), .o (n4988) );
  buffer buf_n4989( .i (n4988), .o (n4989) );
  buffer buf_n4990( .i (n4989), .o (n4990) );
  assign n4991 = n3474 | n4893 ;
  buffer buf_n4863( .i (n4862), .o (n4863) );
  buffer buf_n4864( .i (n4863), .o (n4864) );
  buffer buf_n4865( .i (n4864), .o (n4865) );
  assign n4992 = n4305 | n4879 ;
  buffer buf_n4993( .i (n4992), .o (n4993) );
  buffer buf_n4994( .i (n4993), .o (n4994) );
  buffer buf_n4995( .i (n4994), .o (n4995) );
  assign n4996 = n4776 | n4995 ;
  assign n4997 = ( ~n4475 & n4865 ) | ( ~n4475 & n4996 ) | ( n4865 & n4996 ) ;
  assign n4998 = n4476 | n4997 ;
  assign n4999 = n4991 | n4998 ;
  assign n5000 = ( ~n4294 & n4990 ) | ( ~n4294 & n4999 ) | ( n4990 & n4999 ) ;
  assign n5001 = n4295 | n5000 ;
  buffer buf_n4519( .i (n4518), .o (n4519) );
  buffer buf_n4520( .i (n4519), .o (n4520) );
  assign n5002 = n3919 | n3924 ;
  buffer buf_n5003( .i (n5002), .o (n5003) );
  buffer buf_n5004( .i (n5003), .o (n5004) );
  buffer buf_n5005( .i (n5004), .o (n5005) );
  buffer buf_n5006( .i (n5005), .o (n5006) );
  buffer buf_n5007( .i (n5006), .o (n5007) );
  assign n5008 = n4520 | n5007 ;
  assign n5009 = ( ~n4983 & n5001 ) | ( ~n4983 & n5008 ) | ( n5001 & n5008 ) ;
  assign n5010 = n4984 | n5009 ;
  buffer buf_n4662( .i (n4661), .o (n4662) );
  buffer buf_n225( .i (n224), .o (n225) );
  assign n5011 = ( n225 & n1802 ) | ( n225 & n4855 ) | ( n1802 & n4855 ) ;
  assign n5012 = ~n4857 & n5011 ;
  buffer buf_n5013( .i (n4169), .o (n5013) );
  buffer buf_n5014( .i (n5013), .o (n5014) );
  assign n5015 = ~n4031 & n5014 ;
  buffer buf_n5016( .i (n764), .o (n5016) );
  assign n5017 = ( n5012 & n5015 ) | ( n5012 & n5016 ) | ( n5015 & n5016 ) ;
  assign n5018 = ~n766 & n5017 ;
  assign n5019 = n1350 & n5018 ;
  buffer buf_n5020( .i (n5019), .o (n5020) );
  buffer buf_n5021( .i (n5020), .o (n5021) );
  buffer buf_n5022( .i (n5021), .o (n5022) );
  buffer buf_n5023( .i (n5022), .o (n5023) );
  buffer buf_n5024( .i (n5023), .o (n5024) );
  buffer buf_n5025( .i (n5024), .o (n5025) );
  buffer buf_n5026( .i (n5025), .o (n5026) );
  buffer buf_n4379( .i (n4378), .o (n4379) );
  assign n5027 = n221 & n338 ;
  assign n5028 = ( n4070 & n4073 ) | ( n4070 & n5027 ) | ( n4073 & n5027 ) ;
  assign n5029 = ~n4645 & n5028 ;
  buffer buf_n5030( .i (n5029), .o (n5030) );
  buffer buf_n5031( .i (n5030), .o (n5031) );
  assign n5032 = ( n1858 & n5013 ) | ( n1858 & ~n5030 ) | ( n5013 & ~n5030 ) ;
  assign n5033 = n5031 & n5032 ;
  assign n5034 = ( n4671 & n4672 ) | ( n4671 & n5033 ) | ( n4672 & n5033 ) ;
  assign n5035 = ~n4119 & n5034 ;
  buffer buf_n5036( .i (n5035), .o (n5036) );
  buffer buf_n5037( .i (n5036), .o (n5037) );
  buffer buf_n5038( .i (n5037), .o (n5038) );
  buffer buf_n5039( .i (n5038), .o (n5039) );
  buffer buf_n5040( .i (n5039), .o (n5040) );
  buffer buf_n5041( .i (n5040), .o (n5041) );
  buffer buf_n5042( .i (n5041), .o (n5042) );
  assign n5043 = n4379 | n5042 ;
  assign n5044 = n5026 | n5043 ;
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n5045( .i (n4645), .o (n5045) );
  assign n5046 = n280 & ~n5045 ;
  assign n5047 = ( n486 & n2174 ) | ( n486 & n5046 ) | ( n2174 & n5046 ) ;
  assign n5048 = ~n487 & n5047 ;
  buffer buf_n5049( .i (n5048), .o (n5049) );
  buffer buf_n5050( .i (n5049), .o (n5050) );
  buffer buf_n4079( .i (n4078), .o (n4079) );
  buffer buf_n4080( .i (n4079), .o (n4080) );
  buffer buf_n4081( .i (n4080), .o (n4081) );
  assign n5051 = ( n3972 & n4081 ) | ( n3972 & ~n5049 ) | ( n4081 & ~n5049 ) ;
  assign n5052 = n5050 & n5051 ;
  buffer buf_n5053( .i (n5052), .o (n5053) );
  buffer buf_n5054( .i (n5053), .o (n5054) );
  buffer buf_n5055( .i (n5054), .o (n5055) );
  buffer buf_n5056( .i (n5055), .o (n5056) );
  buffer buf_n5057( .i (n5056), .o (n5057) );
  assign n5058 = n301 & n484 ;
  assign n5059 = ( n4075 & n5045 ) | ( n4075 & n5058 ) | ( n5045 & n5058 ) ;
  assign n5060 = ~n4855 & n5059 ;
  buffer buf_n5061( .i (n5060), .o (n5061) );
  buffer buf_n5062( .i (n5061), .o (n5062) );
  assign n5063 = ( n4080 & n4965 ) | ( n4080 & ~n5061 ) | ( n4965 & ~n5061 ) ;
  assign n5064 = n5062 & n5063 ;
  buffer buf_n5065( .i (n5064), .o (n5065) );
  buffer buf_n5066( .i (n5065), .o (n5066) );
  buffer buf_n5067( .i (n5066), .o (n5067) );
  buffer buf_n5068( .i (n5067), .o (n5068) );
  buffer buf_n5069( .i (n5068), .o (n5069) );
  assign n5070 = n4393 | n5069 ;
  assign n5071 = ( ~n3363 & n5057 ) | ( ~n3363 & n5070 ) | ( n5057 & n5070 ) ;
  assign n5072 = n3364 | n5071 ;
  assign n5073 = n4682 | n5072 ;
  assign n5074 = ( ~n4661 & n5044 ) | ( ~n4661 & n5073 ) | ( n5044 & n5073 ) ;
  assign n5075 = n4662 | n5074 ;
  assign n5076 = n5010 | n5075 ;
  assign n5077 = n4980 | n5076 ;
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  buffer buf_n2129( .i (n2128), .o (n2129) );
  buffer buf_n2130( .i (n2129), .o (n2130) );
  assign n5078 = n1666 | n1703 ;
  assign n5079 = n1639 | n5078 ;
  assign n5080 = n2130 | n5079 ;
  assign n5081 = ( n1757 & ~n2109 ) | ( n1757 & n5080 ) | ( ~n2109 & n5080 ) ;
  assign n5082 = n2110 | n5081 ;
  assign n5083 = n1955 | n2045 ;
  buffer buf_n5084( .i (n5083), .o (n5084) );
  assign n5085 = n2032 | n5084 ;
  assign n5086 = ( ~n1521 & n1927 ) | ( ~n1521 & n5085 ) | ( n1927 & n5085 ) ;
  assign n5087 = n1522 | n5086 ;
  assign n5088 = n1582 | n1976 ;
  assign n5089 = n1568 | n5088 ;
  assign n5090 = n2017 | n5089 ;
  assign n5091 = ( ~n1869 & n5087 ) | ( ~n1869 & n5090 ) | ( n5087 & n5090 ) ;
  assign n5092 = n1870 | n5091 ;
  buffer buf_n1821( .i (n1820), .o (n1821) );
  buffer buf_n1822( .i (n1821), .o (n1822) );
  buffer buf_n1823( .i (n1822), .o (n1823) );
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  assign n5093 = n1787 | n1885 ;
  assign n5094 = n1767 | n5093 ;
  assign n5095 = n1842 | n5094 ;
  assign n5096 = ( n1548 & ~n1823 ) | ( n1548 & n5095 ) | ( ~n1823 & n5095 ) ;
  assign n5097 = n1824 | n5096 ;
  assign n5098 = n5092 | n5097 ;
  assign n5099 = n5082 | n5098 ;
  buffer buf_n5100( .i (n5099), .o (n5100) );
  buffer buf_n5101( .i (n5100), .o (n5101) );
  buffer buf_n5102( .i (n5101), .o (n5102) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n2143( .i (n2142), .o (n2143) );
  buffer buf_n2144( .i (n2143), .o (n2144) );
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  assign n5103 = n2072 | n2092 ;
  assign n5104 = n2148 | n5103 ;
  assign n5105 = n1621 | n2171 ;
  buffer buf_n5106( .i (n5105), .o (n5106) );
  assign n5107 = n1685 | n5106 ;
  assign n5108 = n5104 | n5107 ;
  buffer buf_n5109( .i (n5108), .o (n5109) );
  buffer buf_n5110( .i (n5109), .o (n5110) );
  buffer buf_n5111( .i (n5110), .o (n5111) );
  buffer buf_n5112( .i (n5111), .o (n5112) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  buffer buf_n2197( .i (n2196), .o (n2197) );
  buffer buf_n2198( .i (n2197), .o (n2198) );
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n2184( .i (n2183), .o (n2184) );
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  assign n5113 = n2092 | n2186 ;
  assign n5114 = n2199 | n5113 ;
  buffer buf_n5115( .i (n1684), .o (n5115) );
  assign n5116 = n1735 | n5115 ;
  assign n5117 = n5114 | n5116 ;
  buffer buf_n5118( .i (n5117), .o (n5118) );
  buffer buf_n5119( .i (n5118), .o (n5119) );
  buffer buf_n5120( .i (n5119), .o (n5120) );
  buffer buf_n5121( .i (n5120), .o (n5121) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n370( .i (x12), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n5122( .i (n2808), .o (n5122) );
  assign n5123 = ~n411 & n5122 ;
  assign n5124 = ( n390 & ~n434 ) | ( n390 & n5123 ) | ( ~n434 & n5123 ) ;
  assign n5125 = ~n391 & n5124 ;
  assign n5126 = ~n4030 & n5125 ;
  buffer buf_n5127( .i (n3125), .o (n5127) );
  buffer buf_n5128( .i (n4321), .o (n5128) );
  assign n5129 = ( n5126 & n5127 ) | ( n5126 & ~n5128 ) | ( n5127 & ~n5128 ) ;
  assign n5130 = ~n828 & n5129 ;
  buffer buf_n5131( .i (n4859), .o (n5131) );
  assign n5132 = n5130 & ~n5131 ;
  buffer buf_n5133( .i (n5132), .o (n5133) );
  buffer buf_n5134( .i (n5133), .o (n5134) );
  buffer buf_n5135( .i (n5134), .o (n5135) );
  buffer buf_n5136( .i (n5135), .o (n5136) );
  buffer buf_n5137( .i (n5136), .o (n5137) );
  buffer buf_n5138( .i (n5137), .o (n5138) );
  buffer buf_n5139( .i (n5138), .o (n5139) );
  buffer buf_n5140( .i (n5139), .o (n5140) );
  buffer buf_n5141( .i (n5140), .o (n5141) );
  buffer buf_n5142( .i (n5141), .o (n5142) );
  buffer buf_n5143( .i (n5142), .o (n5143) );
  buffer buf_n5144( .i (n5143), .o (n5144) );
  buffer buf_n5145( .i (n5144), .o (n5145) );
  buffer buf_n3996( .i (n3995), .o (n3996) );
  assign n5146 = n3962 | n3977 ;
  assign n5147 = ( ~n2593 & n3996 ) | ( ~n2593 & n5146 ) | ( n3996 & n5146 ) ;
  assign n5148 = n2594 | n5147 ;
  buffer buf_n5149( .i (n5148), .o (n5149) );
  buffer buf_n5150( .i (n5149), .o (n5150) );
  buffer buf_n5151( .i (n5150), .o (n5151) );
  buffer buf_n5152( .i (n5151), .o (n5152) );
  buffer buf_n5153( .i (n5152), .o (n5153) );
  buffer buf_n5154( .i (n5153), .o (n5154) );
  buffer buf_n2348( .i (n2347), .o (n2348) );
  buffer buf_n2349( .i (n2348), .o (n2349) );
  buffer buf_n2350( .i (n2349), .o (n2350) );
  buffer buf_n2351( .i (n2350), .o (n2351) );
  assign n5155 = n2351 | n2546 ;
  assign n5156 = n2525 | n5155 ;
  assign n5157 = n2330 | n3816 ;
  assign n5158 = n3118 | n5157 ;
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  buffer buf_n2563( .i (n2562), .o (n2563) );
  buffer buf_n2564( .i (n2563), .o (n2564) );
  buffer buf_n5159( .i (n959), .o (n5159) );
  assign n5160 = n2559 & n5159 ;
  buffer buf_n5161( .i (n5160), .o (n5161) );
  buffer buf_n5162( .i (n5161), .o (n5162) );
  buffer buf_n5163( .i (n5162), .o (n5163) );
  buffer buf_n5164( .i (n5163), .o (n5164) );
  assign n5165 = ( ~n1025 & n2564 ) | ( ~n1025 & n5164 ) | ( n2564 & n5164 ) ;
  assign n5166 = n5158 | n5165 ;
  assign n5167 = n5156 | n5166 ;
  buffer buf_n5168( .i (n5167), .o (n5168) );
  buffer buf_n5169( .i (n5168), .o (n5169) );
  buffer buf_n3382( .i (n3381), .o (n3382) );
  buffer buf_n3383( .i (n3382), .o (n3383) );
  buffer buf_n3384( .i (n3383), .o (n3384) );
  buffer buf_n3385( .i (n3384), .o (n3385) );
  buffer buf_n3386( .i (n3385), .o (n3386) );
  buffer buf_n3387( .i (n3386), .o (n3387) );
  buffer buf_n3201( .i (n3200), .o (n3201) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n1585( .i (n1584), .o (n1585) );
  assign n5170 = n1439 | n1476 ;
  assign n5171 = n2935 | n5170 ;
  buffer buf_n5172( .i (n5171), .o (n5172) );
  assign n5173 = ( n1585 & ~n3200 ) | ( n1585 & n5172 ) | ( ~n3200 & n5172 ) ;
  assign n5174 = n3201 | n5173 ;
  buffer buf_n4632( .i (n4631), .o (n4632) );
  buffer buf_n4633( .i (n4632), .o (n4633) );
  buffer buf_n4634( .i (n4633), .o (n4634) );
  buffer buf_n4635( .i (n4634), .o (n4635) );
  buffer buf_n4636( .i (n4635), .o (n4636) );
  buffer buf_n4637( .i (n4636), .o (n4637) );
  buffer buf_n3367( .i (n3366), .o (n3367) );
  buffer buf_n3368( .i (n3367), .o (n3368) );
  buffer buf_n3369( .i (n3368), .o (n3369) );
  buffer buf_n3370( .i (n3369), .o (n3370) );
  assign n5175 = n2863 | n3847 ;
  assign n5176 = n3370 | n5175 ;
  assign n5177 = n4637 | n5176 ;
  assign n5178 = ( ~n3386 & n5174 ) | ( ~n3386 & n5177 ) | ( n5174 & n5177 ) ;
  assign n5179 = n3387 | n5178 ;
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  assign n5180 = n2185 | n3160 ;
  assign n5181 = n2198 | n5180 ;
  buffer buf_n3181( .i (n3180), .o (n3181) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  assign n5182 = n2630 & n4810 ;
  buffer buf_n5183( .i (n5182), .o (n5183) );
  buffer buf_n5184( .i (n5183), .o (n5184) );
  assign n5185 = n1663 | n2632 ;
  assign n5186 = n1729 | n5185 ;
  assign n5187 = n1681 | n5186 ;
  assign n5188 = ( ~n3825 & n5184 ) | ( ~n3825 & n5187 ) | ( n5184 & n5187 ) ;
  assign n5189 = n3826 | n5188 ;
  assign n5190 = n3181 | n5189 ;
  assign n5191 = ( ~n1720 & n5181 ) | ( ~n1720 & n5190 ) | ( n5181 & n5190 ) ;
  assign n5192 = n1721 | n5191 ;
  buffer buf_n2815( .i (n2814), .o (n2815) );
  buffer buf_n2816( .i (n2815), .o (n2816) );
  buffer buf_n2817( .i (n2816), .o (n2817) );
  buffer buf_n2818( .i (n2817), .o (n2818) );
  buffer buf_n3151( .i (n3150), .o (n3151) );
  buffer buf_n3152( .i (n3151), .o (n3152) );
  buffer buf_n3153( .i (n3152), .o (n3153) );
  assign n5193 = ( n893 & n2818 ) | ( n893 & n3153 ) | ( n2818 & n3153 ) ;
  assign n5194 = ~n894 & n5193 ;
  buffer buf_n5195( .i (n5194), .o (n5195) );
  buffer buf_n2853( .i (n2852), .o (n2853) );
  assign n5196 = ( ~n2853 & n3149 ) | ( ~n2853 & n4939 ) | ( n3149 & n4939 ) ;
  assign n5197 = ~n4371 & n5196 ;
  buffer buf_n5198( .i (n5197), .o (n5198) );
  assign n5199 = n1785 | n5198 ;
  buffer buf_n5200( .i (n5199), .o (n5200) );
  assign n5201 = n2825 | n5200 ;
  assign n5202 = n1754 | n5201 ;
  assign n5203 = ( ~n2462 & n5195 ) | ( ~n2462 & n5202 ) | ( n5195 & n5202 ) ;
  assign n5204 = n2463 | n5203 ;
  buffer buf_n2468( .i (n2467), .o (n2468) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  buffer buf_n2470( .i (n2469), .o (n2470) );
  buffer buf_n2471( .i (n2470), .o (n2471) );
  buffer buf_n5205( .i (n4939), .o (n5205) );
  assign n5206 = n2471 & ~n5205 ;
  assign n5207 = ~n4808 & n5206 ;
  buffer buf_n5208( .i (n5207), .o (n5208) );
  buffer buf_n5209( .i (n5208), .o (n5209) );
  buffer buf_n5210( .i (n5209), .o (n5210) );
  assign n5212 = n3582 | n5210 ;
  assign n5213 = n2091 | n5212 ;
  assign n5214 = n3603 | n5213 ;
  assign n5215 = ( ~n2384 & n5204 ) | ( ~n2384 & n5214 ) | ( n5204 & n5214 ) ;
  assign n5216 = n2385 | n5215 ;
  assign n5217 = n5192 | n5216 ;
  assign n5218 = ( ~n5168 & n5179 ) | ( ~n5168 & n5217 ) | ( n5179 & n5217 ) ;
  assign n5219 = n5169 | n5218 ;
  buffer buf_n5220( .i (n5219), .o (n5220) );
  assign n5221 = n4136 | n4762 ;
  buffer buf_n5222( .i (n4134), .o (n5222) );
  assign n5223 = ( n251 & n5221 ) | ( n251 & ~n5222 ) | ( n5221 & ~n5222 ) ;
  assign n5224 = n136 | n5223 ;
  assign n5225 = n4694 | n5224 ;
  assign n5226 = ( n3634 & n5045 ) | ( n3634 & ~n5225 ) | ( n5045 & ~n5225 ) ;
  buffer buf_n5227( .i (n5045), .o (n5227) );
  assign n5228 = n5226 & ~n5227 ;
  assign n5229 = ( n1575 & n5128 ) | ( n1575 & n5228 ) | ( n5128 & n5228 ) ;
  assign n5230 = ~n4939 & n5229 ;
  buffer buf_n5231( .i (n5230), .o (n5231) );
  assign n5238 = n1750 | n5231 ;
  assign n5239 = n3640 | n5238 ;
  assign n5240 = n2474 | n3576 ;
  assign n5241 = ( n2085 & ~n2101 ) | ( n2085 & n5240 ) | ( ~n2101 & n5240 ) ;
  assign n5242 = n2102 | n5241 ;
  assign n5243 = n3763 | n5242 ;
  assign n5244 = ( ~n3746 & n5239 ) | ( ~n3746 & n5243 ) | ( n5239 & n5243 ) ;
  assign n5245 = n3747 | n5244 ;
  buffer buf_n5246( .i (n5245), .o (n5246) );
  buffer buf_n5247( .i (n5246), .o (n5247) );
  assign n5248 = n2150 | n3598 ;
  assign n5249 = ( ~n3509 & n3520 ) | ( ~n3509 & n5248 ) | ( n3520 & n5248 ) ;
  assign n5250 = n3510 | n5249 ;
  assign n5251 = n2068 | n3487 ;
  buffer buf_n5252( .i (n5251), .o (n5252) );
  assign n5255 = n5250 | n5252 ;
  assign n5256 = ( n2201 & ~n5246 ) | ( n2201 & n5255 ) | ( ~n5246 & n5255 ) ;
  assign n5257 = n5247 | n5256 ;
  buffer buf_n5258( .i (n5257), .o (n5258) );
  buffer buf_n5259( .i (n5258), .o (n5259) );
  assign n5260 = n1700 | n3538 ;
  buffer buf_n5261( .i (n5260), .o (n5261) );
  assign n5263 = n2169 | n5261 ;
  assign n5264 = ( ~n1620 & n3554 ) | ( ~n1620 & n5263 ) | ( n3554 & n5263 ) ;
  assign n5265 = n1621 | n5264 ;
  assign n5266 = n4338 | n5265 ;
  assign n5267 = n1735 | n5266 ;
  buffer buf_n2340( .i (n2339), .o (n2340) );
  buffer buf_n2341( .i (n2340), .o (n2341) );
  buffer buf_n2342( .i (n2341), .o (n2342) );
  assign n5268 = n2603 | n3900 ;
  assign n5269 = ( ~n2341 & n2614 ) | ( ~n2341 & n5268 ) | ( n2614 & n5268 ) ;
  assign n5270 = n2342 | n5269 ;
  assign n5271 = n3976 | n5183 ;
  assign n5272 = n3995 | n5271 ;
  assign n5273 = n1683 | n5272 ;
  assign n5274 = n3135 | n5273 ;
  assign n5275 = n5270 | n5274 ;
  assign n5276 = ( ~n5258 & n5267 ) | ( ~n5258 & n5275 ) | ( n5267 & n5275 ) ;
  assign n5277 = n5259 | n5276 ;
  buffer buf_n5278( .i (n5277), .o (n5278) );
  buffer buf_n5279( .i (n5278), .o (n5279) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  assign n5280 = n1904 | n3021 ;
  buffer buf_n5281( .i (n5280), .o (n5281) );
  buffer buf_n5282( .i (n5281), .o (n5282) );
  buffer buf_n5283( .i (n5282), .o (n5283) );
  assign n5284 = n1956 | n3097 ;
  assign n5285 = ( ~n1520 & n3034 ) | ( ~n1520 & n5284 ) | ( n3034 & n5284 ) ;
  assign n5286 = n1521 | n5285 ;
  assign n5287 = n2052 | n5286 ;
  assign n5288 = ( ~n1924 & n5283 ) | ( ~n1924 & n5287 ) | ( n5283 & n5287 ) ;
  assign n5289 = n1925 | n5288 ;
  buffer buf_n5290( .i (n5289), .o (n5290) );
  buffer buf_n5291( .i (n5290), .o (n5291) );
  assign n5292 = n2014 | n2970 ;
  buffer buf_n5293( .i (n5292), .o (n5293) );
  buffer buf_n5294( .i (n5293), .o (n5294) );
  buffer buf_n5295( .i (n5294), .o (n5295) );
  buffer buf_n5296( .i (n5295), .o (n5296) );
  buffer buf_n5297( .i (n5296), .o (n5297) );
  buffer buf_n5298( .i (n5297), .o (n5298) );
  buffer buf_n4550( .i (n4549), .o (n4550) );
  buffer buf_n4551( .i (n4550), .o (n4551) );
  buffer buf_n5299( .i (n2896), .o (n5299) );
  assign n5300 = n1976 | n5299 ;
  buffer buf_n5301( .i (n5300), .o (n5301) );
  assign n5302 = n2936 | n5301 ;
  assign n5303 = ( n1585 & ~n2995 ) | ( n1585 & n5302 ) | ( ~n2995 & n5302 ) ;
  assign n5304 = n2996 | n5303 ;
  assign n5305 = n4551 | n5304 ;
  assign n5306 = ( ~n5290 & n5298 ) | ( ~n5290 & n5305 ) | ( n5298 & n5305 ) ;
  assign n5307 = n5291 | n5306 ;
  buffer buf_n1846( .i (n1845), .o (n1846) );
  assign n5308 = n1547 | n4014 ;
  assign n5309 = ( ~n1823 & n4052 ) | ( ~n1823 & n5308 ) | ( n4052 & n5308 ) ;
  assign n5310 = n1824 | n5309 ;
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n2003), .o (n2004) );
  buffer buf_n2954( .i (n2953), .o (n2954) );
  buffer buf_n2955( .i (n2954), .o (n2955) );
  assign n5311 = n1868 | n2955 ;
  assign n5312 = n2004 | n5311 ;
  assign n5313 = n3303 | n5312 ;
  assign n5314 = ( ~n1845 & n5310 ) | ( ~n1845 & n5313 ) | ( n5310 & n5313 ) ;
  assign n5315 = n1846 | n5314 ;
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  buffer buf_n4444( .i (n4443), .o (n4444) );
  buffer buf_n4445( .i (n4444), .o (n4445) );
  buffer buf_n4446( .i (n4445), .o (n4446) );
  buffer buf_n4082( .i (n4081), .o (n4082) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n4022( .i (n4021), .o (n4022) );
  buffer buf_n4023( .i (n4022), .o (n4023) );
  buffer buf_n4024( .i (n4023), .o (n4024) );
  buffer buf_n5316( .i (n4857), .o (n5316) );
  assign n5317 = ( n257 & n4024 ) | ( n257 & ~n5316 ) | ( n4024 & ~n5316 ) ;
  assign n5318 = ~n258 & n5317 ;
  buffer buf_n5319( .i (n4965), .o (n5319) );
  buffer buf_n5320( .i (n5319), .o (n5320) );
  assign n5321 = ( n4082 & n5318 ) | ( n4082 & n5320 ) | ( n5318 & n5320 ) ;
  assign n5322 = ~n635 & n5321 ;
  assign n5323 = n1352 & n5322 ;
  buffer buf_n5324( .i (n5323), .o (n5324) );
  buffer buf_n5325( .i (n5324), .o (n5325) );
  buffer buf_n5326( .i (n5325), .o (n5326) );
  buffer buf_n5327( .i (n5326), .o (n5327) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n5328( .i (n4645), .o (n5328) );
  assign n5329 = n167 | n5328 ;
  assign n5330 = ( ~n139 & n2174 ) | ( ~n139 & n5329 ) | ( n2174 & n5329 ) ;
  assign n5331 = n140 | n5330 ;
  assign n5332 = n4033 | n5331 ;
  assign n5333 = n5319 | n5332 ;
  assign n5334 = ( n1578 & n3485 ) | ( n1578 & ~n5333 ) | ( n3485 & ~n5333 ) ;
  assign n5335 = ~n2181 & n5334 ;
  buffer buf_n5336( .i (n5335), .o (n5336) );
  buffer buf_n5337( .i (n5336), .o (n5337) );
  buffer buf_n5338( .i (n5337), .o (n5338) );
  assign n5339 = n1886 | n4571 ;
  buffer buf_n5340( .i (n1788), .o (n5340) );
  assign n5341 = ( n5338 & n5339 ) | ( n5338 & ~n5340 ) | ( n5339 & ~n5340 ) ;
  buffer buf_n5342( .i (n5340), .o (n5342) );
  assign n5343 = n5341 | n5342 ;
  assign n5344 = n5327 | n5343 ;
  assign n5345 = ( ~n1771 & n4446 ) | ( ~n1771 & n5344 ) | ( n4446 & n5344 ) ;
  assign n5346 = n1772 | n5345 ;
  assign n5347 = n5315 | n5346 ;
  assign n5348 = ( ~n5278 & n5307 ) | ( ~n5278 & n5347 ) | ( n5307 & n5347 ) ;
  assign n5349 = n5279 | n5348 ;
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n3177( .i (n3176), .o (n3177) );
  assign n5350 = n2637 | n4331 ;
  assign n5351 = n3177 | n5350 ;
  buffer buf_n3812( .i (n3811), .o (n3812) );
  buffer buf_n3813( .i (n3812), .o (n3813) );
  assign n5352 = n1636 | n3131 ;
  assign n5353 = n1681 | n5352 ;
  assign n5354 = n2340 | n5353 ;
  buffer buf_n5355( .i (n3825), .o (n5355) );
  assign n5356 = ( ~n3812 & n5354 ) | ( ~n3812 & n5355 ) | ( n5354 & n5355 ) ;
  assign n5357 = n3813 | n5356 ;
  assign n5358 = n5106 | n5357 ;
  assign n5359 = ( ~n1707 & n5351 ) | ( ~n1707 & n5358 ) | ( n5351 & n5358 ) ;
  assign n5360 = n1708 | n5359 ;
  buffer buf_n5361( .i (n5360), .o (n5361) );
  buffer buf_n5362( .i (n5361), .o (n5362) );
  buffer buf_n3089( .i (n3088), .o (n3089) );
  buffer buf_n3090( .i (n3089), .o (n3090) );
  buffer buf_n3091( .i (n3090), .o (n3091) );
  buffer buf_n3092( .i (n3091), .o (n3092) );
  buffer buf_n3093( .i (n3092), .o (n3093) );
  buffer buf_n3094( .i (n3093), .o (n3094) );
  buffer buf_n3047( .i (n3046), .o (n3047) );
  assign n5363 = ( n433 & ~n1874 ) | ( n433 & n4766 ) | ( ~n1874 & n4766 ) ;
  buffer buf_n5364( .i (n433), .o (n5364) );
  assign n5365 = n5363 & ~n5364 ;
  assign n5366 = ~n3984 & n5365 ;
  assign n5367 = ( ~n4030 & n5013 ) | ( ~n4030 & n5366 ) | ( n5013 & n5366 ) ;
  assign n5368 = ~n5014 & n5367 ;
  buffer buf_n5369( .i (n5128), .o (n5369) );
  assign n5370 = n5368 & ~n5369 ;
  assign n5371 = ~n5131 & n5370 ;
  buffer buf_n5372( .i (n5371), .o (n5372) );
  buffer buf_n5373( .i (n5372), .o (n5373) );
  buffer buf_n5374( .i (n5373), .o (n5374) );
  buffer buf_n5375( .i (n5374), .o (n5375) );
  buffer buf_n5376( .i (n5375), .o (n5376) );
  buffer buf_n5377( .i (n5376), .o (n5377) );
  assign n5378 = ( n430 & n1446 ) | ( n430 & ~n4763 ) | ( n1446 & ~n4763 ) ;
  assign n5379 = ~n431 & n5378 ;
  assign n5380 = ~n698 & n5379 ;
  assign n5381 = ( ~n823 & n5122 ) | ( ~n823 & n5380 ) | ( n5122 & n5380 ) ;
  assign n5382 = ~n4694 & n5381 ;
  buffer buf_n5383( .i (n3718), .o (n5383) );
  assign n5384 = n5382 & ~n5383 ;
  buffer buf_n5385( .i (n4029), .o (n5385) );
  assign n5386 = ( ~n4319 & n5384 ) | ( ~n4319 & n5385 ) | ( n5384 & n5385 ) ;
  buffer buf_n5387( .i (n5385), .o (n5387) );
  assign n5388 = n5386 & ~n5387 ;
  buffer buf_n5389( .i (n5388), .o (n5389) );
  buffer buf_n5390( .i (n5389), .o (n5390) );
  buffer buf_n5391( .i (n5390), .o (n5391) );
  buffer buf_n5392( .i (n5391), .o (n5392) );
  buffer buf_n5393( .i (n5392), .o (n5393) );
  buffer buf_n5394( .i (n5393), .o (n5394) );
  buffer buf_n5395( .i (n5394), .o (n5395) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n5396( .i (n4694), .o (n5396) );
  assign n5397 = n413 & ~n5396 ;
  buffer buf_n5398( .i (n3984), .o (n5398) );
  assign n5399 = ( n436 & n5397 ) | ( n436 & ~n5398 ) | ( n5397 & ~n5398 ) ;
  assign n5400 = ~n437 & n5399 ;
  assign n5401 = ~n5369 & n5400 ;
  buffer buf_n5402( .i (n4671), .o (n5402) );
  assign n5403 = ( ~n5131 & n5401 ) | ( ~n5131 & n5402 ) | ( n5401 & n5402 ) ;
  assign n5404 = ~n2822 & n5403 ;
  buffer buf_n5405( .i (n5404), .o (n5405) );
  buffer buf_n5406( .i (n5405), .o (n5406) );
  buffer buf_n5407( .i (n5406), .o (n5407) );
  buffer buf_n5408( .i (n5407), .o (n5408) );
  assign n5409 = n5395 | n5408 ;
  assign n5410 = ( ~n5138 & n5377 ) | ( ~n5138 & n5409 ) | ( n5377 & n5409 ) ;
  assign n5411 = n5139 | n5410 ;
  buffer buf_n5412( .i (n456), .o (n5412) );
  buffer buf_n5413( .i (n5412), .o (n5413) );
  buffer buf_n5414( .i (n1325), .o (n5414) );
  assign n5415 = ( n223 & n5413 ) | ( n223 & n5414 ) | ( n5413 & n5414 ) ;
  assign n5416 = ~n224 & n5415 ;
  buffer buf_n5417( .i (n5416), .o (n5417) );
  buffer buf_n5418( .i (n5417), .o (n5418) );
  assign n5419 = ( n1970 & n5014 ) | ( n1970 & ~n5417 ) | ( n5014 & ~n5417 ) ;
  assign n5420 = n5418 & n5419 ;
  assign n5421 = ( n4651 & n5402 ) | ( n4651 & n5420 ) | ( n5402 & n5420 ) ;
  assign n5422 = ~n2822 & n5421 ;
  buffer buf_n5423( .i (n5422), .o (n5423) );
  buffer buf_n5424( .i (n5423), .o (n5424) );
  buffer buf_n5425( .i (n5424), .o (n5425) );
  buffer buf_n5426( .i (n5425), .o (n5426) );
  buffer buf_n5427( .i (n5426), .o (n5427) );
  assign n5428 = ( ~n2900 & n5172 ) | ( ~n2900 & n5427 ) | ( n5172 & n5427 ) ;
  assign n5429 = n2901 | n5428 ;
  assign n5430 = n5411 | n5429 ;
  assign n5431 = ( n3047 & ~n3093 ) | ( n3047 & n5430 ) | ( ~n3093 & n5430 ) ;
  assign n5432 = n3094 | n5431 ;
  assign n5433 = n2145 | n3159 ;
  buffer buf_n5434( .i (n5433), .o (n5434) );
  buffer buf_n5435( .i (n5434), .o (n5435) );
  buffer buf_n5436( .i (n5435), .o (n5436) );
  buffer buf_n5211( .i (n5210), .o (n5211) );
  assign n5437 = n2091 | n5211 ;
  assign n5438 = n2130 | n5437 ;
  assign n5439 = n1883 | n5198 ;
  assign n5440 = ( n2722 & ~n4011 ) | ( n2722 & n5439 ) | ( ~n4011 & n5439 ) ;
  assign n5441 = n4012 | n5440 ;
  assign n5442 = n1767 | n5441 ;
  assign n5443 = ( ~n2107 & n5195 ) | ( ~n2107 & n5442 ) | ( n5195 & n5442 ) ;
  assign n5444 = n2108 | n5443 ;
  assign n5445 = n5438 | n5444 ;
  assign n5446 = ( ~n2074 & n5436 ) | ( ~n2074 & n5445 ) | ( n5436 & n5445 ) ;
  assign n5447 = n2075 | n5446 ;
  buffer buf_n4054( .i (n4053), .o (n4054) );
  buffer buf_n4055( .i (n4054), .o (n4055) );
  buffer buf_n4206( .i (n4205), .o (n4206) );
  buffer buf_n4207( .i (n4206), .o (n4207) );
  assign n5448 = n456 & ~n4069 ;
  buffer buf_n5449( .i (n4161), .o (n5449) );
  assign n5450 = ( n222 & n5448 ) | ( n222 & n5449 ) | ( n5448 & n5449 ) ;
  assign n5451 = ~n223 & n5450 ;
  assign n5452 = n3634 & n5451 ;
  assign n5453 = ( n5013 & n5385 ) | ( n5013 & n5452 ) | ( n5385 & n5452 ) ;
  assign n5454 = ~n5387 & n5453 ;
  assign n5455 = n4672 & n5454 ;
  buffer buf_n5456( .i (n5455), .o (n5456) );
  buffer buf_n5457( .i (n5456), .o (n5457) );
  buffer buf_n5458( .i (n5457), .o (n5458) );
  buffer buf_n5459( .i (n5458), .o (n5459) );
  buffer buf_n5460( .i (n5459), .o (n5460) );
  buffer buf_n5461( .i (n5460), .o (n5461) );
  buffer buf_n5462( .i (n4764), .o (n5462) );
  buffer buf_n5463( .i (n5462), .o (n5463) );
  assign n5464 = ~n483 & n5463 ;
  assign n5465 = ( n279 & ~n4074 ) | ( n279 & n5464 ) | ( ~n4074 & n5464 ) ;
  assign n5466 = ~n280 & n5465 ;
  buffer buf_n5467( .i (n5466), .o (n5467) );
  buffer buf_n5468( .i (n5467), .o (n5468) );
  buffer buf_n5469( .i (n1969), .o (n5469) );
  assign n5470 = ( n5014 & ~n5467 ) | ( n5014 & n5469 ) | ( ~n5467 & n5469 ) ;
  assign n5471 = n5468 & n5470 ;
  assign n5472 = ( n3150 & n5205 ) | ( n3150 & n5471 ) | ( n5205 & n5471 ) ;
  buffer buf_n5473( .i (n5205), .o (n5473) );
  assign n5474 = n5472 & ~n5473 ;
  buffer buf_n5475( .i (n5474), .o (n5475) );
  buffer buf_n5476( .i (n5475), .o (n5476) );
  buffer buf_n5477( .i (n5476), .o (n5477) );
  buffer buf_n5478( .i (n482), .o (n5478) );
  assign n5479 = ( n300 & n1325 ) | ( n300 & n5478 ) | ( n1325 & n5478 ) ;
  assign n5480 = ~n301 & n5479 ;
  buffer buf_n5481( .i (n5480), .o (n5481) );
  buffer buf_n5482( .i (n5481), .o (n5482) );
  buffer buf_n5483( .i (n5396), .o (n5483) );
  assign n5484 = ( n1969 & ~n5481 ) | ( n1969 & n5483 ) | ( ~n5481 & n5483 ) ;
  assign n5485 = n5482 & n5484 ;
  assign n5486 = ( n3149 & n5369 ) | ( n3149 & n5485 ) | ( n5369 & n5485 ) ;
  assign n5487 = ~n5205 & n5486 ;
  buffer buf_n5488( .i (n5487), .o (n5488) );
  buffer buf_n5489( .i (n5488), .o (n5489) );
  buffer buf_n5490( .i (n5489), .o (n5490) );
  assign n5491 = n2920 | n5490 ;
  assign n5492 = n5477 | n5491 ;
  assign n5493 = n5461 | n5492 ;
  assign n5494 = ( ~n2974 & n4207 ) | ( ~n2974 & n5493 ) | ( n4207 & n5493 ) ;
  assign n5495 = n2975 | n5494 ;
  buffer buf_n3374( .i (n3373), .o (n3374) );
  buffer buf_n3375( .i (n3374), .o (n3375) );
  assign n5496 = ~n482 & n4161 ;
  assign n5497 = ( n278 & ~n5463 ) | ( n278 & n5496 ) | ( ~n5463 & n5496 ) ;
  assign n5498 = ~n279 & n5497 ;
  buffer buf_n5499( .i (n5498), .o (n5499) );
  buffer buf_n5500( .i (n5499), .o (n5500) );
  assign n5501 = ( n4078 & n5483 ) | ( n4078 & ~n5499 ) | ( n5483 & ~n5499 ) ;
  assign n5502 = n5500 & n5501 ;
  buffer buf_n5503( .i (n5502), .o (n5503) );
  buffer buf_n5504( .i (n5503), .o (n5504) );
  buffer buf_n5505( .i (n5504), .o (n5505) );
  buffer buf_n5506( .i (n5505), .o (n5506) );
  buffer buf_n5507( .i (n5506), .o (n5507) );
  buffer buf_n5508( .i (n5507), .o (n5508) );
  buffer buf_n5509( .i (n5508), .o (n5509) );
  buffer buf_n5510( .i (n5509), .o (n5510) );
  buffer buf_n5511( .i (n481), .o (n5511) );
  assign n5512 = ~n5462 & n5511 ;
  assign n5513 = ( n300 & n5449 ) | ( n300 & n5512 ) | ( n5449 & n5512 ) ;
  assign n5514 = ~n301 & n5513 ;
  buffer buf_n5515( .i (n5514), .o (n5515) );
  buffer buf_n5516( .i (n5515), .o (n5516) );
  assign n5517 = ( n4078 & n5483 ) | ( n4078 & ~n5515 ) | ( n5483 & ~n5515 ) ;
  assign n5518 = n5516 & n5517 ;
  buffer buf_n5519( .i (n5518), .o (n5519) );
  buffer buf_n5520( .i (n5519), .o (n5520) );
  buffer buf_n5521( .i (n5520), .o (n5521) );
  buffer buf_n5522( .i (n5521), .o (n5522) );
  buffer buf_n5523( .i (n5522), .o (n5523) );
  buffer buf_n5524( .i (n5523), .o (n5524) );
  buffer buf_n5525( .i (n5524), .o (n5525) );
  assign n5526 = n2955 | n5525 ;
  assign n5527 = n5510 | n5526 ;
  assign n5528 = n3375 | n5527 ;
  assign n5529 = ( ~n4054 & n5495 ) | ( ~n4054 & n5528 ) | ( n5495 & n5528 ) ;
  assign n5530 = n4055 | n5529 ;
  assign n5531 = n5447 | n5530 ;
  assign n5532 = ( ~n5361 & n5432 ) | ( ~n5361 & n5531 ) | ( n5432 & n5531 ) ;
  assign n5533 = n5362 | n5532 ;
  buffer buf_n4605( .i (n4604), .o (n4605) );
  buffer buf_n4606( .i (n4605), .o (n4606) );
  buffer buf_n4589( .i (n4588), .o (n4589) );
  buffer buf_n4590( .i (n4589), .o (n4590) );
  assign n5534 = n4590 | n5003 ;
  assign n5535 = ( n3891 & ~n4605 ) | ( n3891 & n5534 ) | ( ~n4605 & n5534 ) ;
  assign n5536 = n4606 | n5535 ;
  buffer buf_n5537( .i (n5536), .o (n5537) );
  buffer buf_n5538( .i (n5537), .o (n5538) );
  assign n5539 = n1682 | n5184 ;
  assign n5540 = n3978 | n5539 ;
  assign n5541 = ( n1022 & n2561 ) | ( n1022 & n5161 ) | ( n2561 & n5161 ) ;
  assign n5542 = n2602 | n4361 ;
  assign n5543 = n5541 | n5542 ;
  assign n5544 = n3315 | n5543 ;
  assign n5545 = ( ~n1640 & n5540 ) | ( ~n1640 & n5544 ) | ( n5540 & n5544 ) ;
  assign n5546 = n1641 | n5545 ;
  buffer buf_n4593( .i (n4592), .o (n4593) );
  buffer buf_n4594( .i (n4593), .o (n4594) );
  buffer buf_n4595( .i (n4594), .o (n4595) );
  buffer buf_n5547( .i (n958), .o (n5547) );
  assign n5548 = n2558 & ~n5547 ;
  assign n5549 = ~n1020 & n5548 ;
  assign n5550 = n2542 | n5549 ;
  assign n5551 = n4224 | n5550 ;
  assign n5552 = n4595 | n5551 ;
  assign n5553 = ( ~n3956 & n4218 ) | ( ~n3956 & n5552 ) | ( n4218 & n5552 ) ;
  assign n5554 = n3957 | n5553 ;
  assign n5555 = n1716 | n3173 ;
  assign n5556 = n1731 | n5555 ;
  buffer buf_n5262( .i (n5261), .o (n5262) );
  assign n5557 = n2657 | n4324 ;
  assign n5558 = n3787 | n5557 ;
  assign n5559 = n2632 | n5558 ;
  assign n5560 = ( ~n1664 & n3993 ) | ( ~n1664 & n5559 ) | ( n3993 & n5559 ) ;
  assign n5561 = n1665 | n5560 ;
  assign n5562 = n5262 | n5561 ;
  assign n5563 = ( ~n2688 & n5556 ) | ( ~n2688 & n5562 ) | ( n5556 & n5562 ) ;
  assign n5564 = n2689 | n5563 ;
  assign n5565 = n5554 | n5564 ;
  assign n5566 = ( ~n5537 & n5546 ) | ( ~n5537 & n5565 ) | ( n5546 & n5565 ) ;
  assign n5567 = n5538 | n5566 ;
  buffer buf_n5568( .i (n5567), .o (n5568) );
  buffer buf_n5569( .i (n5568), .o (n5569) );
  buffer buf_n5232( .i (n5231), .o (n5232) );
  buffer buf_n5233( .i (n5232), .o (n5233) );
  buffer buf_n5234( .i (n5233), .o (n5234) );
  buffer buf_n5235( .i (n5234), .o (n5235) );
  buffer buf_n5236( .i (n5235), .o (n5236) );
  buffer buf_n5237( .i (n5236), .o (n5237) );
  assign n5570 = n4276 | n5324 ;
  assign n5571 = ( n5195 & ~n5236 ) | ( n5195 & n5570 ) | ( ~n5236 & n5570 ) ;
  assign n5572 = n5237 | n5571 ;
  assign n5573 = n2104 | n5208 ;
  assign n5574 = n2460 | n5573 ;
  assign n5575 = n2086 | n4249 ;
  assign n5576 = ( ~n2477 & n3579 ) | ( ~n2477 & n5575 ) | ( n3579 & n5575 ) ;
  assign n5577 = n2478 | n5576 ;
  assign n5578 = n4260 | n5577 ;
  assign n5579 = ( ~n4181 & n5574 ) | ( ~n4181 & n5578 ) | ( n5574 & n5578 ) ;
  assign n5580 = n4182 | n5579 ;
  assign n5581 = n2799 | n2836 ;
  assign n5582 = n3641 | n5581 ;
  assign n5583 = n2502 | n5582 ;
  assign n5584 = ( ~n3748 & n3766 ) | ( ~n3748 & n5583 ) | ( n3766 & n5583 ) ;
  assign n5585 = n3749 | n5584 ;
  assign n5586 = n5580 | n5585 ;
  assign n5587 = n5572 | n5586 ;
  buffer buf_n5588( .i (n5587), .o (n5588) );
  buffer buf_n5589( .i (n5588), .o (n5589) );
  buffer buf_n2675( .i (n2674), .o (n2675) );
  buffer buf_n5253( .i (n5252), .o (n5253) );
  buffer buf_n5254( .i (n5253), .o (n5254) );
  assign n5590 = n2675 | n5254 ;
  assign n5591 = ( n2203 & ~n2437 ) | ( n2203 & n5590 ) | ( ~n2437 & n5590 ) ;
  assign n5592 = n2438 | n5591 ;
  assign n5593 = n3624 | n4775 ;
  assign n5594 = ( ~n3510 & n4867 ) | ( ~n3510 & n5593 ) | ( n4867 & n5593 ) ;
  assign n5595 = n3511 | n5594 ;
  assign n5596 = n2128 | n4528 ;
  assign n5597 = n5595 | n5596 ;
  assign n5598 = ( ~n2408 & n5434 ) | ( ~n2408 & n5597 ) | ( n5434 & n5597 ) ;
  assign n5599 = n2409 | n5598 ;
  assign n5600 = n2171 | n4746 ;
  assign n5601 = ( ~n1622 & n2699 ) | ( ~n1622 & n5600 ) | ( n2699 & n5600 ) ;
  assign n5602 = n1623 | n5601 ;
  assign n5603 = n5599 | n5602 ;
  assign n5604 = ( ~n5588 & n5592 ) | ( ~n5588 & n5603 ) | ( n5592 & n5603 ) ;
  assign n5605 = n5589 | n5604 ;
  assign n5606 = n1836 | n3356 ;
  assign n5607 = n4046 | n5606 ;
  assign n5608 = n3297 | n5607 ;
  assign n5609 = ( ~n1865 & n3366 ) | ( ~n1865 & n5608 ) | ( n3366 & n5608 ) ;
  assign n5610 = n1866 | n5609 ;
  buffer buf_n5611( .i (n5610), .o (n5611) );
  buffer buf_n5612( .i (n5611), .o (n5612) );
  assign n5613 = n4011 | n4390 ;
  assign n5614 = ( ~n1820 & n3845 ) | ( ~n1820 & n5613 ) | ( n3845 & n5613 ) ;
  assign n5615 = n1821 | n5614 ;
  assign n5616 = n1997 | n5519 ;
  assign n5617 = n2950 | n5616 ;
  assign n5618 = n5065 | n5617 ;
  assign n5619 = ( ~n4654 & n5053 ) | ( ~n4654 & n5618 ) | ( n5053 & n5618 ) ;
  assign n5620 = n4655 | n5619 ;
  assign n5621 = n3377 | n5503 ;
  assign n5622 = n5456 | n5621 ;
  assign n5623 = n5036 | n5622 ;
  assign n5624 = ( ~n4676 & n5020 ) | ( ~n4676 & n5623 ) | ( n5020 & n5623 ) ;
  assign n5625 = n4677 | n5624 ;
  assign n5626 = n5620 | n5625 ;
  assign n5627 = ( ~n5611 & n5615 ) | ( ~n5611 & n5626 ) | ( n5615 & n5626 ) ;
  assign n5628 = n5612 | n5627 ;
  buffer buf_n5629( .i (n5628), .o (n5629) );
  buffer buf_n5630( .i (n5629), .o (n5630) );
  buffer buf_n1889( .i (n1888), .o (n1889) );
  assign n5631 = n3669 | n4038 ;
  assign n5632 = n3473 | n5631 ;
  assign n5633 = n4125 | n5632 ;
  assign n5634 = ( ~n1888 & n2864 ) | ( ~n1888 & n5633 ) | ( n2864 & n5633 ) ;
  assign n5635 = n1889 | n5634 ;
  assign n5636 = n5200 | n5336 ;
  assign n5637 = n3657 | n4993 ;
  assign n5638 = ( ~n1765 & n2824 ) | ( ~n1765 & n5637 ) | ( n2824 & n5637 ) ;
  assign n5639 = n1766 | n5638 ;
  assign n5640 = n5636 | n5639 ;
  assign n5641 = ( ~n4067 & n4566 ) | ( ~n4067 & n5640 ) | ( n4566 & n5640 ) ;
  assign n5642 = n4068 | n5641 ;
  assign n5643 = n2724 | n4987 ;
  assign n5644 = ( ~n1547 & n4893 ) | ( ~n1547 & n5643 ) | ( n4893 & n5643 ) ;
  assign n5645 = n1548 | n5644 ;
  assign n5646 = n5642 | n5645 ;
  assign n5647 = ( ~n5629 & n5635 ) | ( ~n5629 & n5646 ) | ( n5635 & n5646 ) ;
  assign n5648 = n5630 | n5647 ;
  assign n5649 = n4543 | n4941 ;
  assign n5650 = n5488 | n5649 ;
  assign n5651 = ( ~n4959 & n5475 ) | ( ~n4959 & n5650 ) | ( n5475 & n5650 ) ;
  assign n5652 = n4960 | n5651 ;
  assign n5653 = n5293 | n5652 ;
  assign n5654 = ( ~n4377 & n4635 ) | ( ~n4377 & n5653 ) | ( n4635 & n5653 ) ;
  assign n5655 = n4378 | n5654 ;
  buffer buf_n5656( .i (n5655), .o (n5656) );
  buffer buf_n5657( .i (n5656), .o (n5657) );
  assign n5658 = n1440 | n3273 ;
  assign n5659 = n1431 | n5658 ;
  assign n5660 = n1519 | n3058 ;
  assign n5661 = n3087 | n5660 ;
  buffer buf_n5662( .i (n3033), .o (n5662) );
  assign n5663 = n5084 | n5662 ;
  assign n5664 = n5661 | n5663 ;
  assign n5665 = n3077 | n5664 ;
  assign n5666 = ( ~n1362 & n5659 ) | ( ~n1362 & n5665 ) | ( n5659 & n5665 ) ;
  assign n5667 = n1363 | n5666 ;
  assign n5668 = n2988 | n4701 ;
  assign n5669 = n3259 | n5668 ;
  assign n5670 = n3245 | n5669 ;
  assign n5671 = ( n1581 & ~n2933 ) | ( n1581 & n5670 ) | ( ~n2933 & n5670 ) ;
  assign n5672 = n2934 | n5671 ;
  assign n5673 = n3205 | n5423 ;
  assign n5674 = n4971 | n5673 ;
  assign n5675 = n5672 | n5674 ;
  assign n5676 = ( ~n3199 & n5301 ) | ( ~n3199 & n5675 ) | ( n5301 & n5675 ) ;
  assign n5677 = n3200 | n5676 ;
  buffer buf_n3290( .i (n3289), .o (n3290) );
  buffer buf_n2033( .i (n2032), .o (n2033) );
  assign n5678 = n1921 | n4718 ;
  assign n5679 = n2033 | n5678 ;
  assign n5680 = n797 & n1536 ;
  buffer buf_n5681( .i (n5680), .o (n5681) );
  buffer buf_n5682( .i (n5681), .o (n5682) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  assign n5683 = ( n1803 & n4857 ) | ( n1803 & ~n5681 ) | ( n4857 & ~n5681 ) ;
  assign n5684 = n5682 & n5683 ;
  assign n5685 = n5389 | n5684 ;
  assign n5686 = n3683 | n5685 ;
  assign n5687 = n5372 | n5686 ;
  assign n5688 = ( ~n5134 & n5405 ) | ( ~n5134 & n5687 ) | ( n5405 & n5687 ) ;
  assign n5689 = n5135 | n5688 ;
  assign n5690 = n5281 | n5689 ;
  assign n5691 = ( ~n3289 & n5679 ) | ( ~n3289 & n5690 ) | ( n5679 & n5690 ) ;
  assign n5692 = n3290 | n5691 ;
  assign n5693 = n5677 | n5692 ;
  assign n5694 = ( ~n5656 & n5667 ) | ( ~n5656 & n5693 ) | ( n5667 & n5693 ) ;
  assign n5695 = n5657 | n5694 ;
  assign n5696 = n5648 | n5695 ;
  assign n5697 = ( ~n5568 & n5605 ) | ( ~n5568 & n5696 ) | ( n5605 & n5696 ) ;
  assign n5698 = n5569 | n5697 ;
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  assign n5699 = n637 & n1353 ;
  assign n5700 = ( n538 & n1509 ) | ( n538 & n5699 ) | ( n1509 & n5699 ) ;
  assign n5701 = ~n539 & n5700 ;
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n571( .i (n570), .o (n571) );
  assign n5702 = ~n5320 & n5473 ;
  buffer buf_n5703( .i (n5702), .o (n5703) );
  assign n5704 = ~n928 & n5703 ;
  assign n5705 = n537 & n5704 ;
  assign n5706 = ( n571 & n603 ) | ( n571 & n5705 ) | ( n603 & n5705 ) ;
  assign n5707 = ~n604 & n5706 ;
  assign n5708 = n5701 | n5707 ;
  buffer buf_n5709( .i (n5708), .o (n5709) );
  buffer buf_n5710( .i (n5709), .o (n5710) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  assign n5711 = n775 & n5709 ;
  assign n5712 = ( n679 & n5710 ) | ( n679 & n5711 ) | ( n5710 & n5711 ) ;
  buffer buf_n5713( .i (n5712), .o (n5713) );
  buffer buf_n5714( .i (n5713), .o (n5714) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  assign n5715 = n4029 & ~n5328 ;
  buffer buf_n5716( .i (n5715), .o (n5716) );
  buffer buf_n5717( .i (n5716), .o (n5717) );
  assign n5722 = n368 & n4319 ;
  assign n5723 = ( n799 & ~n5716 ) | ( n799 & n5722 ) | ( ~n5716 & n5722 ) ;
  assign n5724 = n5717 & n5723 ;
  buffer buf_n5725( .i (n5724), .o (n5725) );
  buffer buf_n5726( .i (n5725), .o (n5726) );
  buffer buf_n5727( .i (n5726), .o (n5727) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  assign n5728 = ( n172 & n567 ) | ( n172 & n5725 ) | ( n567 & n5725 ) ;
  assign n5729 = n831 & ~n5728 ;
  assign n5730 = ( n832 & n5727 ) | ( n832 & ~n5729 ) | ( n5727 & ~n5729 ) ;
  assign n5731 = n537 & ~n5730 ;
  buffer buf_n5718( .i (n5717), .o (n5718) );
  buffer buf_n5719( .i (n5718), .o (n5719) );
  buffer buf_n5720( .i (n5719), .o (n5720) );
  buffer buf_n5721( .i (n5720), .o (n5721) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  assign n5732 = ~n172 & n4808 ;
  assign n5733 = n144 & n5732 ;
  assign n5734 = n5721 & n5733 ;
  assign n5735 = n537 | n5734 ;
  assign n5736 = ~n5731 & n5735 ;
  assign n5737 = ~n896 & n5736 ;
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  assign n5738 = n668 & n4671 ;
  assign n5739 = ( ~n228 & n4967 ) | ( ~n228 & n5738 ) | ( n4967 & n5738 ) ;
  assign n5740 = n567 & ~n5739 ;
  buffer buf_n705( .i (n704), .o (n705) );
  assign n5741 = n705 & ~n5402 ;
  assign n5742 = n567 | n5741 ;
  assign n5743 = ~n5740 & n5742 ;
  buffer buf_n5744( .i (n4810), .o (n5744) );
  assign n5745 = ( n536 & n5743 ) | ( n536 & ~n5744 ) | ( n5743 & ~n5744 ) ;
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  assign n5746 = n202 | n829 ;
  assign n5747 = n5227 & ~n5385 ;
  buffer buf_n5748( .i (n5747), .o (n5748) );
  assign n5751 = n5316 & ~n5748 ;
  buffer buf_n5752( .i (n5751), .o (n5752) );
  assign n5753 = ~n5746 & n5752 ;
  buffer buf_n5749( .i (n5748), .o (n5749) );
  buffer buf_n5750( .i (n5749), .o (n5750) );
  assign n5754 = ( n802 & ~n5750 ) | ( n802 & n5752 ) | ( ~n5750 & n5752 ) ;
  assign n5755 = ( ~n860 & n5753 ) | ( ~n860 & n5754 ) | ( n5753 & n5754 ) ;
  assign n5756 = ( n536 & n5744 ) | ( n536 & ~n5755 ) | ( n5744 & ~n5755 ) ;
  assign n5757 = n5745 & ~n5756 ;
  assign n5758 = ~n228 & n5131 ;
  assign n5759 = ~n830 & n5758 ;
  assign n5760 = n535 & n5759 ;
  assign n5761 = ( n569 & n861 ) | ( n569 & n5760 ) | ( n861 & n5760 ) ;
  assign n5762 = ~n862 & n5761 ;
  assign n5763 = n5757 | n5762 ;
  buffer buf_n5764( .i (n895), .o (n5764) );
  assign n5765 = n5763 & n5764 ;
  assign n5766 = n5737 | n5765 ;
  assign n5767 = n606 & n5766 ;
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n5768( .i (n5473), .o (n5768) );
  assign n5769 = ( ~n803 & n860 ) | ( ~n803 & n5768 ) | ( n860 & n5768 ) ;
  buffer buf_n5770( .i (n5769), .o (n5770) );
  assign n5771 = ( n894 & n929 ) | ( n894 & ~n5770 ) | ( n929 & ~n5770 ) ;
  assign n5772 = ( ~n862 & n929 ) | ( ~n862 & n5770 ) | ( n929 & n5770 ) ;
  assign n5773 = n5771 & ~n5772 ;
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  assign n5774 = n570 & ~n1335 ;
  buffer buf_n5775( .i (n5774), .o (n5775) );
  assign n5776 = n5773 & n5775 ;
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n5777( .i (n5402), .o (n5777) );
  buffer buf_n5778( .i (n5777), .o (n5778) );
  assign n5779 = n5768 & ~n5778 ;
  assign n5780 = ( n231 & ~n5744 ) | ( n231 & n5779 ) | ( ~n5744 & n5779 ) ;
  assign n5781 = ~n232 & n5780 ;
  buffer buf_n145( .i (n144), .o (n145) );
  assign n5782 = ( n144 & n1351 ) | ( n144 & n5778 ) | ( n1351 & n5778 ) ;
  assign n5783 = ~n145 & n5782 ;
  assign n5784 = ~n175 & n5783 ;
  assign n5785 = ( ~n176 & n5781 ) | ( ~n176 & n5784 ) | ( n5781 & n5784 ) ;
  assign n5786 = ( ~n1337 & n5775 ) | ( ~n1337 & n5785 ) | ( n5775 & n5785 ) ;
  assign n5787 = ( ~n540 & n5776 ) | ( ~n540 & n5786 ) | ( n5776 & n5786 ) ;
  assign n5788 = n606 | n5787 ;
  assign n5789 = ( ~n607 & n5767 ) | ( ~n607 & n5788 ) | ( n5767 & n5788 ) ;
  assign n5790 = n643 | n5789 ;
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n5791( .i (n5387), .o (n5791) );
  assign n5792 = n227 | n5791 ;
  assign n5793 = n463 | n5792 ;
  buffer buf_n5794( .i (n5793), .o (n5794) );
  buffer buf_n5795( .i (n5794), .o (n5795) );
  assign n5798 = ( n599 & n670 ) | ( n599 & n5777 ) | ( n670 & n5777 ) ;
  assign n5799 = n5794 | n5798 ;
  assign n5800 = ( n861 & ~n5795 ) | ( n861 & n5799 ) | ( ~n5795 & n5799 ) ;
  assign n5801 = n570 & ~n5800 ;
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n5802( .i (n569), .o (n5802) );
  assign n5803 = n1951 | n5802 ;
  assign n5804 = ~n5801 & n5803 ;
  buffer buf_n5805( .i (n5804), .o (n5805) );
  buffer buf_n5806( .i (n5805), .o (n5806) );
  assign n5807 = ( n540 & ~n932 ) | ( n540 & n5805 ) | ( ~n932 & n5805 ) ;
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n5796( .i (n5795), .o (n5796) );
  buffer buf_n5797( .i (n5796), .o (n5797) );
  assign n5808 = ( n571 & n1810 ) | ( n571 & ~n5797 ) | ( n1810 & ~n5797 ) ;
  assign n5809 = ~n572 & n5808 ;
  assign n5810 = n932 & n5809 ;
  assign n5811 = ( n5806 & ~n5807 ) | ( n5806 & n5810 ) | ( ~n5807 & n5810 ) ;
  assign n5812 = ~n899 & n5811 ;
  assign n5813 = n643 & ~n5812 ;
  assign n5814 = n5790 & ~n5813 ;
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  assign n5815 = ~n673 & n709 ;
  buffer buf_n1543( .i (n1542), .o (n1543) );
  assign n5816 = n5473 | n5777 ;
  assign n5817 = n4810 & n5816 ;
  assign n5818 = ( n1543 & n5703 ) | ( n1543 & ~n5817 ) | ( n5703 & ~n5817 ) ;
  assign n5819 = ~n602 & n5818 ;
  assign n5820 = ( n674 & n5815 ) | ( n674 & n5819 ) | ( n5815 & n5819 ) ;
  assign n5821 = ( n115 & n1337 ) | ( n115 & n5820 ) | ( n1337 & n5820 ) ;
  assign n5822 = ~n116 & n5821 ;
  assign n5823 = n1389 | n5822 ;
  assign n5824 = ( ~n1417 & n1464 ) | ( ~n1417 & n5823 ) | ( n1464 & n5823 ) ;
  assign n5825 = n1418 | n5824 ;
  buffer buf_n5826( .i (n5825), .o (n5826) );
  assign n5827 = ( ~n5713 & n5814 ) | ( ~n5713 & n5826 ) | ( n5814 & n5826 ) ;
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  assign n5828 = n83 & ~n5826 ;
  assign n5829 = ( n5714 & n5827 ) | ( n5714 & ~n5828 ) | ( n5827 & ~n5828 ) ;
  assign n5830 = n3862 | n3978 ;
  assign n5831 = ( n2615 & ~n2664 ) | ( n2615 & n5830 ) | ( ~n2664 & n5830 ) ;
  assign n5832 = n2665 | n5831 ;
  buffer buf_n5833( .i (n5832), .o (n5833) );
  buffer buf_n5834( .i (n5833), .o (n5834) );
  buffer buf_n4556( .i (n4555), .o (n4556) );
  buffer buf_n4557( .i (n4556), .o (n4557) );
  buffer buf_n4558( .i (n4557), .o (n4558) );
  buffer buf_n4559( .i (n4558), .o (n4559) );
  assign n5835 = n2919 | n2952 ;
  buffer buf_n5836( .i (n2970), .o (n5836) );
  assign n5837 = ( ~n3299 & n5835 ) | ( ~n3299 & n5836 ) | ( n5835 & n5836 ) ;
  assign n5838 = n3300 | n5837 ;
  assign n5839 = n4051 | n5838 ;
  assign n5840 = ( n2726 & ~n4015 ) | ( n2726 & n5839 ) | ( ~n4015 & n5839 ) ;
  assign n5841 = n4016 | n5840 ;
  buffer buf_n4183( .i (n4182), .o (n4183) );
  assign n5842 = n2837 | n2873 ;
  assign n5843 = ( ~n2801 & n2825 ) | ( ~n2801 & n5842 ) | ( n2825 & n5842 ) ;
  assign n5844 = n2802 | n5843 ;
  assign n5845 = n4150 | n5844 ;
  assign n5846 = ( ~n2505 & n4183 ) | ( ~n2505 & n5845 ) | ( n4183 & n5845 ) ;
  assign n5847 = n2506 | n5846 ;
  assign n5848 = n5841 | n5847 ;
  assign n5849 = ( n4559 & ~n5833 ) | ( n4559 & n5848 ) | ( ~n5833 & n5848 ) ;
  assign n5850 = n5834 | n5849 ;
  buffer buf_n5851( .i (n5850), .o (n5851) );
  buffer buf_n5852( .i (n5851), .o (n5852) );
  buffer buf_n4127( .i (n4126), .o (n4127) );
  buffer buf_n4128( .i (n4127), .o (n4128) );
  buffer buf_n4184( .i (n4183), .o (n4184) );
  buffer buf_n3997( .i (n3996), .o (n3997) );
  assign n5853 = n4971 | n5021 ;
  assign n5854 = ( ~n4039 & n5039 ) | ( ~n4039 & n5853 ) | ( n5039 & n5853 ) ;
  assign n5855 = n4040 | n5854 ;
  assign n5856 = n3997 | n5855 ;
  assign n5857 = ( ~n4127 & n4184 ) | ( ~n4127 & n5856 ) | ( n4184 & n5856 ) ;
  assign n5858 = n4128 | n5857 ;
  buffer buf_n5859( .i (n5858), .o (n5859) );
  buffer buf_n5860( .i (n5859), .o (n5860) );
  buffer buf_n5861( .i (n5860), .o (n5861) );
  buffer buf_n5862( .i (n5861), .o (n5862) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  buffer buf_n1983( .i (n1982), .o (n1983) );
  buffer buf_n1984( .i (n1983), .o (n1984) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n1986( .i (n1985), .o (n1986) );
  buffer buf_n4823( .i (n4822), .o (n4823) );
  buffer buf_n4824( .i (n4823), .o (n4824) );
  buffer buf_n4825( .i (n4824), .o (n4825) );
  buffer buf_n4826( .i (n4825), .o (n4826) );
  buffer buf_n4827( .i (n4826), .o (n4827) );
  buffer buf_n4828( .i (n4827), .o (n4828) );
  assign y0 = n1469 ;
  assign y1 = n1474 ;
  assign y2 = 1'b0 ;
  assign y3 = n1486 ;
  assign y4 = n1492 ;
  assign y5 = n1595 ;
  assign y6 = n2209 ;
  assign y7 = n2219 ;
  assign y8 = n2234 ;
  assign y9 = n2244 ;
  assign y10 = n3108 ;
  assign y11 = n3310 ;
  assign y12 = n3483 ;
  assign y13 = n3801 ;
  assign y14 = n3870 ;
  assign y15 = n4216 ;
  assign y16 = n4345 ;
  assign y17 = n4435 ;
  assign y18 = n4495 ;
  assign y19 = n4585 ;
  assign y20 = n2415 ;
  assign y21 = n2443 ;
  assign y22 = n4839 ;
  assign y23 = n4849 ;
  assign y24 = n4300 ;
  assign y25 = n4904 ;
  assign y26 = n4917 ;
  assign y27 = n4929 ;
  assign y28 = n5077 ;
  assign y29 = n5102 ;
  assign y30 = n5112 ;
  assign y31 = n5121 ;
  assign y32 = n5145 ;
  assign y33 = n5154 ;
  assign y34 = n5220 ;
  assign y35 = n5349 ;
  assign y36 = n5533 ;
  assign y37 = n5698 ;
  assign y38 = n5829 ;
  assign y39 = n5852 ;
  assign y40 = n5862 ;
  assign y41 = n1986 ;
  assign y42 = 1'b0 ;
  assign y43 = n4828 ;
  assign y44 = n4300 ;
endmodule
