module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( N1 , N101 , N106 , N111 , N116 , N121 , N126 , N13 , N130 , N135 , N138 , N143 , N146 , N149 , N152 , N153 , N156 , N159 , N165 , N17 , N171 , N177 , N183 , N189 , N195 , N201 , N207 , N210 , N219 , N228 , N237 , N246 , N255 , N259 , N26 , N260 , N261 , N267 , N268 , N29 , N36 , N42 , N51 , N55 , N59 , N68 , N72 , N73 , N74 , N75 , N8 , N80 , N85 , N86 , N87 , N88 , N89 , N90 , N91 , N96 , N388 , N389 , N390 , N391 , N418 , N419 , N420 , N421 , N422 , N423 , N446 , N447 , N448 , N449 , N450 , N767 , N768 , N850 , N863 , N864 , N865 , N866 , N874 , N878 , N879 , N880 );
  input N1 , N101 , N106 , N111 , N116 , N121 , N126 , N13 , N130 , N135 , N138 , N143 , N146 , N149 , N152 , N153 , N156 , N159 , N165 , N17 , N171 , N177 , N183 , N189 , N195 , N201 , N207 , N210 , N219 , N228 , N237 , N246 , N255 , N259 , N26 , N260 , N261 , N267 , N268 , N29 , N36 , N42 , N51 , N55 , N59 , N68 , N72 , N73 , N74 , N75 , N8 , N80 , N85 , N86 , N87 , N88 , N89 , N90 , N91 , N96 ;
  output N388 , N389 , N390 , N391 , N418 , N419 , N420 , N421 , N422 , N423 , N446 , N447 , N448 , N449 , N450 , N767 , N768 , N850 , N863 , N864 , N865 , N866 , N874 , N878 , N879 , N880 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 ;
  assign n61 = N29 & N75 ;
  buffer buf_n62( .i (n61), .o (n62) );
  assign n63 = N42 & n62 ;
  assign n64 = N29 & N36 ;
  buffer buf_n65( .i (n64), .o (n65) );
  assign n66 = N80 & n65 ;
  assign n67 = N42 & n65 ;
  buffer buf_n68( .i (n67), .o (n68) );
  assign n69 = N85 & N86 ;
  assign n70 = N1 & N8 ;
  buffer buf_n71( .i (n70), .o (n71) );
  assign n72 = N13 & N17 ;
  buffer buf_n73( .i (n72), .o (n73) );
  assign n74 = n71 & n73 ;
  assign n75 = N1 & N26 ;
  buffer buf_n76( .i (n75), .o (n76) );
  assign n77 = n73 & n76 ;
  buffer buf_n78( .i (n77), .o (n78) );
  assign n79 = n68 | ~n78 ;
  assign n80 = N59 & N75 ;
  buffer buf_n81( .i (n80), .o (n81) );
  assign n82 = ~N80 | ~n81 ;
  assign n83 = N36 & N59 ;
  buffer buf_n84( .i (n83), .o (n84) );
  assign n85 = ~N80 | ~n84 ;
  assign n86 = ~N42 | ~n84 ;
  assign n87 = N87 | N88 ;
  buffer buf_n88( .i (n87), .o (n88) );
  assign n89 = N90 & n88 ;
  assign n90 = ~n68 | ~n78 ;
  assign n91 = N51 & n76 ;
  buffer buf_n92( .i (n91), .o (n92) );
  assign n93 = N13 & N55 ;
  assign n94 = n71 & n93 ;
  buffer buf_n95( .i (n94), .o (n95) );
  assign n96 = N29 & N68 ;
  assign n97 = n95 & n96 ;
  assign n98 = N59 & N68 ;
  buffer buf_n99( .i (n98), .o (n99) );
  assign n100 = N74 & n99 ;
  assign n101 = n95 & n100 ;
  assign n102 = N89 & n88 ;
  assign n103 = N130 | N96 ;
  assign n104 = N130 & N96 ;
  assign n105 = n103 & ~n104 ;
  buffer buf_n106( .i (n105), .o (n106) );
  assign n107 = N91 & n106 ;
  assign n108 = N91 | n106 ;
  assign n109 = ~n107 & n108 ;
  buffer buf_n110( .i (n109), .o (n110) );
  assign n111 = N121 | N135 ;
  assign n112 = N121 & N135 ;
  assign n113 = n111 & ~n112 ;
  buffer buf_n114( .i (n113), .o (n114) );
  assign n115 = N126 & ~n114 ;
  assign n116 = ~N126 & n114 ;
  assign n117 = n115 | n116 ;
  buffer buf_n118( .i (n117), .o (n118) );
  assign n119 = N101 & ~N106 ;
  assign n120 = ~N101 & N106 ;
  assign n121 = n119 | n120 ;
  buffer buf_n122( .i (n121), .o (n122) );
  assign n123 = N111 | N116 ;
  assign n124 = N111 & N116 ;
  assign n125 = n123 & ~n124 ;
  buffer buf_n126( .i (n125), .o (n126) );
  assign n127 = n122 | n126 ;
  assign n128 = n122 & n126 ;
  assign n129 = n127 & ~n128 ;
  buffer buf_n130( .i (n129), .o (n130) );
  assign n131 = n118 | n130 ;
  assign n132 = n118 & n130 ;
  assign n133 = n131 & ~n132 ;
  buffer buf_n134( .i (n133), .o (n134) );
  assign n135 = ~n110 & n134 ;
  assign n136 = n110 & ~n134 ;
  assign n137 = n135 | n136 ;
  assign n138 = N159 | N177 ;
  assign n139 = N159 & N177 ;
  assign n140 = n138 & ~n139 ;
  buffer buf_n141( .i (n140), .o (n141) );
  assign n142 = N130 & ~n141 ;
  assign n143 = ~N130 & n141 ;
  assign n144 = n142 | n143 ;
  buffer buf_n145( .i (n144), .o (n145) );
  assign n146 = N189 | N195 ;
  assign n147 = N189 & N195 ;
  assign n148 = n146 & ~n147 ;
  buffer buf_n149( .i (n148), .o (n149) );
  assign n150 = N207 & ~n149 ;
  assign n151 = ~N207 & n149 ;
  assign n152 = n150 | n151 ;
  buffer buf_n153( .i (n152), .o (n153) );
  assign n154 = ~N165 & N201 ;
  assign n155 = N165 & ~N201 ;
  assign n156 = n154 | n155 ;
  buffer buf_n157( .i (n156), .o (n157) );
  assign n158 = N171 & ~N183 ;
  assign n159 = ~N171 & N183 ;
  assign n160 = n158 | n159 ;
  buffer buf_n161( .i (n160), .o (n161) );
  assign n162 = n157 & ~n161 ;
  assign n163 = ~n157 & n161 ;
  assign n164 = n162 | n163 ;
  buffer buf_n165( .i (n164), .o (n165) );
  assign n166 = ~n153 & n165 ;
  assign n167 = n153 & ~n165 ;
  assign n168 = n166 | n167 ;
  buffer buf_n169( .i (n168), .o (n169) );
  assign n170 = n145 & ~n169 ;
  assign n171 = ~n145 & n169 ;
  assign n172 = n170 | n171 ;
  assign n173 = N156 & N59 ;
  buffer buf_n174( .i (n173), .o (n174) );
  assign n175 = n92 & ~n174 ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n177 = N17 & n176 ;
  assign n178 = N1 & ~n177 ;
  buffer buf_n179( .i (n178), .o (n179) );
  assign n180 = N153 & ~n179 ;
  assign n181 = N80 & n62 ;
  assign n182 = n92 & n181 ;
  buffer buf_n183( .i (n182), .o (n183) );
  assign n184 = N55 & n183 ;
  assign n185 = ~N268 & n184 ;
  buffer buf_n186( .i (n185), .o (n186) );
  assign n191 = N17 & ~N42 ;
  assign n192 = ~N17 & N42 ;
  assign n193 = n191 | n192 ;
  assign n194 = n92 & n174 ;
  assign n195 = n193 & n194 ;
  assign n196 = N42 & n81 ;
  assign n197 = N17 & N51 ;
  assign n198 = n71 & n197 ;
  assign n199 = ~n196 & n198 ;
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  assign n202 = n195 | n201 ;
  buffer buf_n203( .i (n202), .o (n203) );
  assign n208 = N126 & n203 ;
  assign n209 = n186 | n208 ;
  assign n210 = n180 | n209 ;
  buffer buf_n211( .i (n210), .o (n211) );
  assign n212 = N201 | n211 ;
  buffer buf_n213( .i (n212), .o (n213) );
  assign n215 = N201 & n211 ;
  buffer buf_n216( .i (n215), .o (n216) );
  assign n217 = n213 & ~n216 ;
  buffer buf_n218( .i (n217), .o (n218) );
  assign n219 = N261 & n218 ;
  buffer buf_n220( .i (n219), .o (n220) );
  assign n221 = N261 | n218 ;
  assign n222 = N219 & n221 ;
  assign n223 = ~n220 & n222 ;
  assign n224 = N228 & n218 ;
  assign n225 = N237 & n216 ;
  assign n226 = N246 & n211 ;
  assign n227 = N42 & N72 ;
  assign n228 = N73 & n227 ;
  assign n229 = n99 & n228 ;
  assign n230 = n95 & n229 ;
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  assign n233 = N201 & n232 ;
  assign n234 = N255 & N267 ;
  assign n235 = N121 & N210 ;
  assign n236 = n234 | n235 ;
  assign n237 = n233 | n236 ;
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  assign n242 = n226 | n241 ;
  buffer buf_n243( .i (n242), .o (n243) );
  assign n244 = n225 | n243 ;
  buffer buf_n245( .i (n244), .o (n245) );
  assign n246 = n224 | n245 ;
  buffer buf_n247( .i (n246), .o (n247) );
  assign n248 = n223 | n247 ;
  assign n249 = N146 & ~n179 ;
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  assign n254 = N116 & n207 ;
  assign n255 = n190 | n254 ;
  assign n256 = n253 | n255 ;
  buffer buf_n257( .i (n256), .o (n257) );
  assign n258 = N189 & n257 ;
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  assign n263 = N189 | n257 ;
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  assign n267 = N149 & ~n179 ;
  buffer buf_n268( .i (n267), .o (n268) );
  assign n269 = N121 & n204 ;
  assign n270 = n187 | n269 ;
  assign n271 = n268 | n270 ;
  buffer buf_n272( .i (n271), .o (n272) );
  assign n273 = N195 & n272 ;
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  assign n278 = N195 | n272 ;
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n282 = N261 | n216 ;
  assign n283 = n214 & n282 ;
  buffer buf_n284( .i (n283), .o (n284) );
  assign n285 = n281 & n284 ;
  assign n286 = n277 | n285 ;
  buffer buf_n287( .i (n286), .o (n287) );
  assign n288 = n266 & n287 ;
  assign n289 = n262 | n288 ;
  buffer buf_n290( .i (n289), .o (n290) );
  assign n291 = N111 & n204 ;
  assign n292 = N143 & ~n179 ;
  assign n293 = n291 | n292 ;
  assign n294 = n188 | n293 ;
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = N183 & n295 ;
  buffer buf_n297( .i (n296), .o (n297) );
  assign n307 = N183 | n295 ;
  buffer buf_n308( .i (n307), .o (n308) );
  assign n317 = ~n297 & n308 ;
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  assign n325 = n290 | n324 ;
  assign n326 = n290 & n324 ;
  assign n327 = n325 & ~n326 ;
  assign n328 = N219 & n327 ;
  assign n329 = N228 & n318 ;
  assign n330 = N237 & n297 ;
  assign n331 = N246 & n295 ;
  assign n332 = N183 & n232 ;
  assign n333 = N106 & N210 ;
  assign n334 = n332 | n333 ;
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  assign n340 = n331 | n339 ;
  buffer buf_n341( .i (n340), .o (n341) );
  assign n342 = n330 | n341 ;
  buffer buf_n343( .i (n342), .o (n343) );
  assign n344 = n329 | n343 ;
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  assign n352 = n328 | n351 ;
  assign n353 = ~n259 & n264 ;
  buffer buf_n354( .i (n353), .o (n354) );
  assign n355 = n287 | n354 ;
  assign n356 = n287 & n354 ;
  assign n357 = n355 & ~n356 ;
  assign n358 = N219 & n357 ;
  assign n359 = N228 & n354 ;
  assign n360 = N237 & n259 ;
  assign n361 = N246 & n257 ;
  assign n362 = N189 & n232 ;
  assign n363 = N111 & N210 ;
  assign n364 = N255 & N259 ;
  assign n365 = n363 | n364 ;
  assign n366 = n362 | n365 ;
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  assign n375 = n361 | n374 ;
  buffer buf_n376( .i (n375), .o (n376) );
  assign n377 = n360 | n376 ;
  buffer buf_n378( .i (n377), .o (n378) );
  assign n379 = n359 | n378 ;
  buffer buf_n380( .i (n379), .o (n380) );
  assign n381 = n358 | n380 ;
  assign n382 = ~n274 & n279 ;
  buffer buf_n383( .i (n382), .o (n383) );
  assign n384 = n284 | n383 ;
  assign n385 = n284 & n383 ;
  assign n386 = n384 & ~n385 ;
  assign n387 = N219 & n386 ;
  assign n388 = N228 & n383 ;
  assign n389 = N237 & n274 ;
  assign n390 = N246 & n272 ;
  assign n391 = N195 & n232 ;
  assign n392 = N255 & N260 ;
  assign n393 = N116 & N210 ;
  assign n394 = n392 | n393 ;
  assign n395 = n391 | n394 ;
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  assign n401 = n390 | n400 ;
  buffer buf_n402( .i (n401), .o (n402) );
  assign n403 = n389 | n402 ;
  buffer buf_n404( .i (n403), .o (n404) );
  assign n405 = n388 | n404 ;
  buffer buf_n406( .i (n405), .o (n406) );
  assign n407 = n387 | n406 ;
  assign n408 = N91 & n204 ;
  assign n409 = N55 & n176 ;
  buffer buf_n410( .i (n409), .o (n410) );
  assign n411 = N143 & n410 ;
  assign n412 = N17 & ~N268 ;
  assign n413 = n183 & n412 ;
  buffer buf_n414( .i (n413), .o (n414) );
  assign n415 = N138 & N8 ;
  assign n416 = n414 | n415 ;
  assign n417 = n411 | n416 ;
  assign n418 = n408 | n417 ;
  buffer buf_n419( .i (n418), .o (n419) );
  assign n420 = N159 & n419 ;
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  assign n444 = N159 | n419 ;
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n203), .o (n467) );
  assign n468 = N96 & n467 ;
  assign n469 = N146 & n410 ;
  assign n470 = N138 & N51 ;
  assign n471 = n414 | n470 ;
  assign n472 = n469 | n471 ;
  assign n473 = n468 | n472 ;
  buffer buf_n474( .i (n473), .o (n474) );
  assign n475 = N165 & n474 ;
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  assign n496 = N165 | n474 ;
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  assign n516 = N101 & n467 ;
  assign n517 = N149 & n410 ;
  assign n518 = N138 & N17 ;
  assign n519 = n414 | n518 ;
  assign n520 = n517 | n519 ;
  assign n521 = n516 | n520 ;
  buffer buf_n522( .i (n521), .o (n522) );
  assign n523 = N171 & n522 ;
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  assign n541 = N171 | n522 ;
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  assign n558 = N106 & n467 ;
  assign n559 = N153 & n410 ;
  assign n560 = N138 & N152 ;
  assign n561 = n414 | n560 ;
  assign n562 = n559 | n561 ;
  assign n563 = n558 | n562 ;
  buffer buf_n564( .i (n563), .o (n564) );
  assign n565 = N177 & n564 ;
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  assign n580 = N177 | n564 ;
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  assign n594 = n290 & n316 ;
  assign n595 = n306 | n594 ;
  buffer buf_n596( .i (n595), .o (n596) );
  assign n597 = n593 & n596 ;
  assign n598 = n579 | n597 ;
  buffer buf_n599( .i (n598), .o (n599) );
  assign n600 = n557 & n599 ;
  assign n601 = n540 | n600 ;
  buffer buf_n602( .i (n601), .o (n602) );
  assign n603 = n515 & n602 ;
  assign n604 = n495 | n603 ;
  buffer buf_n605( .i (n604), .o (n605) );
  assign n606 = n466 & n605 ;
  assign n607 = n443 | n606 ;
  assign n608 = ~n566 & n581 ;
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  assign n622 = N219 & ~n596 ;
  assign n623 = N228 | n622 ;
  assign n624 = n621 & n623 ;
  assign n625 = N219 & ~n609 ;
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  assign n635 = n596 & n634 ;
  assign n636 = N237 & n566 ;
  assign n637 = N246 & n564 ;
  buffer buf_n638( .i (n231), .o (n638) );
  assign n639 = N177 & n638 ;
  assign n640 = N101 & N210 ;
  assign n641 = n639 | n640 ;
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  assign n646 = n637 | n645 ;
  buffer buf_n647( .i (n646), .o (n647) );
  assign n648 = n636 | n647 ;
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  assign n660 = n635 | n659 ;
  buffer buf_n661( .i (n660), .o (n661) );
  assign n662 = n624 | n661 ;
  assign n663 = ~n421 & n445 ;
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  assign n684 = n605 | n683 ;
  buffer buf_n685( .i (n684), .o (n685) );
  assign n686 = n605 & n683 ;
  assign n687 = N219 & ~n686 ;
  assign n688 = n685 & n687 ;
  assign n689 = N228 & n664 ;
  assign n690 = N237 & n421 ;
  assign n691 = N246 & n419 ;
  assign n692 = N159 & n638 ;
  assign n693 = N210 & N268 ;
  assign n694 = n692 | n693 ;
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  assign n699 = n691 | n698 ;
  buffer buf_n700( .i (n699), .o (n700) );
  assign n701 = n690 | n700 ;
  buffer buf_n702( .i (n701), .o (n702) );
  assign n703 = n689 | n702 ;
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  assign n724 = n688 | n723 ;
  assign n725 = ~n476 & n497 ;
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  assign n743 = n602 & n742 ;
  buffer buf_n744( .i (n743), .o (n744) );
  assign n745 = n602 | n742 ;
  assign n746 = N219 & n745 ;
  assign n747 = ~n744 & n746 ;
  assign n748 = N228 & n726 ;
  assign n749 = N237 & n476 ;
  assign n750 = N246 & n474 ;
  assign n751 = N210 & N91 ;
  assign n752 = N165 & n638 ;
  assign n753 = n751 | n752 ;
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = n750 | n757 ;
  buffer buf_n759( .i (n758), .o (n759) );
  assign n760 = n749 | n759 ;
  buffer buf_n761( .i (n760), .o (n761) );
  assign n762 = n748 | n761 ;
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  assign n780 = n747 | n779 ;
  assign n781 = ~n524 & n542 ;
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  assign n796 = n599 & n795 ;
  buffer buf_n797( .i (n796), .o (n797) );
  assign n798 = n599 | n795 ;
  assign n799 = N219 & n798 ;
  assign n800 = ~n797 & n799 ;
  assign n801 = N228 & n782 ;
  assign n802 = N237 & n524 ;
  assign n803 = N246 & n522 ;
  assign n804 = N210 & N96 ;
  assign n805 = N171 & n638 ;
  assign n806 = n804 | n805 ;
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  assign n811 = n803 | n810 ;
  buffer buf_n812( .i (n811), .o (n812) );
  assign n813 = n802 | n812 ;
  buffer buf_n814( .i (n813), .o (n814) );
  assign n815 = n801 | n814 ;
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  assign n830 = n800 | n829 ;
  assign N388 = n63 ;
  assign N389 = n66 ;
  assign N390 = n68 ;
  assign N391 = n69 ;
  assign N418 = n74 ;
  assign N419 = n79 ;
  assign N420 = n82 ;
  assign N421 = n85 ;
  assign N422 = n86 ;
  assign N423 = n89 ;
  assign N446 = n90 ;
  assign N447 = n92 ;
  assign N448 = n97 ;
  assign N449 = n101 ;
  assign N450 = n102 ;
  assign N767 = n137 ;
  assign N768 = n172 ;
  assign N850 = n248 ;
  assign N863 = n352 ;
  assign N864 = n381 ;
  assign N865 = n407 ;
  assign N866 = n607 ;
  assign N874 = n662 ;
  assign N878 = n724 ;
  assign N879 = n780 ;
  assign N880 = n830 ;
endmodule
