module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 );
  input G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 ;
  output G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 ;
  wire n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 ;
  assign n158 = G141 | G142 ;
  assign n159 = G139 | G140 ;
  assign n160 = n158 | n159 ;
  assign n161 = G121 | G2 ;
  assign n162 = G11 | n161 ;
  assign n163 = G115 & ~G74 ;
  assign n164 = G121 | G7 ;
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  assign n167 = G119 | n165 ;
  assign n168 = G147 | n165 ;
  assign n169 = G53 & ~G96 ;
  assign n170 = G43 | G86 ;
  assign n171 = n169 & ~n170 ;
  buffer buf_n172( .i (n171), .o (n172) );
  assign n173 = ~G106 & G32 ;
  assign n174 = G64 | G76 ;
  assign n175 = n173 & ~n174 ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n177 = n172 | n176 ;
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  assign n183 = G147 & ~n176 ;
  assign n184 = G119 & ~n172 ;
  assign n185 = n183 | n184 ;
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  assign n190 = G145 | G146 ;
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  assign n206 = G109 & ~n194 ;
  assign n207 = G79 & ~n194 ;
  assign n208 = n206 | n207 ;
  assign n209 = G89 & ~n194 ;
  buffer buf_n210( .i (n193), .o (n210) );
  assign n211 = G99 & ~n210 ;
  assign n212 = n209 | n211 ;
  assign n213 = n208 | n212 ;
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  assign n236 = G108 | n204 ;
  assign n237 = G98 & ~n204 ;
  assign n238 = n236 & ~n237 ;
  assign n239 = G88 & ~n204 ;
  buffer buf_n240( .i (n203), .o (n240) );
  assign n241 = G78 & ~n240 ;
  assign n242 = n239 | n241 ;
  assign n243 = n238 & ~n242 ;
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  assign n256 = G80 | n210 ;
  assign n257 = G90 & ~n210 ;
  assign n258 = n256 & ~n257 ;
  assign n259 = G100 & ~n210 ;
  buffer buf_n260( .i (n193), .o (n260) );
  assign n261 = G110 & ~n260 ;
  assign n262 = n259 | n261 ;
  assign n263 = n258 & ~n262 ;
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  assign n286 = G117 & ~G36 ;
  assign n287 = G117 & ~G68 ;
  assign n288 = G120 | n287 ;
  assign n289 = n286 & ~n288 ;
  assign n290 = G117 | G120 ;
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  assign n305 = G46 & ~n296 ;
  assign n306 = G57 & ~n296 ;
  assign n307 = n305 | n306 ;
  assign n308 = n289 & ~n307 ;
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  assign n321 = G117 & ~G37 ;
  assign n322 = G117 & ~G69 ;
  assign n323 = G120 | n322 ;
  assign n324 = n321 & ~n323 ;
  assign n325 = G47 & ~n295 ;
  assign n326 = G58 & ~n295 ;
  assign n327 = n325 | n326 ;
  assign n328 = n324 & ~n327 ;
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  assign n342 = G117 & ~G38 ;
  assign n343 = G117 & ~G70 ;
  assign n344 = G120 | n343 ;
  assign n345 = n342 & ~n344 ;
  assign n346 = G48 & ~n295 ;
  buffer buf_n347( .i (n294), .o (n347) );
  assign n348 = G59 & ~n347 ;
  assign n349 = n346 | n348 ;
  assign n350 = n345 & ~n349 ;
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  assign n364 = G117 & ~G31 ;
  assign n365 = G117 & ~G63 ;
  assign n366 = G120 | n365 ;
  assign n367 = n364 & ~n366 ;
  assign n368 = G42 & ~n294 ;
  assign n369 = G52 & ~n294 ;
  assign n370 = n368 | n369 ;
  assign n371 = n367 & ~n370 ;
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  assign n385 = G122 | n384 ;
  assign n386 = G116 | G121 ;
  assign n387 = n186 | n386 ;
  buffer buf_n388( .i (n387), .o (n388) );
  assign n389 = G28 | n388 ;
  assign n390 = G1 & ~G3 ;
  assign n391 = n388 | n390 ;
  assign n392 = G117 | G39 ;
  assign n393 = G117 & ~G71 ;
  assign n394 = G120 | n393 ;
  assign n395 = n392 & ~n394 ;
  buffer buf_n396( .i (n293), .o (n396) );
  assign n397 = G49 & ~n396 ;
  assign n398 = G60 & ~n396 ;
  assign n399 = n397 | n398 ;
  assign n400 = n395 | n399 ;
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  assign n415 = G56 & ~n299 ;
  assign n416 = G117 | G35 ;
  assign n417 = G117 & ~G67 ;
  assign n418 = G120 | n417 ;
  assign n419 = n416 & ~n418 ;
  assign n420 = n415 & ~n419 ;
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  assign n431 = G117 & ~G34 ;
  assign n432 = G117 & ~G66 ;
  assign n433 = G120 | n432 ;
  assign n434 = n431 & ~n433 ;
  assign n435 = G45 & ~n296 ;
  buffer buf_n436( .i (n347), .o (n436) );
  assign n437 = G55 & ~n436 ;
  assign n438 = n435 | n437 ;
  assign n439 = n434 & ~n438 ;
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  assign n452 = G117 & ~G33 ;
  assign n453 = G117 & ~G65 ;
  assign n454 = G120 | n453 ;
  assign n455 = n452 & ~n454 ;
  assign n456 = G44 & ~n436 ;
  assign n457 = G54 & ~n436 ;
  assign n458 = n456 | n457 ;
  assign n459 = n455 & ~n458 ;
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  assign n472 = G117 & ~G40 ;
  assign n473 = G117 & ~G72 ;
  assign n474 = G120 | n473 ;
  assign n475 = n472 & ~n474 ;
  assign n476 = G50 & ~n396 ;
  assign n477 = G61 & ~n396 ;
  assign n478 = n476 | n477 ;
  assign n479 = n475 & ~n478 ;
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  assign n493 = G123 | n490 ;
  assign n494 = G123 & ~n360 ;
  assign n495 = n493 & ~n494 ;
  buffer buf_n496( .i (n495), .o (n496) );
  assign n497 = G123 | n411 ;
  assign n498 = ~G123 & n338 ;
  assign n499 = n497 & ~n498 ;
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  assign n501 = G118 & ~G122 ;
  assign n502 = n492 | n501 ;
  assign n503 = G123 & ~n382 ;
  assign n504 = G118 | G123 ;
  assign n505 = n490 & ~n504 ;
  assign n506 = n503 | n505 ;
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n205( .i (n204), .o (n205) );
  assign n508 = G77 & ~n205 ;
  assign n509 = G97 & ~n205 ;
  assign n510 = n508 & ~n509 ;
  assign n511 = G107 & ~n205 ;
  assign n512 = G87 & ~n205 ;
  assign n513 = n511 | n512 ;
  assign n514 = n510 & ~n513 ;
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  assign n523 = G143 | n522 ;
  assign n524 = G143 & ~n522 ;
  assign n525 = n523 & ~n524 ;
  assign n526 = G144 | n525 ;
  assign n527 = ~G19 & G23 ;
  buffer buf_n528( .i (n240), .o (n528) );
  assign n529 = G75 & ~n528 ;
  assign n530 = G85 & ~n528 ;
  assign n531 = n529 & ~n530 ;
  assign n532 = G95 & ~n528 ;
  assign n533 = G105 & ~n528 ;
  assign n534 = n532 | n533 ;
  assign n535 = n531 & ~n534 ;
  buffer buf_n536( .i (n535), .o (n536) );
  assign n538 = G23 & ~n536 ;
  assign n539 = n527 & ~n538 ;
  assign n540 = G135 & ~n539 ;
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  assign n544 = G12 & ~G13 ;
  assign n545 = G12 & ~n374 ;
  assign n546 = n544 & ~n545 ;
  assign n547 = G125 & ~n546 ;
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  assign n551 = G12 & ~G15 ;
  assign n552 = ~G12 & n330 ;
  assign n553 = n551 & ~n552 ;
  assign n554 = G130 & ~n553 ;
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  assign n558 = n550 | n557 ;
  assign n559 = n543 | n558 ;
  assign n560 = G12 & ~G5 ;
  assign n561 = G12 & ~n352 ;
  assign n562 = n560 & ~n561 ;
  assign n563 = G129 & ~n562 ;
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  assign n566 = ~G21 & G23 ;
  assign n567 = G23 & ~n275 ;
  assign n568 = n566 & ~n567 ;
  assign n569 = G140 & ~n568 ;
  buffer buf_n570( .i (n569), .o (n570) );
  assign n571 = n565 | n570 ;
  assign n572 = G23 & ~G27 ;
  assign n573 = G23 & ~n244 ;
  assign n574 = n572 & ~n573 ;
  assign n575 = G142 & ~n574 ;
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  assign n578 = n541 | n577 ;
  assign n579 = n571 | n578 ;
  assign n580 = G12 & ~G14 ;
  assign n581 = ~G12 & n403 ;
  assign n582 = n580 & ~n581 ;
  assign n583 = G128 & ~n582 ;
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  assign n586 = G12 & ~G4 ;
  assign n587 = G12 & ~n482 ;
  assign n588 = n586 & ~n587 ;
  assign n589 = G126 & ~n588 ;
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  assign n592 = n585 | n591 ;
  assign n593 = G23 & ~G26 ;
  assign n594 = G23 & ~n224 ;
  assign n595 = n593 & ~n594 ;
  assign n596 = G141 & ~n595 ;
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  assign n599 = n570 | n598 ;
  assign n600 = n592 | n599 ;
  assign n601 = n579 | n600 ;
  assign n602 = n559 | n601 ;
  assign n603 = G23 & ~G24 ;
  buffer buf_n604( .i (n240), .o (n604) );
  assign n605 = G93 & ~n604 ;
  assign n606 = G103 & ~n604 ;
  assign n607 = n605 & ~n606 ;
  assign n608 = G113 & ~n604 ;
  assign n609 = G83 & ~n604 ;
  assign n610 = n608 | n609 ;
  assign n611 = n607 & ~n610 ;
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  assign n614 = G23 & ~n613 ;
  assign n615 = n603 & ~n614 ;
  buffer buf_n616( .i (n615), .o (n616) );
  assign n617 = G136 | n616 ;
  assign n618 = G136 & ~n616 ;
  assign n619 = n617 & ~n618 ;
  assign n620 = G12 & ~G16 ;
  assign n621 = G12 & ~n310 ;
  assign n622 = n620 & ~n621 ;
  buffer buf_n623( .i (n622), .o (n623) );
  assign n624 = G131 | n623 ;
  assign n625 = G131 & ~n623 ;
  assign n626 = n624 & ~n625 ;
  assign n627 = ~G20 & G23 ;
  buffer buf_n628( .i (n240), .o (n628) );
  assign n629 = G82 & ~n628 ;
  assign n630 = G102 & ~n628 ;
  assign n631 = n629 & ~n630 ;
  assign n632 = G112 & ~n628 ;
  assign n633 = G92 & ~n628 ;
  assign n634 = n632 | n633 ;
  assign n635 = n631 & ~n634 ;
  buffer buf_n636( .i (n635), .o (n636) );
  assign n639 = G23 & ~n636 ;
  assign n640 = n627 & ~n639 ;
  buffer buf_n641( .i (n640), .o (n641) );
  assign n642 = G138 | n641 ;
  assign n643 = G138 & ~n641 ;
  assign n644 = n642 & ~n643 ;
  assign n645 = n626 | n644 ;
  assign n646 = n619 | n645 ;
  assign n647 = G23 & ~G25 ;
  buffer buf_n648( .i (n203), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  assign n650 = G81 & ~n649 ;
  assign n651 = G101 & ~n649 ;
  assign n652 = n650 & ~n651 ;
  assign n653 = G111 & ~n649 ;
  assign n654 = G91 & ~n649 ;
  assign n655 = n653 | n654 ;
  assign n656 = n652 & ~n655 ;
  assign n657 = G23 & ~n656 ;
  assign n658 = n647 & ~n657 ;
  assign n659 = G139 & ~n658 ;
  buffer buf_n660( .i (n659), .o (n660) );
  assign n661 = n555 | n660 ;
  assign n662 = G12 & ~G18 ;
  assign n663 = G12 & ~n460 ;
  assign n664 = n662 & ~n663 ;
  assign n665 = G134 & ~n664 ;
  buffer buf_n666( .i (n665), .o (n666) );
  assign n667 = n590 | n666 ;
  assign n668 = n661 | n667 ;
  assign n669 = G12 & ~G6 ;
  assign n670 = G12 & ~n440 ;
  assign n671 = n669 & ~n670 ;
  assign n672 = G133 & ~n671 ;
  buffer buf_n673( .i (n672), .o (n673) );
  assign n674 = G23 & ~n516 ;
  assign n675 = ~G22 & G23 ;
  assign n676 = G9 | n675 ;
  assign n677 = n674 | n676 ;
  assign n678 = n673 | n677 ;
  assign n679 = n576 | n673 ;
  assign n680 = n678 | n679 ;
  assign n681 = n668 | n680 ;
  assign n682 = n564 | n597 ;
  assign n683 = n548 | n584 ;
  assign n684 = n682 | n683 ;
  assign n685 = n660 | n666 ;
  assign n686 = G12 & ~G17 ;
  assign n687 = G12 & ~n421 ;
  assign n688 = n686 & ~n687 ;
  assign n689 = G132 & ~n688 ;
  assign n690 = n685 | n689 ;
  assign n691 = n684 | n690 ;
  assign n692 = n681 | n691 ;
  assign n693 = n646 | n692 ;
  assign n694 = n602 | n693 ;
  buffer buf_n695( .i (n694), .o (n695) );
  assign n696 = G117 & ~G41 ;
  assign n697 = G117 & ~G73 ;
  assign n698 = G120 | n697 ;
  assign n699 = n696 & ~n698 ;
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  assign n700 = G51 & ~n304 ;
  assign n701 = G62 & ~n304 ;
  assign n702 = n700 | n701 ;
  assign n703 = n699 & ~n702 ;
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  assign n706 = G122 & ~n705 ;
  assign n707 = G122 | n706 ;
  assign n708 = n246 | n516 ;
  assign n709 = n246 & ~n516 ;
  assign n710 = n708 & ~n709 ;
  buffer buf_n711( .i (n710), .o (n711) );
  assign n712 = n229 | n711 ;
  assign n713 = ~n229 & n711 ;
  assign n714 = n712 & ~n713 ;
  assign n715 = G29 | n714 ;
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  inverter inv_n718( .i (n717), .o (n718) );
  assign n719 = G123 & ~n704 ;
  assign n720 = G123 | n719 ;
  buffer buf_n721( .i (n720), .o (n721) );
  assign n722 = G127 | n264 ;
  buffer buf_n723( .i (n722), .o (n723) );
  assign n724 = G30 | n214 ;
  buffer buf_n725( .i (n724), .o (n725) );
  assign n726 = n723 | n725 ;
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  assign n732 = ~G8 & n729 ;
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  assign n743 = ~G133 & n742 ;
  assign n744 = G8 | n729 ;
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  assign n754 = n446 | n753 ;
  assign n755 = ~G132 & n740 ;
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  assign n756 = G129 & n731 ;
  assign n757 = G140 & ~n731 ;
  assign n758 = n756 & ~n757 ;
  assign n759 = n352 & ~n758 ;
  buffer buf_n760( .i (n759), .o (n760) );
  assign n761 = ~G128 & n728 ;
  assign n762 = G139 & ~n728 ;
  assign n763 = n761 | n762 ;
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  assign n767 = ~n403 & n766 ;
  assign n768 = ~G126 & n728 ;
  buffer buf_n769( .i (n727), .o (n769) );
  assign n770 = G138 & ~n769 ;
  assign n771 = n768 | n770 ;
  buffer buf_n772( .i (n771), .o (n772) );
  assign n773 = n480 | n772 ;
  assign n774 = ~G125 & n729 ;
  buffer buf_n775( .i (n769), .o (n775) );
  assign n776 = G136 & ~n775 ;
  assign n777 = n774 | n776 ;
  assign n778 = ~n372 & n777 ;
  assign n779 = n773 & n778 ;
  assign n780 = n480 & n772 ;
  assign n781 = n401 & n764 ;
  assign n782 = n780 | n781 ;
  assign n783 = n779 | n782 ;
  assign n784 = ~n767 & n783 ;
  assign n785 = n760 | n784 ;
  assign n786 = G8 & ~n329 ;
  assign n787 = G130 & n733 ;
  assign n788 = G141 & ~n745 ;
  assign n789 = n787 & ~n788 ;
  assign n790 = n786 & ~n789 ;
  buffer buf_n791( .i (n790), .o (n791) );
  assign n793 = n760 | n791 ;
  assign n794 = n785 & ~n793 ;
  buffer buf_n792( .i (n791), .o (n792) );
  assign n795 = G8 & ~n309 ;
  assign n796 = G131 & n734 ;
  assign n797 = G142 & ~n746 ;
  assign n798 = n796 & ~n797 ;
  assign n799 = n795 & ~n798 ;
  buffer buf_n800( .i (n799), .o (n800) );
  assign n802 = n792 | n800 ;
  assign n803 = n794 | n802 ;
  buffer buf_n801( .i (n800), .o (n801) );
  assign n804 = n422 & ~n750 ;
  assign n805 = n801 | n804 ;
  assign n806 = n803 & ~n805 ;
  assign n807 = n755 | n806 ;
  assign n808 = n754 & n807 ;
  assign n809 = n743 | n808 ;
  assign n810 = n723 & ~n725 ;
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  assign n823 = G136 | n612 ;
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  assign n827 = n822 & ~n826 ;
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  assign n828 = G138 | n638 ;
  assign n829 = n821 & ~n828 ;
  buffer buf_n830( .i (n829), .o (n830) );
  assign n834 = n827 & ~n830 ;
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n537( .i (n536), .o (n537) );
  assign n836 = G135 | n537 ;
  buffer buf_n837( .i (n836), .o (n837) );
  assign n840 = G134 & ~n463 ;
  assign n841 = n837 & ~n840 ;
  assign n842 = n822 & ~n841 ;
  assign n843 = n830 | n842 ;
  assign n844 = G135 & ~n537 ;
  assign n845 = n824 & ~n844 ;
  assign n846 = n821 & ~n845 ;
  buffer buf_n847( .i (n846), .o (n847) );
  assign n849 = G134 | n463 ;
  assign n850 = n821 & ~n849 ;
  buffer buf_n851( .i (n850), .o (n851) );
  assign n852 = n847 | n851 ;
  assign n853 = n843 | n852 ;
  assign n854 = n835 & ~n853 ;
  assign n855 = n809 & n854 ;
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  assign n856 = n839 & ~n851 ;
  assign n857 = n848 & ~n856 ;
  assign n858 = n835 & ~n857 ;
  assign n859 = n833 | n858 ;
  assign n860 = ~n855 & ~n859 ;
  assign n861 = G10 & ~n186 ;
  assign n862 = n716 & n861 ;
  inverter inv_n863( .i (n862), .o (n863) );
  assign G2531 = G115 ;
  assign G2532 = G115 ;
  assign G2533 = G115 ;
  assign G2534 = G124 ;
  assign G2535 = G124 ;
  assign G2536 = G137 ;
  assign G2537 = G137 ;
  assign G2538 = G137 ;
  assign G2539 = G32 ;
  assign G2540 = G106 ;
  assign G2541 = G64 ;
  assign G2542 = G76 ;
  assign G2543 = G53 ;
  assign G2544 = G96 ;
  assign G2545 = G43 ;
  assign G2546 = G86 ;
  assign G2547 = n160 ;
  assign G2548 = n162 ;
  assign G2549 = G115 ;
  assign G2550 = n163 ;
  assign G2551 = n166 ;
  assign G2552 = n167 ;
  assign G2553 = n168 ;
  assign G2554 = n182 ;
  assign G2555 = n182 ;
  assign G2556 = n189 ;
  assign G2557 = n235 ;
  assign G2558 = n255 ;
  assign G2559 = n285 ;
  assign G2560 = n320 ;
  assign G2561 = n341 ;
  assign G2562 = n363 ;
  assign G2563 = n385 ;
  assign G2564 = n389 ;
  assign G2565 = n391 ;
  assign G2566 = n414 ;
  assign G2567 = n363 ;
  assign G2568 = n341 ;
  assign G2569 = n320 ;
  assign G2570 = n430 ;
  assign G2571 = n451 ;
  assign G2572 = n471 ;
  assign G2573 = n496 ;
  assign G2574 = n496 ;
  assign G2575 = n500 ;
  assign G2576 = n500 ;
  assign G2577 = n502 ;
  assign G2578 = n507 ;
  assign G2579 = n507 ;
  assign G2580 = n526 ;
  assign G2581 = ~G10 ;
  assign G2582 = 1'b0 ;
  assign G2583 = 1'b0 ;
  assign G2584 = n695 ;
  assign G2585 = n695 ;
  assign G2586 = n707 ;
  assign G2587 = n718 ;
  assign G2588 = n721 ;
  assign G2589 = n721 ;
  assign G2590 = 1'b0 ;
  assign G2591 = n860 ;
  assign G2592 = 1'b0 ;
  assign G2593 = n863 ;
  assign G2594 = n863 ;
endmodule
