module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 ;
  wire n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 ;
  buffer buf_n34( .i (x0), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n378( .i (x22), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n274( .i (x16), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n254( .i (x15), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n526( .i (x31), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  assign n535 = ~n256 & n528 ;
  assign n536 = ~n277 & n535 ;
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n56( .i (x1), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n504( .i (x30), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n465( .i (x28), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n529( .i (n528), .o (n529) );
  assign n540 = n468 & ~n529 ;
  assign n541 = n508 & n540 ;
  assign n542 = ( n61 & n537 ) | ( n61 & n541 ) | ( n537 & n541 ) ;
  assign n543 = n384 & ~n542 ;
  assign n544 = ( n385 & n539 ) | ( n385 & ~n543 ) | ( n539 & ~n543 ) ;
  assign n545 = ~n42 & n544 ;
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n112( .i (x4), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n530( .i (x32), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  assign n559 = ( ~n38 & n116 ) | ( ~n38 & n534 ) | ( n116 & n534 ) ;
  buffer buf_n408( .i (x24), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n486( .i (x29), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  assign n560 = n465 & ~n530 ;
  assign n561 = n487 & n560 ;
  assign n562 = n410 & n561 ;
  assign n563 = n59 & n562 ;
  assign n564 = ~n38 & n563 ;
  assign n565 = ( ~n117 & n559 ) | ( ~n117 & n564 ) | ( n559 & n564 ) ;
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n92( .i (x3), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  assign n582 = n111 & ~n484 ;
  assign n583 = ( n54 & ~n524 ) | ( n54 & n582 ) | ( ~n524 & n582 ) ;
  assign n584 = ~n55 & n583 ;
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  assign n585 = ~n480 & n501 ;
  assign n586 = ~n520 & n585 ;
  assign n587 = n51 | n586 ;
  assign n588 = ( n52 & n110 ) | ( n52 & n587 ) | ( n110 & n587 ) ;
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n202( .i (x11), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n218( .i (x12), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  assign n592 = ( n211 & ~n227 ) | ( n211 & n495 ) | ( ~n227 & n495 ) ;
  buffer buf_n183( .i (x10), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  assign n593 = ~n192 & n495 ;
  assign n594 = ( ~n212 & n592 ) | ( ~n212 & n593 ) | ( n592 & n593 ) ;
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n348( .i (x20), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n334( .i (x19), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n364( .i (x21), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  assign n597 = n345 & n375 ;
  assign n598 = ( n360 & ~n595 ) | ( n360 & n597 ) | ( ~n595 & n597 ) ;
  assign n599 = n596 & n598 ;
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n164( .i (x9), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  assign n604 = ~n181 & n602 ;
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  assign n605 = ~n197 & n216 ;
  assign n606 = ( n179 & ~n233 ) | ( n179 & n605 ) | ( ~n233 & n605 ) ;
  assign n607 = ~n180 & n606 ;
  buffer buf_n198( .i (n197), .o (n198) );
  assign n608 = n211 | n227 ;
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n346( .i (n345), .o (n346) );
  assign n613 = ( ~n228 & n358 ) | ( ~n228 & n496 ) | ( n358 & n496 ) ;
  assign n614 = ( n228 & n374 ) | ( n228 & n496 ) | ( n374 & n496 ) ;
  assign n615 = n613 & n614 ;
  assign n616 = n346 & n615 ;
  assign n617 = n215 & ~n616 ;
  assign n618 = n612 & ~n617 ;
  assign n619 = ( ~n179 & n198 ) | ( ~n179 & n618 ) | ( n198 & n618 ) ;
  assign n620 = n374 & ~n496 ;
  assign n621 = ( n229 & ~n375 ) | ( n229 & n620 ) | ( ~n375 & n620 ) ;
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  assign n624 = ( n215 & n231 ) | ( n215 & n622 ) | ( n231 & n622 ) ;
  assign n625 = ( n612 & n623 ) | ( n612 & ~n624 ) | ( n623 & ~n624 ) ;
  assign n626 = ( n179 & n198 ) | ( n179 & ~n625 ) | ( n198 & ~n625 ) ;
  assign n627 = n619 & n626 ;
  assign n628 = n607 | n627 ;
  assign n629 = ( n603 & ~n604 ) | ( n603 & n628 ) | ( ~n604 & n628 ) ;
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n485( .i (n484), .o (n485) );
  assign n632 = ~n52 & n522 ;
  buffer buf_n633( .i (n632), .o (n633) );
  assign n634 = ( n485 & n630 ) | ( n485 & ~n633 ) | ( n630 & ~n633 ) ;
  assign n635 = n631 & ~n634 ;
  buffer buf_n314( .i (x18), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  assign n636 = n189 & ~n208 ;
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  assign n643 = ( n177 & ~n231 ) | ( n177 & n642 ) | ( ~n231 & n642 ) ;
  assign n644 = ~n178 & n643 ;
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n238( .i (x14), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n294( .i (x17), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  assign n647 = n264 & ~n475 ;
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  assign n651 = ( n252 & n308 ) | ( n252 & n650 ) | ( n308 & n650 ) ;
  assign n652 = ~n253 & n651 ;
  assign n653 = ( n520 & ~n645 ) | ( n520 & n652 ) | ( ~n645 & n652 ) ;
  buffer buf_n121( .i (x6), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  assign n654 = ( ~n124 & n257 ) | ( ~n124 & n297 ) | ( n257 & n297 ) ;
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  assign n662 = ~n259 & n655 ;
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n136( .i (x7), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  assign n665 = ( n143 & ~n301 ) | ( n143 & n663 ) | ( ~n301 & n663 ) ;
  assign n666 = ( n658 & n664 ) | ( n658 & n665 ) | ( n664 & n665 ) ;
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  assign n670 = ( ~n248 & n264 ) | ( ~n248 & n667 ) | ( n264 & n667 ) ;
  assign n671 = n305 & ~n670 ;
  assign n672 = ( n306 & n669 ) | ( n306 & ~n671 ) | ( n669 & ~n671 ) ;
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n393( .i (x23), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  assign n675 = n68 & n477 ;
  buffer buf_n676( .i (n675), .o (n676) );
  assign n677 = ( n407 & ~n673 ) | ( n407 & n676 ) | ( ~n673 & n676 ) ;
  assign n678 = n674 & n677 ;
  assign n679 = n520 & n678 ;
  assign n680 = ( n646 & n653 ) | ( n646 & n679 ) | ( n653 & n679 ) ;
  assign n681 = ~n292 & n680 ;
  assign n682 = ( n53 & ~n333 ) | ( n53 & n681 ) | ( ~n333 & n681 ) ;
  assign n683 = ~n54 & n682 ;
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  assign n685 = n208 | n471 ;
  buffer buf_n686( .i (n685), .o (n686) );
  assign n693 = n226 | n686 ;
  assign n694 = ~n171 & n190 ;
  buffer buf_n695( .i (n694), .o (n695) );
  assign n701 = ~n693 & n695 ;
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  assign n705 = ( n67 & n404 ) | ( n67 & n702 ) | ( n404 & n702 ) ;
  assign n706 = n477 & ~n705 ;
  assign n707 = ( n478 & n704 ) | ( n478 & ~n706 ) | ( n704 & ~n706 ) ;
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  assign n710 = n287 & n327 ;
  assign n711 = n307 & ~n327 ;
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  assign n712 = n133 | n286 ;
  assign n713 = n307 & n712 ;
  assign n714 = ( n710 & n711 ) | ( n710 & ~n713 ) | ( n711 & ~n713 ) ;
  assign n715 = ( n519 & ~n708 ) | ( n519 & n714 ) | ( ~n708 & n714 ) ;
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  assign n716 = ~n295 & n315 ;
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n153( .i (x8), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  assign n721 = n317 & ~n717 ;
  assign n722 = ~n157 & n721 ;
  assign n723 = ( n299 & n719 ) | ( n299 & ~n722 ) | ( n719 & ~n722 ) ;
  assign n724 = ( ~n127 & n720 ) | ( ~n127 & n723 ) | ( n720 & n723 ) ;
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  assign n727 = ~n281 & n400 ;
  assign n728 = ( ~n473 & n725 ) | ( ~n473 & n727 ) | ( n725 & n727 ) ;
  assign n729 = ~n726 & n728 ;
  assign n730 = n228 & n729 ;
  assign n731 = ( n194 & n213 ) | ( n194 & n730 ) | ( n213 & n730 ) ;
  assign n732 = ~n195 & n731 ;
  assign n733 = ~n177 & n732 ;
  assign n734 = n70 & n733 ;
  assign n735 = n519 & n734 ;
  assign n736 = ( n709 & n715 ) | ( n709 & n735 ) | ( n715 & n735 ) ;
  assign n737 = ~n51 & n736 ;
  assign n738 = ~n272 & n737 ;
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  assign n742 = n208 & n224 ;
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  assign n748 = ( n174 & n193 ) | ( n174 & ~n475 ) | ( n193 & ~n475 ) ;
  assign n749 = n746 & n748 ;
  assign n750 = ( n477 & n747 ) | ( n477 & ~n749 ) | ( n747 & ~n749 ) ;
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  assign n753 = ~n327 & n391 ;
  assign n754 = ( n268 & ~n751 ) | ( n268 & n753 ) | ( ~n751 & n753 ) ;
  assign n755 = n752 & n754 ;
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  assign n758 = ( n73 & n521 ) | ( n73 & ~n756 ) | ( n521 & ~n756 ) ;
  assign n759 = ( n67 & n389 ) | ( n67 & n702 ) | ( n389 & n702 ) ;
  buffer buf_n760( .i (n476), .o (n760) );
  assign n761 = ~n759 & n760 ;
  assign n762 = ( n478 & n704 ) | ( n478 & ~n761 ) | ( n704 & ~n761 ) ;
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  assign n765 = ~n48 & n328 ;
  assign n766 = ( n269 & n763 ) | ( n269 & ~n765 ) | ( n763 & ~n765 ) ;
  assign n767 = n764 & ~n766 ;
  assign n768 = n521 & n767 ;
  assign n769 = ( n757 & n758 ) | ( n757 & n768 ) | ( n758 & n768 ) ;
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  assign n772 = ( n53 & n293 ) | ( n53 & ~n313 ) | ( n293 & ~n313 ) ;
  assign n773 = n770 & ~n772 ;
  assign n774 = ( n55 & n771 ) | ( n55 & ~n773 ) | ( n771 & ~n773 ) ;
  assign n775 = n283 & ~n303 ;
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n392( .i (n391), .o (n392) );
  assign n781 = n392 & n479 ;
  assign n782 = ( ~n289 & n780 ) | ( ~n289 & n781 ) | ( n780 & n781 ) ;
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  assign n785 = ( n73 & n521 ) | ( n73 & ~n783 ) | ( n521 & ~n783 ) ;
  assign n786 = n282 & n386 ;
  assign n787 = ( n303 & n744 ) | ( n303 & n786 ) | ( n744 & n786 ) ;
  assign n788 = ~n304 & n787 ;
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  assign n791 = n65 & ~n192 ;
  assign n792 = ( n131 & n163 ) | ( n131 & n791 ) | ( n163 & n791 ) ;
  assign n793 = ~n132 & n792 ;
  assign n794 = ( n46 & n789 ) | ( n46 & ~n793 ) | ( n789 & ~n793 ) ;
  assign n795 = ~n226 & n637 ;
  buffer buf_n796( .i (n795), .o (n796) );
  assign n800 = ~n282 & n302 ;
  buffer buf_n801( .i (n800), .o (n801) );
  assign n811 = ( n248 & n796 ) | ( n248 & n801 ) | ( n796 & n801 ) ;
  assign n812 = ~n249 & n811 ;
  assign n813 = ~n46 & n812 ;
  assign n814 = ( n790 & ~n794 ) | ( n790 & n813 ) | ( ~n794 & n813 ) ;
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  assign n817 = n227 | n303 ;
  assign n818 = ( ~n212 & n284 ) | ( ~n212 & n817 ) | ( n284 & n817 ) ;
  assign n819 = n213 | n818 ;
  assign n820 = n195 & ~n819 ;
  assign n821 = ( n134 & n149 ) | ( n134 & n820 ) | ( n149 & n820 ) ;
  assign n822 = ~n135 & n821 ;
  assign n823 = ~n815 & n822 ;
  assign n824 = n178 | n479 ;
  buffer buf_n825( .i (n824), .o (n825) );
  assign n826 = ( n816 & n823 ) | ( n816 & ~n825 ) | ( n823 & ~n825 ) ;
  buffer buf_n827( .i (n519), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  assign n829 = n826 & n828 ;
  assign n830 = ( n784 & n785 ) | ( n784 & n829 ) | ( n785 & n829 ) ;
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n273( .i (n272), .o (n273) );
  assign n833 = ( n53 & n273 ) | ( n53 & ~n333 ) | ( n273 & ~n333 ) ;
  assign n834 = n831 & ~n833 ;
  assign n835 = ( n55 & n832 ) | ( n55 & ~n834 ) | ( n832 & ~n834 ) ;
  assign n836 = n306 & n648 ;
  assign n837 = ~n231 & n836 ;
  assign n838 = ~n252 & n837 ;
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  assign n841 = ( n48 & ~n216 ) | ( n48 & n700 ) | ( ~n216 & n700 ) ;
  assign n842 = ~n49 & n841 ;
  assign n843 = ( n827 & ~n839 ) | ( n827 & n842 ) | ( ~n839 & n842 ) ;
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  assign n844 = ( n248 & n264 ) | ( n248 & ~n304 ) | ( n264 & ~n304 ) ;
  assign n845 = n661 & ~n844 ;
  assign n846 = ~n126 & n141 ;
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  assign n849 = ~n302 & n848 ;
  assign n850 = n263 & n849 ;
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  assign n853 = n45 & ~n851 ;
  assign n854 = ( n845 & n852 ) | ( n845 & ~n853 ) | ( n852 & ~n853 ) ;
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  assign n857 = ( n392 & n676 ) | ( n392 & ~n855 ) | ( n676 & ~n855 ) ;
  assign n858 = n856 & n857 ;
  assign n859 = n827 & n858 ;
  assign n860 = ( n840 & n843 ) | ( n840 & n859 ) | ( n843 & n859 ) ;
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  assign n863 = n50 & n152 ;
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  assign n868 = ( n292 & n332 ) | ( n292 & ~n864 ) | ( n332 & ~n864 ) ;
  assign n869 = n861 & n868 ;
  assign n870 = ( n862 & n866 ) | ( n862 & ~n869 ) | ( n866 & ~n869 ) ;
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  assign n872 = n123 & ~n276 ;
  assign n873 = ( n123 & n155 ) | ( n123 & n276 ) | ( n155 & n276 ) ;
  assign n874 = ~n256 & n276 ;
  assign n875 = ( n872 & n873 ) | ( n872 & ~n874 ) | ( n873 & ~n874 ) ;
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  assign n878 = ( n39 & n470 ) | ( n39 & n876 ) | ( n470 & n876 ) ;
  assign n879 = n139 & ~n257 ;
  assign n880 = ~n278 & n879 ;
  assign n881 = ~n470 & n880 ;
  assign n882 = ( n877 & ~n878 ) | ( n877 & n881 ) | ( ~n878 & n881 ) ;
  assign n883 = n225 & n882 ;
  assign n884 = ( n191 & n210 ) | ( n191 & n883 ) | ( n210 & n883 ) ;
  assign n885 = ~n192 & n884 ;
  assign n886 = ( n174 & ~n324 ) | ( n174 & n885 ) | ( ~n324 & n885 ) ;
  assign n887 = n261 & n472 ;
  assign n888 = ( n282 & n848 ) | ( n282 & n887 ) | ( n848 & n887 ) ;
  assign n889 = ~n283 & n888 ;
  assign n890 = ~n324 & n889 ;
  assign n891 = ( ~n175 & n886 ) | ( ~n175 & n890 ) | ( n886 & n890 ) ;
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  assign n894 = n42 | n262 ;
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  assign n898 = n284 & n475 ;
  assign n899 = ( n325 & n896 ) | ( n325 & n898 ) | ( n896 & n898 ) ;
  assign n900 = ~n897 & n899 ;
  assign n901 = ~n892 & n900 ;
  assign n902 = n69 & n391 ;
  assign n903 = ( n893 & n901 ) | ( n893 & n902 ) | ( n901 & n902 ) ;
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  assign n907 = n259 & ~n319 ;
  buffer buf_n908( .i (n907), .o (n908) );
  assign n917 = ( n281 & n847 ) | ( n281 & n908 ) | ( n847 & n908 ) ;
  buffer buf_n918( .i (n281), .o (n918) );
  assign n919 = n917 & ~n918 ;
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  assign n923 = ( n284 & ~n895 ) | ( n284 & n920 ) | ( ~n895 & n920 ) ;
  assign n924 = n325 & ~n923 ;
  assign n925 = ( n326 & n922 ) | ( n326 & ~n924 ) | ( n922 & ~n924 ) ;
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  assign n928 = ( n232 & n692 ) | ( n232 & n926 ) | ( n692 & n926 ) ;
  assign n929 = n927 & ~n928 ;
  assign n930 = ( ~n180 & n904 ) | ( ~n180 & n929 ) | ( n904 & n929 ) ;
  assign n931 = n200 & ~n930 ;
  assign n932 = ( n201 & n906 ) | ( n201 & ~n931 ) | ( n906 & ~n931 ) ;
  assign n933 = ( ~n313 & n865 ) | ( ~n313 & n932 ) | ( n865 & n932 ) ;
  assign n934 = n524 & ~n933 ;
  assign n935 = ( n525 & n867 ) | ( n525 & ~n934 ) | ( n867 & ~n934 ) ;
  assign n936 = ( n288 & n308 ) | ( n288 & n407 ) | ( n308 & n407 ) ;
  assign n937 = ( n288 & n308 ) | ( n288 & ~n479 ) | ( n308 & ~n479 ) ;
  assign n938 = n936 & ~n937 ;
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  assign n939 = ~n476 & n776 ;
  assign n940 = ( n176 & n798 ) | ( n176 & ~n939 ) | ( n798 & ~n939 ) ;
  assign n941 = n225 & n400 ;
  assign n942 = ( n302 & n918 ) | ( n302 & n941 ) | ( n918 & n941 ) ;
  assign n943 = ~n283 & n942 ;
  assign n944 = n65 & n211 ;
  assign n945 = ( n193 & n943 ) | ( n193 & n944 ) | ( n943 & n944 ) ;
  assign n946 = ~n194 & n945 ;
  assign n947 = ~n176 & n946 ;
  assign n948 = ( n799 & ~n940 ) | ( n799 & n947 ) | ( ~n940 & n947 ) ;
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  assign n951 = n71 | n949 ;
  assign n952 = ( n938 & n950 ) | ( n938 & n951 ) | ( n950 & n951 ) ;
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  assign n955 = ~n271 & n828 ;
  assign n956 = ( n332 & ~n953 ) | ( n332 & n955 ) | ( ~n953 & n955 ) ;
  assign n957 = n954 & n956 ;
  assign n958 = ~n54 & n957 ;
  assign n959 = ( n55 & ~n867 ) | ( n55 & n958 ) | ( ~n867 & n958 ) ;
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n960( .i (n478), .o (n960) );
  assign n961 = n407 & n960 ;
  assign n962 = ( ~n269 & n916 ) | ( ~n269 & n961 ) | ( n916 & n961 ) ;
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  assign n965 = ( n73 & n828 ) | ( n73 & ~n963 ) | ( n828 & ~n963 ) ;
  assign n966 = n62 & ~n159 ;
  assign n967 = ~n190 & n966 ;
  assign n968 = n401 & n967 ;
  assign n969 = ( n323 & ~n744 ) | ( n323 & n968 ) | ( ~n744 & n968 ) ;
  assign n970 = n745 & n969 ;
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n191), .o (n973) );
  buffer buf_n974( .i (n226), .o (n974) );
  assign n975 = n973 & ~n974 ;
  assign n976 = ( n212 & ~n324 ) | ( n212 & n975 ) | ( ~n324 & n975 ) ;
  assign n977 = ~n213 & n976 ;
  assign n978 = ~n971 & n977 ;
  assign n979 = n133 | n266 ;
  assign n980 = ( n972 & n978 ) | ( n972 & ~n979 ) | ( n978 & ~n979 ) ;
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  assign n983 = ~n326 & n798 ;
  assign n984 = ( n251 & n267 ) | ( n251 & n983 ) | ( n267 & n983 ) ;
  assign n985 = ~n252 & n984 ;
  assign n986 = ~n981 & n985 ;
  assign n987 = ( ~n825 & n982 ) | ( ~n825 & n986 ) | ( n982 & n986 ) ;
  assign n988 = n828 & n987 ;
  assign n989 = ( n964 & n965 ) | ( n964 & n988 ) | ( n965 & n988 ) ;
  assign n990 = n810 & n989 ;
  buffer buf_n991( .i (n52), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  assign n993 = n990 & ~n992 ;
  buffer buf_n994( .i (n992), .o (n994) );
  assign n995 = ( ~n867 & n993 ) | ( ~n867 & n994 ) | ( n993 & n994 ) ;
  assign n996 = ( n34 & n408 ) | ( n34 & n486 ) | ( n408 & n486 ) ;
  buffer buf_n423( .i (x25), .o (n423) );
  assign n997 = n423 & n486 ;
  assign n998 = ( ~n35 & n996 ) | ( ~n35 & n997 ) | ( n996 & n997 ) ;
  assign n999 = ( n36 & n58 ) | ( n36 & n998 ) | ( n58 & n998 ) ;
  assign n1000 = n468 & ~n999 ;
  assign n1001 = ( n38 & n469 ) | ( n38 & ~n1000 ) | ( n469 & ~n1000 ) ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n236( .i (x13), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  assign n1019 = n56 & ~n378 ;
  assign n1020 = ( n35 & n237 ) | ( n35 & n1019 ) | ( n237 & n1019 ) ;
  assign n1021 = ~n36 & n1020 ;
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n411( .i (n410), .o (n411) );
  assign n1024 = n411 & n489 ;
  assign n1025 = ( n469 & ~n1022 ) | ( n469 & n1024 ) | ( ~n1022 & n1024 ) ;
  assign n1026 = n1023 & n1025 ;
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  assign n1043 = ( n48 & n422 ) | ( n48 & n676 ) | ( n422 & n676 ) ;
  assign n1044 = ~n49 & n1043 ;
  assign n1045 = n502 & n1044 ;
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n118( .i (x5), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  assign n1051 = ( n118 & n378 ) | ( n118 & n465 ) | ( n378 & n465 ) ;
  assign n1052 = n505 & ~n1051 ;
  assign n1053 = ( n120 & n506 ) | ( n120 & ~n1052 ) | ( n506 & ~n1052 ) ;
  assign n1054 = ~n37 & n1053 ;
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n444( .i (x27), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  assign n1073 = ~n229 & n515 ;
  assign n1074 = ( n214 & ~n760 ) | ( n214 & n1073 ) | ( ~n760 & n1073 ) ;
  assign n1075 = ~n215 & n1074 ;
  buffer buf_n1076( .i (n47), .o (n1076) );
  assign n1077 = ( n700 & n1075 ) | ( n700 & n1076 ) | ( n1075 & n1076 ) ;
  assign n1078 = ~n49 & n1077 ;
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  assign n1082 = ( n111 & n463 ) | ( n111 & ~n1081 ) | ( n463 & ~n1081 ) ;
  buffer buf_n424( .i (x26), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  assign n1083 = n443 | n1081 ;
  assign n1084 = ( n464 & ~n1082 ) | ( n464 & n1083 ) | ( ~n1082 & n1083 ) ;
  assign n1085 = n994 | n1084 ;
  assign n1086 = ( ~n109 & n461 ) | ( ~n109 & n1079 ) | ( n461 & n1079 ) ;
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  assign n1089 = ( n110 & n442 ) | ( n110 & n1080 ) | ( n442 & n1080 ) ;
  assign n1090 = n1087 | n1089 ;
  assign n1091 = ( ~n464 & n1088 ) | ( ~n464 & n1090 ) | ( n1088 & n1090 ) ;
  assign n1092 = n994 | n1091 ;
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n217( .i (n216), .o (n217) );
  assign n1093 = ( n198 & ~n217 ) | ( n198 & n600 ) | ( ~n217 & n600 ) ;
  assign n1094 = n234 & ~n1093 ;
  assign n1095 = ( n235 & n602 ) | ( n235 & ~n1094 ) | ( n602 & ~n1094 ) ;
  buffer buf_n1096( .i (n225), .o (n1096) );
  assign n1097 = ( n342 & n356 ) | ( n342 & ~n1096 ) | ( n356 & ~n1096 ) ;
  assign n1098 = ( n342 & n372 ) | ( n342 & n1096 ) | ( n372 & n1096 ) ;
  assign n1099 = n1097 & n1098 ;
  assign n1100 = n174 & ~n1099 ;
  assign n1101 = n373 & n974 ;
  buffer buf_n1102( .i (n173), .o (n1102) );
  assign n1103 = n1101 | n1102 ;
  assign n1104 = ~n1100 & n1103 ;
  assign n1105 = n498 & n1104 ;
  assign n1106 = n196 & ~n1105 ;
  assign n1107 = n176 | n230 ;
  assign n1108 = ~n196 & n1107 ;
  assign n1109 = n1106 | n1108 ;
  assign n1110 = n217 & ~n1109 ;
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  assign n1113 = n181 | n1111 ;
  assign n1114 = ( n1095 & n1112 ) | ( n1095 & n1113 ) | ( n1112 & n1113 ) ;
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  assign n1117 = ( n485 & ~n633 ) | ( n485 & n1115 ) | ( ~n633 & n1115 ) ;
  assign n1118 = n1116 & ~n1117 ;
  buffer buf_n74( .i (x2), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n1119( .i (n827), .o (n1119) );
  assign n1120 = ( n91 & n503 ) | ( n91 & ~n1119 ) | ( n503 & ~n1119 ) ;
  assign n1121 = ( n109 & n503 ) | ( n109 & n1119 ) | ( n503 & n1119 ) ;
  assign n1122 = n1120 & ~n1121 ;
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n1125( .i (n495), .o (n1125) );
  assign n1126 = n374 & n1125 ;
  buffer buf_n1127( .i (n210), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  assign n1130 = ( ~n609 & n1126 ) | ( ~n609 & n1129 ) | ( n1126 & n1129 ) ;
  assign n1131 = n360 & n1130 ;
  assign n1132 = ( n196 & n347 ) | ( n196 & n1131 ) | ( n347 & n1131 ) ;
  assign n1133 = ~n197 & n1132 ;
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n1136( .i (n974), .o (n1136) );
  assign n1137 = ( ~n193 & n1128 ) | ( ~n193 & n1136 ) | ( n1128 & n1136 ) ;
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  assign n1142 = n230 & ~n1138 ;
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  assign n1145 = n345 & n497 ;
  buffer buf_n1146( .i (n1145), .o (n1146) );
  assign n1149 = n377 & n1146 ;
  assign n1150 = ( n216 & n1143 ) | ( n216 & n1149 ) | ( n1143 & n1149 ) ;
  assign n1151 = ( ~n1141 & n1144 ) | ( ~n1141 & n1150 ) | ( n1144 & n1150 ) ;
  assign n1152 = n1125 & n1136 ;
  assign n1153 = n375 & n1152 ;
  assign n1154 = n214 & n1153 ;
  buffer buf_n1155( .i (n195), .o (n1155) );
  assign n1156 = ( n177 & n1154 ) | ( n177 & n1155 ) | ( n1154 & n1155 ) ;
  assign n1157 = ~n178 & n1156 ;
  buffer buf_n1158( .i (n1157), .o (n1158) );
  assign n1159 = ( ~n1134 & n1151 ) | ( ~n1134 & n1158 ) | ( n1151 & n1158 ) ;
  assign n1160 = n180 | n1158 ;
  assign n1161 = ( n1135 & n1159 ) | ( n1135 & n1160 ) | ( n1159 & n1160 ) ;
  assign n1162 = n522 & ~n1161 ;
  assign n1163 = n109 & ~n503 ;
  assign n1164 = n522 | n1163 ;
  assign n1165 = ~n1162 & n1164 ;
  assign n1166 = ( n992 & ~n1123 ) | ( n992 & n1165 ) | ( ~n1123 & n1165 ) ;
  assign n1167 = n485 & ~n992 ;
  assign n1168 = ( n1124 & n1166 ) | ( n1124 & ~n1167 ) | ( n1166 & ~n1167 ) ;
  assign n1169 = ( n111 & ~n484 ) | ( n111 & n523 ) | ( ~n484 & n523 ) ;
  buffer buf_n182( .i (n181), .o (n182) );
  assign n1170 = n354 & n492 ;
  assign n1171 = n371 & n1170 ;
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  assign n1174 = n172 & n342 ;
  assign n1175 = ( n974 & ~n1172 ) | ( n974 & n1174 ) | ( ~n1172 & n1174 ) ;
  assign n1176 = n1173 & n1175 ;
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n175), .o (n1180) );
  assign n1181 = ( n230 & ~n1177 ) | ( n230 & n1180 ) | ( ~n1177 & n1180 ) ;
  buffer buf_n1182( .i (n214), .o (n1182) );
  assign n1183 = n1181 & n1182 ;
  buffer buf_n1184( .i (n1182), .o (n1184) );
  assign n1185 = ( n1179 & ~n1183 ) | ( n1179 & n1184 ) | ( ~n1183 & n1184 ) ;
  buffer buf_n1186( .i (n197), .o (n1186) );
  assign n1187 = n1185 & ~n1186 ;
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  assign n1190 = ~n210 & n1096 ;
  buffer buf_n1191( .i (n1190), .o (n1191) );
  assign n1194 = n1136 & ~n1191 ;
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n194), .o (n1196) );
  assign n1197 = n1195 & n1196 ;
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  assign n1198 = ( n376 & ~n1193 ) | ( n376 & n1195 ) | ( ~n1193 & n1195 ) ;
  assign n1199 = ( ~n1182 & n1197 ) | ( ~n1182 & n1198 ) | ( n1197 & n1198 ) ;
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  assign n1202 = ( n363 & n1148 ) | ( n363 & ~n1200 ) | ( n1148 & ~n1200 ) ;
  assign n1203 = n1201 & n1202 ;
  assign n1204 = n1188 | n1203 ;
  assign n1205 = ( n182 & n1189 ) | ( n182 & n1204 ) | ( n1189 & n1204 ) ;
  assign n1206 = ( n484 & n523 ) | ( n484 & ~n1205 ) | ( n523 & ~n1205 ) ;
  assign n1207 = n1169 & ~n1206 ;
  assign n1208 = ~n994 & n1207 ;
  assign n1209 = n173 & n1127 ;
  buffer buf_n1210( .i (n973), .o (n1210) );
  assign n1211 = ( n44 & n1209 ) | ( n44 & n1210 ) | ( n1209 & n1210 ) ;
  assign n1212 = ~n45 & n1211 ;
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n229), .o (n1215) );
  assign n1216 = n360 & n1215 ;
  assign n1217 = ( n347 & ~n1213 ) | ( n347 & n1216 ) | ( ~n1213 & n1216 ) ;
  assign n1218 = n1214 & n1217 ;
  buffer buf_n1219( .i (n518), .o (n1219) );
  assign n1220 = n1218 & n1219 ;
  assign n1221 = ( n481 & n502 ) | ( n481 & n1220 ) | ( n502 & n1220 ) ;
  assign n1222 = ~n482 & n1221 ;
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  assign y0 = n558 ;
  assign y1 = n581 ;
  assign y2 = n584 ;
  assign y3 = n591 ;
  assign y4 = n635 ;
  assign y5 = n684 ;
  assign y6 = n741 ;
  assign y7 = n774 ;
  assign y8 = n835 ;
  assign y9 = n871 ;
  assign y10 = n935 ;
  assign y11 = n959 ;
  assign y12 = n995 ;
  assign y13 = n1018 ;
  assign y14 = n1042 ;
  assign y15 = n1050 ;
  assign y16 = n1072 ;
  assign y17 = n1085 ;
  assign y18 = n1092 ;
  assign y19 = n1118 ;
  assign y20 = n1168 ;
  assign y21 = n1208 ;
  assign y22 = n1226 ;
endmodule
