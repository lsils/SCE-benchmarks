module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( in_6_ , in_15_ , in_13_ , in_14_ , in_2_ , in_10_ , in_24_ , in_8_ , in_22_ , in_20_ , in_7_ , in_25_ , in_5_ , in_4_ , in_23_ , in_27_ , in_1_ , in_0_ , in_16_ , in_30_ , in_26_ , in_12_ , in_11_ , in_17_ , in_19_ , in_18_ , in_21_ , in_31_ , in_29_ , in_28_ , in_9_ , in_3_ , out_2_ , out_1_ , out_3_ , out_0_ , out_5_ , out_4_ );
  input in_6_ , in_15_ , in_13_ , in_14_ , in_2_ , in_10_ , in_24_ , in_8_ , in_22_ , in_20_ , in_7_ , in_25_ , in_5_ , in_4_ , in_23_ , in_27_ , in_1_ , in_0_ , in_16_ , in_30_ , in_26_ , in_12_ , in_11_ , in_17_ , in_19_ , in_18_ , in_21_ , in_31_ , in_29_ , in_28_ , in_9_ , in_3_ ;
  output out_2_ , out_1_ , out_3_ , out_0_ , out_5_ , out_4_ ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 ;
  assign n33 = in_29_ | in_28_ ;
  buffer buf_n34( .i (n33), .o (n34) );
  assign n37 = in_20_ | in_21_ ;
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  assign n41 = in_16_ | in_17_ ;
  buffer buf_n42( .i (n41), .o (n42) );
  assign n43 = in_19_ & in_18_ ;
  buffer buf_n44( .i (n43), .o (n44) );
  assign n45 = ( n38 & n42 ) | ( n38 & n44 ) | ( n42 & n44 ) ;
  buffer buf_n46( .i (n45), .o (n46) );
  assign n51 = ( ~n38 & n42 ) | ( ~n38 & n44 ) | ( n42 & n44 ) ;
  buffer buf_n52( .i (n51), .o (n52) );
  assign n53 = ( n40 & ~n46 ) | ( n40 & n52 ) | ( ~n46 & n52 ) ;
  buffer buf_n54( .i (n53), .o (n54) );
  assign n55 = in_27_ & in_26_ ;
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  assign n59 = in_22_ & in_23_ ;
  buffer buf_n60( .i (n59), .o (n60) );
  assign n61 = in_24_ | in_25_ ;
  buffer buf_n62( .i (n61), .o (n62) );
  assign n63 = ( n56 & n60 ) | ( n56 & n62 ) | ( n60 & n62 ) ;
  buffer buf_n64( .i (n63), .o (n64) );
  assign n69 = ( ~n56 & n60 ) | ( ~n56 & n62 ) | ( n60 & n62 ) ;
  buffer buf_n70( .i (n69), .o (n70) );
  assign n71 = ( n58 & ~n64 ) | ( n58 & n70 ) | ( ~n64 & n70 ) ;
  buffer buf_n72( .i (n71), .o (n72) );
  assign n73 = ( n34 & n54 ) | ( n34 & n72 ) | ( n54 & n72 ) ;
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  assign n77 = ( n50 & n68 ) | ( n50 & n74 ) | ( n68 & n74 ) ;
  buffer buf_n78( .i (n77), .o (n78) );
  assign n83 = ( n50 & n68 ) | ( n50 & ~n74 ) | ( n68 & ~n74 ) ;
  buffer buf_n84( .i (n83), .o (n84) );
  assign n85 = ( n76 & ~n78 ) | ( n76 & n84 ) | ( ~n78 & n84 ) ;
  buffer buf_n86( .i (n85), .o (n86) );
  assign n87 = in_30_ & in_31_ ;
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  assign n89 = ( ~n34 & n54 ) | ( ~n34 & n72 ) | ( n54 & n72 ) ;
  buffer buf_n90( .i (n89), .o (n90) );
  assign n91 = ( n36 & ~n74 ) | ( n36 & n90 ) | ( ~n74 & n90 ) ;
  buffer buf_n92( .i (n91), .o (n92) );
  assign n93 = n88 & n92 ;
  buffer buf_n94( .i (n93), .o (n94) );
  assign n95 = n86 & n94 ;
  buffer buf_n96( .i (n95), .o (n96) );
  assign n97 = n86 | n94 ;
  buffer buf_n98( .i (n97), .o (n98) );
  assign n99 = ~n96 & n98 ;
  buffer buf_n100( .i (n99), .o (n100) );
  assign n101 = in_13_ | in_12_ ;
  buffer buf_n102( .i (n101), .o (n102) );
  assign n105 = in_5_ | in_4_ ;
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  assign n109 = in_1_ | in_0_ ;
  buffer buf_n110( .i (n109), .o (n110) );
  assign n111 = in_2_ & in_3_ ;
  buffer buf_n112( .i (n111), .o (n112) );
  assign n113 = ( n106 & n110 ) | ( n106 & n112 ) | ( n110 & n112 ) ;
  buffer buf_n114( .i (n113), .o (n114) );
  assign n119 = ( ~n106 & n110 ) | ( ~n106 & n112 ) | ( n110 & n112 ) ;
  buffer buf_n120( .i (n119), .o (n120) );
  assign n121 = ( n108 & ~n114 ) | ( n108 & n120 ) | ( ~n114 & n120 ) ;
  buffer buf_n122( .i (n121), .o (n122) );
  assign n123 = in_10_ & in_11_ ;
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  assign n127 = in_6_ & in_7_ ;
  buffer buf_n128( .i (n127), .o (n128) );
  assign n129 = in_8_ | in_9_ ;
  buffer buf_n130( .i (n129), .o (n130) );
  assign n131 = ( n124 & n128 ) | ( n124 & n130 ) | ( n128 & n130 ) ;
  buffer buf_n132( .i (n131), .o (n132) );
  assign n137 = ( ~n124 & n128 ) | ( ~n124 & n130 ) | ( n128 & n130 ) ;
  buffer buf_n138( .i (n137), .o (n138) );
  assign n139 = ( n126 & ~n132 ) | ( n126 & n138 ) | ( ~n132 & n138 ) ;
  buffer buf_n140( .i (n139), .o (n140) );
  assign n141 = ( n102 & n122 ) | ( n102 & n140 ) | ( n122 & n140 ) ;
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  assign n145 = ( n118 & n136 ) | ( n118 & n142 ) | ( n136 & n142 ) ;
  buffer buf_n146( .i (n145), .o (n146) );
  assign n151 = ( n118 & n136 ) | ( n118 & ~n142 ) | ( n136 & ~n142 ) ;
  buffer buf_n152( .i (n151), .o (n152) );
  assign n153 = ( n144 & ~n146 ) | ( n144 & n152 ) | ( ~n146 & n152 ) ;
  buffer buf_n154( .i (n153), .o (n154) );
  assign n155 = in_15_ & in_14_ ;
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  assign n157 = ( ~n102 & n122 ) | ( ~n102 & n140 ) | ( n122 & n140 ) ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n159 = ( n104 & ~n142 ) | ( n104 & n158 ) | ( ~n142 & n158 ) ;
  buffer buf_n160( .i (n159), .o (n160) );
  assign n161 = n156 & n160 ;
  buffer buf_n162( .i (n161), .o (n162) );
  assign n163 = n154 & n162 ;
  buffer buf_n164( .i (n163), .o (n164) );
  assign n165 = n154 | n162 ;
  buffer buf_n166( .i (n165), .o (n166) );
  assign n167 = ~n164 & n166 ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = n100 & n168 ;
  assign n170 = n100 | n168 ;
  assign n171 = ~n169 & n170 ;
  buffer buf_n172( .i (n171), .o (n172) );
  assign n173 = n88 | n92 ;
  buffer buf_n174( .i (n173), .o (n174) );
  assign n175 = ~n94 & n174 ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n177 = n156 | n160 ;
  buffer buf_n178( .i (n177), .o (n178) );
  assign n179 = ~n162 & n178 ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = n176 & n180 ;
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  assign n186 = n172 & n185 ;
  assign n187 = n172 | n185 ;
  assign n188 = ~n186 & n187 ;
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  assign n191 = n176 | n180 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = ~n182 & n192 ;
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  assign n200 = n82 & n96 ;
  buffer buf_n201( .i (n200), .o (n201) );
  assign n206 = n82 | n96 ;
  buffer buf_n207( .i (n206), .o (n207) );
  assign n208 = ~n201 & n207 ;
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  assign n210 = n150 & n164 ;
  buffer buf_n211( .i (n210), .o (n211) );
  assign n216 = n150 | n164 ;
  buffer buf_n217( .i (n216), .o (n217) );
  assign n218 = ~n211 & n217 ;
  buffer buf_n219( .i (n218), .o (n219) );
  assign n220 = n209 & n219 ;
  assign n221 = n209 | n219 ;
  assign n222 = ~n220 & n221 ;
  buffer buf_n223( .i (n222), .o (n223) );
  assign n224 = ( n100 & n168 ) | ( n100 & n182 ) | ( n168 & n182 ) ;
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  assign n229 = n223 & n228 ;
  assign n230 = n223 | n228 ;
  assign n231 = ~n229 & n230 ;
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  assign n232 = ( n209 & n219 ) | ( n209 & n225 ) | ( n219 & n225 ) ;
  buffer buf_n233( .i (n232), .o (n233) );
  assign n234 = ( n205 & n215 ) | ( n205 & n233 ) | ( n215 & n233 ) ;
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  assign n237 = n201 | n211 ;
  assign n238 = n201 & n211 ;
  assign n239 = n237 & ~n238 ;
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  assign n242 = n233 & n241 ;
  assign n243 = n233 | n241 ;
  assign n244 = ~n242 & n243 ;
  buffer buf_n245( .i (n244), .o (n245) );
  assign out_2_ = n190 ;
  assign out_1_ = n199 ;
  assign out_3_ = n231 ;
  assign out_0_ = 1'b0 ;
  assign out_5_ = n236 ;
  assign out_4_ = n245 ;
endmodule
