module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( N1 , N102 , N105 , N108 , N11 , N112 , N115 , N14 , N17 , N21 , N24 , N27 , N30 , N34 , N37 , N4 , N40 , N43 , N47 , N50 , N53 , N56 , N60 , N63 , N66 , N69 , N73 , N76 , N79 , N8 , N82 , N86 , N89 , N92 , N95 , N99 , N223 , N329 , N370 , N421 , N430 , N431 , N432 );
  input N1 , N102 , N105 , N108 , N11 , N112 , N115 , N14 , N17 , N21 , N24 , N27 , N30 , N34 , N37 , N4 , N40 , N43 , N47 , N50 , N53 , N56 , N60 , N63 , N66 , N69 , N73 , N76 , N79 , N8 , N82 , N86 , N89 , N92 , N95 , N99 ;
  output N223 , N329 , N370 , N421 , N430 , N431 , N432 ;
  wire n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 ;
  assign n37 = ~N24 & N30 ;
  buffer buf_n38( .i (n37), .o (n38) );
  assign n44 = ~N102 & N108 ;
  assign n45 = n38 | n44 ;
  assign n46 = ~N1 & N4 ;
  assign n47 = ~N89 & N95 ;
  assign n48 = ~N76 & N82 ;
  assign n49 = n47 | n48 ;
  assign n50 = n46 | n49 ;
  assign n51 = ~N63 & N69 ;
  buffer buf_n52( .i (n51), .o (n52) );
  assign n59 = ~N37 & N43 ;
  assign n60 = n52 | n59 ;
  assign n61 = ~N50 & N56 ;
  assign n62 = ~N11 & N17 ;
  assign n63 = n61 | n62 ;
  assign n64 = n60 | n63 ;
  assign n65 = n50 | n64 ;
  assign n66 = n45 | n65 ;
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n120( .i (n67), .o (n120) );
  buffer buf_n68( .i (n67), .o (n68) );
  assign n69 = N102 & n68 ;
  assign n70 = N108 & ~n69 ;
  buffer buf_n71( .i (n70), .o (n71) );
  assign n79 = ~N112 & n71 ;
  assign n80 = N76 & n68 ;
  assign n81 = N82 & ~n80 ;
  buffer buf_n82( .i (n81), .o (n82) );
  assign n91 = ~N86 & n82 ;
  assign n92 = n79 | n91 ;
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  assign n93 = N30 & ~n68 ;
  assign n94 = n43 | n93 ;
  buffer buf_n95( .i (n94), .o (n95) );
  assign n105 = ~N34 & n95 ;
  assign n106 = N11 & n68 ;
  assign n107 = N17 & ~n106 ;
  buffer buf_n108( .i (n107), .o (n108) );
  assign n117 = ~N21 & n108 ;
  assign n118 = n105 | n117 ;
  assign n119 = n92 | n118 ;
  assign n121 = N1 & n120 ;
  assign n122 = N4 & ~n121 ;
  buffer buf_n123( .i (n122), .o (n123) );
  assign n132 = ~N8 & n123 ;
  assign n133 = N89 & n120 ;
  assign n134 = N95 & ~n133 ;
  buffer buf_n135( .i (n134), .o (n135) );
  assign n144 = ~N99 & n135 ;
  assign n145 = n132 | n144 ;
  assign n146 = N50 & n120 ;
  assign n147 = N56 & ~n146 ;
  buffer buf_n148( .i (n147), .o (n148) );
  assign n155 = ~N60 & n148 ;
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  assign n156 = N69 & ~n67 ;
  assign n157 = n58 | n156 ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n167 = ~N73 & n158 ;
  assign n168 = N37 & n67 ;
  assign n169 = N43 & ~n168 ;
  buffer buf_n170( .i (n169), .o (n170) );
  assign n179 = ~N47 & n170 ;
  assign n180 = n167 | n179 ;
  assign n181 = n155 | n180 ;
  assign n182 = n145 | n181 ;
  assign n183 = n119 | n182 ;
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  assign n188 = N34 & n187 ;
  assign n189 = n104 & ~n188 ;
  buffer buf_n190( .i (n189), .o (n190) );
  assign n197 = ~N40 & n190 ;
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  assign n198 = N99 & n186 ;
  assign n199 = n143 & ~n198 ;
  buffer buf_n200( .i (n199), .o (n200) );
  assign n209 = ~N105 & n200 ;
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  assign n210 = N21 & n186 ;
  assign n211 = n116 & ~n210 ;
  buffer buf_n212( .i (n211), .o (n212) );
  assign n220 = ~N27 & n212 ;
  assign n221 = n209 | n220 ;
  assign n222 = n197 | n221 ;
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  assign n223 = N8 & n186 ;
  assign n224 = n131 & ~n223 ;
  buffer buf_n225( .i (n224), .o (n225) );
  assign n239 = ~N14 & n225 ;
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n240( .i (n185), .o (n240) );
  assign n241 = N86 & n240 ;
  assign n242 = n90 & ~n241 ;
  buffer buf_n243( .i (n242), .o (n243) );
  assign n252 = ~N92 & n243 ;
  assign n253 = n239 | n252 ;
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  assign n254 = N73 & n185 ;
  assign n255 = n166 & ~n254 ;
  buffer buf_n256( .i (n255), .o (n256) );
  assign n266 = ~N79 & n256 ;
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  assign n267 = N60 & n184 ;
  assign n268 = n154 & ~n267 ;
  buffer buf_n269( .i (n268), .o (n269) );
  assign n279 = ~N66 & n269 ;
  buffer buf_n280( .i (n279), .o (n280) );
  assign n289 = n266 | n280 ;
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  assign n290 = N47 & n185 ;
  assign n291 = n178 & ~n290 ;
  buffer buf_n292( .i (n291), .o (n292) );
  assign n301 = ~N53 & n292 ;
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n302( .i (n184), .o (n302) );
  assign n303 = N112 & n302 ;
  assign n304 = n78 & ~n303 ;
  buffer buf_n305( .i (n304), .o (n305) );
  assign n317 = ~N115 & n305 ;
  assign n318 = n301 | n317 ;
  assign n319 = n289 | n318 ;
  assign n320 = n253 | n319 ;
  assign n321 = n222 | n320 ;
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n323( .i (n322), .o (n323) );
  assign n330 = N40 & n323 ;
  assign n331 = n196 & ~n330 ;
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  assign n337 = N27 & n323 ;
  assign n338 = n219 & ~n337 ;
  buffer buf_n339( .i (n338), .o (n339) );
  assign n345 = n332 | n339 ;
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  assign n349 = N53 & n323 ;
  assign n350 = n300 & ~n349 ;
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n324( .i (n323), .o (n324) );
  assign n354 = n278 & ~n324 ;
  assign n355 = n288 | n354 ;
  assign n356 = n351 | n355 ;
  buffer buf_n357( .i (n356), .o (n357) );
  assign n359 = n346 | n357 ;
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  assign n361 = N92 & n324 ;
  assign n362 = n251 & ~n361 ;
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  assign n364 = N79 & n324 ;
  assign n365 = n265 & ~n364 ;
  buffer buf_n366( .i (n365), .o (n366) );
  assign n368 = n363 | n366 ;
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n370( .i (n322), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  assign n372 = N105 & n371 ;
  assign n373 = n208 & ~n372 ;
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  assign n376 = N115 & n326 ;
  assign n377 = n316 & ~n376 ;
  assign n378 = n375 | n377 ;
  assign n379 = n369 | n378 ;
  assign n380 = n360 | n379 ;
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  assign n381 = N14 & n329 ;
  assign n382 = n238 & ~n381 ;
  assign n383 = n380 & ~n382 ;
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n358( .i (n357), .o (n358) );
  assign n384 = ~n358 & n369 ;
  assign n385 = n348 | n384 ;
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n367( .i (n366), .o (n367) );
  assign n386 = ~n357 & n367 ;
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  assign n387 = ~n363 & n374 ;
  assign n388 = n353 | n387 ;
  assign n389 = n386 | n388 ;
  assign n390 = ~n336 & n389 ;
  assign n391 = n344 | n390 ;
  assign N223 = n120 ;
  assign N329 = n184 ;
  assign N370 = n322 ;
  assign N421 = n383 ;
  assign N430 = n360 ;
  assign N431 = n385 ;
  assign N432 = n391 ;
endmodule
