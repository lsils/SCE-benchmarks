module top( in_15_ , in_0_ , in_4_ , in_29_ , in_38_ , in_53_ , in_42_ , in_11_ , in_59_ , in_48_ , in_54_ , in_16_ , in_43_ , in_37_ , in_61_ , in_14_ , in_62_ , in_60_ , in_40_ , in_5_ , in_28_ , in_7_ , in_6_ , in_34_ , in_57_ , in_3_ , in_56_ , in_45_ , in_10_ , in_27_ , in_21_ , in_25_ , in_22_ , in_12_ , in_58_ , in_36_ , in_51_ , in_18_ , in_9_ , in_39_ , in_24_ , in_26_ , in_8_ , in_41_ , in_55_ , in_2_ , in_49_ , in_19_ , in_35_ , in_50_ , in_32_ , in_30_ , in_33_ , in_17_ , in_31_ , in_44_ , in_1_ , in_23_ , in_52_ , in_20_ , in_46_ , in_13_ , in_63_ , in_47_ , out_1_ , out_3_ , out_6_ , out_2_ , out_0_ , out_4_ , out_5_ );
  input in_15_ , in_0_ , in_4_ , in_29_ , in_38_ , in_53_ , in_42_ , in_11_ , in_59_ , in_48_ , in_54_ , in_16_ , in_43_ , in_37_ , in_61_ , in_14_ , in_62_ , in_60_ , in_40_ , in_5_ , in_28_ , in_7_ , in_6_ , in_34_ , in_57_ , in_3_ , in_56_ , in_45_ , in_10_ , in_27_ , in_21_ , in_25_ , in_22_ , in_12_ , in_58_ , in_36_ , in_51_ , in_18_ , in_9_ , in_39_ , in_24_ , in_26_ , in_8_ , in_41_ , in_55_ , in_2_ , in_49_ , in_19_ , in_35_ , in_50_ , in_32_ , in_30_ , in_33_ , in_17_ , in_31_ , in_44_ , in_1_ , in_23_ , in_52_ , in_20_ , in_46_ , in_13_ , in_63_ , in_47_ ;
  output out_1_ , out_3_ , out_6_ , out_2_ , out_0_ , out_4_ , out_5_ ;
  wire n65 , n75 , n83 , n87 , n89 , n91 , n97 , n99 , n101 , n105 , n107 , n109 , n115 , n117 , n119 , n123 , n125 , n127 , n129 , n131 , n133 , n143 , n151 , n155 , n157 , n159 , n165 , n167 , n169 , n173 , n175 , n177 , n183 , n185 , n187 , n191 , n193 , n195 , n197 , n199 , n201 , n206 , n208 , n210 , n220 , n228 , n232 , n234 , n236 , n242 , n244 , n246 , n250 , n252 , n254 , n260 , n262 , n264 , n268 , n270 , n272 , n274 , n276 , n278 , n288 , n296 , n300 , n302 , n304 , n310 , n312 , n314 , n318 , n320 , n322 , n328 , n330 , n332 , n336 , n338 , n340 , n342 , n344 , n346 , n351 , n353 , n355 , n362 , n364 , n374 , n380 , n382 , n384 , n386 , n392 , n394 , n396 , n402 , n404 , n406 , n408 , n414 , n416 , n418 , n419 , n420 , n422 , n424 , n426 , n428 , n430 , n435 , n436 , n437 , n439 , n445 , n447 , n449 , n451 , n457 , n459 , n461 , n467 , n469 , n471 , n473 , n479 , n481 , n483 , n484 , n485 , n487 , n489 , n491 , n493 , n495 , n500 , n501 , n502 , n504 , n505 , n506 , n508 , n509 , n510 , n512 , n513 , n514 , n516 , n517 , n518 , n520 , n521 , n522 , n524 , n529 , n530 , n531 , n533 , n535 , n543 , n545 , n553 , n554 , n555 , n557 , n558 , n559 , n564 , n565 , n566 , n568 , n569 , n570 , n575 , n577 , n579 , n581 , n582 , n583 , n585 , n586 , n587 , n591 , n592 , n593 , n595 , n596 , n597 , n600 , n601 , n602 , n604 , n605 , n606 ;
  assign n65 = in_15_ & in_14_ ;
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  assign n75 = in_12_ | in_13_ ;
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  assign n83 = in_4_ | in_5_ ;
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  assign n87 = in_0_ | in_1_ ;
  buffer buf_n88( .i (n87), .o (n88) );
  assign n89 = in_3_ & in_2_ ;
  buffer buf_n90( .i (n89), .o (n90) );
  assign n91 = ( n84 & n88 ) | ( n84 & n90 ) | ( n88 & n90 ) ;
  buffer buf_n92( .i (n91), .o (n92) );
  assign n97 = ( ~n84 & n88 ) | ( ~n84 & n90 ) | ( n88 & n90 ) ;
  buffer buf_n98( .i (n97), .o (n98) );
  assign n99 = ( n86 & ~n92 ) | ( n86 & n98 ) | ( ~n92 & n98 ) ;
  buffer buf_n100( .i (n99), .o (n100) );
  assign n101 = in_11_ & in_10_ ;
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  assign n105 = in_7_ & in_6_ ;
  buffer buf_n106( .i (n105), .o (n106) );
  assign n107 = in_9_ | in_8_ ;
  buffer buf_n108( .i (n107), .o (n108) );
  assign n109 = ( n102 & n106 ) | ( n102 & n108 ) | ( n106 & n108 ) ;
  buffer buf_n110( .i (n109), .o (n110) );
  assign n115 = ( ~n102 & n106 ) | ( ~n102 & n108 ) | ( n106 & n108 ) ;
  buffer buf_n116( .i (n115), .o (n116) );
  assign n117 = ( n104 & ~n110 ) | ( n104 & n116 ) | ( ~n110 & n116 ) ;
  buffer buf_n118( .i (n117), .o (n118) );
  assign n119 = ( n80 & n100 ) | ( n80 & n118 ) | ( n100 & n118 ) ;
  buffer buf_n120( .i (n119), .o (n120) );
  assign n123 = ( ~n80 & n100 ) | ( ~n80 & n118 ) | ( n100 & n118 ) ;
  buffer buf_n124( .i (n123), .o (n124) );
  assign n125 = ( n82 & ~n120 ) | ( n82 & n124 ) | ( ~n120 & n124 ) ;
  buffer buf_n126( .i (n125), .o (n126) );
  assign n127 = n74 & n126 ;
  buffer buf_n128( .i (n127), .o (n128) );
  assign n129 = n74 | n126 ;
  buffer buf_n130( .i (n129), .o (n130) );
  assign n131 = ~n128 & n130 ;
  buffer buf_n132( .i (n131), .o (n132) );
  assign n133 = in_30_ & in_31_ ;
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  assign n143 = in_29_ | in_28_ ;
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  assign n151 = in_21_ | in_20_ ;
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  assign n155 = in_16_ | in_17_ ;
  buffer buf_n156( .i (n155), .o (n156) );
  assign n157 = in_18_ & in_19_ ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n159 = ( n152 & n156 ) | ( n152 & n158 ) | ( n156 & n158 ) ;
  buffer buf_n160( .i (n159), .o (n160) );
  assign n165 = ( ~n152 & n156 ) | ( ~n152 & n158 ) | ( n156 & n158 ) ;
  buffer buf_n166( .i (n165), .o (n166) );
  assign n167 = ( n154 & ~n160 ) | ( n154 & n166 ) | ( ~n160 & n166 ) ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = in_27_ & in_26_ ;
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  assign n173 = in_22_ & in_23_ ;
  buffer buf_n174( .i (n173), .o (n174) );
  assign n175 = in_25_ | in_24_ ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n177 = ( n170 & n174 ) | ( n170 & n176 ) | ( n174 & n176 ) ;
  buffer buf_n178( .i (n177), .o (n178) );
  assign n183 = ( ~n170 & n174 ) | ( ~n170 & n176 ) | ( n174 & n176 ) ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n185 = ( n172 & ~n178 ) | ( n172 & n184 ) | ( ~n178 & n184 ) ;
  buffer buf_n186( .i (n185), .o (n186) );
  assign n187 = ( n148 & n168 ) | ( n148 & n186 ) | ( n168 & n186 ) ;
  buffer buf_n188( .i (n187), .o (n188) );
  assign n191 = ( ~n148 & n168 ) | ( ~n148 & n186 ) | ( n168 & n186 ) ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = ( n150 & ~n188 ) | ( n150 & n192 ) | ( ~n188 & n192 ) ;
  buffer buf_n194( .i (n193), .o (n194) );
  assign n195 = n142 & n194 ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n197 = n142 | n194 ;
  buffer buf_n198( .i (n197), .o (n198) );
  assign n199 = ~n196 & n198 ;
  buffer buf_n200( .i (n199), .o (n200) );
  assign n201 = n132 & n200 ;
  buffer buf_n202( .i (n201), .o (n202) );
  assign n206 = n132 | n200 ;
  buffer buf_n207( .i (n206), .o (n207) );
  assign n208 = ~n202 & n207 ;
  buffer buf_n209( .i (n208), .o (n209) );
  assign n210 = in_46_ & in_47_ ;
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  assign n220 = in_45_ | in_44_ ;
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  assign n228 = in_37_ | in_36_ ;
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  assign n232 = in_32_ | in_33_ ;
  buffer buf_n233( .i (n232), .o (n233) );
  assign n234 = in_34_ & in_35_ ;
  buffer buf_n235( .i (n234), .o (n235) );
  assign n236 = ( n229 & n233 ) | ( n229 & n235 ) | ( n233 & n235 ) ;
  buffer buf_n237( .i (n236), .o (n237) );
  assign n242 = ( ~n229 & n233 ) | ( ~n229 & n235 ) | ( n233 & n235 ) ;
  buffer buf_n243( .i (n242), .o (n243) );
  assign n244 = ( n231 & ~n237 ) | ( n231 & n243 ) | ( ~n237 & n243 ) ;
  buffer buf_n245( .i (n244), .o (n245) );
  assign n246 = in_42_ & in_43_ ;
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  assign n250 = in_38_ & in_39_ ;
  buffer buf_n251( .i (n250), .o (n251) );
  assign n252 = in_40_ | in_41_ ;
  buffer buf_n253( .i (n252), .o (n253) );
  assign n254 = ( n247 & n251 ) | ( n247 & n253 ) | ( n251 & n253 ) ;
  buffer buf_n255( .i (n254), .o (n255) );
  assign n260 = ( ~n247 & n251 ) | ( ~n247 & n253 ) | ( n251 & n253 ) ;
  buffer buf_n261( .i (n260), .o (n261) );
  assign n262 = ( n249 & ~n255 ) | ( n249 & n261 ) | ( ~n255 & n261 ) ;
  buffer buf_n263( .i (n262), .o (n263) );
  assign n264 = ( n225 & n245 ) | ( n225 & n263 ) | ( n245 & n263 ) ;
  buffer buf_n265( .i (n264), .o (n265) );
  assign n268 = ( ~n225 & n245 ) | ( ~n225 & n263 ) | ( n245 & n263 ) ;
  buffer buf_n269( .i (n268), .o (n269) );
  assign n270 = ( n227 & ~n265 ) | ( n227 & n269 ) | ( ~n265 & n269 ) ;
  buffer buf_n271( .i (n270), .o (n271) );
  assign n272 = n219 & n271 ;
  buffer buf_n273( .i (n272), .o (n273) );
  assign n274 = n219 | n271 ;
  buffer buf_n275( .i (n274), .o (n275) );
  assign n276 = ~n273 & n275 ;
  buffer buf_n277( .i (n276), .o (n277) );
  assign n278 = in_62_ & in_63_ ;
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  assign n288 = in_61_ | in_60_ ;
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = in_53_ | in_52_ ;
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  assign n300 = in_48_ | in_49_ ;
  buffer buf_n301( .i (n300), .o (n301) );
  assign n302 = in_51_ & in_50_ ;
  buffer buf_n303( .i (n302), .o (n303) );
  assign n304 = ( n297 & n301 ) | ( n297 & n303 ) | ( n301 & n303 ) ;
  buffer buf_n305( .i (n304), .o (n305) );
  assign n310 = ( ~n297 & n301 ) | ( ~n297 & n303 ) | ( n301 & n303 ) ;
  buffer buf_n311( .i (n310), .o (n311) );
  assign n312 = ( n299 & ~n305 ) | ( n299 & n311 ) | ( ~n305 & n311 ) ;
  buffer buf_n313( .i (n312), .o (n313) );
  assign n314 = in_59_ & in_58_ ;
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  assign n318 = in_54_ & in_55_ ;
  buffer buf_n319( .i (n318), .o (n319) );
  assign n320 = in_57_ | in_56_ ;
  buffer buf_n321( .i (n320), .o (n321) );
  assign n322 = ( n315 & n319 ) | ( n315 & n321 ) | ( n319 & n321 ) ;
  buffer buf_n323( .i (n322), .o (n323) );
  assign n328 = ( ~n315 & n319 ) | ( ~n315 & n321 ) | ( n319 & n321 ) ;
  buffer buf_n329( .i (n328), .o (n329) );
  assign n330 = ( n317 & ~n323 ) | ( n317 & n329 ) | ( ~n323 & n329 ) ;
  buffer buf_n331( .i (n330), .o (n331) );
  assign n332 = ( n293 & n313 ) | ( n293 & n331 ) | ( n313 & n331 ) ;
  buffer buf_n333( .i (n332), .o (n333) );
  assign n336 = ( ~n293 & n313 ) | ( ~n293 & n331 ) | ( n313 & n331 ) ;
  buffer buf_n337( .i (n336), .o (n337) );
  assign n338 = ( n295 & ~n333 ) | ( n295 & n337 ) | ( ~n333 & n337 ) ;
  buffer buf_n339( .i (n338), .o (n339) );
  assign n340 = n287 | n339 ;
  buffer buf_n341( .i (n340), .o (n341) );
  assign n342 = n287 & n339 ;
  buffer buf_n343( .i (n342), .o (n343) );
  assign n344 = n341 & ~n343 ;
  buffer buf_n345( .i (n344), .o (n345) );
  assign n346 = n277 & n345 ;
  buffer buf_n347( .i (n346), .o (n347) );
  assign n351 = n277 | n345 ;
  buffer buf_n352( .i (n351), .o (n352) );
  assign n353 = ~n347 & n352 ;
  buffer buf_n354( .i (n353), .o (n354) );
  assign n355 = n209 & n354 ;
  buffer buf_n356( .i (n355), .o (n356) );
  assign n362 = n209 | n354 ;
  buffer buf_n363( .i (n362), .o (n363) );
  assign n364 = ~n356 & n363 ;
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  assign n374 = ( n96 & n114 ) | ( n96 & n120 ) | ( n114 & n120 ) ;
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  assign n380 = ( n96 & n114 ) | ( n96 & ~n120 ) | ( n114 & ~n120 ) ;
  buffer buf_n381( .i (n380), .o (n381) );
  assign n382 = ( n122 & ~n375 ) | ( n122 & n381 ) | ( ~n375 & n381 ) ;
  buffer buf_n383( .i (n382), .o (n383) );
  assign n384 = n128 & n383 ;
  buffer buf_n385( .i (n384), .o (n385) );
  assign n386 = n379 & n385 ;
  buffer buf_n387( .i (n386), .o (n387) );
  assign n392 = n379 | n385 ;
  buffer buf_n393( .i (n392), .o (n393) );
  assign n394 = ~n387 & n393 ;
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  assign n396 = ( n164 & n182 ) | ( n164 & n188 ) | ( n182 & n188 ) ;
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  assign n402 = ( n164 & n182 ) | ( n164 & ~n188 ) | ( n182 & ~n188 ) ;
  buffer buf_n403( .i (n402), .o (n403) );
  assign n404 = ( n190 & ~n397 ) | ( n190 & n403 ) | ( ~n397 & n403 ) ;
  buffer buf_n405( .i (n404), .o (n405) );
  assign n406 = n196 & n405 ;
  buffer buf_n407( .i (n406), .o (n407) );
  assign n408 = n401 & n407 ;
  buffer buf_n409( .i (n408), .o (n409) );
  assign n414 = n401 | n407 ;
  buffer buf_n415( .i (n414), .o (n415) );
  assign n416 = ~n409 & n415 ;
  buffer buf_n417( .i (n416), .o (n417) );
  assign n418 = n395 & n417 ;
  assign n419 = n395 | n417 ;
  assign n420 = ~n418 & n419 ;
  buffer buf_n421( .i (n420), .o (n421) );
  assign n422 = n128 | n383 ;
  buffer buf_n423( .i (n422), .o (n423) );
  assign n424 = ~n385 & n423 ;
  buffer buf_n425( .i (n424), .o (n425) );
  assign n426 = n196 | n405 ;
  buffer buf_n427( .i (n426), .o (n427) );
  assign n428 = ~n407 & n427 ;
  buffer buf_n429( .i (n428), .o (n429) );
  assign n430 = ( n202 & n425 ) | ( n202 & n429 ) | ( n425 & n429 ) ;
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  assign n435 = n421 & n434 ;
  assign n436 = n421 | n434 ;
  assign n437 = ~n435 & n436 ;
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  assign n439 = ( n241 & n259 ) | ( n241 & n265 ) | ( n259 & n265 ) ;
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  assign n445 = ( n241 & n259 ) | ( n241 & ~n265 ) | ( n259 & ~n265 ) ;
  buffer buf_n446( .i (n445), .o (n446) );
  assign n447 = ( n267 & ~n440 ) | ( n267 & n446 ) | ( ~n440 & n446 ) ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = n273 & n448 ;
  buffer buf_n450( .i (n449), .o (n450) );
  assign n451 = n444 & n450 ;
  buffer buf_n452( .i (n451), .o (n452) );
  assign n457 = n444 | n450 ;
  buffer buf_n458( .i (n457), .o (n458) );
  assign n459 = ~n452 & n458 ;
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  assign n461 = ( n309 & n327 ) | ( n309 & n333 ) | ( n327 & n333 ) ;
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  assign n467 = ( n309 & n327 ) | ( n309 & ~n333 ) | ( n327 & ~n333 ) ;
  buffer buf_n468( .i (n467), .o (n468) );
  assign n469 = ( n335 & ~n462 ) | ( n335 & n468 ) | ( ~n462 & n468 ) ;
  buffer buf_n470( .i (n469), .o (n470) );
  assign n471 = n343 & n470 ;
  buffer buf_n472( .i (n471), .o (n472) );
  assign n473 = n466 & n472 ;
  buffer buf_n474( .i (n473), .o (n474) );
  assign n479 = n466 | n472 ;
  buffer buf_n480( .i (n479), .o (n480) );
  assign n481 = ~n474 & n480 ;
  buffer buf_n482( .i (n481), .o (n482) );
  assign n483 = n460 & n482 ;
  assign n484 = n460 | n482 ;
  assign n485 = ~n483 & n484 ;
  buffer buf_n486( .i (n485), .o (n486) );
  assign n487 = n273 | n448 ;
  buffer buf_n488( .i (n487), .o (n488) );
  assign n489 = ~n450 & n488 ;
  buffer buf_n490( .i (n489), .o (n490) );
  assign n491 = n343 | n470 ;
  buffer buf_n492( .i (n491), .o (n492) );
  assign n493 = ~n472 & n492 ;
  buffer buf_n494( .i (n493), .o (n494) );
  assign n495 = ( n347 & n490 ) | ( n347 & n494 ) | ( n490 & n494 ) ;
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  assign n500 = n486 & n499 ;
  assign n501 = n486 | n499 ;
  assign n502 = ~n500 & n501 ;
  buffer buf_n503( .i (n502), .o (n503) );
  assign n504 = n438 & n503 ;
  assign n505 = n438 | n503 ;
  assign n506 = ~n504 & n505 ;
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  assign n508 = n425 & n429 ;
  assign n509 = n425 | n429 ;
  assign n510 = ~n508 & n509 ;
  buffer buf_n511( .i (n510), .o (n511) );
  assign n512 = n205 & n511 ;
  assign n513 = n205 | n511 ;
  assign n514 = ~n512 & n513 ;
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  assign n516 = n490 & n494 ;
  assign n517 = n490 | n494 ;
  assign n518 = ~n516 & n517 ;
  buffer buf_n519( .i (n518), .o (n519) );
  assign n520 = n350 & n519 ;
  assign n521 = n350 | n519 ;
  assign n522 = ~n520 & n521 ;
  buffer buf_n523( .i (n522), .o (n523) );
  assign n524 = ( n358 & n515 ) | ( n358 & n523 ) | ( n515 & n523 ) ;
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  assign n529 = n507 & n528 ;
  assign n530 = n507 | n528 ;
  assign n531 = ~n529 & n530 ;
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  assign n533 = ( n395 & n417 ) | ( n395 & n431 ) | ( n417 & n431 ) ;
  buffer buf_n534( .i (n533), .o (n534) );
  assign n535 = ( n391 & n413 ) | ( n391 & n534 ) | ( n413 & n534 ) ;
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  assign n543 = ( n460 & n482 ) | ( n460 & n496 ) | ( n482 & n496 ) ;
  buffer buf_n544( .i (n543), .o (n544) );
  assign n545 = ( n456 & n478 ) | ( n456 & n544 ) | ( n478 & n544 ) ;
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  assign n553 = n388 & n410 ;
  assign n554 = n388 | n410 ;
  assign n555 = ~n553 & n554 ;
  buffer buf_n556( .i (n555), .o (n556) );
  assign n557 = n534 & n556 ;
  assign n558 = n534 | n556 ;
  assign n559 = ~n557 & n558 ;
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  assign n564 = n453 & n475 ;
  assign n565 = n453 | n475 ;
  assign n566 = ~n564 & n565 ;
  buffer buf_n567( .i (n566), .o (n567) );
  assign n568 = n544 & n567 ;
  assign n569 = n544 | n567 ;
  assign n570 = ~n568 & n569 ;
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  assign n575 = ( n438 & n503 ) | ( n438 & n525 ) | ( n503 & n525 ) ;
  buffer buf_n576( .i (n575), .o (n576) );
  assign n577 = ( n563 & n574 ) | ( n563 & n576 ) | ( n574 & n576 ) ;
  buffer buf_n578( .i (n577), .o (n578) );
  assign n579 = ( n542 & n552 ) | ( n542 & n578 ) | ( n552 & n578 ) ;
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  assign n581 = n515 & n523 ;
  assign n582 = n515 | n523 ;
  assign n583 = ~n581 & n582 ;
  buffer buf_n584( .i (n583), .o (n584) );
  assign n585 = n361 & n584 ;
  assign n586 = n361 | n584 ;
  assign n587 = ~n585 & n586 ;
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  assign n591 = n560 & n571 ;
  assign n592 = n560 | n571 ;
  assign n593 = ~n591 & n592 ;
  buffer buf_n594( .i (n593), .o (n594) );
  assign n595 = n576 & n594 ;
  assign n596 = n576 | n594 ;
  assign n597 = ~n595 & n596 ;
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  assign n600 = n539 & n549 ;
  assign n601 = n539 | n549 ;
  assign n602 = ~n600 & n601 ;
  buffer buf_n603( .i (n602), .o (n603) );
  assign n604 = n578 & n603 ;
  assign n605 = n578 | n603 ;
  assign n606 = ~n604 & n605 ;
  assign out_1_ = n373 ;
  assign out_3_ = n532 ;
  assign out_6_ = n580 ;
  assign out_2_ = n590 ;
  assign out_0_ = 1'b0 ;
  assign out_4_ = n599 ;
  assign out_5_ = n606 ;
endmodule
