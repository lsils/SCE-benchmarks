module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 ;
  buffer buf_n17( .i (x1), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n29( .i (x2), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n67( .i (x5), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  assign n115 = n31 | n69 ;
  buffer buf_n116( .i (n115), .o (n116) );
  assign n122 = n21 | n116 ;
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n42( .i (x3), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n104( .i (x8), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  assign n126 = ~n44 & n106 ;
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n54( .i (x4), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  assign n132 = n4 | n56 ;
  buffer buf_n133( .i (n132), .o (n133) );
  assign n141 = n127 & ~n133 ;
  buffer buf_n142( .i (n141), .o (n142) );
  assign n145 = ~n123 & n142 ;
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n93( .i (x7), .o (n93) );
  assign n153 = n93 & ~n104 ;
  buffer buf_n154( .i (n153), .o (n154) );
  assign n161 = ~n93 & n104 ;
  buffer buf_n162( .i (n161), .o (n162) );
  assign n170 = n154 | n162 ;
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  assign n181 = n18 | n30 ;
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  assign n191 = n12 & n52 ;
  assign n192 = ( n13 & n190 ) | ( n13 & n191 ) | ( n190 & n191 ) ;
  buffer buf_n193( .i (n192), .o (n193) );
  assign n195 = n180 & ~n193 ;
  assign n196 = ~n152 & n195 ;
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  assign n197 = n95 & n106 ;
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n70( .i (n69), .o (n70) );
  assign n204 = ~n45 & n70 ;
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  assign n209 = ~n101 & n208 ;
  assign n210 = n203 | n209 ;
  assign n211 = ~n44 & n56 ;
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n71( .i (n70), .o (n71) );
  assign n217 = ~n19 & n31 ;
  buffer buf_n218( .i (n217), .o (n218) );
  assign n223 = n71 & n218 ;
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  assign n226 = ~n215 & n225 ;
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n57( .i (n56), .o (n57) );
  assign n228 = n32 & n57 ;
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  assign n234 = n19 & ~n44 ;
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n241( .i (n43), .o (n241) );
  assign n242 = n31 & n241 ;
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  assign n247 = n236 | n244 ;
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  assign n250 = n232 | n249 ;
  assign n251 = n227 | n250 ;
  assign n252 = n210 & ~n251 ;
  buffer buf_n80( .i (x6), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  assign n253 = n43 | n81 ;
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n260( .i (n30), .o (n260) );
  assign n261 = ~n56 & n260 ;
  buffer buf_n262( .i (n261), .o (n262) );
  assign n268 = ~n255 & n262 ;
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  assign n273 = n43 | n55 ;
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  assign n279 = n166 & n277 ;
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n219( .i (n218), .o (n219) );
  assign n281 = ~n98 & n219 ;
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  assign n284 = n280 | n283 ;
  assign n285 = n272 | n284 ;
  buffer buf_n286( .i (n55), .o (n286) );
  assign n287 = n19 | n286 ;
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  assign n292 = n32 | n96 ;
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n296( .i (n42), .o (n296) );
  assign n297 = n55 & n296 ;
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  assign n304 = n294 | n301 ;
  assign n305 = n291 & ~n304 ;
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  assign n308 = n106 | n241 ;
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n82( .i (n81), .o (n82) );
  assign n314 = n69 & n82 ;
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n319( .i (n54), .o (n319) );
  assign n320 = n105 | n319 ;
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  assign n329 = n317 | n324 ;
  assign n330 = n312 & n329 ;
  buffer buf_n331( .i (n330), .o (n331) );
  assign n332 = n306 | n331 ;
  assign n333 = ( n285 & n307 ) | ( n285 & n332 ) | ( n307 & n332 ) ;
  assign n334 = n252 | n333 ;
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  assign n336 = ~n114 & n189 ;
  assign n337 = n7 | n98 ;
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  assign n343 = n336 | n342 ;
  buffer buf_n344( .i (n343), .o (n344) );
  assign n345 = n335 & ~n344 ;
  buffer buf_n346( .i (n18), .o (n346) );
  assign n347 = n4 | n346 ;
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  assign n357 = n32 & ~n96 ;
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  assign n362 = n202 | n361 ;
  assign n363 = ( n203 & ~n331 ) | ( n203 & n362 ) | ( ~n331 & n362 ) ;
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  assign n366 = ~n356 & n365 ;
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  assign n367 = n69 & n286 ;
  buffer buf_n368( .i (n367), .o (n368) );
  assign n372 = n84 & n368 ;
  buffer buf_n373( .i (n372), .o (n373) );
  assign n377 = n129 & ~n373 ;
  buffer buf_n378( .i (n377), .o (n378) );
  assign n379 = n18 & ~n30 ;
  buffer buf_n380( .i (n379), .o (n380) );
  assign n388 = ~n5 & n380 ;
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  assign n394 = n378 & n392 ;
  buffer buf_n395( .i (n17), .o (n395) );
  assign n396 = ~n3 & n395 ;
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n408( .i (n260), .o (n408) );
  assign n409 = n397 & n408 ;
  buffer buf_n410( .i (n409), .o (n410) );
  assign n415 = n3 & ~n296 ;
  buffer buf_n416( .i (n415), .o (n416) );
  assign n422 = ~n182 & n416 ;
  buffer buf_n423( .i (n422), .o (n423) );
  assign n429 = n410 | n423 ;
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n433( .i (n68), .o (n433) );
  assign n434 = n4 | n433 ;
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  assign n440 = n213 | n436 ;
  buffer buf_n441( .i (n440), .o (n441) );
  assign n442 = n174 & n441 ;
  assign n443 = n431 & n442 ;
  assign n444 = n394 | n443 ;
  buffer buf_n445( .i (n444), .o (n445) );
  assign n446 = n6 | n183 ;
  buffer buf_n447( .i (n446), .o (n447) );
  assign n450 = ~n171 & n255 ;
  buffer buf_n451( .i (n450), .o (n451) );
  assign n454 = ~n447 & n451 ;
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  assign n458 = n174 & n258 ;
  buffer buf_n459( .i (n458), .o (n459) );
  assign n460 = n414 & n459 ;
  assign n461 = n457 | n460 ;
  assign n462 = n445 | n461 ;
  buffer buf_n463( .i (n462), .o (n463) );
  assign n464 = n366 | n463 ;
  assign n465 = n345 | n464 ;
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n466( .i (n105), .o (n466) );
  assign n467 = n433 & ~n466 ;
  buffer buf_n468( .i (n467), .o (n468) );
  assign n473 = ~n58 & n468 ;
  buffer buf_n474( .i (n473), .o (n474) );
  assign n477 = n82 & n286 ;
  buffer buf_n478( .i (n477), .o (n478) );
  assign n484 = n433 & n466 ;
  buffer buf_n485( .i (n484), .o (n485) );
  assign n490 = n478 & n485 ;
  buffer buf_n491( .i (n490), .o (n491) );
  assign n494 = n474 | n491 ;
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  assign n497 = n26 & ~n496 ;
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  assign n500 = n46 & n108 ;
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  assign n504 = n45 & ~n83 ;
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  assign n508 = n95 & ~n433 ;
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  assign n514 = n506 & n511 ;
  buffer buf_n515( .i (n514), .o (n515) );
  assign n518 = n503 | n515 ;
  assign n519 = n38 & n518 ;
  buffer buf_n520( .i (n519), .o (n520) );
  assign n521 = ~n241 & n260 ;
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  assign n529 = n58 & n156 ;
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  assign n535 = ~n528 & n534 ;
  assign n536 = ~n520 & n535 ;
  assign n537 = n94 & ~n296 ;
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  assign n545 = ~n82 & n260 ;
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  assign n550 = ~n60 & n548 ;
  buffer buf_n551( .i (n550), .o (n551) );
  assign n552 = n543 & n551 ;
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n68), .o (n554) );
  buffer buf_n555( .i (n81), .o (n555) );
  assign n556 = n554 | n555 ;
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n563( .i (n29), .o (n563) );
  assign n564 = n296 & ~n563 ;
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  assign n573 = ~n559 & n568 ;
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  assign n576 = n37 & n131 ;
  assign n577 = n575 | n576 ;
  assign n578 = n553 | n577 ;
  assign n579 = n498 & n578 ;
  assign n580 = ( n499 & n536 ) | ( n499 & n579 ) | ( n536 & n579 ) ;
  assign n581 = n335 | n580 ;
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n398( .i (n397), .o (n398) );
  assign n582 = n398 & n566 ;
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  assign n586 = n425 | n584 ;
  assign n587 = n175 & n586 ;
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  assign n590 = n286 | n554 ;
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  assign n599 = n99 | n593 ;
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n42), .o (n602) );
  assign n603 = n81 & n602 ;
  buffer buf_n604( .i (n603), .o (n604) );
  assign n610 = n254 & ~n604 ;
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n3), .o (n615) );
  buffer buf_n616( .i (n563), .o (n616) );
  assign n617 = n615 | n616 ;
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  assign n626 = n466 & n555 ;
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  assign n634 = n621 | n630 ;
  assign n635 = n614 & ~n634 ;
  assign n636 = ~n601 & n635 ;
  buffer buf_n393( .i (n392), .o (n393) );
  assign n637 = n393 & n496 ;
  assign n638 = n636 | n637 ;
  assign n639 = n589 | n638 ;
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  assign n642 = n15 & ~n640 ;
  assign n643 = ( n581 & n641 ) | ( n581 & ~n642 ) | ( n641 & ~n642 ) ;
  assign n644 = n48 & ~n200 ;
  buffer buf_n645( .i (n644), .o (n645) );
  assign n646 = ~n83 & n96 ;
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  assign n652 = n301 & ~n648 ;
  buffer buf_n653( .i (n652), .o (n653) );
  assign n654 = n645 | n653 ;
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n655( .i (n319), .o (n655) );
  assign n656 = ~n616 & n655 ;
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  assign n662 = n472 & n661 ;
  assign n663 = n654 & ~n662 ;
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  assign n665 = n110 & ~n370 ;
  buffer buf_n666( .i (n665), .o (n666) );
  assign n667 = n661 | n666 ;
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  assign n669 = ( n50 & ~n101 ) | ( n50 & n120 ) | ( ~n101 & n120 ) ;
  assign n670 = n121 & ~n669 ;
  assign n671 = ( ~n52 & n668 ) | ( ~n52 & n670 ) | ( n668 & n670 ) ;
  assign n672 = n664 | n671 ;
  assign n673 = ~n368 & n591 ;
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  assign n679 = n46 & n97 ;
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  assign n683 = ~n37 & n682 ;
  assign n684 = n677 & n683 ;
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  assign n685 = n466 | n554 ;
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  assign n691 = n547 & ~n687 ;
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  assign n694 = ~n62 & n693 ;
  assign n695 = n26 & ~n694 ;
  assign n696 = ~n684 & n695 ;
  assign n697 = ~n520 & n696 ;
  assign n698 = n672 & n697 ;
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n313( .i (n312), .o (n313) );
  assign n699 = ~n101 & n313 ;
  assign n700 = n596 & n699 ;
  assign n701 = ~n166 & n311 ;
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n371( .i (n370), .o (n371) );
  assign n703 = n95 | n241 ;
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  assign n710 = ~n371 & n707 ;
  assign n711 = ~n702 & n710 ;
  buffer buf_n712( .i (n711), .o (n712) );
  assign n713 = n700 | n712 ;
  assign n714 = ~n625 & n713 ;
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n715( .i (n2), .o (n715) );
  assign n716 = n563 & ~n715 ;
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  assign n723 = n215 & n721 ;
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  assign n726 = n203 | n403 ;
  assign n727 = ( n404 & n725 ) | ( n404 & n726 ) | ( n725 & n726 ) ;
  assign n728 = n94 | n105 ;
  buffer buf_n729( .i (n728), .o (n729) );
  assign n735 = n57 | n729 ;
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  assign n741 = ~n436 & n523 ;
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  assign n745 = ~n740 & n744 ;
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  assign n746 = n112 & ~n513 ;
  assign n747 = ~n615 & n655 ;
  buffer buf_n748( .i (n747), .o (n748) );
  assign n753 = n243 & n748 ;
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = ~n746 & n757 ;
  assign n759 = n745 | n758 ;
  assign n760 = n727 | n759 ;
  assign n761 = n714 | n760 ;
  assign n762 = ~n698 & n761 ;
  buffer buf_n763( .i (n94), .o (n763) );
  assign n764 = n554 & n763 ;
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n769( .i (n68), .o (n769) );
  assign n770 = n763 | n769 ;
  buffer buf_n771( .i (n770), .o (n771) );
  assign n776 = ~n765 & n771 ;
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  assign n782 = ~n267 & n527 ;
  assign n783 = ~n781 & n782 ;
  assign n784 = n346 & n616 ;
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n602), .o (n790) );
  assign n791 = ~n763 & n790 ;
  buffer buf_n792( .i (n791), .o (n792) );
  assign n796 = ~n108 & n792 ;
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  assign n800 = ~n789 & n799 ;
  assign n801 = n202 & n208 ;
  assign n802 = n800 | n801 ;
  buffer buf_n803( .i (n802), .o (n803) );
  assign n804 = n783 | n803 ;
  assign n805 = ~n23 & n118 ;
  assign n806 = ~n225 & n805 ;
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  assign n809 = n23 & ~n60 ;
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  assign n812 = ~n6 & n84 ;
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  assign n817 = ~n811 & n816 ;
  assign n818 = ~n808 & n817 ;
  buffer buf_n819( .i (n818), .o (n819) );
  assign n820 = n804 & n819 ;
  assign n821 = ~n655 & n763 ;
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  assign n828 = n47 & n719 ;
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  assign n831 = n826 & n830 ;
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  assign n835 = ~n317 & n824 ;
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  assign n840 = n177 & n428 ;
  assign n841 = ~n839 & n840 ;
  assign n842 = n834 | n841 ;
  assign n843 = n820 | n842 ;
  assign n844 = n762 | n843 ;
  assign n845 = ~n555 & n655 ;
  buffer buf_n846( .i (n845), .o (n846) );
  assign n851 = ~n309 & n846 ;
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n100), .o (n855) );
  assign n856 = n854 & n855 ;
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  assign n859 = n20 & n57 ;
  buffer buf_n860( .i (n859), .o (n860) );
  assign n865 = n289 & ~n860 ;
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  assign n870 = ~n485 & n686 ;
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n875( .i (n319), .o (n875) );
  buffer buf_n876( .i (n93), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  assign n878 = n875 & ~n877 ;
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  assign n884 = ~n86 & n881 ;
  assign n885 = n872 & n884 ;
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  assign n888 = n869 | n887 ;
  assign n889 = ~n769 & n790 ;
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  assign n895 = n541 | n892 ;
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n877), .o (n898) );
  assign n899 = n70 & ~n898 ;
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n906( .i (n104), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  assign n908 = n555 | n907 ;
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  assign n916 = n215 | n912 ;
  assign n917 = n903 & n916 ;
  assign n918 = n897 | n917 ;
  assign n919 = ~n857 & n918 ;
  assign n920 = ( n858 & n888 ) | ( n858 & ~n919 ) | ( n888 & ~n919 ) ;
  assign n921 = ~n319 & n602 ;
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n928( .i (n80), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  assign n930 = n907 & ~n929 ;
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  assign n937 = n510 & n932 ;
  buffer buf_n938( .i (n937), .o (n938) );
  assign n940 = n926 & n938 ;
  assign n941 = n183 & ~n785 ;
  buffer buf_n942( .i (n941), .o (n942) );
  assign n943 = n166 & n942 ;
  buffer buf_n944( .i (n943), .o (n944) );
  assign n945 = n940 | n944 ;
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  assign n946 = n47 & ~n184 ;
  buffer buf_n947( .i (n946), .o (n947) );
  assign n948 = n159 & n947 ;
  buffer buf_n933( .i (n932), .o (n933) );
  assign n949 = n21 & ~n71 ;
  buffer buf_n950( .i (n949), .o (n950) );
  assign n953 = n933 | n950 ;
  buffer buf_n954( .i (n875), .o (n954) );
  assign n955 = n408 | n954 ;
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  assign n959 = n99 & ~n957 ;
  assign n960 = n953 & n959 ;
  assign n961 = n948 | n960 ;
  assign n962 = n945 | n961 ;
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  assign n965 = n40 | n963 ;
  assign n966 = ( n920 & n964 ) | ( n920 & n965 ) | ( n964 & n965 ) ;
  assign n967 = ~n15 & n966 ;
  buffer buf_n968( .i (n54), .o (n968) );
  assign n969 = n906 & n968 ;
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  assign n977 = n158 & n264 ;
  buffer buf_n766( .i (n765), .o (n766) );
  assign n978 = n658 & n766 ;
  buffer buf_n979( .i (n67), .o (n979) );
  assign n980 = ~n968 & n979 ;
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  assign n988 = ~n97 & n982 ;
  buffer buf_n989( .i (n988), .o (n989) );
  assign n994 = n978 | n989 ;
  assign n995 = n977 | n994 ;
  buffer buf_n996( .i (n995), .o (n996) );
  assign n997 = n976 | n996 ;
  buffer buf_n998( .i (n997), .o (n998) );
  assign n999 = n875 & n877 ;
  buffer buf_n1000( .i (n999), .o (n1000) );
  assign n1005 = n875 | n877 ;
  buffer buf_n1006( .i (n1005), .o (n1006) );
  assign n1011 = ~n1000 & n1006 ;
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  assign n1016 = n395 | n602 ;
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  assign n1023 = ~n616 & n907 ;
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  assign n1027 = n1020 | n1026 ;
  buffer buf_n1028( .i (n1027), .o (n1028) );
  assign n1029 = ( n1014 & n1022 ) | ( n1014 & n1028 ) | ( n1022 & n1028 ) ;
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  assign n1032 = n12 & ~n1030 ;
  assign n1033 = ( n998 & n1031 ) | ( n998 & ~n1032 ) | ( n1031 & ~n1032 ) ;
  assign n1034 = n720 & n797 ;
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  assign n1037 = n677 & n1036 ;
  assign n1038 = ~n71 & n718 ;
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n134( .i (n133), .o (n134) );
  assign n1042 = ~n134 & n199 ;
  buffer buf_n1043( .i (n1042), .o (n1043) );
  assign n1044 = n1040 & n1043 ;
  buffer buf_n1045( .i (n1044), .o (n1045) );
  assign n1046 = n26 & ~n1045 ;
  assign n1047 = ~n1037 & n1046 ;
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  assign n1048 = n60 | n487 ;
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  assign n1049 = ~n620 & n773 ;
  assign n1050 = ~n1048 & n1049 ;
  assign n1051 = n58 & ~n435 ;
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  assign n1054 = ~n346 & n790 ;
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  assign n1059 = n732 & n1057 ;
  assign n1060 = ( ~n1053 & n1058 ) | ( ~n1053 & n1059 ) | ( n1058 & n1059 ) ;
  assign n1061 = ~n1050 & n1060 ;
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  assign n1064 = ~n107 & n954 ;
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  assign n1072 = ~n621 & n1067 ;
  assign n1073 = n144 | n1072 ;
  assign n1074 = ~n897 & n1073 ;
  assign n1075 = ~n1062 & n1074 ;
  assign n1076 = ( n1047 & n1063 ) | ( n1047 & ~n1075 ) | ( n1063 & ~n1075 ) ;
  assign n1077 = n1033 & ~n1076 ;
  assign n1078 = n35 & ~n901 ;
  buffer buf_n1079( .i (n1078), .o (n1079) );
  assign n1081 = n25 | n1079 ;
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  assign n1082 = n361 & n952 ;
  assign n1083 = n1081 & ~n1082 ;
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n135( .i (n134), .o (n135) );
  assign n1084 = ~n907 & n929 ;
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  assign n1094 = ~n135 & n1087 ;
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  assign n1097 = ~n544 & n1096 ;
  assign n1098 = ~n1083 & n1097 ;
  assign n1099 = n85 & n165 ;
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  assign n1103 = n426 & n1101 ;
  buffer buf_n847( .i (n846), .o (n847) );
  assign n1104 = ~n70 & n107 ;
  buffer buf_n1105( .i (n1104), .o (n1105) );
  assign n1110 = n847 & n1105 ;
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  assign n1113 = n836 | n1112 ;
  assign n1114 = ( n427 & n1103 ) | ( n427 & n1113 ) | ( n1103 & n1113 ) ;
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  assign n1115 = ~n348 & n522 ;
  buffer buf_n1116( .i (n1115), .o (n1116) );
  assign n1119 = n629 & n1116 ;
  buffer buf_n1120( .i (n1119), .o (n1120) );
  assign n1121 = n75 & n1120 ;
  buffer buf_n479( .i (n478), .o (n479) );
  assign n1122 = n479 & ~n510 ;
  buffer buf_n1123( .i (n1122), .o (n1123) );
  assign n1125 = n391 & n1123 ;
  assign n1126 = ~n615 & n790 ;
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  assign n1133 = n1065 & n1128 ;
  buffer buf_n1134( .i (n1133), .o (n1134) );
  assign n1135 = n548 & n950 ;
  assign n1136 = n1134 & n1135 ;
  assign n1137 = n1125 | n1136 ;
  assign n1138 = n1121 | n1137 ;
  assign n1139 = n1114 | n1138 ;
  assign n1140 = n1098 | n1139 ;
  assign n1141 = n83 | n954 ;
  buffer buf_n1142( .i (n1141), .o (n1142) );
  assign n1147 = ~n479 & n1142 ;
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n432( .i (n431), .o (n432) );
  assign n1152 = n208 | n743 ;
  assign n1153 = ( n432 & n744 ) | ( n432 & n1152 ) | ( n744 & n1152 ) ;
  assign n1154 = ~n1151 & n1153 ;
  assign n1155 = ~n509 & n718 ;
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  assign n1160 = n203 & n1159 ;
  buffer buf_n1161( .i (n1160), .o (n1161) );
  assign n1162 = n687 & n719 ;
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  assign n1167 = n177 & ~n1166 ;
  assign n1168 = ( n1154 & n1161 ) | ( n1154 & n1167 ) | ( n1161 & n1167 ) ;
  assign n1169 = n1140 | n1168 ;
  assign n1170 = n1077 | n1169 ;
  assign n1171 = n967 | n1170 ;
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n1172( .i (n769), .o (n1172) );
  assign n1173 = n45 & n1172 ;
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  assign n1178 = ~n98 & n658 ;
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  assign n1181 = n1177 & n1180 ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  assign n1184 = n968 & ~n979 ;
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  assign n1190 = n501 & n1188 ;
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  assign n1193 = n38 & n1192 ;
  assign n1194 = n517 | n1193 ;
  assign n1195 = n1183 | n1194 ;
  assign n1196 = n406 & n1195 ;
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  assign n1197 = ~n315 & n557 ;
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  assign n1203 = n544 & n1201 ;
  assign n1204 = n408 & ~n1172 ;
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  assign n1210 = n88 & ~n208 ;
  assign n1211 = ~n1209 & n1210 ;
  assign n1212 = n1203 | n1211 ;
  assign n1213 = n1071 & n1212 ;
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  assign n1214 = ~n34 & n510 ;
  buffer buf_n1215( .i (n1214), .o (n1215) );
  assign n1216 = ~n325 & n1215 ;
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n507( .i (n506), .o (n507) );
  assign n1219 = n507 & n902 ;
  buffer buf_n1220( .i (n1219), .o (n1220) );
  assign n1221 = n85 & n891 ;
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  assign n1225 = n1220 | n1224 ;
  assign n1226 = ( ~n328 & n1218 ) | ( ~n328 & n1225 ) | ( n1218 & n1225 ) ;
  buffer buf_n1227( .i (n1226), .o (n1227) );
  assign n1228 = n1213 | n1227 ;
  assign n1229 = ( n407 & n1196 ) | ( n407 & n1228 ) | ( n1196 & n1228 ) ;
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  assign n1230 = ~n184 & n891 ;
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  assign n1233 = n526 | n1232 ;
  assign n1234 = ~n86 & n158 ;
  assign n1235 = n1100 | n1234 ;
  buffer buf_n1236( .i (n1235), .o (n1236) );
  assign n1237 = n1233 & n1236 ;
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  assign n1238 = ~n125 & n1089 ;
  assign n1239 = ~n627 & n909 ;
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1245( .i (n1172), .o (n1245) );
  assign n1246 = ~n21 & n1245 ;
  buffer buf_n1247( .i (n1246), .o (n1247) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  assign n1250 = n525 & n1248 ;
  assign n1251 = ~n1242 & n1250 ;
  assign n1252 = n1238 | n1251 ;
  assign n1253 = n1237 | n1252 ;
  assign n1254 = ~n140 & n1253 ;
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  assign n1255 = ~n200 & n750 ;
  buffer buf_n1256( .i (n1255), .o (n1256) );
  assign n1257 = n46 | n183 ;
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  assign n1260 = n778 | n1259 ;
  assign n1261 = n1256 & ~n1260 ;
  assign n1262 = n8 | n173 ;
  buffer buf_n1263( .i (n1262), .o (n1263) );
  assign n1266 = n107 & ~n954 ;
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  assign n1272 = n911 & ~n1268 ;
  assign n1273 = n225 & n1272 ;
  assign n1274 = ~n1263 & n1273 ;
  assign n1275 = n1261 | n1274 ;
  assign n1276 = ~n633 & n1275 ;
  buffer buf_n1277( .i (n59), .o (n1277) );
  assign n1278 = n548 | n1277 ;
  buffer buf_n1279( .i (n1278), .o (n1279) );
  assign n1280 = n199 | n505 ;
  buffer buf_n1281( .i (n1280), .o (n1281) );
  assign n1283 = n99 & n1175 ;
  assign n1284 = n1281 | n1283 ;
  assign n1285 = ~n1279 & n1284 ;
  buffer buf_n1286( .i (n876), .o (n1286) );
  assign n1287 = n929 | n1286 ;
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  assign n1292 = ~n110 & n1290 ;
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  assign n1295 = n902 | n1107 ;
  assign n1296 = n1293 | n1295 ;
  assign n1297 = ~n1285 & n1296 ;
  assign n1298 = n219 & n1128 ;
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  assign n1303 = n201 | n351 ;
  assign n1304 = n690 & ~n1303 ;
  assign n1305 = n1301 | n1304 ;
  assign n1306 = ~n1297 & n1305 ;
  assign n1307 = n1276 | n1306 ;
  assign n1308 = n1254 | n1307 ;
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  assign n1309 = n607 & n777 ;
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n547), .o (n1311) );
  assign n1312 = n206 & ~n1311 ;
  buffer buf_n1313( .i (n1312), .o (n1313) );
  assign n1314 = n1310 | n1313 ;
  buffer buf_n1315( .i (n1314), .o (n1315) );
  assign n1316 = n267 & n403 ;
  assign n1317 = n1315 & n1316 ;
  assign n1318 = n346 & ~n1286 ;
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  assign n1325 = ~n9 & n1322 ;
  buffer buf_n1326( .i (n1325), .o (n1326) );
  assign n1327 = n274 & ~n298 ;
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1331( .i (n563), .o (n1331) );
  buffer buf_n1332( .i (n906), .o (n1332) );
  assign n1333 = n1331 & n1332 ;
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  assign n1338 = ~n1329 & n1336 ;
  buffer buf_n1339( .i (n1338), .o (n1339) );
  assign n1341 = n300 | n687 ;
  buffer buf_n1342( .i (n1341), .o (n1342) );
  assign n1344 = n86 | n264 ;
  assign n1345 = n1342 | n1344 ;
  assign n1346 = ~n1339 & n1345 ;
  assign n1347 = n1326 & ~n1346 ;
  assign n1348 = n769 & ~n929 ;
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1353( .i (n968), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  assign n1356 = n1349 & n1355 ;
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  assign n1359 = n310 | n349 ;
  buffer buf_n1360( .i (n1359), .o (n1360) );
  assign n1362 = n1358 & ~n1360 ;
  buffer buf_n1363( .i (n1362), .o (n1363) );
  assign n1364 = ~n715 & n876 ;
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  assign n1371 = n316 & n1367 ;
  buffer buf_n1372( .i (n1371), .o (n1372) );
  assign n1373 = n947 & n1372 ;
  assign n1374 = n658 | n1019 ;
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  assign n1377 = ~n688 & n1368 ;
  assign n1378 = ~n1375 & n1377 ;
  assign n1379 = n1373 | n1378 ;
  assign n1380 = n1363 | n1379 ;
  assign n1381 = n1347 | n1380 ;
  assign n1382 = n1317 | n1381 ;
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  assign n1383 = n59 & n469 ;
  assign n1384 = n1002 | n1383 ;
  buffer buf_n1385( .i (n1384), .o (n1385) );
  assign n1388 = ~n7 & n1056 ;
  buffer buf_n1389( .i (n1388), .o (n1389) );
  assign n1391 = ~n1163 & n1389 ;
  assign n1392 = n1385 & n1391 ;
  assign n1393 = ~n348 & n1245 ;
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  assign n1396 = n1331 & ~n1332 ;
  buffer buf_n1397( .i (n1396), .o (n1397) );
  assign n1404 = n164 | n1397 ;
  assign n1405 = ~n276 & n1404 ;
  buffer buf_n1406( .i (n1405), .o (n1406) );
  assign n1407 = n1395 & n1406 ;
  buffer buf_n1408( .i (n1407), .o (n1408) );
  assign n1409 = n1392 | n1408 ;
  assign n1410 = n321 & ~n970 ;
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  assign n1417 = n424 & n1351 ;
  buffer buf_n1418( .i (n1417), .o (n1418) );
  assign n1420 = ~n1414 & n1418 ;
  assign n1421 = n165 | n647 ;
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n979), .o (n1424) );
  assign n1425 = ~n1331 & n1424 ;
  buffer buf_n1426( .i (n1425), .o (n1426) );
  assign n1429 = n5 & ~n20 ;
  assign n1430 = n1426 & n1429 ;
  buffer buf_n1431( .i (n1430), .o (n1431) );
  assign n1436 = n214 & n1431 ;
  buffer buf_n1437( .i (n1436), .o (n1437) );
  assign n1439 = n1423 & n1437 ;
  assign n1440 = n1420 | n1439 ;
  assign n1441 = n1409 | n1440 ;
  assign n1442 = n200 & ~n1198 ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n245( .i (n244), .o (n245) );
  assign n1446 = ~n245 & n400 ;
  buffer buf_n1447( .i (n1446), .o (n1447) );
  assign n1448 = n1443 & n1447 ;
  buffer buf_n1041( .i (n1040), .o (n1041) );
  assign n1449 = ~n20 & n1354 ;
  buffer buf_n1450( .i (n1449), .o (n1450) );
  assign n1454 = n1289 & ~n1450 ;
  assign n1455 = n129 & ~n1454 ;
  buffer buf_n1456( .i (n1455), .o (n1456) );
  assign n1459 = n1041 & n1456 ;
  assign n1460 = n1448 | n1459 ;
  assign n1461 = n116 | n288 ;
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  assign n1465 = ~n158 & n419 ;
  assign n1466 = ~n1100 & n1465 ;
  assign n1467 = ~n1464 & n1466 ;
  buffer buf_n1468( .i (n928), .o (n1468) );
  assign n1469 = n1286 & n1468 ;
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  assign n1477 = n424 & n1188 ;
  buffer buf_n1478( .i (n1477), .o (n1478) );
  assign n1479 = n1474 & n1478 ;
  assign n1480 = n1467 | n1479 ;
  assign n1481 = n1460 | n1480 ;
  assign n1482 = n1441 | n1481 ;
  assign n1483 = n1382 | n1482 ;
  assign n1484 = n1308 | n1483 ;
  assign n1485 = n1229 | n1484 ;
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  assign n1486 = n110 & ~n773 ;
  buffer buf_n1487( .i (n1486), .o (n1487) );
  assign n1488 = n316 & n1267 ;
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  assign n1491 = n1487 | n1490 ;
  assign n1492 = n571 & n1491 ;
  assign n1493 = ( n572 & n887 ) | ( n572 & n1492 ) | ( n887 & n1492 ) ;
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  assign n1494 = n85 | n705 ;
  buffer buf_n1495( .i (n1494), .o (n1495) );
  assign n1497 = n509 & n1355 ;
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  assign n1501 = n1495 & ~n1499 ;
  assign n1502 = n1401 & ~n1501 ;
  buffer buf_n1189( .i (n1188), .o (n1189) );
  assign n1503 = n567 & n932 ;
  buffer buf_n1504( .i (n1503), .o (n1504) );
  assign n1505 = n1189 & n1504 ;
  assign n1506 = n25 | n1505 ;
  assign n1507 = n1502 | n1506 ;
  assign n1508 = n900 & n972 ;
  buffer buf_n1509( .i (n1508), .o (n1509) );
  assign n1511 = n525 & n1509 ;
  assign n1512 = ( n526 & n1443 ) | ( n526 & n1511 ) | ( n1443 & n1511 ) ;
  assign n1513 = n523 | n567 ;
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  assign n1516 = ~n173 & n373 ;
  buffer buf_n1517( .i (n1516), .o (n1517) );
  assign n1518 = ~n1515 & n1517 ;
  assign n1519 = n1512 | n1518 ;
  assign n1520 = n1507 | n1519 ;
  assign n1521 = n1493 | n1520 ;
  buffer buf_n89( .i (n88), .o (n89) );
  assign n1522 = n1206 & ~n1329 ;
  assign n1523 = n214 & ~n1206 ;
  assign n1524 = n1522 | n1523 ;
  buffer buf_n1525( .i (n1524), .o (n1525) );
  assign n1526 = ~n89 & n1525 ;
  buffer buf_n1527( .i (n84), .o (n1527) );
  assign n1528 = ~n592 & n1527 ;
  buffer buf_n1529( .i (n1528), .o (n1529) );
  assign n1532 = n1358 | n1529 ;
  assign n1533 = n36 & ~n681 ;
  assign n1534 = n1532 & ~n1533 ;
  assign n1535 = ~n113 & n1534 ;
  assign n1536 = ( ~n114 & n1526 ) | ( ~n114 & n1535 ) | ( n1526 & n1535 ) ;
  assign n1537 = n487 & ~n524 ;
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  assign n1540 = n361 & ~n1149 ;
  assign n1541 = n1539 & n1540 ;
  assign n1542 = ~n37 & n1223 ;
  buffer buf_n1543( .i (n42), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1468), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  assign n1549 = ~n1546 & n1548 ;
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1553( .i (n199), .o (n1553) );
  assign n1554 = n1550 & n1553 ;
  buffer buf_n1555( .i (n1554), .o (n1555) );
  assign n1556 = n25 & ~n1555 ;
  assign n1557 = ~n1542 & n1556 ;
  assign n1558 = ~n1541 & n1557 ;
  assign n1559 = ~n1536 & n1558 ;
  assign n1560 = n1521 & ~n1559 ;
  assign n1561 = ~n898 & n1547 ;
  buffer buf_n1562( .i (n1561), .o (n1562) );
  assign n1568 = n47 & n1562 ;
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  assign n1572 = n62 | n1022 ;
  assign n1573 = ~n1571 & n1572 ;
  buffer buf_n1415( .i (n1414), .o (n1415) );
  assign n1574 = n1209 & n1415 ;
  assign n1575 = ~n1573 & n1574 ;
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  assign n1576 = n187 | n614 ;
  buffer buf_n1577( .i (n1576), .o (n1577) );
  assign n1579 = n993 & ~n1577 ;
  assign n1580 = n1575 | n1579 ;
  assign n1581 = ~n14 & n1580 ;
  assign n1582 = ( ~n15 & n1560 ) | ( ~n15 & n1581 ) | ( n1560 & n1581 ) ;
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  assign n1583 = n400 & n674 ;
  assign n1584 = n1514 & n1583 ;
  buffer buf_n1585( .i (n1584), .o (n1585) );
  assign n1587 = n1324 & n1585 ;
  buffer buf_n1243( .i (n1242), .o (n1243) );
  assign n1588 = n981 & ~n1017 ;
  buffer buf_n1589( .i (n1588), .o (n1589) );
  assign n1593 = n7 & n1589 ;
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1596( .i (n182), .o (n1596) );
  assign n1597 = n97 & ~n1596 ;
  buffer buf_n1598( .i (n1597), .o (n1598) );
  assign n1602 = ~n1087 & n1598 ;
  assign n1603 = n1594 & n1602 ;
  buffer buf_n1604( .i (n1603), .o (n1604) );
  assign n1605 = n1243 & ~n1604 ;
  assign n1606 = ~n1587 & n1605 ;
  buffer buf_n1607( .i (n395), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  assign n1609 = n1172 | n1608 ;
  buffer buf_n1610( .i (n1609), .o (n1610) );
  assign n1611 = ~n1174 & n1610 ;
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  assign n1615 = n431 & n1014 ;
  assign n1616 = n719 & n1001 ;
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  assign n1619 = ~n1613 & n1618 ;
  assign n1620 = ( ~n1614 & n1615 ) | ( ~n1614 & n1619 ) | ( n1615 & n1619 ) ;
  buffer buf_n1621( .i (n1424), .o (n1621) );
  assign n1622 = ~n5 & n1621 ;
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  assign n1630 = n391 | n1625 ;
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  assign n1633 = ~n135 & n794 ;
  buffer buf_n1634( .i (n1633), .o (n1634) );
  buffer buf_n1635( .i (n1634), .o (n1635) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  assign n1636 = n222 & n1634 ;
  assign n1637 = ( ~n1631 & n1635 ) | ( ~n1631 & n1636 ) | ( n1635 & n1636 ) ;
  assign n1638 = n1620 | n1637 ;
  assign n1639 = n1606 & ~n1638 ;
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  assign n1640 = n212 & ~n1596 ;
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  assign n1645 = ~n775 & n1643 ;
  buffer buf_n585( .i (n584), .o (n585) );
  assign n1646 = n585 & ~n600 ;
  assign n1647 = n1645 | n1646 ;
  assign n1648 = ~n182 & n538 ;
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  assign n1651 = ~n135 & n1650 ;
  buffer buf_n1652( .i (n1651), .o (n1652) );
  assign n1653 = n615 | n1544 ;
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n1658( .i (n898), .o (n1658) );
  assign n1659 = n368 & n1658 ;
  buffer buf_n1660( .i (n1659), .o (n1660) );
  assign n1662 = ~n1656 & n1660 ;
  buffer buf_n1663( .i (n1662), .o (n1663) );
  assign n1664 = n1652 | n1663 ;
  buffer buf_n1665( .i (n1664), .o (n1665) );
  assign n1666 = n1647 | n1665 ;
  assign n1667 = n300 & n389 ;
  buffer buf_n1668( .i (n1667), .o (n1668) );
  assign n1670 = n1473 & n1668 ;
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  assign n1673 = n424 & n1002 ;
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  assign n1677 = n1243 | n1675 ;
  assign n1678 = n1672 | n1677 ;
  assign n1679 = n1666 | n1678 ;
  assign n1680 = ~n1639 & n1679 ;
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  assign n1681 = n90 & n1586 ;
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1682( .i (n1658), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n423), .o (n1684) );
  assign n1685 = ~n1683 & n1684 ;
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  assign n1689 = n1202 | n1688 ;
  assign n1690 = n100 & n1299 ;
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  assign n1693 = n1202 & ~n1692 ;
  assign n1694 = ( n1681 & n1689 ) | ( n1681 & ~n1693 ) | ( n1689 & ~n1693 ) ;
  buffer buf_n939( .i (n938), .o (n939) );
  assign n1695 = n756 & n939 ;
  assign n1696 = n24 & ~n1067 ;
  assign n1697 = n33 | n1546 ;
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  assign n1702 = n688 & n1368 ;
  assign n1703 = ~n1699 & n1702 ;
  assign n1704 = ~n1696 & n1703 ;
  assign n1705 = n1695 | n1704 ;
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  assign n1708 = n65 & ~n1706 ;
  assign n1709 = ( n1694 & n1707 ) | ( n1694 & ~n1708 ) | ( n1707 & ~n1708 ) ;
  assign n1710 = n1680 | n1709 ;
  assign n1711 = n1582 | n1710 ;
  assign n1712 = n108 & ~n243 ;
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  assign n1716 = n862 | n1489 ;
  assign n1717 = n1715 & n1716 ;
  buffer buf_n848( .i (n847), .o (n848) );
  assign n1718 = n848 & ~n1698 ;
  buffer buf_n1719( .i (n1718), .o (n1719) );
  assign n1720 = ~n75 & n1719 ;
  assign n1721 = n1717 | n1720 ;
  assign n1722 = ~n12 & n1721 ;
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n608( .i (n607), .o (n608) );
  assign n1723 = ~n608 & n1148 ;
  assign n1724 = n222 & ~n1723 ;
  assign n1725 = n408 & n1547 ;
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  assign n1730 = n1545 & n1608 ;
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  assign n1736 = ~n848 & n1732 ;
  assign n1737 = ~n1728 & n1736 ;
  assign n1738 = n1108 & n1737 ;
  assign n1739 = ( n1109 & n1724 ) | ( n1109 & n1738 ) | ( n1724 & n1738 ) ;
  buffer buf_n1740( .i (n1332), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  assign n1742 = n1546 & ~n1741 ;
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  assign n1746 = ~n568 & n593 ;
  buffer buf_n1747( .i (n1746), .o (n1747) );
  assign n1748 = n1745 & n1747 ;
  assign n1749 = n974 & n1058 ;
  assign n1750 = n1200 & n1749 ;
  assign n1751 = ( n1201 & n1748 ) | ( n1201 & n1750 ) | ( n1748 & n1750 ) ;
  assign n1752 = n1739 | n1751 ;
  assign n1753 = ( ~n13 & n1722 ) | ( ~n13 & n1752 ) | ( n1722 & n1752 ) ;
  buffer buf_n102( .i (n101), .o (n102) );
  assign n1754 = n102 & ~n1363 ;
  buffer buf_n1755( .i (n1754), .o (n1755) );
  assign n1756 = n349 | n1527 ;
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1546), .o (n1759) );
  assign n1760 = ~n592 & n1759 ;
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  assign n1763 = ~n1758 & n1762 ;
  buffer buf_n1764( .i (n1763), .o (n1764) );
  assign n1765 = ~n1019 & n1025 ;
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  assign n1768 = ~n62 & n1767 ;
  assign n1769 = n23 & n73 ;
  buffer buf_n1770( .i (n1769), .o (n1770) );
  assign n1772 = n1095 & n1770 ;
  assign n1773 = n1768 | n1772 ;
  assign n1774 = n1764 | n1773 ;
  assign n1775 = n1755 & ~n1774 ;
  assign n1776 = ~n1753 & n1775 ;
  buffer buf_n1302( .i (n1301), .o (n1302) );
  assign n1777 = n88 | n472 ;
  assign n1778 = n1415 & ~n1777 ;
  assign n1779 = ~n1302 & n1778 ;
  assign n1780 = n72 & n229 ;
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  assign n1783 = n1490 | n1782 ;
  buffer buf_n1784( .i (n1783), .o (n1784) );
  assign n1785 = ~n354 & n1784 ;
  assign n1786 = ( ~n355 & n1779 ) | ( ~n355 & n1785 ) | ( n1779 & n1785 ) ;
  buffer buf_n1787( .i (n54), .o (n1787) );
  assign n1788 = n928 & ~n1787 ;
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n381( .i (n380), .o (n381) );
  assign n1797 = n381 & ~n1654 ;
  buffer buf_n1798( .i (n1797), .o (n1798) );
  assign n1801 = n688 & n1798 ;
  buffer buf_n1802( .i (n1801), .o (n1802) );
  assign n1803 = ~n1794 & n1802 ;
  buffer buf_n1804( .i (n1803), .o (n1804) );
  assign n1805 = n787 & n1624 ;
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n849( .i (n848), .o (n849) );
  assign n1807 = n278 & ~n849 ;
  assign n1808 = n1806 & n1807 ;
  buffer buf_n437( .i (n436), .o (n437) );
  assign n1809 = n214 & ~n437 ;
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  assign n1811 = n111 | n384 ;
  assign n1812 = n1810 & ~n1811 ;
  assign n1813 = n1808 | n1812 ;
  assign n1814 = ( ~n1796 & n1804 ) | ( ~n1796 & n1813 ) | ( n1804 & n1813 ) ;
  assign n1815 = n975 & n1300 ;
  assign n1816 = n102 | n1815 ;
  assign n1817 = ~n348 & n1024 ;
  buffer buf_n1818( .i (n1817), .o (n1818) );
  assign n1823 = n1357 & n1818 ;
  buffer buf_n1824( .i (n1823), .o (n1824) );
  assign n1825 = ~n1547 & n1608 ;
  buffer buf_n1826( .i (n1825), .o (n1826) );
  assign n1830 = ~n34 & n1826 ;
  buffer buf_n1831( .i (n1830), .o (n1831) );
  assign n1832 = ~n441 & n1831 ;
  assign n1833 = n1824 | n1832 ;
  buffer buf_n1834( .i (n1833), .o (n1834) );
  assign n1835 = n1816 | n1834 ;
  assign n1836 = n1814 | n1835 ;
  assign n1837 = n1786 | n1836 ;
  assign n1838 = ~n1776 & n1837 ;
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  assign n1839 = n455 & n986 ;
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  assign n1842 = n989 | n1002 ;
  buffer buf_n1843( .i (n1842), .o (n1843) );
  assign n1845 = n1800 & n1843 ;
  buffer buf_n1846( .i (n22), .o (n1846) );
  assign n1847 = ~n881 & n1846 ;
  assign n1848 = n742 & n1847 ;
  assign n1849 = n1242 | n1848 ;
  assign n1850 = n1845 | n1849 ;
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  assign n1851 = n399 & n891 ;
  buffer buf_n1852( .i (n1851), .o (n1852) );
  assign n1854 = n425 | n1852 ;
  assign n1855 = n883 & n1854 ;
  assign n1856 = ~n749 & n1649 ;
  buffer buf_n1857( .i (n1856), .o (n1857) );
  assign n1859 = n74 & n1857 ;
  buffer buf_n1860( .i (n1859), .o (n1860) );
  assign n1861 = n1855 | n1860 ;
  assign n1862 = n1850 | n1861 ;
  assign n1863 = n1841 | n1862 ;
  assign n1864 = n398 & n522 ;
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  assign n1869 = n903 | n1500 ;
  assign n1870 = n1868 & ~n1869 ;
  assign n1871 = n391 | n1299 ;
  assign n1872 = n1500 & n1871 ;
  buffer buf_n1129( .i (n1128), .o (n1129) );
  assign n1873 = n419 | n1129 ;
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  assign n1876 = n59 | n184 ;
  buffer buf_n1877( .i (n1876), .o (n1877) );
  assign n1883 = n768 | n1877 ;
  assign n1884 = n1874 & ~n1883 ;
  assign n1885 = n1872 | n1884 ;
  assign n1886 = n1870 | n1885 ;
  assign n1887 = n583 & n984 ;
  buffer buf_n1888( .i (n1887), .o (n1888) );
  assign n1890 = n1437 | n1888 ;
  assign n1891 = n102 & n1890 ;
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  assign n1892 = n294 & ~n1156 ;
  buffer buf_n1893( .i (n1892), .o (n1893) );
  assign n1896 = n1592 & ~n1893 ;
  assign n1897 = ~n133 & n235 ;
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  assign n1900 = ~n774 & n1899 ;
  assign n1901 = n1242 & ~n1900 ;
  assign n1902 = ~n1896 & n1901 ;
  assign n1903 = ~n1891 & n1902 ;
  assign n1904 = ~n1886 & n1903 ;
  assign n1905 = n1863 & ~n1904 ;
  buffer buf_n1853( .i (n1852), .o (n1853) );
  assign n1906 = n661 & n1853 ;
  buffer buf_n1907( .i (n1906), .o (n1907) );
  buffer buf_n1908( .i (n1907), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  assign n1911 = n1905 | n1910 ;
  assign n1912 = n1838 | n1911 ;
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  assign n1913 = ~n541 & n720 ;
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n1915( .i (n1914), .o (n1915) );
  buffer buf_n1916( .i (n1915), .o (n1916) );
  buffer buf_n1917( .i (n1916), .o (n1917) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  assign n1918 = n869 & ~n905 ;
  assign n1919 = n1917 & n1918 ;
  buffer buf_n1676( .i (n1675), .o (n1676) );
  assign n1920 = n1091 & n1676 ;
  buffer buf_n1921( .i (n1920), .o (n1921) );
  assign n1922 = ( n1093 & n1919 ) | ( n1093 & n1921 ) | ( n1919 & n1921 ) ;
  assign n1923 = n289 & ~n1759 ;
  assign n1924 = n1247 | n1923 ;
  buffer buf_n1925( .i (n1924), .o (n1925) );
  assign n1926 = ~n1331 & n1468 ;
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1934( .i (n1608), .o (n1934) );
  assign n1935 = n1927 & ~n1934 ;
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  assign n1938 = ~n134 & n165 ;
  buffer buf_n1939( .i (n1938), .o (n1939) );
  assign n1941 = n1937 & n1939 ;
  assign n1942 = n1925 & ~n1941 ;
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  assign n1945 = n911 & n1039 ;
  buffer buf_n1946( .i (n1945), .o (n1946) );
  assign n1947 = n1288 & ~n1470 ;
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  assign n1954 = n1389 & ~n1949 ;
  assign n1955 = n1946 & n1954 ;
  buffer buf_n1352( .i (n1351), .o (n1352) );
  assign n1956 = ~n738 & n1352 ;
  assign n1957 = n1800 & n1956 ;
  assign n1958 = n1955 | n1957 ;
  buffer buf_n1959( .i (n1958), .o (n1959) );
  assign n1960 = ~n1944 & n1959 ;
  assign n1961 = n430 & ~n1612 ;
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  assign n1964 = ~n612 & n1624 ;
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  assign n1967 = ~n137 & n561 ;
  assign n1968 = n1966 | n1967 ;
  assign n1969 = n1963 | n1968 ;
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n1970( .i (n36), .o (n1970) );
  buffer buf_n1971( .i (n207), .o (n1971) );
  assign n1972 = ( n88 & ~n1970 ) | ( n88 & n1971 ) | ( ~n1970 & n1971 ) ;
  assign n1973 = ~n864 & n1972 ;
  assign n1974 = n1057 & ~n1683 ;
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  assign n1977 = n73 & n787 ;
  buffer buf_n1978( .i (n1977), .o (n1978) );
  assign n1980 = n175 & ~n1978 ;
  assign n1981 = ~n1976 & n1980 ;
  assign n1982 = ~n1973 & n1981 ;
  assign n1983 = n1969 & n1982 ;
  assign n1984 = n1960 | n1983 ;
  assign n1985 = n1922 | n1984 ;
  assign n1986 = n1245 & ~n1397 ;
  buffer buf_n1987( .i (n1986), .o (n1987) );
  assign n1989 = n22 & ~n1142 ;
  assign n1990 = ~n1987 & n1989 ;
  buffer buf_n1991( .i (n1990), .o (n1991) );
  buffer buf_n480( .i (n479), .o (n480) );
  assign n1992 = n1548 & ~n1934 ;
  buffer buf_n1993( .i (n1992), .o (n1993) );
  assign n1997 = n480 | n1993 ;
  assign n1998 = n1781 | n1997 ;
  assign n1999 = n1991 | n1998 ;
  assign n2000 = n359 | n1993 ;
  assign n2001 = ~n985 & n2000 ;
  buffer buf_n2002( .i (n157), .o (n2002) );
  assign n2003 = n1129 & ~n2002 ;
  buffer buf_n2004( .i (n2003), .o (n2004) );
  assign n2008 = ~n2001 & n2004 ;
  assign n2009 = n1999 & n2008 ;
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  assign n2010 = n755 & n1322 ;
  assign n2011 = ~n922 & n1365 ;
  buffer buf_n2012( .i (n2011), .o (n2012) );
  assign n2016 = n380 & n1789 ;
  buffer buf_n2017( .i (n2016), .o (n2017) );
  assign n2020 = n2012 & n2017 ;
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  assign n2023 = n2010 | n2022 ;
  assign n2024 = n874 & n2023 ;
  assign n2025 = n2009 | n2024 ;
  assign n2026 = ~n558 & n1759 ;
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2028( .i (n2027), .o (n2028) );
  assign n2029 = n910 & ~n1759 ;
  buffer buf_n2030( .i (n2029), .o (n2030) );
  assign n2032 = n1199 & n2030 ;
  assign n2033 = n2028 | n2032 ;
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  assign n2034 = n912 & ~n1009 ;
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  assign n2035 = n448 | n1003 ;
  assign n2036 = n2034 | n2035 ;
  assign n2037 = n2033 & ~n2036 ;
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  assign n2038 = n493 | n1310 ;
  assign n2039 = n393 & n2038 ;
  assign n2040 = n2037 | n2039 ;
  assign n2041 = n2025 | n2040 ;
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  assign n2042 = n1451 & n1929 ;
  buffer buf_n2043( .i (n2042), .o (n2043) );
  assign n2046 = n378 & n2043 ;
  assign n2047 = n1332 | n1607 ;
  buffer buf_n2048( .i (n2047), .o (n2048) );
  assign n2055 = n718 & ~n2048 ;
  buffer buf_n2056( .i (n2055), .o (n2056) );
  buffer buf_n2057( .i (n2056), .o (n2057) );
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  assign n2059 = n774 | n1330 ;
  assign n2060 = n2058 & ~n2059 ;
  assign n2061 = n2046 | n2060 ;
  assign n2062 = n1553 & n1865 ;
  assign n2063 = n423 & ~n736 ;
  buffer buf_n2064( .i (n2063), .o (n2064) );
  assign n2067 = n2062 | n2064 ;
  buffer buf_n2068( .i (n2067), .o (n2068) );
  assign n2069 = ~n255 & n822 ;
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  assign n2073 = n1003 | n2071 ;
  buffer buf_n2074( .i (n390), .o (n2074) );
  assign n2075 = ~n872 & n2074 ;
  assign n2076 = n2073 & n2075 ;
  assign n2077 = n2068 | n2076 ;
  assign n2078 = n2061 | n2077 ;
  assign n2079 = ~n704 & n1085 ;
  buffer buf_n2080( .i (n2079), .o (n2080) );
  assign n2083 = n1052 & n2080 ;
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  assign n2086 = ~n1427 & n1562 ;
  assign n2087 = n1898 & n2086 ;
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2089( .i (n890), .o (n2089) );
  assign n2090 = n1826 & ~n2089 ;
  buffer buf_n2091( .i (n2090), .o (n2091) );
  assign n2092 = n1617 & n2091 ;
  assign n2093 = n2088 | n2092 ;
  assign n2094 = n2085 | n2093 ;
  assign n2095 = n813 | n1008 ;
  assign n2096 = n1259 | n2095 ;
  assign n2097 = n873 & ~n2096 ;
  assign n2098 = n1604 | n2097 ;
  assign n2099 = n2094 | n2098 ;
  assign n2100 = n2078 | n2099 ;
  assign n2101 = n2041 | n2100 ;
  assign n2102 = n1024 & n1366 ;
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  assign n2106 = n1925 | n2105 ;
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  assign n2109 = ~n1943 & n2107 ;
  assign n2110 = ( n1959 & n2108 ) | ( n1959 & n2109 ) | ( n2108 & n2109 ) ;
  buffer buf_n2005( .i (n2004), .o (n2005) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n2007( .i (n2006), .o (n2007) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n2111( .i (n87), .o (n2111) );
  assign n2112 = n1361 & ~n2111 ;
  assign n2113 = ~n350 & n1087 ;
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  assign n2116 = n2112 | n2115 ;
  buffer buf_n1249( .i (n1248), .o (n1249) );
  assign n2117 = n952 | n1249 ;
  assign n2118 = n724 & ~n2117 ;
  assign n2119 = n2116 & n2118 ;
  buffer buf_n733( .i (n732), .o (n733) );
  assign n2120 = n24 | n733 ;
  assign n2121 = n1279 & ~n2120 ;
  assign n2122 = n206 & n720 ;
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  assign n2125 = n629 & n1683 ;
  buffer buf_n2126( .i (n2125), .o (n2126) );
  assign n2127 = n2123 & n2126 ;
  assign n2128 = ( n2121 & n2124 ) | ( n2121 & n2127 ) | ( n2124 & n2127 ) ;
  assign n2129 = ~n2006 & n2128 ;
  assign n2130 = ( ~n2007 & n2119 ) | ( ~n2007 & n2129 ) | ( n2119 & n2129 ) ;
  assign n2131 = n2110 | n2130 ;
  assign n2132 = n2101 | n2131 ;
  assign n2133 = n1985 | n2132 ;
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n237( .i (n236), .o (n237) );
  assign n2134 = n237 & ~n871 ;
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  buffer buf_n2137( .i (n2136), .o (n2137) );
  buffer buf_n233( .i (n232), .o (n233) );
  assign n2138 = ~n11 & n233 ;
  assign n2139 = n2137 & n2138 ;
  buffer buf_n1390( .i (n1389), .o (n1390) );
  assign n2140 = n325 & n1207 ;
  assign n2141 = n1390 & n2140 ;
  buffer buf_n2142( .i (n2141), .o (n2142) );
  assign n2143 = n90 & n2142 ;
  assign n2144 = ( n91 & n2139 ) | ( n91 & n2143 ) | ( n2139 & n2143 ) ;
  assign n2145 = n546 & n1934 ;
  buffer buf_n2146( .i (n2145), .o (n2146) );
  assign n2148 = n1936 | n2146 ;
  buffer buf_n2149( .i (n2148), .o (n2149) );
  assign n2150 = n325 & n1176 ;
  assign n2151 = n2149 & n2150 ;
  assign n2152 = n146 | n855 ;
  assign n2153 = n2151 | n2152 ;
  assign n2154 = n985 | n1111 ;
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2155( .i (n1607), .o (n2155) );
  assign n2156 = n1740 & n2155 ;
  buffer buf_n2157( .i (n2156), .o (n2157) );
  assign n2160 = n2049 & ~n2157 ;
  buffer buf_n2161( .i (n2160), .o (n2161) );
  assign n2163 = n549 & ~n2161 ;
  assign n2164 = n2154 & n2163 ;
  assign n2165 = n675 | n926 ;
  assign n2166 = n2114 & ~n2165 ;
  assign n2167 = n2164 | n2166 ;
  assign n2168 = n2153 | n2167 ;
  assign n2169 = n925 & n1727 ;
  buffer buf_n2170( .i (n2169), .o (n2170) );
  buffer buf_n2171( .i (n24), .o (n2171) );
  assign n2172 = n2170 & n2171 ;
  assign n2173 = ~n257 & n1188 ;
  buffer buf_n2174( .i (n2173), .o (n2174) );
  assign n2177 = ~n112 & n2174 ;
  assign n2178 = ( ~n113 & n2172 ) | ( ~n113 & n2177 ) | ( n2172 & n2177 ) ;
  assign n2179 = ~n1268 & n1846 ;
  buffer buf_n2180( .i (n2179), .o (n2180) );
  assign n2181 = n574 & ~n2180 ;
  assign n2182 = ~n436 & n1025 ;
  buffer buf_n2183( .i (n2182), .o (n2183) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  assign n2185 = n1827 | n1993 ;
  assign n2186 = n2183 & ~n2185 ;
  assign n2187 = n1055 & n1349 ;
  buffer buf_n2188( .i (n2187), .o (n2188) );
  assign n2191 = ~n324 & n2188 ;
  buffer buf_n2192( .i (n2191), .o (n2192) );
  assign n2193 = n2186 | n2192 ;
  assign n2194 = n2181 | n2193 ;
  assign n2195 = n2178 | n2194 ;
  assign n2196 = n2168 | n2195 ;
  assign n2197 = n2144 | n2196 ;
  assign n2198 = n1198 & n1277 ;
  buffer buf_n2199( .i (n2198), .o (n2199) );
  assign n2201 = n612 & n942 ;
  buffer buf_n2202( .i (n2201), .o (n2202) );
  assign n2203 = n2199 & n2202 ;
  assign n2204 = n972 & n1350 ;
  buffer buf_n2205( .i (n2204), .o (n2205) );
  assign n2206 = n942 | n1656 ;
  assign n2207 = n2205 & ~n2206 ;
  buffer buf_n2208( .i (n2207), .o (n2208) );
  assign n2210 = n2203 | n2208 ;
  assign n2211 = n235 | n1055 ;
  buffer buf_n2212( .i (n2211), .o (n2212) );
  assign n2215 = n35 & n2212 ;
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n1994( .i (n1993), .o (n1994) );
  assign n2219 = n675 | n1994 ;
  assign n2220 = n2216 & ~n2219 ;
  assign n2221 = n1108 & n2149 ;
  assign n2222 = n2220 | n2221 ;
  assign n2223 = n2210 | n2222 ;
  buffer buf_n2224( .i (n1846), .o (n2224) );
  assign n2225 = ( n36 & n926 ) | ( n36 & ~n2224 ) | ( n926 & ~n2224 ) ;
  assign n2226 = n1793 | n2224 ;
  assign n2227 = ~n2225 & n2226 ;
  buffer buf_n2189( .i (n2188), .o (n2189) );
  buffer buf_n2190( .i (n2189), .o (n2190) );
  assign n2228 = ~n301 & n470 ;
  assign n2229 = ~n849 & n2228 ;
  assign n2230 = ~n2190 & n2229 ;
  assign n2231 = ~n2227 & n2230 ;
  assign n2232 = n985 & n1504 ;
  buffer buf_n2233( .i (n2232), .o (n2233) );
  assign n2234 = n692 & ~n1330 ;
  assign n2235 = n855 & ~n2234 ;
  assign n2236 = ~n2233 & n2235 ;
  assign n2237 = ~n2231 & n2236 ;
  assign n2238 = ~n2223 & n2237 ;
  assign n2239 = n14 | n2238 ;
  assign n2240 = n2197 & ~n2239 ;
  buffer buf_n2175( .i (n2174), .o (n2175) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  buffer buf_n987( .i (n986), .o (n987) );
  assign n2241 = n51 & n987 ;
  assign n2242 = n2176 | n2241 ;
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  assign n2243 = n387 & ~n1265 ;
  assign n2244 = n2242 & n2243 ;
  buffer buf_n1416( .i (n1415), .o (n1416) );
  assign n2245 = n1649 & n1791 ;
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  assign n2249 = n1691 | n2248 ;
  assign n2250 = n1416 & n2249 ;
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n2251( .i (n657), .o (n2251) );
  assign n2252 = n1007 & ~n2251 ;
  assign n2253 = ~n1727 & n2252 ;
  buffer buf_n2254( .i (n2253), .o (n2254) );
  assign n2256 = n1004 | n2254 ;
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  assign n2259 = n426 | n1118 ;
  assign n2260 = n936 & n2259 ;
  assign n2261 = ~n2257 & n2260 ;
  assign n2262 = n2250 | n2261 ;
  assign n2263 = n2244 | n2262 ;
  assign n2264 = n164 & ~n1355 ;
  buffer buf_n2265( .i (n2264), .o (n2265) );
  assign n2269 = n2002 | n2265 ;
  buffer buf_n2270( .i (n2269), .o (n2270) );
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  assign n2273 = n50 | n1149 ;
  buffer buf_n2274( .i (n2273), .o (n2274) );
  assign n2275 = n2272 & ~n2274 ;
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  assign n2276 = n393 & ~n483 ;
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  assign n2277 = ( n160 & ~n1145 ) | ( n160 & n1800 ) | ( ~n1145 & n1800 ) ;
  buffer buf_n2278( .i (n2277), .o (n2278) );
  assign n2279 = n2276 & n2278 ;
  assign n2280 = ~n2275 & n2279 ;
  assign n2281 = n431 & n1517 ;
  assign n2282 = n539 | n618 ;
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2285( .i (n1545), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  assign n2287 = n479 & ~n2286 ;
  assign n2288 = ~n2283 & n2287 ;
  buffer buf_n2289( .i (n2288), .o (n2289) );
  assign n2291 = ~n2135 & n2289 ;
  assign n2292 = n2281 | n2291 ;
  assign n2293 = ~n119 & n1088 ;
  assign n2294 = n1674 & n2293 ;
  buffer buf_n2184( .i (n2183), .o (n2184) );
  assign n2295 = n48 & n848 ;
  assign n2296 = n2071 | n2295 ;
  assign n2297 = n2184 & n2296 ;
  assign n2298 = n2294 | n2297 ;
  assign n2299 = n2292 | n2298 ;
  buffer buf_n2018( .i (n2017), .o (n2018) );
  buffer buf_n2019( .i (n2018), .o (n2019) );
  buffer buf_n2300( .i (n164), .o (n2300) );
  assign n2301 = n1128 & n2300 ;
  buffer buf_n2302( .i (n2301), .o (n2302) );
  assign n2303 = n2019 & n2302 ;
  assign n2304 = n1865 & n2070 ;
  buffer buf_n2305( .i (n2304), .o (n2305) );
  assign n2308 = n2303 | n2305 ;
  assign n2309 = n852 & n1431 ;
  buffer buf_n2310( .i (n2309), .o (n2310) );
  assign n2311 = n35 & n317 ;
  assign n2312 = n143 & n2311 ;
  assign n2313 = n2310 | n2312 ;
  assign n2314 = n2308 | n2313 ;
  assign n2315 = n1671 | n2068 ;
  assign n2316 = n2314 | n2315 ;
  assign n2317 = n2299 | n2316 ;
  assign n2318 = n2280 | n2317 ;
  assign n2319 = n2263 | n2318 ;
  assign n2320 = n2240 | n2319 ;
  assign n2321 = n156 | n1334 ;
  assign n2322 = ( n157 & ~n1328 ) | ( n157 & n2321 ) | ( ~n1328 & n2321 ) ;
  buffer buf_n2323( .i (n2322), .o (n2323) );
  assign n2326 = n1406 & ~n2323 ;
  assign n2327 = n230 & n1553 ;
  assign n2328 = n156 & n923 ;
  buffer buf_n2329( .i (n2328), .o (n2329) );
  assign n2330 = n1846 | n2329 ;
  assign n2331 = n2327 | n2330 ;
  assign n2332 = n2326 | n2331 ;
  buffer buf_n2333( .i (n2332), .o (n2333) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  assign n2335 = n230 | n1713 ;
  assign n2336 = n212 | n1741 ;
  buffer buf_n2337( .i (n2336), .o (n2337) );
  assign n2340 = n1286 & ~n1607 ;
  buffer buf_n2341( .i (n2340), .o (n2341) );
  assign n2345 = n1319 | n2341 ;
  buffer buf_n2346( .i (n2345), .o (n2346) );
  assign n2348 = n2337 & ~n2346 ;
  assign n2349 = ~n2335 & n2348 ;
  buffer buf_n2350( .i (n2349), .o (n2350) );
  buffer buf_n2351( .i (n2350), .o (n2351) );
  buffer buf_n2352( .i (n2351), .o (n2352) );
  assign n2353 = ( n109 & n293 ) | ( n109 & ~n2286 ) | ( n293 & ~n2286 ) ;
  buffer buf_n2354( .i (n2353), .o (n2354) );
  assign n2356 = n1277 | n1743 ;
  assign n2357 = n2354 | n2356 ;
  assign n2358 = n230 & n1743 ;
  assign n2359 = n127 & n879 ;
  buffer buf_n2360( .i (n2359), .o (n2360) );
  buffer buf_n2362( .i (n22), .o (n2362) );
  assign n2363 = ~n2360 & n2362 ;
  assign n2364 = ~n2358 & n2363 ;
  assign n2365 = n2357 & n2364 ;
  assign n2366 = ~n2350 & n2365 ;
  buffer buf_n2367( .i (n2366), .o (n2367) );
  assign n2368 = ( n2334 & n2352 ) | ( n2334 & ~n2367 ) | ( n2352 & ~n2367 ) ;
  buffer buf_n2369( .i (n11), .o (n2369) );
  assign n2370 = ( n1202 & n2351 ) | ( n1202 & n2369 ) | ( n2351 & n2369 ) ;
  assign n2371 = ( n1202 & n2333 ) | ( n1202 & n2369 ) | ( n2333 & n2369 ) ;
  assign n2372 = ( ~n2367 & n2370 ) | ( ~n2367 & n2371 ) | ( n2370 & n2371 ) ;
  assign n2373 = n2368 & ~n2372 ;
  assign n2374 = ~n942 & n1792 ;
  buffer buf_n2375( .i (n2374), .o (n2375) );
  assign n2376 = n100 & ~n207 ;
  assign n2377 = n2375 & n2376 ;
  assign n2378 = n777 & n1277 ;
  buffer buf_n2379( .i (n2378), .o (n2379) );
  assign n2381 = ~n825 & n1831 ;
  assign n2382 = ~n2379 & n2381 ;
  assign n2383 = n2377 | n2382 ;
  assign n2384 = ~n114 & n2383 ;
  assign n2385 = n471 | n951 ;
  assign n2386 = n2184 | n2385 ;
  buffer buf_n216( .i (n215), .o (n216) );
  assign n2387 = n216 & n1474 ;
  assign n2388 = n2386 & n2387 ;
  assign n2389 = n283 & n1456 ;
  assign n2390 = n793 & n1726 ;
  buffer buf_n2391( .i (n2390), .o (n2391) );
  assign n2392 = n1215 | n2391 ;
  buffer buf_n1269( .i (n1268), .o (n1269) );
  assign n2393 = n1269 & n2224 ;
  assign n2394 = n2392 & n2393 ;
  assign n2395 = n2389 | n2394 ;
  assign n2396 = n2388 | n2395 ;
  assign n2397 = n2384 | n2396 ;
  buffer buf_n1930( .i (n1929), .o (n1930) );
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  assign n2398 = n901 & n1412 ;
  buffer buf_n2399( .i (n198), .o (n2399) );
  assign n2400 = n2286 & n2399 ;
  assign n2401 = ~n984 & n2400 ;
  assign n2402 = n2398 | n2401 ;
  buffer buf_n2403( .i (n2402), .o (n2403) );
  buffer buf_n2404( .i (n2171), .o (n2404) );
  assign n2405 = n2403 & ~n2404 ;
  buffer buf_n2406( .i (n2300), .o (n2406) );
  assign n2407 = ~n48 & n2406 ;
  buffer buf_n2408( .i (n2407), .o (n2408) );
  assign n2411 = n594 & n2224 ;
  assign n2412 = n2408 & ~n2411 ;
  assign n2413 = n984 & n2002 ;
  buffer buf_n2414( .i (n2413), .o (n2414) );
  assign n2415 = n1931 & n2414 ;
  assign n2416 = ( n1932 & n2412 ) | ( n1932 & n2415 ) | ( n2412 & n2415 ) ;
  assign n2417 = ( n1933 & n2405 ) | ( n1933 & n2416 ) | ( n2405 & n2416 ) ;
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  assign n2418 = n109 | n1471 ;
  assign n2419 = ~n593 & n2418 ;
  buffer buf_n2420( .i (n2419), .o (n2420) );
  assign n2421 = n475 | n1422 ;
  assign n2422 = ( n476 & n2420 ) | ( n476 & n2421 ) | ( n2420 & n2421 ) ;
  assign n2423 = n886 | n2422 ;
  assign n2424 = n766 & ~n1267 ;
  assign n2425 = n612 & n2424 ;
  buffer buf_n2426( .i (n2425), .o (n2426) );
  assign n2427 = ~n867 & n2426 ;
  assign n2428 = n38 & n2427 ;
  assign n2429 = n705 & n1019 ;
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  assign n2432 = n866 & n2430 ;
  assign n2433 = ( ~n2426 & n2431 ) | ( ~n2426 & n2432 ) | ( n2431 & n2432 ) ;
  buffer buf_n2434( .i (n1970), .o (n2434) );
  assign n2435 = ~n2433 & n2434 ;
  assign n2436 = ( n2423 & n2428 ) | ( n2423 & n2435 ) | ( n2428 & n2435 ) ;
  assign n2437 = n2417 | n2436 ;
  assign n2438 = n2397 | n2437 ;
  assign n2439 = ( ~n15 & n2373 ) | ( ~n15 & n2438 ) | ( n2373 & n2438 ) ;
  assign n2440 = ~n112 & n676 ;
  assign n2441 = n432 & n2440 ;
  assign n2442 = ~n2274 & n2441 ;
  assign n2443 = n867 & n935 ;
  buffer buf_n2444( .i (n1934), .o (n2444) );
  assign n2445 = n1065 & n2444 ;
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n2448( .i (n2447), .o (n2448) );
  assign n2449 = n2443 | n2448 ;
  assign n2450 = ~n120 & n815 ;
  buffer buf_n722( .i (n721), .o (n722) );
  assign n2451 = n722 & n1177 ;
  assign n2452 = n2450 | n2451 ;
  assign n2453 = n2449 & n2452 ;
  assign n2454 = n2442 | n2453 ;
  buffer buf_n2081( .i (n2080), .o (n2081) );
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  assign n2455 = n1432 & n2081 ;
  buffer buf_n438( .i (n437), .o (n438) );
  assign n2456 = n384 & ~n438 ;
  assign n2457 = ( n2082 & n2455 ) | ( n2082 & n2456 ) | ( n2455 & n2456 ) ;
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  assign n2460 = n421 & n1600 ;
  buffer buf_n2461( .i (n2460), .o (n2461) );
  assign n2462 = n1201 | n1415 ;
  assign n2463 = n2461 & ~n2462 ;
  assign n2464 = n2459 | n2463 ;
  assign n2465 = n2454 | n2464 ;
  buffer buf_n2466( .i (n2286), .o (n2466) );
  assign n2467 = ~n2002 & n2466 ;
  buffer buf_n2468( .i (n983), .o (n2468) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  assign n2470 = ~n2467 & n2469 ;
  buffer buf_n2471( .i (n1355), .o (n2471) );
  buffer buf_n2472( .i (n2471), .o (n2472) );
  assign n2473 = ~n767 & n2472 ;
  assign n2474 = ~n1757 & n2473 ;
  assign n2475 = ( ~n1758 & n2470 ) | ( ~n1758 & n2474 ) | ( n2470 & n2474 ) ;
  buffer buf_n2476( .i (n2475), .o (n2476) );
  assign n2477 = n50 & n175 ;
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n2478( .i (n174), .o (n2478) );
  assign n2479 = n894 | n2478 ;
  assign n2480 = ( n2434 & ~n2477 ) | ( n2434 & n2479 ) | ( ~n2477 & n2479 ) ;
  assign n2481 = n2476 & n2480 ;
  buffer buf_n2482( .i (n2481), .o (n2482) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  assign n2483 = n173 & n1394 ;
  buffer buf_n2484( .i (n2483), .o (n2484) );
  buffer buf_n2485( .i (n2484), .o (n2485) );
  assign n2486 = ~n1701 & n2485 ;
  assign n2487 = n2476 | n2486 ;
  buffer buf_n2488( .i (n2487), .o (n2488) );
  assign n2489 = n2482 & ~n2488 ;
  buffer buf_n2209( .i (n2208), .o (n2209) );
  assign n2490 = n881 & n892 ;
  buffer buf_n2491( .i (n2490), .o (n2491) );
  assign n2492 = n2058 & n2491 ;
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  assign n2493 = ~n689 & n1564 ;
  assign n2494 = n1300 & n2493 ;
  assign n2495 = n2492 | n2494 ;
  assign n2496 = n2209 | n2495 ;
  assign n2497 = ~n872 & n2246 ;
  buffer buf_n2498( .i (n2497), .o (n2498) );
  buffer buf_n2499( .i (n2498), .o (n2499) );
  buffer buf_n488( .i (n487), .o (n488) );
  assign n2500 = n488 & n2074 ;
  buffer buf_n2501( .i (n2500), .o (n2501) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  assign n2502 = n49 & n882 ;
  assign n2503 = n2072 | n2502 ;
  assign n2504 = n2501 & n2503 ;
  assign n2505 = n2499 | n2504 ;
  assign n2506 = n2496 | n2505 ;
  assign n2507 = ( ~n2482 & n2488 ) | ( ~n2482 & n2506 ) | ( n2488 & n2506 ) ;
  assign n2508 = ( n2465 & ~n2489 ) | ( n2465 & n2507 ) | ( ~n2489 & n2507 ) ;
  assign n2509 = n2439 | n2508 ;
  assign n2510 = n1700 & ~n2190 ;
  buffer buf_n2511( .i (n61), .o (n2511) );
  assign n2512 = n187 & ~n2511 ;
  assign n2513 = ~n2510 & n2512 ;
  assign n2514 = ~n177 & n2513 ;
  buffer buf_n850( .i (n849), .o (n850) );
  assign n2515 = n10 | n850 ;
  buffer buf_n2213( .i (n2212), .o (n2213) );
  buffer buf_n2214( .i (n2213), .o (n2214) );
  assign n2516 = n74 | n221 ;
  assign n2517 = n2214 | n2516 ;
  assign n2518 = n2515 & ~n2517 ;
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  assign n2519 = n527 & n1531 ;
  assign n2520 = n2518 | n2519 ;
  assign n2521 = ( ~n178 & n2514 ) | ( ~n178 & n2520 ) | ( n2514 & n2520 ) ;
  buffer buf_n2306( .i (n2305), .o (n2306) );
  buffer buf_n2307( .i (n2306), .o (n2307) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  assign n2522 = n1644 & n1951 ;
  assign n2523 = n2307 | n2522 ;
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  assign n2524 = n259 | n1626 ;
  assign n2525 = n187 & n883 ;
  assign n2526 = ( n1601 & ~n2524 ) | ( n1601 & n2525 ) | ( ~n2524 & n2525 ) ;
  assign n2527 = n222 & n1474 ;
  assign n2528 = n874 & n2527 ;
  assign n2529 = n2526 | n2528 ;
  assign n2530 = n2523 | n2529 ;
  assign n2531 = n2521 | n2530 ;
  assign n2532 = ~n435 & n1055 ;
  buffer buf_n2533( .i (n2532), .o (n2533) );
  assign n2540 = n2406 & n2533 ;
  buffer buf_n2541( .i (n2540), .o (n2541) );
  buffer buf_n2542( .i (n2541), .o (n2542) );
  assign n2543 = ~n2434 & n2542 ;
  assign n2544 = n160 & n1118 ;
  assign n2545 = n1150 & n2544 ;
  assign n2546 = ( n1151 & n2543 ) | ( n1151 & n2545 ) | ( n2543 & n2545 ) ;
  assign n2547 = n1021 & ~n1728 ;
  assign n2548 = ~n2202 & n2547 ;
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  assign n2549 = n168 & ~n1747 ;
  assign n2550 = ~n2548 & n2549 ;
  assign n2551 = n647 & ~n956 ;
  buffer buf_n2552( .i (n2551), .o (n2552) );
  assign n2553 = n236 & ~n263 ;
  buffer buf_n2554( .i (n2553), .o (n2554) );
  assign n2556 = n2552 | n2554 ;
  assign n2557 = n476 & n2556 ;
  assign n2558 = n1311 & ~n1553 ;
  assign n2559 = n1591 & n2558 ;
  assign n2560 = n2192 | n2559 ;
  assign n2561 = n2557 | n2560 ;
  assign n2562 = n2550 | n2561 ;
  assign n2563 = n2546 | n2562 ;
  assign n2564 = ~n14 & n2563 ;
  buffer buf_n1878( .i (n1877), .o (n1878) );
  buffer buf_n1879( .i (n1878), .o (n1879) );
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n2565( .i (n13), .o (n2565) );
  assign n2566 = n1882 & n2565 ;
  assign n2567 = ( n2531 & n2564 ) | ( n2531 & ~n2566 ) | ( n2564 & ~n2566 ) ;
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  assign n2568 = ~n1416 & n2461 ;
  buffer buf_n2569( .i (n2285), .o (n2569) );
  assign n2570 = n289 & n2569 ;
  assign n2571 = n2103 & n2570 ;
  buffer buf_n2572( .i (n2571), .o (n2572) );
  buffer buf_n2573( .i (n2572), .o (n2573) );
  buffer buf_n2574( .i (n2573), .o (n2574) );
  assign n2575 = ~n77 & n2574 ;
  assign n2576 = ( ~n78 & n2568 ) | ( ~n78 & n2575 ) | ( n2568 & n2575 ) ;
  buffer buf_n2290( .i (n2289), .o (n2290) );
  assign n2577 = n76 | n2290 ;
  assign n2578 = n398 & n546 ;
  buffer buf_n2579( .i (n2578), .o (n2579) );
  buffer buf_n2580( .i (n2579), .o (n2580) );
  buffer buf_n2581( .i (n2580), .o (n2581) );
  assign n2582 = ~n645 & n2581 ;
  assign n2583 = n2302 & n2391 ;
  buffer buf_n2584( .i (n2583), .o (n2584) );
  assign n2585 = n2582 | n2584 ;
  assign n2586 = n2577 | n2585 ;
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  assign n2587 = n1129 & ~n2050 ;
  buffer buf_n2588( .i (n2587), .o (n2588) );
  buffer buf_n2589( .i (n2588), .o (n2589) );
  assign n2590 = n2255 & n2589 ;
  assign n2591 = n411 | n1650 ;
  buffer buf_n2592( .i (n2591), .o (n2592) );
  assign n2593 = n1256 & n2592 ;
  buffer buf_n2594( .i (n2593), .o (n2594) );
  assign n2595 = n2590 | n2594 ;
  assign n2596 = n2586 | n2595 ;
  assign n2597 = n2576 | n2596 ;
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n2598( .i (n880), .o (n2598) );
  assign n2599 = ~n311 & n2598 ;
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2158( .i (n2157), .o (n2158) );
  buffer buf_n2159( .i (n2158), .o (n2159) );
  assign n2601 = n925 & n2406 ;
  assign n2602 = n2159 | n2601 ;
  assign n2603 = n2600 | n2602 ;
  assign n2604 = n1340 | n2603 ;
  assign n2605 = n280 & n789 ;
  assign n2606 = n816 & ~n2605 ;
  assign n2607 = n2604 & n2606 ;
  buffer buf_n2608( .i (n2607), .o (n2608) );
  buffer buf_n2361( .i (n2360), .o (n2361) );
  assign n2609 = n2361 & n2580 ;
  assign n2610 = n75 & ~n2609 ;
  assign n2611 = n1134 & n1930 ;
  buffer buf_n2612( .i (n2155), .o (n2612) );
  assign n2613 = ~n1741 & n2612 ;
  buffer buf_n2614( .i (n2613), .o (n2614) );
  assign n2617 = ~n256 & n1367 ;
  assign n2618 = n2614 & n2617 ;
  buffer buf_n2619( .i (n2618), .o (n2619) );
  assign n2620 = n2611 | n2619 ;
  assign n2621 = n2610 & ~n2620 ;
  assign n2622 = n1035 & ~n2111 ;
  assign n2623 = n631 & n1674 ;
  assign n2624 = n2622 | n2623 ;
  assign n2625 = n2621 & ~n2624 ;
  buffer buf_n2626( .i (n847), .o (n2626) );
  assign n2627 = n568 & n2626 ;
  buffer buf_n2628( .i (n2627), .o (n2628) );
  assign n2629 = n2375 | n2628 ;
  assign n2630 = ~n1264 & n2629 ;
  assign n2631 = n2458 | n2630 ;
  assign n2632 = n2625 & ~n2631 ;
  assign n2633 = ~n2608 & n2632 ;
  assign n2634 = n2597 & ~n2633 ;
  assign n2635 = n2567 | n2634 ;
  assign n2636 = n1106 | n1683 ;
  buffer buf_n2637( .i (n2636), .o (n2637) );
  assign n2638 = n653 & n2637 ;
  buffer buf_n2639( .i (n157), .o (n2639) );
  assign n2640 = ~n1143 & n2639 ;
  buffer buf_n2641( .i (n2640), .o (n2641) );
  assign n2642 = n894 & n2641 ;
  assign n2643 = n2638 | n2642 ;
  assign n2644 = ~n39 & n2643 ;
  buffer buf_n2645( .i (n1527), .o (n2645) );
  assign n2646 = n1020 & n2645 ;
  buffer buf_n2647( .i (n2646), .o (n2647) );
  buffer buf_n2648( .i (n2647), .o (n2648) );
  buffer buf_n2649( .i (n111), .o (n2649) );
  assign n2650 = n896 & n2649 ;
  assign n2651 = n2648 & n2650 ;
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  assign n2652 = n239 & ~n690 ;
  assign n2653 = ~n827 & n2652 ;
  assign n2654 = n2651 | n2653 ;
  assign n2655 = ( ~n40 & n2644 ) | ( ~n40 & n2654 ) | ( n2644 & n2654 ) ;
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n2656( .i (n2362), .o (n2656) );
  assign n2657 = ~n302 & n2656 ;
  assign n2658 = n1729 & n2657 ;
  assign n2659 = ~n176 & n2658 ;
  assign n2660 = ~n1386 & n2233 ;
  assign n2661 = ( ~n1387 & n2659 ) | ( ~n1387 & n2660 ) | ( n2659 & n2660 ) ;
  assign n2662 = n565 & n1185 ;
  buffer buf_n2663( .i (n2662), .o (n2663) );
  assign n2668 = n924 | n2663 ;
  buffer buf_n2669( .i (n2668), .o (n2669) );
  assign n2672 = n474 & ~n524 ;
  assign n2673 = n474 & n524 ;
  assign n2674 = ( n2669 & ~n2672 ) | ( n2669 & n2673 ) | ( ~n2672 & n2673 ) ;
  buffer buf_n2675( .i (n2674), .o (n2675) );
  buffer buf_n2676( .i (n2675), .o (n2676) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  assign n2677 = n1566 & ~n2404 ;
  assign n2678 = n2676 & n2677 ;
  assign n2679 = n2661 | n2678 ;
  assign n2680 = n2655 | n2679 ;
  buffer buf_n2681( .i (n2565), .o (n2681) );
  assign n2682 = n2680 & ~n2681 ;
  buffer buf_n1979( .i (n1978), .o (n1979) );
  assign n2683 = n807 | n1979 ;
  assign n2684 = n543 & ~n1149 ;
  assign n2685 = n8 & n185 ;
  buffer buf_n2686( .i (n2685), .o (n2686) );
  assign n2688 = n1414 & ~n2686 ;
  assign n2689 = n2684 & n2688 ;
  assign n2690 = n2683 & n2689 ;
  buffer buf_n2691( .i (n1086), .o (n2691) );
  assign n2692 = n437 & n2691 ;
  buffer buf_n2693( .i (n2692), .o (n2693) );
  assign n2694 = n1618 & n2693 ;
  assign n2695 = n1478 | n2088 ;
  assign n2696 = n2694 | n2695 ;
  assign n2697 = n358 & ~n369 ;
  buffer buf_n2698( .i (n2697), .o (n2698) );
  buffer buf_n2699( .i (n2698), .o (n2699) );
  assign n2700 = n1120 & ~n2699 ;
  buffer buf_n2701( .i (n1354), .o (n2701) );
  assign n2702 = ~n686 & n2701 ;
  buffer buf_n2703( .i (n2702), .o (n2703) );
  buffer buf_n2704( .i (n2703), .o (n2704) );
  buffer buf_n2705( .i (n2704), .o (n2705) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  assign n2706 = n1527 | n2444 ;
  buffer buf_n2707( .i (n2706), .o (n2707) );
  assign n2709 = n2284 | n2707 ;
  assign n2710 = n2705 & ~n2709 ;
  assign n2711 = n2700 | n2710 ;
  assign n2712 = n2696 | n2711 ;
  assign n2713 = n2690 | n2712 ;
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n2162( .i (n2161), .o (n2162) );
  assign n2714 = n609 | n2162 ;
  assign n2715 = n1012 | n2362 ;
  buffer buf_n2716( .i (n2715), .o (n2716) );
  assign n2718 = n237 & n2626 ;
  buffer buf_n2719( .i (n2718), .o (n2719) );
  assign n2720 = n2716 & ~n2719 ;
  assign n2721 = n2714 & n2720 ;
  assign n2722 = ~n111 & n1495 ;
  assign n2723 = ~n2716 & n2722 ;
  assign n2724 = n73 & ~n620 ;
  buffer buf_n2725( .i (n2724), .o (n2725) );
  buffer buf_n2342( .i (n2341), .o (n2342) );
  buffer buf_n2343( .i (n2342), .o (n2343) );
  buffer buf_n2344( .i (n2343), .o (n2344) );
  assign n2728 = n130 & ~n2344 ;
  assign n2729 = n2725 & ~n2728 ;
  assign n2730 = ~n2723 & n2729 ;
  assign n2731 = ~n2721 & n2730 ;
  assign n2732 = n142 | n2579 ;
  assign n2733 = n512 & n2732 ;
  buffer buf_n2734( .i (n2733), .o (n2734) );
  buffer buf_n2735( .i (n611), .o (n2735) );
  buffer buf_n2736( .i (n1001), .o (n2736) );
  assign n2737 = n2735 | n2736 ;
  buffer buf_n2738( .i (n2737), .o (n2738) );
  assign n2740 = n2057 & ~n2698 ;
  assign n2741 = ~n2738 & n2740 ;
  assign n2742 = n2734 | n2741 ;
  assign n2743 = ~n495 & n1686 ;
  buffer buf_n439( .i (n438), .o (n439) );
  assign n2744 = ~n439 & n2247 ;
  assign n2745 = n2743 | n2744 ;
  assign n2746 = n2742 | n2745 ;
  assign n2747 = n2731 | n2746 ;
  assign n2748 = n2713 | n2747 ;
  buffer buf_n2749( .i (n717), .o (n2749) );
  buffer buf_n2750( .i (n2749), .o (n2750) );
  buffer buf_n2751( .i (n2750), .o (n2751) );
  assign n2752 = n933 & n2751 ;
  buffer buf_n2753( .i (n2752), .o (n2753) );
  buffer buf_n2754( .i (n2753), .o (n2754) );
  buffer buf_n2755( .i (n2754), .o (n2755) );
  buffer buf_n2756( .i (n2755), .o (n2756) );
  assign n2757 = n903 | n1975 ;
  assign n2758 = n1175 & ~n2362 ;
  buffer buf_n2759( .i (n2758), .o (n2759) );
  assign n2760 = n2511 | n2759 ;
  assign n2761 = n2757 & ~n2760 ;
  buffer buf_n1661( .i (n1660), .o (n1661) );
  assign n2762 = n862 | n1661 ;
  buffer buf_n2763( .i (n2762), .o (n2763) );
  buffer buf_n2764( .i (n2763), .o (n2764) );
  assign n2765 = n2761 | n2764 ;
  buffer buf_n2380( .i (n2379), .o (n2380) );
  assign n2766 = ( ~n51 & n2380 ) | ( ~n51 & n2754 ) | ( n2380 & n2754 ) ;
  assign n2767 = n52 & n2766 ;
  assign n2768 = ( n2756 & n2765 ) | ( n2756 & n2767 ) | ( n2765 & n2767 ) ;
  buffer buf_n2347( .i (n2346), .o (n2347) );
  assign n2769 = n1949 & ~n2347 ;
  buffer buf_n2770( .i (n2769), .o (n2770) );
  buffer buf_n2771( .i (n2770), .o (n2771) );
  assign n2772 = ~n229 & n956 ;
  buffer buf_n2773( .i (n2772), .o (n2773) );
  buffer buf_n2774( .i (n2773), .o (n2774) );
  buffer buf_n2775( .i (n2774), .o (n2775) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  assign n2776 = n1829 | n2431 ;
  assign n2777 = n2775 & ~n2776 ;
  assign n2778 = ~n2771 & n2777 ;
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n2779 = ~n61 & n1130 ;
  assign n2780 = ~n649 & n1625 ;
  assign n2781 = ( ~n650 & n2779 ) | ( ~n650 & n2780 ) | ( n2779 & n2780 ) ;
  buffer buf_n2782( .i (n2781), .o (n2782) );
  buffer buf_n2783( .i (n2782), .o (n2783) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n958( .i (n957), .o (n958) );
  assign n2784 = ~n958 & n1564 ;
  assign n2785 = ~n231 & n1625 ;
  assign n2786 = ~n2784 & n2785 ;
  assign n2787 = n1735 & ~n2786 ;
  assign n2788 = n2782 & n2787 ;
  assign n2789 = ( n2778 & n2783 ) | ( n2778 & n2788 ) | ( n2783 & n2788 ) ;
  assign n2790 = n2768 | n2789 ;
  assign n2791 = n2748 | n2790 ;
  assign n2792 = n2682 | n2791 ;
  assign n2793 = n794 | n2736 ;
  buffer buf_n2794( .i (n2793), .o (n2794) );
  buffer buf_n2795( .i (n2794), .o (n2795) );
  assign n2796 = n113 & n2795 ;
  buffer buf_n1102( .i (n1101), .o (n1102) );
  assign n2797 = n987 | n1102 ;
  assign n2798 = n2796 | n2797 ;
  assign n2799 = n89 & n1701 ;
  assign n2800 = n768 | n1473 ;
  assign n2801 = n1447 & ~n2800 ;
  buffer buf_n2802( .i (n2801), .o (n2802) );
  assign n2803 = ~n2799 & n2802 ;
  assign n2804 = n2798 & n2803 ;
  assign n2805 = ~n731 & n1623 ;
  buffer buf_n2806( .i (n2805), .o (n2806) );
  buffer buf_n2807( .i (n2806), .o (n2807) );
  buffer buf_n2808( .i (n2807), .o (n2808) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  assign n2809 = n1376 & ~n2170 ;
  assign n2810 = n2628 & n2807 ;
  assign n2811 = ( n2808 & ~n2809 ) | ( n2808 & n2810 ) | ( ~n2809 & n2810 ) ;
  buffer buf_n2812( .i (n2811), .o (n2812) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n2687( .i (n2686), .o (n2687) );
  buffer buf_n449( .i (n448), .o (n449) );
  assign n2813 = n449 & ~n1515 ;
  assign n2814 = ~n2687 & n2813 ;
  assign n2815 = n1445 & n2814 ;
  assign n2816 = n2812 | n2815 ;
  assign n2817 = n2804 | n2816 ;
  buffer buf_n2818( .i (n34), .o (n2818) );
  assign n2819 = n1792 & ~n2818 ;
  buffer buf_n2820( .i (n2819), .o (n2820) );
  assign n2824 = n1719 | n2820 ;
  buffer buf_n2825( .i (n72), .o (n2825) );
  assign n2826 = n2639 & n2825 ;
  buffer buf_n2827( .i (n2826), .o (n2827) );
  buffer buf_n2828( .i (n2827), .o (n2828) );
  buffer buf_n2829( .i (n925), .o (n2829) );
  assign n2830 = n1728 & ~n2829 ;
  assign n2831 = n2827 & n2830 ;
  assign n2832 = ( n2824 & n2828 ) | ( n2824 & n2831 ) | ( n2828 & n2831 ) ;
  assign n2833 = n1762 & n2126 ;
  buffer buf_n913( .i (n912), .o (n913) );
  assign n2834 = n360 | n594 ;
  assign n2835 = n913 | n2834 ;
  assign n2836 = ~n2833 & n2835 ;
  assign n2837 = ~n2832 & n2836 ;
  assign n2838 = n405 & ~n2837 ;
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  assign n2839 = n739 | n1079 ;
  buffer buf_n2840( .i (n33), .o (n2840) );
  assign n2841 = n2399 & ~n2840 ;
  buffer buf_n2842( .i (n2841), .o (n2842) );
  buffer buf_n2843( .i (n2842), .o (n2843) );
  assign n2844 = n986 | n2843 ;
  assign n2845 = ( n1080 & n2839 ) | ( n1080 & ~n2844 ) | ( n2839 & ~n2844 ) ;
  assign n2846 = ~n27 & n2845 ;
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  assign n2847 = n118 & ~n2406 ;
  buffer buf_n2848( .i (n2847), .o (n2848) );
  assign n2849 = n2180 & n2848 ;
  assign n2850 = n1132 & ~n2849 ;
  assign n2851 = n810 & ~n2848 ;
  assign n2852 = n159 | n265 ;
  assign n2853 = n676 & ~n2852 ;
  assign n2854 = n2851 | n2853 ;
  assign n2855 = n2850 & ~n2854 ;
  assign n2856 = ~n2846 & n2855 ;
  assign n2857 = n2838 | n2856 ;
  assign n2858 = n2817 | n2857 ;
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n2670( .i (n2669), .o (n2670) );
  buffer buf_n2671( .i (n2670), .o (n2671) );
  assign n2859 = n1015 & n2671 ;
  assign n2860 = n49 & ~n902 ;
  assign n2861 = n232 & ~n2860 ;
  assign n2862 = ~n914 & n2861 ;
  assign n2863 = ( ~n915 & n2859 ) | ( ~n915 & n2862 ) | ( n2859 & n2862 ) ;
  assign n2864 = n1487 | n2420 ;
  buffer buf_n2865( .i (n2864), .o (n2865) );
  assign n2866 = ( ~n232 & n526 ) | ( ~n232 & n1555 ) | ( n526 & n1555 ) ;
  assign n2867 = n233 & n2866 ;
  assign n2868 = ( n528 & n2865 ) | ( n528 & n2867 ) | ( n2865 & n2867 ) ;
  assign n2869 = n2863 | n2868 ;
  assign n2870 = ~n356 & n2869 ;
  buffer buf_n2065( .i (n2064), .o (n2065) );
  buffer buf_n2066( .i (n2065), .o (n2066) );
  assign n2871 = ~n76 & n2066 ;
  assign n2872 = n130 & n1179 ;
  assign n2873 = n1965 & n2872 ;
  buffer buf_n1858( .i (n1857), .o (n1858) );
  assign n2874 = ~n690 & n1858 ;
  assign n2875 = n2873 | n2874 ;
  assign n2876 = n2871 | n2875 ;
  assign n2877 = n236 & ~n1411 ;
  buffer buf_n2878( .i (n2877), .o (n2878) );
  buffer buf_n2879( .i (n2878), .o (n2879) );
  assign n2880 = n2725 & n2879 ;
  buffer buf_n1940( .i (n1939), .o (n1940) );
  assign n2881 = n525 & ~n1994 ;
  assign n2882 = n1940 & n2881 ;
  assign n2883 = n2880 | n2882 ;
  assign n2884 = ~n530 & n1684 ;
  buffer buf_n2885( .i (n2884), .o (n2885) );
  assign n2888 = n276 & ~n2300 ;
  buffer buf_n2889( .i (n2888), .o (n2889) );
  assign n2890 = n689 & n2889 ;
  assign n2891 = n2885 & n2890 ;
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  assign n2892 = n361 & n1552 ;
  assign n2893 = n400 & n2703 ;
  buffer buf_n2894( .i (n2893), .o (n2894) );
  buffer buf_n2895( .i (n360), .o (n2895) );
  assign n2896 = ( n1552 & n2894 ) | ( n1552 & n2895 ) | ( n2894 & n2895 ) ;
  assign n2897 = ( n2891 & ~n2892 ) | ( n2891 & n2896 ) | ( ~n2892 & n2896 ) ;
  assign n2898 = n2883 | n2897 ;
  assign n2899 = n2876 | n2898 ;
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  buffer buf_n1821( .i (n1820), .o (n1821) );
  buffer buf_n1822( .i (n1821), .o (n1822) );
  assign n2900 = n778 | n1148 ;
  assign n2901 = ~n608 & n778 ;
  assign n2902 = ( n2174 & n2900 ) | ( n2174 & ~n2901 ) | ( n2900 & ~n2901 ) ;
  buffer buf_n2903( .i (n2902), .o (n2903) );
  assign n2904 = n1822 & n2903 ;
  assign n2905 = ~n186 & n207 ;
  assign n2906 = ~n850 & n2905 ;
  assign n2907 = n205 | n2089 ;
  buffer buf_n2908( .i (n2907), .o (n2908) );
  buffer buf_n2909( .i (n2908), .o (n2909) );
  assign n2911 = n258 & n721 ;
  assign n2912 = ~n2909 & n2911 ;
  assign n2913 = n2906 | n2912 ;
  buffer buf_n2914( .i (n6), .o (n2914) );
  assign n2915 = n2471 & n2914 ;
  buffer buf_n2916( .i (n2915), .o (n2916) );
  buffer buf_n2917( .i (n2916), .o (n2917) );
  assign n2918 = ~n238 & n1144 ;
  assign n2919 = n9 & ~n2916 ;
  assign n2920 = ( ~n2917 & n2918 ) | ( ~n2917 & n2919 ) | ( n2918 & n2919 ) ;
  assign n2921 = n176 & ~n2920 ;
  assign n2922 = n2913 & n2921 ;
  assign n2923 = n2904 | n2922 ;
  assign n2924 = n2899 | n2923 ;
  assign n2925 = n2870 | n2924 ;
  assign n2926 = n2858 | n2925 ;
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n2927( .i (n186), .o (n2927) );
  buffer buf_n2928( .i (n1241), .o (n2928) );
  assign n2929 = n2927 | n2928 ;
  assign n2930 = n1875 & ~n2929 ;
  assign n2931 = n588 | n2930 ;
  assign n2932 = ~n598 & n2931 ;
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  buffer buf_n651( .i (n650), .o (n651) );
  assign n2933 = ~n2343 & n2645 ;
  buffer buf_n2934( .i (n2933), .o (n2934) );
  buffer buf_n2935( .i (n2934), .o (n2935) );
  assign n2936 = n651 | n2935 ;
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n2937( .i (n49), .o (n2937) );
  assign n2938 = n734 & n2937 ;
  assign n2939 = n2935 & n2938 ;
  assign n2940 = ( ~n2054 & n2936 ) | ( ~n2054 & n2939 ) | ( n2936 & n2939 ) ;
  buffer buf_n678( .i (n677), .o (n678) );
  assign n2941 = n138 & ~n393 ;
  assign n2942 = n678 | n2941 ;
  assign n2943 = n2940 & ~n2942 ;
  assign n2944 = n2932 | n2943 ;
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  assign n2945 = ( ~n681 & n2159 ) | ( ~n681 & n2656 ) | ( n2159 & n2656 ) ;
  assign n2946 = n453 | n2945 ;
  assign n2947 = n237 & ~n2639 ;
  buffer buf_n2948( .i (n2444), .o (n2948) );
  assign n2949 = n607 & n2948 ;
  assign n2950 = n2947 | n2949 ;
  assign n2951 = ~n168 & n2950 ;
  assign n2952 = n2946 & ~n2951 ;
  buffer buf_n2953( .i (n2952), .o (n2953) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  assign n2954 = n263 & n1623 ;
  buffer buf_n2955( .i (n2954), .o (n2955) );
  buffer buf_n2956( .i (n2955), .o (n2956) );
  buffer buf_n2957( .i (n2956), .o (n2957) );
  assign n2958 = ~n2589 & n2957 ;
  assign n2959 = ~n1458 & n2958 ;
  assign n2960 = ~n2953 & n2959 ;
  assign n2961 = n754 & n1351 ;
  buffer buf_n2962( .i (n2961), .o (n2962) );
  buffer buf_n2963( .i (n2962), .o (n2963) );
  assign n2964 = n2171 & n2962 ;
  assign n2965 = ( ~n2403 & n2963 ) | ( ~n2403 & n2964 ) | ( n2963 & n2964 ) ;
  buffer buf_n2966( .i (n2965), .o (n2966) );
  buffer buf_n2967( .i (n2966), .o (n2967) );
  assign n2968 = n2960 | n2967 ;
  assign n2969 = n2944 | n2968 ;
  assign n2970 = n618 | n1741 ;
  buffer buf_n2971( .i (n2970), .o (n2971) );
  assign n2975 = n1175 & ~n2971 ;
  buffer buf_n2976( .i (n2975), .o (n2976) );
  assign n2978 = n810 & n2976 ;
  assign n2979 = n146 | n2310 ;
  assign n2980 = n2978 | n2979 ;
  buffer buf_n2981( .i (n1727), .o (n2981) );
  assign n2982 = n1699 & ~n2981 ;
  assign n2983 = n2894 & n2982 ;
  assign n2984 = n269 & n2056 ;
  assign n2985 = n2021 | n2984 ;
  buffer buf_n2986( .i (n2985), .o (n2986) );
  assign n2987 = n2983 | n2986 ;
  assign n2988 = n2980 | n2987 ;
  assign n2989 = n213 & n1289 ;
  buffer buf_n2990( .i (n2989), .o (n2990) );
  assign n2992 = n2806 & n2990 ;
  assign n2993 = ~n619 & n847 ;
  buffer buf_n2994( .i (n2993), .o (n2994) );
  assign n2995 = n1245 | n2285 ;
  buffer buf_n2996( .i (n2995), .o (n2996) );
  assign n2999 = ~n732 & n2996 ;
  assign n3000 = n2994 & n2999 ;
  assign n3001 = n2992 | n3000 ;
  assign n3002 = n2466 & n2614 ;
  assign n3003 = n1372 & n3002 ;
  assign n3004 = n629 & ~n2598 ;
  assign n3005 = n1866 & n3004 ;
  assign n3006 = n3003 | n3005 ;
  assign n3007 = n3001 | n3006 ;
  assign n3008 = n1840 | n3007 ;
  assign n3009 = n2988 | n3008 ;
  assign n3010 = n1451 & ~n1563 ;
  assign n3011 = ~n1199 & n3010 ;
  assign n3012 = n1914 & n3011 ;
  buffer buf_n318( .i (n317), .o (n318) );
  assign n3013 = n318 | n1111 ;
  assign n3014 = n426 & n3013 ;
  assign n3015 = n3012 | n3014 ;
  assign n3016 = n772 | n2914 ;
  buffer buf_n3017( .i (n3016), .o (n3017) );
  buffer buf_n3018( .i (n3017), .o (n3018) );
  assign n3019 = ~n2161 & n2981 ;
  assign n3020 = ~n3018 & n3019 ;
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  assign n3021 = ~n1258 & n2691 ;
  buffer buf_n3022( .i (n3021), .o (n3022) );
  assign n3023 = n752 & n3022 ;
  assign n3024 = n3020 | n3023 ;
  assign n3025 = n3015 | n3024 ;
  assign n3026 = n1231 | n1831 ;
  assign n3027 = n749 & n2399 ;
  buffer buf_n3028( .i (n3027), .o (n3028) );
  buffer buf_n3029( .i (n3028), .o (n3029) );
  assign n3030 = n3026 & n3029 ;
  assign n3031 = n1991 & n2753 ;
  assign n3032 = n3030 | n3031 ;
  assign n3033 = n338 | n594 ;
  buffer buf_n3034( .i (n109), .o (n3034) );
  buffer buf_n3035( .i (n3034), .o (n3035) );
  assign n3036 = ( ~n87 & n951 ) | ( ~n87 & n3035 ) | ( n951 & n3035 ) ;
  assign n3037 = ~n3033 & n3036 ;
  buffer buf_n3038( .i (n235), .o (n3038) );
  assign n3039 = n72 & n3038 ;
  buffer buf_n3040( .i (n3039), .o (n3040) );
  buffer buf_n3041( .i (n3040), .o (n3041) );
  buffer buf_n3043( .i (n1682), .o (n3043) );
  buffer buf_n3044( .i (n3043), .o (n3044) );
  assign n3045 = n2994 & n3044 ;
  assign n3046 = n3041 & n3045 ;
  assign n3047 = n3037 | n3046 ;
  assign n3048 = n3032 | n3047 ;
  assign n3049 = n3025 | n3048 ;
  assign n3050 = n3009 | n3049 ;
  buffer buf_n1578( .i (n1577), .o (n1578) );
  assign n3051 = ~n542 & n2469 ;
  buffer buf_n3052( .i (n3051), .o (n3052) );
  buffer buf_n3053( .i (n3052), .o (n3053) );
  assign n3054 = ~n2903 & n3053 ;
  assign n3055 = ~n1578 & n3054 ;
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  buffer buf_n3056( .i (n1740), .o (n3056) );
  buffer buf_n3057( .i (n3056), .o (n3057) );
  assign n3058 = ~n2444 & n3057 ;
  buffer buf_n3059( .i (n3058), .o (n3059) );
  buffer buf_n3060( .i (n3059), .o (n3060) );
  assign n3061 = n439 & ~n3060 ;
  buffer buf_n2991( .i (n2990), .o (n2991) );
  assign n3062 = ~n2895 & n2991 ;
  assign n3063 = ~n3061 & n3062 ;
  assign n3064 = ~n1895 & n3063 ;
  assign n3065 = n816 & n2734 ;
  assign n3066 = n1200 & n2588 ;
  assign n3067 = n996 & n3066 ;
  assign n3068 = n3065 | n3067 ;
  assign n3069 = n3064 | n3068 ;
  assign n3070 = n3055 | n3069 ;
  assign n3071 = n3050 | n3070 ;
  assign n3072 = n2969 | n3071 ;
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n2664( .i (n2663), .o (n2664) );
  assign n3073 = n1428 | n2664 ;
  buffer buf_n3074( .i (n3073), .o (n3074) );
  buffer buf_n3075( .i (n3074), .o (n3075) );
  buffer buf_n3076( .i (n3075), .o (n3076) );
  assign n3077 = n1950 & n2759 ;
  assign n3078 = ~n774 & n1828 ;
  assign n3079 = n2408 | n3078 ;
  assign n3080 = n3077 | n3079 ;
  assign n3081 = n3076 & ~n3080 ;
  assign n3082 = n125 & ~n1978 ;
  assign n3083 = n1236 & ~n3082 ;
  buffer buf_n1291( .i (n1290), .o (n1291) );
  assign n3084 = n225 & ~n1291 ;
  buffer buf_n3085( .i (n3084), .o (n3085) );
  assign n3086 = ~n118 & n797 ;
  buffer buf_n3087( .i (n3086), .o (n3087) );
  assign n3090 = ~n294 & n506 ;
  assign n3091 = n61 | n3090 ;
  assign n3092 = n3087 | n3091 ;
  assign n3093 = n3085 | n3092 ;
  assign n3094 = n3083 | n3093 ;
  assign n3095 = ~n3081 & n3094 ;
  buffer buf_n1567( .i (n1566), .o (n1567) );
  assign n3096 = n1232 & ~n2928 ;
  assign n3097 = ~n542 & n788 ;
  assign n3098 = n1108 & n3097 ;
  assign n3099 = n3096 | n3098 ;
  assign n3100 = ~n1567 & n3099 ;
  buffer buf_n3042( .i (n3041), .o (n3042) );
  buffer buf_n2355( .i (n2354), .o (n2355) );
  assign n3101 = ~n631 & n2355 ;
  assign n3102 = n3042 & ~n3101 ;
  buffer buf_n2910( .i (n2909), .o (n2910) );
  assign n3103 = n1200 & n2058 ;
  assign n3104 = n2910 & n3103 ;
  assign n3105 = n3102 | n3104 ;
  assign n3106 = n3100 | n3105 ;
  assign n3107 = n3095 | n3106 ;
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  assign n3108 = ~n1022 & n2111 ;
  assign n3109 = n76 & n3108 ;
  assign n3110 = ( n77 & n2218 ) | ( n77 & n3109 ) | ( n2218 & n3109 ) ;
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n2997( .i (n2996), .o (n2997) );
  buffer buf_n2998( .i (n2997), .o (n2998) );
  buffer buf_n3111( .i (n2818), .o (n3111) );
  assign n3112 = ~n649 & n3111 ;
  assign n3113 = n2998 & ~n3112 ;
  assign n3114 = n2770 | n3113 ;
  assign n3115 = ~n1403 & n3114 ;
  assign n3116 = ~n3110 & n3115 ;
  buffer buf_n1282( .i (n1281), .o (n1282) );
  assign n3117 = ~n1282 & n1770 ;
  assign n3118 = ~n1951 & n3117 ;
  assign n3119 = n159 & n1248 ;
  assign n3120 = n614 & n3119 ;
  assign n3121 = n63 & ~n3120 ;
  assign n3122 = ~n3118 & n3121 ;
  buffer buf_n3123( .i (n2369), .o (n3123) );
  assign n3124 = n3122 | n3123 ;
  assign n3125 = ( n2565 & ~n3116 ) | ( n2565 & n3124 ) | ( ~n3116 & n3124 ) ;
  assign n3126 = n3107 & ~n3125 ;
  assign n3127 = n2058 & n2174 ;
  assign n3128 = n1247 & n1368 ;
  buffer buf_n3129( .i (n3128), .o (n3129) );
  assign n3130 = n2170 & n3129 ;
  assign n3131 = n3127 | n3130 ;
  assign n3132 = n1672 | n3131 ;
  buffer buf_n3133( .i (n1127), .o (n3133) );
  buffer buf_n3134( .i (n3133), .o (n3134) );
  assign n3135 = n1498 & n3134 ;
  buffer buf_n3136( .i (n3135), .o (n3136) );
  assign n3137 = n789 & n3136 ;
  buffer buf_n3138( .i (n3137), .o (n3138) );
  buffer buf_n1889( .i (n1888), .o (n1889) );
  assign n3139 = ~n1090 & n1889 ;
  assign n3140 = n3138 | n3139 ;
  assign n3141 = n3132 | n3140 ;
  buffer buf_n2886( .i (n2885), .o (n2886) );
  buffer buf_n2887( .i (n2886), .o (n2887) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  assign n3142 = n2267 | n2414 ;
  buffer buf_n3143( .i (n592), .o (n3143) );
  buffer buf_n3144( .i (n3143), .o (n3144) );
  assign n3145 = n1564 & n3144 ;
  assign n3146 = ~n560 & n733 ;
  assign n3147 = n3145 | n3146 ;
  assign n3148 = n3142 | n3147 ;
  assign n3149 = n2887 & ~n3148 ;
  assign n3150 = n350 | n2466 ;
  buffer buf_n3151( .i (n3150), .o (n3151) );
  assign n3152 = n855 & ~n3151 ;
  assign n3153 = n1326 | n3152 ;
  assign n3154 = n1931 & n2600 ;
  assign n3155 = n1398 & n1791 ;
  buffer buf_n3156( .i (n3155), .o (n3156) );
  assign n3157 = n2552 | n3156 ;
  buffer buf_n3158( .i (n3157), .o (n3158) );
  assign n3159 = n3154 | n3158 ;
  assign n3160 = n3153 & n3159 ;
  assign n3161 = n3149 | n3160 ;
  assign n3162 = n3141 | n3161 ;
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2325( .i (n2324), .o (n2325) );
  buffer buf_n2013( .i (n2012), .o (n2013) );
  buffer buf_n2014( .i (n2013), .o (n2014) );
  buffer buf_n2015( .i (n2014), .o (n2015) );
  assign n3163 = n1395 & ~n2014 ;
  assign n3164 = ( n1437 & ~n2015 ) | ( n1437 & n3163 ) | ( ~n2015 & n3163 ) ;
  assign n3165 = n2325 & n3164 ;
  buffer buf_n3166( .i (n3165), .o (n3166) );
  buffer buf_n3167( .i (n3166), .o (n3167) );
  buffer buf_n3168( .i (n74), .o (n3168) );
  assign n3169 = n810 | n3168 ;
  buffer buf_n2972( .i (n2971), .o (n2972) );
  buffer buf_n2973( .i (n2972), .o (n2973) );
  assign n3170 = n682 & ~n2973 ;
  assign n3171 = n3169 & n3170 ;
  buffer buf_n3172( .i (n117), .o (n3172) );
  buffer buf_n3173( .i (n1367), .o (n3173) );
  assign n3174 = ~n3172 & n3173 ;
  assign n3175 = n2878 & n3174 ;
  buffer buf_n3176( .i (n3175), .o (n3176) );
  buffer buf_n3177( .i (n3176), .o (n3177) );
  assign n3178 = n3171 | n3177 ;
  assign n3179 = ~n63 & n2542 ;
  buffer buf_n2974( .i (n2973), .o (n2974) );
  buffer buf_n3180( .i (n901), .o (n3180) );
  assign n3181 = n481 & n3180 ;
  assign n3182 = n1592 | n3181 ;
  assign n3183 = ~n2974 & n3182 ;
  assign n3184 = n3179 | n3183 ;
  assign n3185 = n3178 | n3184 ;
  assign n3186 = n3167 | n3185 ;
  assign n3187 = n3162 | n3186 ;
  assign n3188 = n3126 | n3187 ;
  buffer buf_n795( .i (n794), .o (n795) );
  assign n3189 = n768 | n795 ;
  assign n3190 = n1794 & ~n3189 ;
  assign n3191 = n2491 & n2649 ;
  buffer buf_n3192( .i (n2649), .o (n3192) );
  assign n3193 = ( n3190 & n3191 ) | ( n3190 & n3192 ) | ( n3191 & n3192 ) ;
  buffer buf_n3194( .i (n3180), .o (n3194) );
  assign n3195 = ~n913 & n3194 ;
  buffer buf_n1124( .i (n1123), .o (n1124) );
  assign n3196 = ~n313 & n1124 ;
  assign n3197 = n3195 | n3196 ;
  assign n3198 = n3193 | n3197 ;
  assign n3199 = n405 & n3198 ;
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  assign n3200 = n1489 | n1761 ;
  assign n3201 = ~n352 & n3200 ;
  assign n3202 = ~n129 & n750 ;
  buffer buf_n3203( .i (n777), .o (n3203) );
  assign n3204 = n3202 & n3203 ;
  assign n3205 = n2162 & n3204 ;
  assign n3206 = n3201 | n3205 ;
  assign n3207 = ~n1476 & n3206 ;
  buffer buf_n3208( .i (n172), .o (n3208) );
  buffer buf_n3209( .i (n3208), .o (n3209) );
  assign n3210 = n1241 & n3209 ;
  assign n3211 = ~n3151 & n3210 ;
  assign n3212 = n399 & n2399 ;
  buffer buf_n3213( .i (n3212), .o (n3213) );
  assign n3215 = n2091 & n3213 ;
  assign n3216 = n1970 & ~n3215 ;
  assign n3217 = ~n3211 & n3216 ;
  assign n3218 = n399 & ~n731 ;
  buffer buf_n3219( .i (n3218), .o (n3219) );
  buffer buf_n3221( .i (n2472), .o (n3221) );
  assign n3222 = n3219 & ~n3221 ;
  assign n3223 = n608 & n3028 ;
  assign n3224 = ( n609 & n3222 ) | ( n609 & n3223 ) | ( n3222 & n3223 ) ;
  assign n3225 = n1965 & n2414 ;
  assign n3226 = n3224 | n3225 ;
  assign n3227 = n3217 & ~n3226 ;
  assign n3228 = ~n3207 & n3227 ;
  assign n3229 = ~n3199 & n3228 ;
  buffer buf_n1844( .i (n1843), .o (n1844) );
  assign n3230 = n1844 & n2589 ;
  assign n3231 = n1970 | n2084 ;
  assign n3232 = n3176 | n3231 ;
  assign n3233 = n3230 | n3232 ;
  buffer buf_n3220( .i (n3219), .o (n3220) );
  assign n3234 = n87 | n2469 ;
  assign n3235 = n3220 & ~n3234 ;
  assign n3236 = n680 & ~n3034 ;
  buffer buf_n3237( .i (n397), .o (n3237) );
  buffer buf_n3238( .i (n3237), .o (n3238) );
  buffer buf_n3239( .i (n3238), .o (n3239) );
  assign n3240 = n2468 & n3239 ;
  assign n3241 = n3236 & n3240 ;
  assign n3242 = n257 & n1247 ;
  assign n3243 = n1043 & n3242 ;
  assign n3244 = n3241 | n3243 ;
  assign n3245 = n3235 | n3244 ;
  assign n3246 = ~n704 & n931 ;
  buffer buf_n3247( .i (n3246), .o (n3247) );
  assign n3250 = ~n1462 & n3247 ;
  buffer buf_n3251( .i (n3250), .o (n3251) );
  assign n3252 = n1222 & n3213 ;
  assign n3253 = n3251 | n3252 ;
  assign n3254 = n900 & n1450 ;
  buffer buf_n3255( .i (n3254), .o (n3255) );
  assign n3258 = n2302 & n3255 ;
  buffer buf_n3259( .i (n1548), .o (n3259) );
  assign n3260 = ~n1610 & n3259 ;
  buffer buf_n3261( .i (n3260), .o (n3261) );
  assign n3263 = n1939 & n3261 ;
  assign n3264 = n3258 | n3263 ;
  assign n3265 = n3253 | n3264 ;
  assign n3266 = n3245 | n3265 ;
  assign n3267 = n3233 | n3266 ;
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  assign n3268 = n1595 | n1663 ;
  assign n3269 = n751 & n3040 ;
  assign n3270 = n3136 | n3269 ;
  assign n3271 = n3268 | n3270 ;
  assign n3272 = ~n1244 & n3271 ;
  assign n3273 = n401 & n3035 ;
  buffer buf_n3274( .i (n3273), .o (n3274) );
  assign n3275 = n613 & n1003 ;
  buffer buf_n3276( .i (n3275), .o (n3276) );
  assign n3277 = n3274 & n3276 ;
  assign n3278 = ( n3052 & n3274 ) | ( n3052 & n3276 ) | ( n3274 & n3276 ) ;
  assign n3279 = ( ~n2903 & n3277 ) | ( ~n2903 & n3278 ) | ( n3277 & n3278 ) ;
  assign n3280 = n3272 | n3279 ;
  assign n3281 = n3267 | n3280 ;
  assign n3282 = ~n3229 & n3281 ;
  assign n3283 = ~n351 & n3044 ;
  buffer buf_n3284( .i (n3283), .o (n3284) );
  assign n3285 = n266 | n1313 ;
  assign n3286 = n3284 & ~n3285 ;
  assign n3287 = n421 & n595 ;
  assign n3288 = n1601 & n3287 ;
  assign n3289 = n3286 | n3288 ;
  assign n3290 = n1427 & ~n1791 ;
  buffer buf_n3291( .i (n3290), .o (n3291) );
  buffer buf_n3292( .i (n3291), .o (n3292) );
  buffer buf_n3293( .i (n3292), .o (n3293) );
  assign n3294 = ~n894 & n2111 ;
  assign n3295 = ~n3293 & n3294 ;
  buffer buf_n2665( .i (n2664), .o (n2665) );
  buffer buf_n2666( .i (n2665), .o (n2666) );
  buffer buf_n2667( .i (n2666), .o (n2667) );
  buffer buf_n3296( .i (n3111), .o (n3296) );
  assign n3297 = ~n259 & n3296 ;
  assign n3298 = n2667 | n3297 ;
  assign n3299 = n3295 | n3298 ;
  assign n3300 = n3289 & n3299 ;
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  buffer buf_n2977( .i (n2976), .o (n2977) );
  assign n3301 = n868 & n2977 ;
  assign n3302 = n487 & n1641 ;
  buffer buf_n3303( .i (n3302), .o (n3303) );
  buffer buf_n3304( .i (n3303), .o (n3304) );
  assign n3305 = n392 & n1191 ;
  assign n3306 = n3304 | n3305 ;
  assign n3307 = n3301 | n3306 ;
  assign n3308 = n1953 & n3307 ;
  assign n3309 = n3300 | n3308 ;
  buffer buf_n3088( .i (n3087), .o (n3088) );
  buffer buf_n3089( .i (n3088), .o (n3089) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  assign n3310 = n353 | n1146 ;
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  assign n3311 = n121 & ~n709 ;
  assign n3312 = ( n3089 & ~n3310 ) | ( n3089 & n3311 ) | ( ~n3310 & n3311 ) ;
  assign n3313 = n2966 | n3312 ;
  buffer buf_n562( .i (n561), .o (n562) );
  assign n3314 = ~n562 & n1015 ;
  buffer buf_n3315( .i (n3314), .o (n3315) );
  assign n3316 = n445 & n3315 ;
  assign n3317 = n3313 | n3316 ;
  assign n3318 = n3309 | n3317 ;
  assign n3319 = n3282 | n3318 ;
  buffer buf_n2534( .i (n2533), .o (n2534) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  buffer buf_n2536( .i (n2535), .o (n2536) );
  buffer buf_n2537( .i (n2536), .o (n2537) );
  buffer buf_n2538( .i (n2537), .o (n2538) );
  buffer buf_n2539( .i (n2538), .o (n2539) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n2821( .i (n2820), .o (n2821) );
  buffer buf_n2822( .i (n2821), .o (n2822) );
  buffer buf_n2823( .i (n2822), .o (n2823) );
  assign n3320 = n39 | n2822 ;
  assign n3321 = ( n2258 & n2823 ) | ( n2258 & n3320 ) | ( n2823 & n3320 ) ;
  assign n3322 = n2539 & n3321 ;
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n295( .i (n294), .o (n295) );
  assign n3323 = n295 & ~n1744 ;
  assign n3324 = n130 & ~n2829 ;
  assign n3325 = ( n927 & n3323 ) | ( n927 & ~n3324 ) | ( n3323 & ~n3324 ) ;
  buffer buf_n3326( .i (n3325), .o (n3326) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n3327( .i (n2645), .o (n3327) );
  buffer buf_n3328( .i (n3327), .o (n3328) );
  assign n3329 = n2927 & ~n3328 ;
  assign n3330 = ~n1271 & n3329 ;
  assign n3331 = n3326 & n3330 ;
  assign n3332 = ~n1794 & n2649 ;
  assign n3333 = n384 & n795 ;
  buffer buf_n3334( .i (n3333), .o (n3334) );
  assign n3335 = ~n3332 & n3334 ;
  assign n3336 = n1628 & n3335 ;
  assign n3337 = ( n1629 & n3331 ) | ( n1629 & n3336 ) | ( n3331 & n3336 ) ;
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  assign n3338 = n1370 & n2928 ;
  buffer buf_n3339( .i (n3338), .o (n3339) );
  buffer buf_n3340( .i (n3339), .o (n3340) );
  assign n3341 = n233 & ~n1525 ;
  buffer buf_n3342( .i (n3341), .o (n3342) );
  assign n3343 = ~n620 & n2212 ;
  buffer buf_n3344( .i (n3343), .o (n3344) );
  buffer buf_n3345( .i (n3344), .o (n3345) );
  assign n3346 = n595 | n789 ;
  assign n3347 = n3345 | n3346 ;
  assign n3348 = n3339 & ~n3347 ;
  assign n3349 = ( n3340 & n3342 ) | ( n3340 & n3348 ) | ( n3342 & n3348 ) ;
  assign n3350 = n3337 | n3349 ;
  assign n3351 = n3322 | n3350 ;
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  assign n3352 = ~n1434 & n1951 ;
  assign n3353 = ( n1435 & n1632 ) | ( n1435 & ~n3352 ) | ( n1632 & ~n3352 ) ;
  buffer buf_n2726( .i (n2725), .o (n2726) );
  buffer buf_n2727( .i (n2726), .o (n2727) );
  assign n3354 = n2274 | n2727 ;
  assign n3355 = n3353 & ~n3354 ;
  buffer buf_n3356( .i (n1793), .o (n3356) );
  assign n3357 = n2541 & ~n3356 ;
  assign n3358 = n2986 | n3357 ;
  assign n3359 = n266 & n2484 ;
  buffer buf_n3360( .i (n924), .o (n3360) );
  assign n3361 = ~n1948 & n3360 ;
  buffer buf_n3362( .i (n3361), .o (n3362) );
  assign n3363 = n1853 & n3362 ;
  assign n3364 = n3359 | n3363 ;
  assign n3365 = n3358 | n3364 ;
  assign n3366 = ~n682 & n2928 ;
  assign n3367 = ~n649 & n1053 ;
  assign n3368 = n1281 | n1799 ;
  assign n3369 = n3367 & ~n3368 ;
  assign n3370 = ~n3366 & n3369 ;
  assign n3371 = n1179 & n1852 ;
  assign n3372 = n1824 | n3371 ;
  buffer buf_n3373( .i (n591), .o (n3373) );
  assign n3374 = n647 & ~n3373 ;
  buffer buf_n3375( .i (n3374), .o (n3375) );
  assign n3378 = n1866 & n3375 ;
  assign n3379 = ~n1360 & n1781 ;
  assign n3380 = n3378 | n3379 ;
  assign n3381 = n3372 | n3380 ;
  assign n3382 = n3370 | n3381 ;
  assign n3383 = n3365 | n3382 ;
  assign n3384 = n3355 | n3383 ;
  assign n3385 = n1271 & n1962 ;
  assign n3386 = n3034 | n3143 ;
  buffer buf_n3387( .i (n3386), .o (n3387) );
  assign n3388 = n3344 & ~n3387 ;
  assign n3389 = n1053 | n1642 ;
  buffer buf_n1657( .i (n1656), .o (n1657) );
  assign n3390 = n1657 & n3059 ;
  assign n3391 = n3389 & n3390 ;
  assign n3392 = n3388 | n3391 ;
  assign n3393 = n3385 | n3392 ;
  assign n3394 = n1953 & n3393 ;
  buffer buf_n2555( .i (n2554), .o (n2555) );
  assign n3395 = n2555 | n3328 ;
  assign n3396 = n401 | n1766 ;
  assign n3397 = ~n481 & n768 ;
  assign n3398 = n3396 & n3397 ;
  assign n3399 = n3395 & n3398 ;
  buffer buf_n2031( .i (n2030), .o (n2031) );
  buffer buf_n3400( .i (n628), .o (n3400) );
  assign n3401 = n2468 & ~n3400 ;
  assign n3402 = ~n448 & n3401 ;
  assign n3403 = ~n2031 & n3402 ;
  assign n3404 = ~n459 & n3403 ;
  assign n3405 = n3399 | n3404 ;
  assign n3406 = n1131 | n1802 ;
  assign n3407 = n1949 & n2446 ;
  assign n3408 = ~n2976 & n3407 ;
  assign n3409 = n3406 & n3408 ;
  assign n3410 = n659 | n1732 ;
  assign n3411 = ~n3017 & n3410 ;
  assign n3412 = n8 & ~n511 ;
  assign n3413 = ~n1877 & n3412 ;
  assign n3414 = n3411 | n3413 ;
  buffer buf_n3415( .i (n1241), .o (n3415) );
  assign n3416 = ~n570 & n3415 ;
  assign n3417 = n3414 & n3416 ;
  assign n3418 = n3409 | n3417 ;
  assign n3419 = n3405 | n3418 ;
  assign n3420 = n3394 | n3419 ;
  assign n3421 = n3384 | n3420 ;
  assign n3422 = n3351 | n3421 ;
  buffer buf_n2200( .i (n2199), .o (n2200) );
  buffer buf_n3423( .i (n2057), .o (n3423) );
  assign n3424 = ~n708 & n3423 ;
  assign n3425 = ~n2200 & n3424 ;
  assign n3426 = n3059 | n3327 ;
  assign n3427 = n221 & n3035 ;
  assign n3428 = n3426 & ~n3427 ;
  buffer buf_n2615( .i (n2614), .o (n2615) );
  assign n3429 = n549 | n2615 ;
  assign n3430 = n1810 & ~n3429 ;
  assign n3431 = ~n3428 & n3430 ;
  assign n3432 = n3425 | n3431 ;
  assign n3433 = n1806 & n3362 ;
  buffer buf_n3434( .i (n3433), .o (n3434) );
  assign n3435 = n650 | n2082 ;
  buffer buf_n1343( .i (n1342), .o (n1343) );
  assign n3436 = n622 | n1343 ;
  assign n3437 = n3435 & ~n3436 ;
  assign n3438 = n3434 | n3437 ;
  assign n3439 = n3432 | n3438 ;
  assign n3440 = ~n1150 & n2501 ;
  assign n3441 = n1004 | n1112 ;
  assign n3442 = n427 & n3441 ;
  assign n3443 = n3440 | n3442 ;
  assign n3444 = n542 | n1569 ;
  buffer buf_n3445( .i (n3444), .o (n3445) );
  assign n3446 = ~n449 & n666 ;
  assign n3447 = n3445 & n3446 ;
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  assign n3448 = n376 & n1691 ;
  assign n3449 = n3447 | n3448 ;
  assign n3450 = n3443 | n3449 ;
  assign n3451 = n3439 | n3450 ;
  buffer buf_n1438( .i (n1437), .o (n1438) );
  assign n3452 = n138 & ~n1438 ;
  buffer buf_n3453( .i (n3452), .o (n3453) );
  assign n3454 = n1205 & n3038 ;
  buffer buf_n3455( .i (n3454), .o (n3455) );
  buffer buf_n3456( .i (n3455), .o (n3456) );
  buffer buf_n3457( .i (n3456), .o (n3457) );
  assign n3458 = n1243 & n3457 ;
  assign n3459 = n588 | n3458 ;
  assign n3460 = ~n3453 & n3459 ;
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  assign n3461 = n266 | n1453 ;
  assign n3462 = n1627 & ~n3461 ;
  assign n3463 = n2410 & n3462 ;
  assign n3464 = n873 & ~n3328 ;
  assign n3465 = ~n1014 & n1118 ;
  assign n3466 = n3464 & n3465 ;
  buffer buf_n2717( .i (n2716), .o (n2717) );
  assign n3467 = n693 & n830 ;
  assign n3468 = ~n2717 & n3467 ;
  assign n3469 = n3466 | n3468 ;
  assign n3470 = n3463 | n3469 ;
  assign n3471 = n3460 | n3470 ;
  assign n3472 = n3451 | n3471 ;
  buffer buf_n3473( .i (n3168), .o (n3473) );
  assign n3474 = ( n51 & n3192 ) | ( n51 & ~n3473 ) | ( n3192 & ~n3473 ) ;
  buffer buf_n3475( .i (n3035), .o (n3475) );
  assign n3476 = ( n2937 & ~n3328 ) | ( n2937 & n3475 ) | ( ~n3328 & n3475 ) ;
  assign n3477 = n3284 & ~n3476 ;
  assign n3478 = n3474 & n3477 ;
  buffer buf_n3479( .i (n1013), .o (n3479) );
  assign n3480 = n595 & n3479 ;
  buffer buf_n3481( .i (n430), .o (n3481) );
  assign n3482 = n2693 & n3481 ;
  assign n3483 = ~n3480 & n3482 ;
  buffer buf_n2616( .i (n2615), .o (n2616) );
  assign n3484 = n1946 & n2616 ;
  assign n3485 = n3445 & n3484 ;
  assign n3486 = n3483 | n3485 ;
  assign n3487 = n3478 | n3486 ;
  buffer buf_n3488( .i (n607), .o (n3488) );
  assign n3489 = n958 | n3488 ;
  assign n3490 = n3129 & ~n3489 ;
  assign n3491 = n1117 & n2205 ;
  assign n3492 = n628 & ~n1731 ;
  buffer buf_n3493( .i (n3492), .o (n3493) );
  assign n3495 = n2955 & n3493 ;
  assign n3496 = n3491 | n3495 ;
  assign n3497 = n3490 | n3496 ;
  buffer buf_n1669( .i (n1668), .o (n1669) );
  assign n3498 = n1565 & n1669 ;
  assign n3499 = n853 & n1866 ;
  assign n3500 = n829 & n938 ;
  assign n3501 = n3499 | n3500 ;
  assign n3502 = n3498 | n3501 ;
  assign n3503 = n3497 | n3502 ;
  assign n3504 = n651 & n1860 ;
  assign n3505 = n1352 & ~n3209 ;
  assign n3506 = n2699 | n3505 ;
  buffer buf_n3494( .i (n3493), .o (n3494) );
  assign n3507 = n302 & n401 ;
  assign n3508 = ( n402 & n3494 ) | ( n402 & n3507 ) | ( n3494 & n3507 ) ;
  assign n3509 = n3506 & n3508 ;
  assign n3510 = n3504 | n3509 ;
  assign n3511 = n3503 | n3510 ;
  assign n3512 = n3487 | n3511 ;
  buffer buf_n489( .i (n488), .o (n489) );
  assign n3513 = n489 & ~n2774 ;
  assign n3514 = n551 & n2171 ;
  assign n3515 = ( n2404 & n3513 ) | ( n2404 & n3514 ) | ( n3513 & n3514 ) ;
  buffer buf_n3516( .i (n1199), .o (n3516) );
  assign n3517 = n3296 | n3516 ;
  buffer buf_n3518( .i (n2656), .o (n3518) );
  assign n3519 = ( ~n1089 & n3296 ) | ( ~n1089 & n3518 ) | ( n3296 & n3518 ) ;
  assign n3520 = n3517 & ~n3519 ;
  assign n3521 = n3515 | n3520 ;
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  assign n3522 = ~n935 & n1131 ;
  assign n3523 = ~n1096 & n3522 ;
  assign n3524 = ~n2045 & n3523 ;
  assign n3525 = n3521 & n3524 ;
  buffer buf_n3256( .i (n3255), .o (n3256) );
  buffer buf_n3257( .i (n3256), .o (n3257) );
  assign n3526 = ~n614 & n3475 ;
  assign n3527 = n3257 & ~n3526 ;
  assign n3528 = n167 & n238 ;
  assign n3529 = ( n239 & ~n3387 ) | ( n239 & n3528 ) | ( ~n3387 & n3528 ) ;
  assign n3530 = n894 & n2267 ;
  assign n3531 = n3529 | n3530 ;
  assign n3532 = n3527 | n3531 ;
  assign n3533 = ~n625 & n3532 ;
  assign n3534 = n3525 | n3533 ;
  assign n3535 = n3512 | n3534 ;
  assign n3536 = n3472 | n3535 ;
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  assign n3537 = n2339 & ~n2879 ;
  buffer buf_n3538( .i (n3537), .o (n3538) );
  buffer buf_n2739( .i (n2738), .o (n2739) );
  assign n3539 = n1914 & n2934 ;
  assign n3540 = n2739 & n3539 ;
  assign n3541 = ~n3538 & n3540 ;
  buffer buf_n3376( .i (n3375), .o (n3376) );
  buffer buf_n3377( .i (n3376), .o (n3377) );
  assign n3542 = n427 & ~n3377 ;
  buffer buf_n1294( .i (n1293), .o (n1294) );
  assign n3543 = n371 | n849 ;
  buffer buf_n3544( .i (n3543), .o (n3544) );
  assign n3545 = n1294 | n3544 ;
  buffer buf_n169( .i (n168), .o (n169) );
  assign n3546 = ~n169 & n3544 ;
  assign n3547 = ( n3542 & ~n3545 ) | ( n3542 & n3546 ) | ( ~n3545 & n3546 ) ;
  assign n3548 = n3541 | n3547 ;
  buffer buf_n3214( .i (n3213), .o (n3214) );
  assign n3549 = ~n2511 & n3214 ;
  assign n3550 = n167 & ~n351 ;
  assign n3551 = n482 & n3550 ;
  assign n3552 = n3549 | n3551 ;
  assign n3553 = n572 & n3552 ;
  assign n3554 = n1118 | n1669 ;
  buffer buf_n3555( .i (n3554), .o (n3555) );
  buffer buf_n3556( .i (n3044), .o (n3556) );
  assign n3557 = ~n676 & n3556 ;
  buffer buf_n3558( .i (n3415), .o (n3558) );
  assign n3559 = n3557 & ~n3558 ;
  assign n3560 = n3555 & n3559 ;
  assign n3561 = n3553 | n3560 ;
  assign n3562 = n3548 | n3561 ;
  assign n3563 = n233 & ~n1614 ;
  assign n3564 = ~n1265 & n3563 ;
  assign n3565 = ~n2953 & n3564 ;
  buffer buf_n1010( .i (n1009), .o (n1010) );
  assign n3566 = ~n1010 & n1867 ;
  buffer buf_n3567( .i (n1726), .o (n3567) );
  assign n3568 = n3360 & ~n3567 ;
  assign n3569 = n3219 & n3568 ;
  assign n3570 = n3028 & n3455 ;
  assign n3571 = n3569 | n3570 ;
  assign n3572 = n3566 | n3571 ;
  buffer buf_n3573( .i (n224), .o (n3573) );
  assign n3574 = n143 & n3573 ;
  assign n3575 = n3251 | n3574 ;
  assign n3576 = n2498 | n3575 ;
  assign n3577 = n3572 | n3576 ;
  assign n3578 = n1232 | n1719 ;
  assign n3579 = n1066 | n1106 ;
  assign n3580 = n1369 & ~n3579 ;
  assign n3581 = n2619 | n3580 ;
  assign n3582 = n3578 & n3581 ;
  assign n3583 = n2414 & ~n2927 ;
  assign n3584 = n1966 & n3583 ;
  assign n3585 = n3582 | n3584 ;
  assign n3586 = n3577 | n3585 ;
  assign n3587 = n3565 | n3586 ;
  assign n3588 = n3562 | n3587 ;
  buffer buf_n3589( .i (n686), .o (n3589) );
  buffer buf_n3590( .i (n3589), .o (n3590) );
  assign n3591 = n3043 & ~n3590 ;
  assign n3592 = ( ~n167 & n1761 ) | ( ~n167 & n3591 ) | ( n1761 & n3591 ) ;
  assign n3593 = ~n216 & n3592 ;
  buffer buf_n1988( .i (n1987), .o (n1988) );
  assign n3594 = n1988 & n2338 ;
  assign n3595 = ~n1538 & n3594 ;
  assign n3596 = ( ~n1539 & n3593 ) | ( ~n1539 & n3595 ) | ( n3593 & n3595 ) ;
  assign n3597 = ( n188 & n1192 ) | ( n188 & n2404 ) | ( n1192 & n2404 ) ;
  assign n3598 = n3596 | n3597 ;
  assign n3599 = n532 & n1729 ;
  assign n3600 = ~n779 & n2820 ;
  assign n3601 = ( ~n780 & n3599 ) | ( ~n780 & n3600 ) | ( n3599 & n3600 ) ;
  buffer buf_n1995( .i (n1994), .o (n1995) );
  buffer buf_n1996( .i (n1995), .o (n1996) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  buffer buf_n3602( .i (n893), .o (n3602) );
  assign n3603 = n1995 | n3602 ;
  assign n3604 = ( n1996 & n2268 ) | ( n1996 & n3603 ) | ( n2268 & n3603 ) ;
  assign n3605 = n3601 | n3604 ;
  assign n3606 = n3598 & n3605 ;
  assign n3607 = n986 & n1515 ;
  assign n3608 = ~n2675 & n3607 ;
  assign n3609 = n2216 & ~n3387 ;
  assign n3610 = n1761 & n2159 ;
  assign n3611 = n3303 | n3610 ;
  assign n3612 = n3609 | n3611 ;
  assign n3613 = n3608 | n3612 ;
  assign n3614 = ~n1953 & n3613 ;
  assign n3615 = n3606 | n3614 ;
  assign n3616 = n493 | n3602 ;
  assign n3617 = n385 & ~n2637 ;
  assign n3618 = n3616 & n3617 ;
  assign n3619 = n2344 | n3221 ;
  buffer buf_n1337( .i (n1336), .o (n1337) );
  assign n3620 = n1337 & n2027 ;
  assign n3621 = n3619 & n3620 ;
  assign n3622 = n1013 | n1248 ;
  assign n3623 = ~n767 & n2691 ;
  assign n3624 = ~n1699 & n3623 ;
  assign n3625 = n3622 & n3624 ;
  assign n3626 = n3621 | n3625 ;
  assign n3627 = n3618 | n3626 ;
  assign n3628 = n481 & n2842 ;
  assign n3629 = n359 & n2691 ;
  assign n3630 = ~n1148 & n3629 ;
  assign n3631 = n3628 | n3630 ;
  buffer buf_n2147( .i (n2146), .o (n2147) );
  assign n3632 = n2147 & ~n2908 ;
  assign n3633 = n2270 & n3632 ;
  assign n3634 = ( ~n2910 & n3631 ) | ( ~n2910 & n3633 ) | ( n3631 & n3633 ) ;
  assign n3635 = n282 & n3156 ;
  assign n3636 = ~n290 & n1026 ;
  buffer buf_n3637( .i (n1948), .o (n3637) );
  assign n3638 = n3636 & ~n3637 ;
  assign n3639 = n3635 | n3638 ;
  buffer buf_n3640( .i (n2937), .o (n3640) );
  assign n3641 = n3639 & n3640 ;
  assign n3642 = n3634 | n3641 ;
  assign n3643 = n3627 | n3642 ;
  assign n3644 = ~n2565 & n3643 ;
  assign n3645 = ( ~n2681 & n3615 ) | ( ~n2681 & n3644 ) | ( n3615 & n3644 ) ;
  assign n3646 = n3588 | n3645 ;
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  assign n3647 = n1510 & n2719 ;
  assign n3648 = ~n2338 & n3291 ;
  assign n3649 = ~n1020 & n1311 ;
  assign n3650 = n2889 & n3649 ;
  assign n3651 = n3648 | n3650 ;
  assign n3652 = n3647 | n3651 ;
  buffer buf_n3653( .i (n1187), .o (n3653) );
  assign n3654 = ~n506 & n3653 ;
  assign n3655 = n248 & n3654 ;
  assign n3656 = n702 & n3655 ;
  assign n3657 = ~n311 & n950 ;
  assign n3658 = n2773 & n3657 ;
  assign n3659 = n3022 | n3658 ;
  assign n3660 = n3656 | n3659 ;
  assign n3661 = n3652 | n3660 ;
  assign n3662 = ~n3123 & n3661 ;
  assign n3663 = n2379 & ~n3041 ;
  assign n3664 = n227 | n3663 ;
  buffer buf_n240( .i (n239), .o (n240) );
  assign n3665 = n238 & ~n630 ;
  buffer buf_n3666( .i (n3038), .o (n3666) );
  buffer buf_n3667( .i (n3666), .o (n3667) );
  assign n3668 = ( n630 & n2469 ) | ( n630 & ~n3667 ) | ( n2469 & ~n3667 ) ;
  assign n3669 = ( n2794 & ~n3665 ) | ( n2794 & n3668 ) | ( ~n3665 & n3668 ) ;
  assign n3670 = n240 & n3669 ;
  assign n3671 = ( n633 & n3664 ) | ( n633 & n3670 ) | ( n3664 & n3670 ) ;
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n3672( .i (n1240), .o (n3672) );
  assign n3673 = n2889 & n3672 ;
  buffer buf_n3674( .i (n3673), .o (n3674) );
  assign n3675 = ( n527 & n1771 ) | ( n527 & n3674 ) | ( n1771 & n3674 ) ;
  buffer buf_n3676( .i (n523), .o (n3676) );
  buffer buf_n3677( .i (n3676), .o (n3677) );
  buffer buf_n3678( .i (n3677), .o (n3678) );
  buffer buf_n3679( .i (n3678), .o (n3679) );
  assign n3680 = ( n267 & n3674 ) | ( n267 & n3679 ) | ( n3674 & n3679 ) ;
  assign n3681 = n3675 & ~n3680 ;
  assign n3682 = n3671 | n3681 ;
  buffer buf_n3683( .i (n3123), .o (n3683) );
  assign n3684 = ( n3662 & n3682 ) | ( n3662 & ~n3683 ) | ( n3682 & ~n3683 ) ;
  assign n3685 = n571 & ~n1220 ;
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  assign n3686 = ~n1496 & n1800 ;
  assign n3687 = n1419 | n3686 ;
  assign n3688 = n3685 | n3687 ;
  buffer buf_n3689( .i (n3518), .o (n3689) );
  assign n3690 = n1475 & n3689 ;
  buffer buf_n3262( .i (n3261), .o (n3262) );
  assign n3691 = n1270 & ~n3262 ;
  buffer buf_n3692( .i (n3691), .o (n3692) );
  assign n3693 = ~n3690 & n3692 ;
  assign n3694 = n3688 & n3693 ;
  buffer buf_n303( .i (n302), .o (n303) );
  assign n3695 = n303 | n2895 ;
  buffer buf_n2708( .i (n2707), .o (n2708) );
  buffer buf_n246( .i (n245), .o (n246) );
  assign n3696 = ~n246 & n1107 ;
  assign n3697 = n2708 & n3696 ;
  assign n3698 = n3695 & n3697 ;
  buffer buf_n3699( .i (n2825), .o (n3699) );
  assign n3700 = ( n825 & ~n3667 ) | ( n825 & n3699 ) | ( ~n3667 & n3699 ) ;
  assign n3701 = ( n549 & n3667 ) | ( n549 & ~n3699 ) | ( n3667 & ~n3699 ) ;
  assign n3702 = n3700 & n3701 ;
  buffer buf_n3248( .i (n3247), .o (n3248) );
  buffer buf_n3249( .i (n3248), .o (n3249) );
  assign n3703 = ~n912 & n2916 ;
  assign n3704 = ( n2917 & n3249 ) | ( n2917 & n3703 ) | ( n3249 & n3703 ) ;
  assign n3705 = n3702 | n3704 ;
  assign n3706 = n3698 | n3705 ;
  assign n3707 = n933 & n1057 ;
  assign n3708 = n9 | n3707 ;
  assign n3709 = n2572 | n3708 ;
  assign n3710 = n779 & n3479 ;
  assign n3711 = n3709 & n3710 ;
  buffer buf_n3712( .i (n619), .o (n3712) );
  assign n3713 = ~n3034 & n3712 ;
  assign n3714 = ~n675 & n3713 ;
  assign n3715 = ~n2647 & n3714 ;
  buffer buf_n3716( .i (n911), .o (n3716) );
  assign n3717 = n1899 & ~n3716 ;
  assign n3718 = n1652 | n3717 ;
  assign n3719 = n3715 | n3718 ;
  assign n3720 = n3711 | n3719 ;
  assign n3721 = n3706 | n3720 ;
  assign n3722 = n3694 | n3721 ;
  assign n3723 = n3684 | n3722 ;
  assign n3724 = ~n194 & n3723 ;
  assign y0 = n196 ;
  assign y1 = n465 ;
  assign y2 = n643 ;
  assign y3 = n844 ;
  assign y4 = n1171 ;
  assign y5 = n1485 ;
  assign y6 = n1711 ;
  assign y7 = n1912 ;
  assign y8 = n2133 ;
  assign y9 = n2320 ;
  assign y10 = n2509 ;
  assign y11 = n2635 ;
  assign y12 = n2792 ;
  assign y13 = n2926 ;
  assign y14 = n3072 ;
  assign y15 = n3188 ;
  assign y16 = n3319 ;
  assign y17 = n3422 ;
  assign y18 = n3536 ;
  assign y19 = n3646 ;
  assign y20 = n3724 ;
endmodule
