module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 );
  input G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 ;
  output G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 ;
  wire n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 ;
  buffer buf_n172( .i (G115), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n225( .i (G124), .o (n225) );
  buffer buf_n287( .i (G137), .o (n287) );
  buffer buf_n332( .i (G32), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n162( .i (G106), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n362( .i (G64), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (G76), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n352( .i (G53), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n397( .i (G96), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n342( .i (G43), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n387( .i (G86), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n312( .i (G141), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n317( .i (G142), .o (n317) );
  assign n407 = n313 | n317 ;
  buffer buf_n298( .i (G139), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n306( .i (G140), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  assign n408 = n302 | n307 ;
  assign n409 = n407 | n408 ;
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n218( .i (G121), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  assign n420 = G2 | n220 ;
  assign n421 = G11 | n420 ;
  assign n422 = ~G74 & n172 ;
  assign n423 = G7 | n219 ;
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n192( .i (G119), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  assign n426 = n197 | n424 ;
  buffer buf_n322( .i (G147), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  assign n427 = n327 | n424 ;
  assign n428 = n352 & ~n397 ;
  assign n429 = n342 | n387 ;
  assign n430 = n428 & ~n429 ;
  buffer buf_n431( .i (n430), .o (n431) );
  assign n432 = ~n162 & n332 ;
  assign n433 = n362 | n372 ;
  assign n434 = n432 & ~n433 ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n436 = n431 | n435 ;
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  assign n442 = n322 & ~n435 ;
  assign n443 = n192 & ~n431 ;
  assign n444 = n442 | n443 ;
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = G145 | G146 ;
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  assign n465 = G109 & ~n453 ;
  assign n466 = G79 & ~n453 ;
  assign n467 = n465 | n466 ;
  assign n468 = G89 & ~n453 ;
  buffer buf_n469( .i (n452), .o (n469) );
  assign n470 = G99 & ~n469 ;
  assign n471 = n468 | n470 ;
  assign n472 = n467 | n471 ;
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  assign n495 = G108 | n463 ;
  assign n496 = G98 & ~n463 ;
  assign n497 = n495 & ~n496 ;
  assign n498 = G88 & ~n463 ;
  buffer buf_n499( .i (n462), .o (n499) );
  assign n500 = G78 & ~n499 ;
  assign n501 = n498 | n500 ;
  assign n502 = n497 & ~n501 ;
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  assign n515 = G80 | n469 ;
  assign n516 = G90 & ~n469 ;
  assign n517 = n515 & ~n516 ;
  assign n518 = G100 & ~n469 ;
  buffer buf_n519( .i (n452), .o (n519) );
  assign n520 = G110 & ~n519 ;
  assign n521 = n518 | n520 ;
  assign n522 = n517 & ~n521 ;
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n174( .i (G117), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  assign n545 = ~G36 & n181 ;
  buffer buf_n203( .i (G120), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  assign n546 = ~G68 & n180 ;
  assign n547 = n210 | n546 ;
  assign n548 = n545 & ~n547 ;
  assign n549 = n174 | n203 ;
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  assign n563 = G46 & ~n555 ;
  assign n564 = G57 & ~n555 ;
  assign n565 = n563 | n564 ;
  assign n566 = n548 & ~n565 ;
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  assign n579 = ~G37 & n180 ;
  assign n580 = ~G69 & n179 ;
  assign n581 = n209 | n580 ;
  assign n582 = n579 & ~n581 ;
  assign n583 = G47 & ~n554 ;
  assign n584 = G58 & ~n554 ;
  assign n585 = n583 | n584 ;
  assign n586 = n582 & ~n585 ;
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  assign n600 = ~G38 & n180 ;
  assign n601 = ~G70 & n179 ;
  assign n602 = n209 | n601 ;
  assign n603 = n600 & ~n602 ;
  assign n604 = G48 & ~n554 ;
  buffer buf_n605( .i (n553), .o (n605) );
  assign n606 = G59 & ~n605 ;
  assign n607 = n604 | n606 ;
  assign n608 = n603 & ~n607 ;
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n221( .i (G122), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  assign n622 = ~G31 & n179 ;
  assign n623 = ~G63 & n178 ;
  assign n624 = n208 | n623 ;
  assign n625 = n622 & ~n624 ;
  assign n626 = G42 & ~n553 ;
  assign n627 = G52 & ~n553 ;
  assign n628 = n626 | n627 ;
  assign n629 = n625 & ~n628 ;
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  assign n643 = n222 | n642 ;
  assign n644 = G116 | n218 ;
  assign n645 = n445 | n644 ;
  buffer buf_n646( .i (n645), .o (n646) );
  assign n647 = G28 | n646 ;
  assign n648 = G1 & ~G3 ;
  assign n649 = n646 | n648 ;
  buffer buf_n650( .i (n178), .o (n650) );
  assign n651 = G39 | n650 ;
  assign n652 = ~G71 & n178 ;
  assign n653 = n208 | n652 ;
  assign n654 = n651 & ~n653 ;
  buffer buf_n655( .i (n552), .o (n655) );
  assign n656 = G49 & ~n655 ;
  assign n657 = G60 & ~n655 ;
  assign n658 = n656 | n657 ;
  assign n659 = n654 | n658 ;
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  assign n674 = G56 & ~n558 ;
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  assign n675 = G35 | n183 ;
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  assign n676 = ~G67 & n182 ;
  assign n677 = n212 | n676 ;
  assign n678 = n675 & ~n677 ;
  assign n679 = n674 & ~n678 ;
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  assign n690 = ~G34 & n181 ;
  buffer buf_n691( .i (n650), .o (n691) );
  assign n692 = ~G66 & n691 ;
  assign n693 = n210 | n692 ;
  assign n694 = n690 & ~n693 ;
  assign n695 = G45 & ~n555 ;
  buffer buf_n696( .i (n605), .o (n696) );
  assign n697 = G55 & ~n696 ;
  assign n698 = n695 | n697 ;
  assign n699 = n694 & ~n698 ;
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  assign n712 = ~G33 & n181 ;
  assign n713 = ~G65 & n691 ;
  assign n714 = n210 | n713 ;
  assign n715 = n712 & ~n714 ;
  assign n716 = G44 & ~n696 ;
  assign n717 = G54 & ~n696 ;
  assign n718 = n716 | n717 ;
  assign n719 = n715 & ~n718 ;
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n223( .i (G123), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  assign n732 = ~G40 & n650 ;
  buffer buf_n733( .i (n177), .o (n733) );
  assign n734 = ~G72 & n733 ;
  assign n735 = n208 | n734 ;
  assign n736 = n732 & ~n735 ;
  assign n737 = G50 & ~n655 ;
  assign n738 = G61 & ~n655 ;
  assign n739 = n737 | n738 ;
  assign n740 = n736 & ~n739 ;
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  assign n754 = n224 | n751 ;
  assign n755 = n224 & ~n618 ;
  assign n756 = n754 & ~n755 ;
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = n224 | n670 ;
  assign n759 = ~n224 & n596 ;
  assign n760 = n758 & ~n759 ;
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n189( .i (G118), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  assign n762 = n191 & ~n221 ;
  assign n763 = n753 | n762 ;
  buffer buf_n764( .i (n223), .o (n764) );
  assign n765 = ~n640 & n764 ;
  assign n766 = n189 | n223 ;
  assign n767 = n751 & ~n766 ;
  assign n768 = n765 | n767 ;
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n321( .i (G143), .o (n321) );
  buffer buf_n464( .i (n463), .o (n464) );
  assign n770 = G77 & ~n464 ;
  assign n771 = G97 & ~n464 ;
  assign n772 = n770 & ~n771 ;
  assign n773 = G107 & ~n464 ;
  assign n774 = G87 & ~n464 ;
  assign n775 = n773 | n774 ;
  assign n776 = n772 & ~n775 ;
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  assign n785 = n321 | n784 ;
  assign n786 = n321 & ~n784 ;
  assign n787 = n785 & ~n786 ;
  assign n788 = G144 | n787 ;
  buffer buf_n158( .i (G10), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  inverter inv_n161( .i (n160), .o (n161) );
  buffer buf_n275( .i (G135), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n328( .i (G23), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  assign n789 = ~G19 & n330 ;
  buffer buf_n790( .i (n499), .o (n790) );
  assign n791 = G75 & ~n790 ;
  assign n792 = G85 & ~n790 ;
  assign n793 = n791 & ~n792 ;
  assign n794 = G95 & ~n790 ;
  assign n795 = G105 & ~n790 ;
  assign n796 = n794 | n795 ;
  assign n797 = n793 & ~n796 ;
  buffer buf_n798( .i (n797), .o (n798) );
  assign n800 = n330 & ~n798 ;
  assign n801 = n789 & ~n800 ;
  assign n802 = n276 & ~n801 ;
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n226( .i (G125), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n198( .i (G12), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  assign n806 = ~G13 & n200 ;
  assign n807 = n200 & ~n632 ;
  assign n808 = n806 & ~n807 ;
  assign n809 = n232 & ~n808 ;
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n254( .i (G130), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  assign n813 = ~G15 & n200 ;
  buffer buf_n814( .i (n199), .o (n814) );
  assign n815 = n588 & ~n814 ;
  assign n816 = n813 & ~n815 ;
  assign n817 = n258 & ~n816 ;
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  assign n821 = n812 | n820 ;
  assign n822 = n805 | n821 ;
  buffer buf_n249( .i (G129), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  assign n823 = ~G5 & n814 ;
  assign n824 = ~n610 & n814 ;
  assign n825 = n823 & ~n824 ;
  assign n826 = n253 & ~n825 ;
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  assign n829 = ~G21 & n330 ;
  buffer buf_n830( .i (n329), .o (n830) );
  assign n831 = ~n534 & n830 ;
  assign n832 = n829 & ~n831 ;
  assign n833 = n311 & ~n832 ;
  buffer buf_n834( .i (n833), .o (n834) );
  assign n835 = n828 | n834 ;
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  assign n836 = ~G27 & n329 ;
  assign n837 = n329 & ~n503 ;
  assign n838 = n836 & ~n837 ;
  assign n839 = n320 & ~n838 ;
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  assign n842 = n803 | n841 ;
  assign n843 = n835 | n842 ;
  buffer buf_n241( .i (G128), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  assign n844 = ~G14 & n814 ;
  buffer buf_n845( .i (n199), .o (n845) );
  assign n846 = n662 & ~n845 ;
  assign n847 = n844 & ~n846 ;
  assign n848 = n248 & ~n847 ;
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n233( .i (G126), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  assign n851 = ~G4 & n845 ;
  assign n852 = ~n743 & n845 ;
  assign n853 = n851 & ~n852 ;
  assign n854 = n240 & ~n853 ;
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  assign n857 = n850 | n856 ;
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n858( .i (n328), .o (n858) );
  assign n859 = ~G26 & n858 ;
  assign n860 = ~n483 & n858 ;
  assign n861 = n859 & ~n860 ;
  assign n862 = n316 & ~n861 ;
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  assign n865 = n834 | n864 ;
  assign n866 = n857 | n865 ;
  assign n867 = n843 | n866 ;
  assign n868 = n822 | n867 ;
  buffer buf_n277( .i (G136), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n331( .i (n330), .o (n331) );
  assign n869 = ~G24 & n331 ;
  buffer buf_n870( .i (n499), .o (n870) );
  assign n871 = G93 & ~n870 ;
  assign n872 = G103 & ~n870 ;
  assign n873 = n871 & ~n872 ;
  assign n874 = G113 & ~n870 ;
  assign n875 = G83 & ~n870 ;
  assign n876 = n874 | n875 ;
  assign n877 = n873 & ~n876 ;
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  assign n880 = n331 & ~n879 ;
  assign n881 = n869 & ~n880 ;
  buffer buf_n882( .i (n881), .o (n882) );
  assign n883 = n286 | n882 ;
  assign n884 = n286 & ~n882 ;
  assign n885 = n883 & ~n884 ;
  buffer buf_n259( .i (G131), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n201( .i (n200), .o (n201) );
  assign n886 = ~G16 & n201 ;
  assign n887 = n201 & ~n568 ;
  assign n888 = n886 & ~n887 ;
  buffer buf_n889( .i (n888), .o (n889) );
  assign n890 = n264 | n889 ;
  assign n891 = n264 & ~n889 ;
  assign n892 = n890 & ~n891 ;
  buffer buf_n288( .i (G138), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  assign n893 = ~G20 & n830 ;
  buffer buf_n894( .i (n499), .o (n894) );
  assign n895 = G82 & ~n894 ;
  assign n896 = G102 & ~n894 ;
  assign n897 = n895 & ~n896 ;
  assign n898 = G112 & ~n894 ;
  assign n899 = G92 & ~n894 ;
  assign n900 = n898 | n899 ;
  assign n901 = n897 & ~n900 ;
  buffer buf_n902( .i (n901), .o (n902) );
  assign n905 = n830 & ~n902 ;
  assign n906 = n893 & ~n905 ;
  buffer buf_n907( .i (n906), .o (n907) );
  assign n908 = n297 | n907 ;
  assign n909 = n297 & ~n907 ;
  assign n910 = n908 & ~n909 ;
  assign n911 = n892 | n910 ;
  assign n912 = n885 | n911 ;
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  assign n913 = ~G25 & n858 ;
  buffer buf_n914( .i (n462), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  assign n916 = G81 & ~n915 ;
  assign n917 = G101 & ~n915 ;
  assign n918 = n916 & ~n917 ;
  assign n919 = G111 & ~n915 ;
  assign n920 = G91 & ~n915 ;
  assign n921 = n919 | n920 ;
  assign n922 = n918 & ~n921 ;
  assign n923 = n858 & ~n922 ;
  assign n924 = n913 & ~n923 ;
  assign n925 = n305 & ~n924 ;
  buffer buf_n926( .i (n925), .o (n926) );
  assign n927 = n818 | n926 ;
  buffer buf_n273( .i (G134), .o (n273) );
  assign n928 = ~G18 & n845 ;
  buffer buf_n929( .i (n199), .o (n929) );
  assign n930 = ~n720 & n929 ;
  assign n931 = n928 & ~n930 ;
  assign n932 = n273 & ~n931 ;
  buffer buf_n933( .i (n932), .o (n933) );
  assign n934 = n855 | n933 ;
  assign n935 = n927 | n934 ;
  buffer buf_n267( .i (G133), .o (n267) );
  assign n936 = ~G6 & n929 ;
  assign n937 = ~n700 & n929 ;
  assign n938 = n936 & ~n937 ;
  assign n939 = n267 & ~n938 ;
  buffer buf_n940( .i (n939), .o (n940) );
  assign n941 = n331 & ~n778 ;
  assign n942 = ~G22 & n830 ;
  assign n943 = G9 | n942 ;
  assign n944 = n941 | n943 ;
  assign n945 = n940 | n944 ;
  assign n946 = n840 | n940 ;
  assign n947 = n945 | n946 ;
  assign n948 = n935 | n947 ;
  assign n949 = n827 | n863 ;
  assign n950 = n810 | n849 ;
  assign n951 = n949 | n950 ;
  assign n952 = n926 | n933 ;
  buffer buf_n265( .i (G132), .o (n265) );
  buffer buf_n202( .i (n201), .o (n202) );
  assign n953 = ~G17 & n202 ;
  assign n954 = n202 & ~n680 ;
  assign n955 = n953 & ~n954 ;
  assign n956 = n265 & ~n955 ;
  assign n957 = n952 | n956 ;
  assign n958 = n951 | n957 ;
  assign n959 = n948 | n958 ;
  assign n960 = n912 | n959 ;
  assign n961 = n868 | n960 ;
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  assign n963 = ~G41 & n188 ;
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  assign n964 = ~G73 & n187 ;
  assign n965 = n217 | n964 ;
  assign n966 = n963 & ~n965 ;
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  assign n967 = G51 & ~n562 ;
  assign n968 = G62 & ~n562 ;
  assign n969 = n967 | n968 ;
  assign n970 = n966 & ~n969 ;
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  assign n974 = n221 & ~n973 ;
  assign n975 = n222 | n974 ;
  assign n976 = n505 | n778 ;
  assign n977 = n505 & ~n778 ;
  assign n978 = n976 & ~n977 ;
  buffer buf_n979( .i (n978), .o (n979) );
  assign n980 = n488 | n979 ;
  assign n981 = ~n488 & n979 ;
  assign n982 = n980 & ~n981 ;
  assign n983 = G29 | n982 ;
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  inverter inv_n986( .i (n985), .o (n986) );
  assign n987 = n223 & ~n971 ;
  assign n988 = n764 | n987 ;
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n382( .i (G8), .o (n382) );
  assign n991 = G127 | n523 ;
  buffer buf_n992( .i (n991), .o (n992) );
  assign n993 = G30 | n473 ;
  buffer buf_n994( .i (n993), .o (n994) );
  assign n995 = n992 | n994 ;
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  assign n1001 = ~n382 & n998 ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  assign n1012 = ~n272 & n1011 ;
  assign n1013 = n382 | n998 ;
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  assign n1023 = n706 | n1022 ;
  buffer buf_n266( .i (n265), .o (n266) );
  assign n1024 = ~n266 & n1009 ;
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  assign n1025 = n249 & n1000 ;
  assign n1026 = n306 & ~n1000 ;
  assign n1027 = n1025 & ~n1026 ;
  assign n1028 = n610 & ~n1027 ;
  buffer buf_n1029( .i (n1028), .o (n1029) );
  assign n1030 = ~n241 & n997 ;
  assign n1031 = n298 & ~n997 ;
  assign n1032 = n1030 | n1031 ;
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  assign n1036 = ~n662 & n1035 ;
  assign n1037 = ~n233 & n997 ;
  buffer buf_n1038( .i (n996), .o (n1038) );
  assign n1039 = n288 & ~n1038 ;
  assign n1040 = n1037 | n1039 ;
  buffer buf_n1041( .i (n1040), .o (n1041) );
  assign n1042 = n741 | n1041 ;
  assign n1043 = ~n226 & n998 ;
  buffer buf_n1044( .i (n1038), .o (n1044) );
  assign n1045 = n277 & ~n1044 ;
  assign n1046 = n1043 | n1045 ;
  assign n1047 = ~n630 & n1046 ;
  assign n1048 = n1042 & n1047 ;
  assign n1049 = n741 & n1041 ;
  assign n1050 = n660 & n1033 ;
  assign n1051 = n1049 | n1050 ;
  assign n1052 = n1048 | n1051 ;
  assign n1053 = ~n1036 & n1052 ;
  assign n1054 = n1029 | n1053 ;
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  assign n1055 = n385 & ~n587 ;
  assign n1056 = n254 & n1002 ;
  assign n1057 = n312 & ~n1014 ;
  assign n1058 = n1056 & ~n1057 ;
  assign n1059 = n1055 & ~n1058 ;
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1062 = n1029 | n1060 ;
  assign n1063 = n1054 & ~n1062 ;
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n386( .i (n385), .o (n386) );
  assign n1064 = n386 & ~n567 ;
  assign n1065 = n259 & n1003 ;
  assign n1066 = n317 & ~n1015 ;
  assign n1067 = n1065 & ~n1066 ;
  assign n1068 = n1064 & ~n1067 ;
  buffer buf_n1069( .i (n1068), .o (n1069) );
  assign n1071 = n1061 | n1069 ;
  assign n1072 = n1063 | n1071 ;
  buffer buf_n1070( .i (n1069), .o (n1070) );
  assign n1073 = n681 & ~n1019 ;
  assign n1074 = n1070 | n1073 ;
  assign n1075 = n1072 & ~n1074 ;
  assign n1076 = n1024 | n1075 ;
  assign n1077 = n1023 & n1076 ;
  assign n1078 = n1012 | n1077 ;
  assign n1079 = n992 & ~n994 ;
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  assign n1092 = n282 | n878 ;
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  assign n1096 = n1091 & ~n1095 ;
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  assign n1097 = n296 | n904 ;
  assign n1098 = n1090 & ~n1097 ;
  buffer buf_n1099( .i (n1098), .o (n1099) );
  assign n1103 = n1096 & ~n1099 ;
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n799( .i (n798), .o (n799) );
  assign n1105 = n275 | n799 ;
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n274( .i (n273), .o (n274) );
  assign n1109 = n274 & ~n723 ;
  assign n1110 = n1106 & ~n1109 ;
  assign n1111 = n1091 & ~n1110 ;
  assign n1112 = n1099 | n1111 ;
  assign n1113 = n275 & ~n799 ;
  assign n1114 = n1093 & ~n1113 ;
  assign n1115 = n1090 & ~n1114 ;
  buffer buf_n1116( .i (n1115), .o (n1116) );
  assign n1118 = n274 | n723 ;
  assign n1119 = n1090 & ~n1118 ;
  buffer buf_n1120( .i (n1119), .o (n1120) );
  assign n1121 = n1116 | n1120 ;
  assign n1122 = n1112 | n1121 ;
  assign n1123 = n1104 & ~n1122 ;
  assign n1124 = n1078 & n1123 ;
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  assign n1125 = n1108 & ~n1120 ;
  assign n1126 = n1117 & ~n1125 ;
  assign n1127 = n1104 & ~n1126 ;
  assign n1128 = n1102 | n1127 ;
  assign n1129 = ~n1124 & ~n1128 ;
  assign n1130 = n158 & ~n445 ;
  assign n1131 = n984 & n1130 ;
  inverter inv_n1132( .i (n1131), .o (n1132) );
  assign G2531 = n173 ;
  assign G2532 = n173 ;
  assign G2533 = n173 ;
  assign G2534 = n225 ;
  assign G2535 = n225 ;
  assign G2536 = n287 ;
  assign G2537 = n287 ;
  assign G2538 = n287 ;
  assign G2539 = n341 ;
  assign G2540 = n171 ;
  assign G2541 = n371 ;
  assign G2542 = n381 ;
  assign G2543 = n361 ;
  assign G2544 = n406 ;
  assign G2545 = n351 ;
  assign G2546 = n396 ;
  assign G2547 = n419 ;
  assign G2548 = n421 ;
  assign G2549 = n173 ;
  assign G2550 = n422 ;
  assign G2551 = n425 ;
  assign G2552 = n426 ;
  assign G2553 = n427 ;
  assign G2554 = n441 ;
  assign G2555 = n441 ;
  assign G2556 = n448 ;
  assign G2557 = n494 ;
  assign G2558 = n514 ;
  assign G2559 = n544 ;
  assign G2560 = n578 ;
  assign G2561 = n599 ;
  assign G2562 = n621 ;
  assign G2563 = n643 ;
  assign G2564 = n647 ;
  assign G2565 = n649 ;
  assign G2566 = n673 ;
  assign G2567 = n621 ;
  assign G2568 = n599 ;
  assign G2569 = n578 ;
  assign G2570 = n689 ;
  assign G2571 = n711 ;
  assign G2572 = n731 ;
  assign G2573 = n757 ;
  assign G2574 = n757 ;
  assign G2575 = n761 ;
  assign G2576 = n761 ;
  assign G2577 = n763 ;
  assign G2578 = n769 ;
  assign G2579 = n769 ;
  assign G2580 = n788 ;
  assign G2581 = n161 ;
  assign G2582 = 1'b0 ;
  assign G2583 = 1'b0 ;
  assign G2584 = n962 ;
  assign G2585 = n962 ;
  assign G2586 = n975 ;
  assign G2587 = n986 ;
  assign G2588 = n990 ;
  assign G2589 = n990 ;
  assign G2590 = 1'b0 ;
  assign G2591 = n1129 ;
  assign G2592 = 1'b0 ;
  assign G2593 = n1132 ;
  assign G2594 = n1132 ;
endmodule
