module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( N1 , N101 , N105 , N109 , N113 , N117 , N121 , N125 , N129 , N13 , N130 , N131 , N132 , N133 , N134 , N135 , N136 , N137 , N17 , N21 , N25 , N29 , N33 , N37 , N41 , N45 , N49 , N5 , N53 , N57 , N61 , N65 , N69 , N73 , N77 , N81 , N85 , N89 , N9 , N93 , N97 , N724 , N725 , N726 , N727 , N728 , N729 , N730 , N731 , N732 , N733 , N734 , N735 , N736 , N737 , N738 , N739 , N740 , N741 , N742 , N743 , N744 , N745 , N746 , N747 , N748 , N749 , N750 , N751 , N752 , N753 , N754 , N755 );
  input N1 , N101 , N105 , N109 , N113 , N117 , N121 , N125 , N129 , N13 , N130 , N131 , N132 , N133 , N134 , N135 , N136 , N137 , N17 , N21 , N25 , N29 , N33 , N37 , N41 , N45 , N49 , N5 , N53 , N57 , N61 , N65 , N69 , N73 , N77 , N81 , N85 , N89 , N9 , N93 , N97 ;
  output N724 , N725 , N726 , N727 , N728 , N729 , N730 , N731 , N732 , N733 , N734 , N735 , N736 , N737 , N738 , N739 , N740 , N741 , N742 , N743 , N744 , N745 , N746 , N747 , N748 , N749 , N750 , N751 , N752 , N753 , N754 , N755 ;
  wire n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 ;
  assign n42 = N33 & ~N49 ;
  assign n43 = ~N33 & N49 ;
  assign n44 = n42 | n43 ;
  buffer buf_n45( .i (n44), .o (n45) );
  assign n46 = N129 & N137 ;
  buffer buf_n47( .i (n46), .o (n47) );
  assign n48 = N1 & ~N17 ;
  assign n49 = ~N1 & N17 ;
  assign n50 = n48 | n49 ;
  buffer buf_n51( .i (n50), .o (n51) );
  assign n52 = n47 & ~n51 ;
  assign n53 = ~n47 & n51 ;
  assign n54 = n52 | n53 ;
  buffer buf_n55( .i (n54), .o (n55) );
  assign n56 = n45 | n55 ;
  assign n57 = n45 & n55 ;
  assign n58 = n56 & ~n57 ;
  buffer buf_n59( .i (n58), .o (n59) );
  assign n60 = N73 | N77 ;
  assign n61 = N73 & N77 ;
  assign n62 = n60 & ~n61 ;
  buffer buf_n63( .i (n62), .o (n63) );
  assign n64 = N65 & ~N69 ;
  assign n65 = ~N65 & N69 ;
  assign n66 = n64 | n65 ;
  buffer buf_n67( .i (n66), .o (n67) );
  assign n68 = ~n63 & n67 ;
  assign n69 = n63 & ~n67 ;
  assign n70 = n68 | n69 ;
  buffer buf_n71( .i (n70), .o (n71) );
  assign n73 = N89 | N93 ;
  assign n74 = N89 & N93 ;
  assign n75 = n73 & ~n74 ;
  buffer buf_n76( .i (n75), .o (n76) );
  assign n77 = N81 & ~N85 ;
  assign n78 = ~N81 & N85 ;
  assign n79 = n77 | n78 ;
  buffer buf_n80( .i (n79), .o (n80) );
  assign n81 = ~n76 & n80 ;
  assign n82 = n76 & ~n80 ;
  assign n83 = n81 | n82 ;
  buffer buf_n84( .i (n83), .o (n84) );
  assign n86 = n71 & n84 ;
  assign n87 = n71 | n84 ;
  assign n88 = ~n86 & n87 ;
  buffer buf_n89( .i (n88), .o (n89) );
  assign n90 = ~n59 & n89 ;
  assign n91 = n59 & ~n89 ;
  assign n92 = n90 | n91 ;
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  assign n106 = N135 & N137 ;
  buffer buf_n107( .i (n106), .o (n107) );
  assign n108 = N105 & ~N121 ;
  assign n109 = ~N105 & N121 ;
  assign n110 = n108 | n109 ;
  buffer buf_n111( .i (n110), .o (n111) );
  assign n112 = N73 & ~N89 ;
  assign n113 = ~N73 & N89 ;
  assign n114 = n112 | n113 ;
  buffer buf_n115( .i (n114), .o (n115) );
  assign n116 = ~n111 & n115 ;
  assign n117 = n111 & ~n115 ;
  assign n118 = n116 | n117 ;
  buffer buf_n119( .i (n118), .o (n119) );
  assign n120 = n107 & n119 ;
  assign n121 = n107 | n119 ;
  assign n122 = ~n120 & n121 ;
  buffer buf_n123( .i (n122), .o (n123) );
  assign n124 = N13 | N9 ;
  assign n125 = N13 & N9 ;
  assign n126 = n124 & ~n125 ;
  buffer buf_n127( .i (n126), .o (n127) );
  assign n128 = N1 & ~N5 ;
  assign n129 = ~N1 & N5 ;
  assign n130 = n128 | n129 ;
  buffer buf_n131( .i (n130), .o (n131) );
  assign n132 = ~n127 & n131 ;
  assign n133 = n127 & ~n131 ;
  assign n134 = n132 | n133 ;
  buffer buf_n135( .i (n134), .o (n135) );
  assign n136 = N41 | N45 ;
  assign n137 = N41 & N45 ;
  assign n138 = n136 & ~n137 ;
  buffer buf_n139( .i (n138), .o (n139) );
  assign n140 = N33 & ~N37 ;
  assign n141 = ~N33 & N37 ;
  assign n142 = n140 | n141 ;
  buffer buf_n143( .i (n142), .o (n143) );
  assign n144 = ~n139 & n143 ;
  assign n145 = n139 & ~n143 ;
  assign n146 = n144 | n145 ;
  buffer buf_n147( .i (n146), .o (n147) );
  assign n148 = n135 & n147 ;
  assign n149 = n135 | n147 ;
  assign n150 = ~n148 & n149 ;
  buffer buf_n151( .i (n150), .o (n151) );
  assign n152 = ~n123 & n151 ;
  assign n153 = n123 & ~n151 ;
  assign n154 = n152 | n153 ;
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  assign n167 = N136 & N137 ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = N109 & ~N125 ;
  assign n170 = ~N109 & N125 ;
  assign n171 = n169 | n170 ;
  buffer buf_n172( .i (n171), .o (n172) );
  assign n173 = N77 & ~N93 ;
  assign n174 = ~N77 & N93 ;
  assign n175 = n173 | n174 ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n177 = ~n172 & n176 ;
  assign n178 = n172 & ~n176 ;
  assign n179 = n177 | n178 ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = n168 & n180 ;
  assign n182 = n168 | n180 ;
  assign n183 = ~n181 & n182 ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n185 = N25 | N29 ;
  assign n186 = N25 & N29 ;
  assign n187 = n185 & ~n186 ;
  buffer buf_n188( .i (n187), .o (n188) );
  assign n189 = N17 & ~N21 ;
  assign n190 = ~N17 & N21 ;
  assign n191 = n189 | n190 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = ~n188 & n192 ;
  assign n194 = n188 & ~n192 ;
  assign n195 = n193 | n194 ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n197 = N57 | N61 ;
  assign n198 = N57 & N61 ;
  assign n199 = n197 & ~n198 ;
  buffer buf_n200( .i (n199), .o (n200) );
  assign n201 = N49 & ~N53 ;
  assign n202 = ~N49 & N53 ;
  assign n203 = n201 | n202 ;
  buffer buf_n204( .i (n203), .o (n204) );
  assign n205 = ~n200 & n204 ;
  assign n206 = n200 & ~n204 ;
  assign n207 = n205 | n206 ;
  buffer buf_n208( .i (n207), .o (n208) );
  assign n209 = n196 & n208 ;
  assign n210 = n196 | n208 ;
  assign n211 = ~n209 & n210 ;
  buffer buf_n212( .i (n211), .o (n212) );
  assign n213 = ~n184 & n212 ;
  assign n214 = n184 & ~n212 ;
  assign n215 = n213 | n214 ;
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  assign n228 = n156 & ~n217 ;
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  assign n236 = N131 & N137 ;
  buffer buf_n237( .i (n236), .o (n237) );
  assign n238 = N41 & ~N57 ;
  assign n239 = ~N41 & N57 ;
  assign n240 = n238 | n239 ;
  buffer buf_n241( .i (n240), .o (n241) );
  assign n242 = ~N25 & N9 ;
  assign n243 = N25 & ~N9 ;
  assign n244 = n242 | n243 ;
  buffer buf_n245( .i (n244), .o (n245) );
  assign n246 = ~n241 & n245 ;
  assign n247 = n241 & ~n245 ;
  assign n248 = n246 | n247 ;
  buffer buf_n249( .i (n248), .o (n249) );
  assign n250 = n237 & n249 ;
  assign n251 = n237 | n249 ;
  assign n252 = ~n250 & n251 ;
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n72( .i (n71), .o (n72) );
  assign n254 = N105 | N109 ;
  assign n255 = N105 & N109 ;
  assign n256 = n254 & ~n255 ;
  buffer buf_n257( .i (n256), .o (n257) );
  assign n258 = ~N101 & N97 ;
  assign n259 = N101 & ~N97 ;
  assign n260 = n258 | n259 ;
  buffer buf_n261( .i (n260), .o (n261) );
  assign n262 = ~n257 & n261 ;
  assign n263 = n257 & ~n261 ;
  assign n264 = n262 | n263 ;
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  assign n267 = n72 & n266 ;
  assign n268 = n72 | n266 ;
  assign n269 = ~n267 & n268 ;
  buffer buf_n270( .i (n269), .o (n270) );
  assign n271 = ~n253 & n270 ;
  assign n272 = n253 & ~n270 ;
  assign n273 = n271 | n272 ;
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  assign n286 = N37 & ~N53 ;
  assign n287 = ~N37 & N53 ;
  assign n288 = n286 | n287 ;
  buffer buf_n289( .i (n288), .o (n289) );
  assign n290 = N130 & N137 ;
  buffer buf_n291( .i (n290), .o (n291) );
  assign n292 = ~N21 & N5 ;
  assign n293 = N21 & ~N5 ;
  assign n294 = n292 | n293 ;
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = n291 & ~n295 ;
  assign n297 = ~n291 & n295 ;
  assign n298 = n296 | n297 ;
  buffer buf_n299( .i (n298), .o (n299) );
  assign n300 = n289 | n299 ;
  assign n301 = n289 & n299 ;
  assign n302 = n300 & ~n301 ;
  buffer buf_n303( .i (n302), .o (n303) );
  assign n304 = N121 | N125 ;
  assign n305 = N121 & N125 ;
  assign n306 = n304 & ~n305 ;
  buffer buf_n307( .i (n306), .o (n307) );
  assign n308 = N113 & ~N117 ;
  assign n309 = ~N113 & N117 ;
  assign n310 = n308 | n309 ;
  buffer buf_n311( .i (n310), .o (n311) );
  assign n312 = ~n307 & n311 ;
  assign n313 = n307 & ~n311 ;
  assign n314 = n312 | n313 ;
  buffer buf_n315( .i (n314), .o (n315) );
  assign n317 = n265 & n315 ;
  assign n318 = n265 | n315 ;
  assign n319 = ~n317 & n318 ;
  buffer buf_n320( .i (n319), .o (n320) );
  assign n321 = ~n303 & n320 ;
  assign n322 = n303 & ~n320 ;
  assign n323 = n321 | n322 ;
  buffer buf_n324( .i (n323), .o (n324) );
  assign n337 = ~n93 & n324 ;
  buffer buf_n338( .i (n337), .o (n338) );
  assign n347 = ~n275 & n338 ;
  buffer buf_n348( .i (n347), .o (n348) );
  assign n355 = n93 & ~n324 ;
  buffer buf_n356( .i (n355), .o (n356) );
  assign n365 = ~n275 & n356 ;
  buffer buf_n366( .i (n365), .o (n366) );
  assign n373 = n348 | n366 ;
  assign n374 = N132 & N137 ;
  buffer buf_n375( .i (n374), .o (n375) );
  assign n376 = N45 & ~N61 ;
  assign n377 = ~N45 & N61 ;
  assign n378 = n376 | n377 ;
  buffer buf_n379( .i (n378), .o (n379) );
  assign n380 = N13 & ~N29 ;
  assign n381 = ~N13 & N29 ;
  assign n382 = n380 | n381 ;
  buffer buf_n383( .i (n382), .o (n383) );
  assign n384 = ~n379 & n383 ;
  assign n385 = n379 & ~n383 ;
  assign n386 = n384 | n385 ;
  buffer buf_n387( .i (n386), .o (n387) );
  assign n388 = n375 & n387 ;
  assign n389 = n375 | n387 ;
  assign n390 = ~n388 & n389 ;
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n316( .i (n315), .o (n316) );
  assign n392 = n85 & n316 ;
  assign n393 = n85 | n316 ;
  assign n394 = ~n392 & n393 ;
  buffer buf_n395( .i (n394), .o (n395) );
  assign n396 = ~n391 & n395 ;
  assign n397 = n391 & ~n395 ;
  assign n398 = n396 | n397 ;
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  assign n411 = n373 & ~n403 ;
  assign n412 = n275 & ~n400 ;
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n276( .i (n275), .o (n276) );
  assign n418 = ~n276 & n401 ;
  assign n419 = n413 | n418 ;
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  assign n420 = n97 | n328 ;
  assign n421 = n419 & ~n420 ;
  assign n422 = n411 | n421 ;
  buffer buf_n423( .i (n422), .o (n423) );
  assign n424 = ~N113 & N97 ;
  assign n425 = N113 & ~N97 ;
  assign n426 = n424 | n425 ;
  buffer buf_n427( .i (n426), .o (n427) );
  assign n428 = N133 & N137 ;
  buffer buf_n429( .i (n428), .o (n429) );
  assign n430 = N65 & ~N81 ;
  assign n431 = ~N65 & N81 ;
  assign n432 = n430 | n431 ;
  buffer buf_n433( .i (n432), .o (n433) );
  assign n434 = n429 & ~n433 ;
  assign n435 = ~n429 & n433 ;
  assign n436 = n434 | n435 ;
  buffer buf_n437( .i (n436), .o (n437) );
  assign n438 = n427 | n437 ;
  assign n439 = n427 & n437 ;
  assign n440 = n438 & ~n439 ;
  buffer buf_n441( .i (n440), .o (n441) );
  assign n442 = n135 & n196 ;
  assign n443 = n135 | n196 ;
  assign n444 = ~n442 & n443 ;
  buffer buf_n445( .i (n444), .o (n445) );
  assign n446 = ~n441 & n445 ;
  assign n447 = n441 & ~n445 ;
  assign n448 = n446 | n447 ;
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  assign n461 = N101 & ~N117 ;
  assign n462 = ~N101 & N117 ;
  assign n463 = n461 | n462 ;
  buffer buf_n464( .i (n463), .o (n464) );
  assign n465 = N134 & N137 ;
  buffer buf_n466( .i (n465), .o (n466) );
  assign n467 = N69 & ~N85 ;
  assign n468 = ~N69 & N85 ;
  assign n469 = n467 | n468 ;
  buffer buf_n470( .i (n469), .o (n470) );
  assign n471 = n466 & ~n470 ;
  assign n472 = ~n466 & n470 ;
  assign n473 = n471 | n472 ;
  buffer buf_n474( .i (n473), .o (n474) );
  assign n475 = n464 | n474 ;
  assign n476 = n464 & n474 ;
  assign n477 = n475 & ~n476 ;
  buffer buf_n478( .i (n477), .o (n478) );
  assign n479 = n147 & n208 ;
  assign n480 = n147 | n208 ;
  assign n481 = ~n479 & n480 ;
  buffer buf_n482( .i (n481), .o (n482) );
  assign n483 = ~n478 & n482 ;
  assign n484 = n478 & ~n482 ;
  assign n485 = n483 | n484 ;
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  assign n498 = n450 & ~n487 ;
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  assign n504 = n423 & n503 ;
  buffer buf_n505( .i (n504), .o (n505) );
  assign n506 = n235 & n505 ;
  buffer buf_n507( .i (n506), .o (n507) );
  assign n508 = n105 & n507 ;
  buffer buf_n509( .i (n508), .o (n509) );
  assign n510 = N1 | n509 ;
  assign n511 = N1 & n509 ;
  assign n512 = n510 & ~n511 ;
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  assign n513 = n336 & n507 ;
  buffer buf_n514( .i (n513), .o (n514) );
  assign n515 = N5 | n514 ;
  assign n516 = N5 & n514 ;
  assign n517 = n515 & ~n516 ;
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  assign n518 = n285 & n507 ;
  buffer buf_n519( .i (n518), .o (n519) );
  assign n520 = N9 & n519 ;
  assign n521 = N9 | n519 ;
  assign n522 = ~n520 & n521 ;
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  assign n523 = n410 & n507 ;
  buffer buf_n524( .i (n523), .o (n524) );
  assign n525 = ~N13 & n524 ;
  assign n526 = N13 & ~n524 ;
  assign n527 = n525 | n526 ;
  assign n528 = ~n156 & n217 ;
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  assign n536 = n505 & n535 ;
  buffer buf_n537( .i (n536), .o (n537) );
  assign n538 = n105 & n537 ;
  buffer buf_n539( .i (n538), .o (n539) );
  assign n540 = N17 | n539 ;
  assign n541 = N17 & n539 ;
  assign n542 = n540 & ~n541 ;
  assign n543 = n336 & n537 ;
  buffer buf_n544( .i (n543), .o (n544) );
  assign n545 = N21 | n544 ;
  assign n546 = N21 & n544 ;
  assign n547 = n545 & ~n546 ;
  assign n548 = n285 & n537 ;
  buffer buf_n549( .i (n548), .o (n549) );
  assign n550 = N25 & n549 ;
  assign n551 = N25 | n549 ;
  assign n552 = ~n550 & n551 ;
  assign n553 = n410 & n537 ;
  buffer buf_n554( .i (n553), .o (n554) );
  assign n555 = ~N29 & n554 ;
  assign n556 = N29 & ~n554 ;
  assign n557 = n555 | n556 ;
  assign n558 = ~n450 & n487 ;
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  assign n564 = n423 & n563 ;
  buffer buf_n565( .i (n564), .o (n565) );
  assign n566 = n235 & n565 ;
  buffer buf_n567( .i (n566), .o (n567) );
  assign n568 = n105 & n567 ;
  buffer buf_n569( .i (n568), .o (n569) );
  assign n570 = N33 | n569 ;
  assign n571 = N33 & n569 ;
  assign n572 = n570 & ~n571 ;
  assign n573 = n336 & n567 ;
  buffer buf_n574( .i (n573), .o (n574) );
  assign n575 = N37 | n574 ;
  assign n576 = N37 & n574 ;
  assign n577 = n575 & ~n576 ;
  assign n578 = n285 & n567 ;
  buffer buf_n579( .i (n578), .o (n579) );
  assign n580 = N41 & n579 ;
  assign n581 = N41 | n579 ;
  assign n582 = ~n580 & n581 ;
  assign n583 = n410 & n567 ;
  buffer buf_n584( .i (n583), .o (n584) );
  assign n585 = N45 | n584 ;
  assign n586 = N45 & n584 ;
  assign n587 = n585 & ~n586 ;
  assign n588 = n535 & n565 ;
  buffer buf_n589( .i (n588), .o (n589) );
  assign n590 = n105 & n589 ;
  buffer buf_n591( .i (n590), .o (n591) );
  assign n592 = N49 | n591 ;
  assign n593 = N49 & n591 ;
  assign n594 = n592 & ~n593 ;
  assign n595 = n336 & n589 ;
  buffer buf_n596( .i (n595), .o (n596) );
  assign n597 = N53 | n596 ;
  assign n598 = N53 & n596 ;
  assign n599 = n597 & ~n598 ;
  assign n600 = n285 & n589 ;
  buffer buf_n601( .i (n600), .o (n601) );
  assign n602 = N57 & n601 ;
  assign n603 = N57 | n601 ;
  assign n604 = ~n602 & n603 ;
  assign n605 = n410 & n589 ;
  buffer buf_n606( .i (n605), .o (n606) );
  assign n607 = N61 & n606 ;
  assign n608 = N61 | n606 ;
  assign n609 = ~n607 & n608 ;
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  assign n610 = n499 | n559 ;
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  assign n611 = n158 | n219 ;
  assign n612 = n610 & ~n611 ;
  assign n613 = n229 | n529 ;
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  assign n614 = n452 | n489 ;
  assign n615 = n613 & ~n614 ;
  assign n616 = n612 | n615 ;
  buffer buf_n617( .i (n616), .o (n617) );
  assign n618 = n417 & n617 ;
  buffer buf_n619( .i (n618), .o (n619) );
  assign n620 = n364 & n619 ;
  buffer buf_n621( .i (n620), .o (n621) );
  assign n622 = n460 & n621 ;
  buffer buf_n623( .i (n622), .o (n623) );
  assign n624 = N65 | n623 ;
  assign n625 = N65 & n623 ;
  assign n626 = n624 & ~n625 ;
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  assign n627 = n497 & n621 ;
  buffer buf_n628( .i (n627), .o (n628) );
  assign n629 = N69 | n628 ;
  assign n630 = N69 & n628 ;
  assign n631 = n629 & ~n630 ;
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  assign n632 = n166 & n621 ;
  buffer buf_n633( .i (n632), .o (n633) );
  assign n634 = ~N73 & n633 ;
  assign n635 = N73 & ~n633 ;
  assign n636 = n634 | n635 ;
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  assign n637 = n227 & n621 ;
  buffer buf_n638( .i (n637), .o (n638) );
  assign n639 = N77 & n638 ;
  assign n640 = N77 | n638 ;
  assign n641 = ~n639 & n640 ;
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  assign n642 = n406 & n617 ;
  buffer buf_n643( .i (n642), .o (n643) );
  assign n644 = n372 & n643 ;
  buffer buf_n645( .i (n644), .o (n645) );
  assign n646 = n460 & n645 ;
  buffer buf_n647( .i (n646), .o (n647) );
  assign n648 = N81 | n647 ;
  assign n649 = N81 & n647 ;
  assign n650 = n648 & ~n649 ;
  assign n651 = n497 & n645 ;
  buffer buf_n652( .i (n651), .o (n652) );
  assign n653 = N85 | n652 ;
  assign n654 = N85 & n652 ;
  assign n655 = n653 & ~n654 ;
  assign n656 = n166 & n645 ;
  buffer buf_n657( .i (n656), .o (n657) );
  assign n658 = N89 & n657 ;
  assign n659 = N89 | n657 ;
  assign n660 = ~n658 & n659 ;
  assign n661 = n227 & n645 ;
  buffer buf_n662( .i (n661), .o (n662) );
  assign n663 = N93 | n662 ;
  assign n664 = N93 & n662 ;
  assign n665 = n663 & ~n664 ;
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  assign n666 = n346 & n619 ;
  buffer buf_n667( .i (n666), .o (n667) );
  assign n668 = n460 & n667 ;
  buffer buf_n669( .i (n668), .o (n669) );
  assign n670 = N97 | n669 ;
  assign n671 = N97 & n669 ;
  assign n672 = n670 & ~n671 ;
  assign n673 = n497 & n667 ;
  buffer buf_n674( .i (n673), .o (n674) );
  assign n675 = N101 | n674 ;
  assign n676 = N101 & n674 ;
  assign n677 = n675 & ~n676 ;
  assign n678 = n166 & n667 ;
  buffer buf_n679( .i (n678), .o (n679) );
  assign n680 = ~N105 & n679 ;
  assign n681 = N105 & ~n679 ;
  assign n682 = n680 | n681 ;
  assign n683 = n227 & n667 ;
  buffer buf_n684( .i (n683), .o (n684) );
  assign n685 = N109 & n684 ;
  assign n686 = N109 | n684 ;
  assign n687 = ~n685 & n686 ;
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  assign n688 = n354 & n643 ;
  buffer buf_n689( .i (n688), .o (n689) );
  assign n690 = n460 & n689 ;
  buffer buf_n691( .i (n690), .o (n691) );
  assign n692 = N113 | n691 ;
  assign n693 = N113 & n691 ;
  assign n694 = n692 & ~n693 ;
  assign n695 = n497 & n689 ;
  buffer buf_n696( .i (n695), .o (n696) );
  assign n697 = N117 | n696 ;
  assign n698 = N117 & n696 ;
  assign n699 = n697 & ~n698 ;
  assign n700 = n166 & n689 ;
  buffer buf_n701( .i (n700), .o (n701) );
  assign n702 = N121 & n701 ;
  assign n703 = N121 | n701 ;
  assign n704 = ~n702 & n703 ;
  assign n705 = n227 & n689 ;
  buffer buf_n706( .i (n705), .o (n706) );
  assign n707 = N125 | n706 ;
  assign n708 = N125 & n706 ;
  assign n709 = n707 & ~n708 ;
  assign N724 = n512 ;
  assign N725 = n517 ;
  assign N726 = n522 ;
  assign N727 = n527 ;
  assign N728 = n542 ;
  assign N729 = n547 ;
  assign N730 = n552 ;
  assign N731 = n557 ;
  assign N732 = n572 ;
  assign N733 = n577 ;
  assign N734 = n582 ;
  assign N735 = n587 ;
  assign N736 = n594 ;
  assign N737 = n599 ;
  assign N738 = n604 ;
  assign N739 = n609 ;
  assign N740 = n626 ;
  assign N741 = n631 ;
  assign N742 = n636 ;
  assign N743 = n641 ;
  assign N744 = n650 ;
  assign N745 = n655 ;
  assign N746 = n660 ;
  assign N747 = n665 ;
  assign N748 = n672 ;
  assign N749 = n677 ;
  assign N750 = n682 ;
  assign N751 = n687 ;
  assign N752 = n694 ;
  assign N753 = n699 ;
  assign N754 = n704 ;
  assign N755 = n709 ;
endmodule
