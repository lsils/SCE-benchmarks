module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( in_18_ , in_1_ , in_7_ , in_109_ , in_13_ , in_106_ , in_54_ , in_118_ , in_101_ , in_3_ , in_0_ , in_113_ , in_56_ , in_30_ , in_89_ , in_35_ , in_70_ , in_38_ , in_100_ , in_105_ , in_28_ , in_10_ , in_9_ , in_78_ , in_29_ , in_60_ , in_94_ , in_108_ , in_117_ , in_103_ , in_67_ , in_44_ , in_57_ , in_76_ , in_47_ , in_20_ , in_84_ , in_17_ , in_72_ , in_116_ , in_16_ , in_120_ , in_104_ , in_64_ , in_125_ , in_58_ , in_42_ , in_40_ , in_81_ , in_115_ , in_88_ , in_24_ , in_33_ , in_123_ , in_61_ , in_79_ , in_31_ , in_36_ , in_82_ , in_111_ , in_68_ , in_2_ , in_87_ , in_74_ , in_114_ , in_53_ , in_83_ , in_86_ , in_65_ , in_102_ , in_6_ , in_75_ , in_4_ , in_93_ , in_45_ , in_90_ , in_80_ , in_73_ , in_46_ , in_25_ , in_107_ , in_37_ , in_85_ , in_49_ , in_39_ , in_63_ , in_12_ , in_112_ , in_32_ , in_119_ , in_77_ , in_34_ , in_41_ , in_122_ , in_124_ , in_48_ , in_92_ , in_15_ , in_55_ , in_50_ , in_5_ , in_127_ , in_96_ , in_22_ , in_43_ , in_52_ , in_51_ , in_21_ , in_95_ , in_59_ , in_69_ , in_121_ , in_97_ , in_11_ , in_98_ , in_126_ , in_14_ , in_91_ , in_26_ , in_99_ , in_27_ , in_71_ , in_8_ , in_23_ , in_110_ , in_62_ , in_66_ , in_19_ , out_3_ , out_2_ , out_5_ , out_1_ , out_0_ , out_7_ , out_4_ , out_6_ );
  input in_18_ , in_1_ , in_7_ , in_109_ , in_13_ , in_106_ , in_54_ , in_118_ , in_101_ , in_3_ , in_0_ , in_113_ , in_56_ , in_30_ , in_89_ , in_35_ , in_70_ , in_38_ , in_100_ , in_105_ , in_28_ , in_10_ , in_9_ , in_78_ , in_29_ , in_60_ , in_94_ , in_108_ , in_117_ , in_103_ , in_67_ , in_44_ , in_57_ , in_76_ , in_47_ , in_20_ , in_84_ , in_17_ , in_72_ , in_116_ , in_16_ , in_120_ , in_104_ , in_64_ , in_125_ , in_58_ , in_42_ , in_40_ , in_81_ , in_115_ , in_88_ , in_24_ , in_33_ , in_123_ , in_61_ , in_79_ , in_31_ , in_36_ , in_82_ , in_111_ , in_68_ , in_2_ , in_87_ , in_74_ , in_114_ , in_53_ , in_83_ , in_86_ , in_65_ , in_102_ , in_6_ , in_75_ , in_4_ , in_93_ , in_45_ , in_90_ , in_80_ , in_73_ , in_46_ , in_25_ , in_107_ , in_37_ , in_85_ , in_49_ , in_39_ , in_63_ , in_12_ , in_112_ , in_32_ , in_119_ , in_77_ , in_34_ , in_41_ , in_122_ , in_124_ , in_48_ , in_92_ , in_15_ , in_55_ , in_50_ , in_5_ , in_127_ , in_96_ , in_22_ , in_43_ , in_52_ , in_51_ , in_21_ , in_95_ , in_59_ , in_69_ , in_121_ , in_97_ , in_11_ , in_98_ , in_126_ , in_14_ , in_91_ , in_26_ , in_99_ , in_27_ , in_71_ , in_8_ , in_23_ , in_110_ , in_62_ , in_66_ , in_19_ ;
  output out_3_ , out_2_ , out_5_ , out_1_ , out_0_ , out_7_ , out_4_ , out_6_ ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 ;
  assign n129 = in_127_ & in_126_ ;
  buffer buf_n130( .i (n129), .o (n130) );
  assign n131 = in_125_ | in_124_ ;
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  assign n135 = in_117_ | in_116_ ;
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  assign n139 = in_113_ | in_112_ ;
  buffer buf_n140( .i (n139), .o (n140) );
  assign n141 = in_115_ & in_114_ ;
  buffer buf_n142( .i (n141), .o (n142) );
  assign n143 = ( n136 & n140 ) | ( n136 & n142 ) | ( n140 & n142 ) ;
  buffer buf_n144( .i (n143), .o (n144) );
  assign n149 = ( ~n136 & n140 ) | ( ~n136 & n142 ) | ( n140 & n142 ) ;
  buffer buf_n150( .i (n149), .o (n150) );
  assign n151 = ( n138 & ~n144 ) | ( n138 & n150 ) | ( ~n144 & n150 ) ;
  buffer buf_n152( .i (n151), .o (n152) );
  assign n153 = in_123_ & in_122_ ;
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  assign n157 = in_118_ & in_119_ ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n159 = in_120_ | in_121_ ;
  buffer buf_n160( .i (n159), .o (n160) );
  assign n161 = ( n154 & n158 ) | ( n154 & n160 ) | ( n158 & n160 ) ;
  buffer buf_n162( .i (n161), .o (n162) );
  assign n167 = ( ~n154 & n158 ) | ( ~n154 & n160 ) | ( n158 & n160 ) ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = ( n156 & ~n162 ) | ( n156 & n168 ) | ( ~n162 & n168 ) ;
  buffer buf_n170( .i (n169), .o (n170) );
  assign n171 = ( n132 & n152 ) | ( n132 & n170 ) | ( n152 & n170 ) ;
  buffer buf_n172( .i (n171), .o (n172) );
  assign n175 = ( ~n132 & n152 ) | ( ~n132 & n170 ) | ( n152 & n170 ) ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n177 = ( n134 & ~n172 ) | ( n134 & n176 ) | ( ~n172 & n176 ) ;
  buffer buf_n178( .i (n177), .o (n178) );
  assign n179 = n130 & n178 ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = n130 | n178 ;
  buffer buf_n182( .i (n181), .o (n182) );
  assign n183 = ~n180 & n182 ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n185 = in_111_ & in_110_ ;
  buffer buf_n186( .i (n185), .o (n186) );
  assign n187 = in_109_ | in_108_ ;
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  assign n191 = in_101_ | in_100_ ;
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  assign n195 = in_96_ | in_97_ ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n197 = in_98_ & in_99_ ;
  buffer buf_n198( .i (n197), .o (n198) );
  assign n199 = ( ~n192 & n196 ) | ( ~n192 & n198 ) | ( n196 & n198 ) ;
  buffer buf_n200( .i (n199), .o (n200) );
  assign n201 = ( n192 & n196 ) | ( n192 & n198 ) | ( n196 & n198 ) ;
  buffer buf_n202( .i (n201), .o (n202) );
  assign n207 = ( n194 & n200 ) | ( n194 & ~n202 ) | ( n200 & ~n202 ) ;
  buffer buf_n208( .i (n207), .o (n208) );
  assign n209 = in_106_ & in_107_ ;
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  assign n213 = in_103_ & in_102_ ;
  buffer buf_n214( .i (n213), .o (n214) );
  assign n215 = in_105_ | in_104_ ;
  buffer buf_n216( .i (n215), .o (n216) );
  assign n217 = ( n210 & n214 ) | ( n210 & n216 ) | ( n214 & n216 ) ;
  buffer buf_n218( .i (n217), .o (n218) );
  assign n223 = ( ~n210 & n214 ) | ( ~n210 & n216 ) | ( n214 & n216 ) ;
  buffer buf_n224( .i (n223), .o (n224) );
  assign n225 = ( n212 & ~n218 ) | ( n212 & n224 ) | ( ~n218 & n224 ) ;
  buffer buf_n226( .i (n225), .o (n226) );
  assign n227 = ( n188 & n208 ) | ( n188 & n226 ) | ( n208 & n226 ) ;
  buffer buf_n228( .i (n227), .o (n228) );
  assign n231 = ( ~n188 & n208 ) | ( ~n188 & n226 ) | ( n208 & n226 ) ;
  buffer buf_n232( .i (n231), .o (n232) );
  assign n233 = ( n190 & ~n228 ) | ( n190 & n232 ) | ( ~n228 & n232 ) ;
  buffer buf_n234( .i (n233), .o (n234) );
  assign n235 = n186 & n234 ;
  buffer buf_n236( .i (n235), .o (n236) );
  assign n237 = n186 | n234 ;
  buffer buf_n238( .i (n237), .o (n238) );
  assign n239 = ~n236 & n238 ;
  buffer buf_n240( .i (n239), .o (n240) );
  assign n241 = n184 & n240 ;
  buffer buf_n242( .i (n241), .o (n242) );
  assign n246 = n184 | n240 ;
  buffer buf_n247( .i (n246), .o (n247) );
  assign n248 = ~n242 & n247 ;
  buffer buf_n249( .i (n248), .o (n249) );
  assign n250 = in_94_ & in_95_ ;
  buffer buf_n251( .i (n250), .o (n251) );
  assign n252 = in_93_ | in_92_ ;
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  assign n256 = in_84_ | in_85_ ;
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  assign n260 = in_81_ | in_80_ ;
  buffer buf_n261( .i (n260), .o (n261) );
  assign n262 = in_82_ & in_83_ ;
  buffer buf_n263( .i (n262), .o (n263) );
  assign n264 = ( n257 & n261 ) | ( n257 & n263 ) | ( n261 & n263 ) ;
  buffer buf_n265( .i (n264), .o (n265) );
  assign n270 = ( ~n257 & n261 ) | ( ~n257 & n263 ) | ( n261 & n263 ) ;
  buffer buf_n271( .i (n270), .o (n271) );
  assign n272 = ( n259 & ~n265 ) | ( n259 & n271 ) | ( ~n265 & n271 ) ;
  buffer buf_n273( .i (n272), .o (n273) );
  assign n274 = in_90_ & in_91_ ;
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  assign n278 = in_87_ & in_86_ ;
  buffer buf_n279( .i (n278), .o (n279) );
  assign n280 = in_89_ | in_88_ ;
  buffer buf_n281( .i (n280), .o (n281) );
  assign n282 = ( n275 & n279 ) | ( n275 & n281 ) | ( n279 & n281 ) ;
  buffer buf_n283( .i (n282), .o (n283) );
  assign n288 = ( ~n275 & n279 ) | ( ~n275 & n281 ) | ( n279 & n281 ) ;
  buffer buf_n289( .i (n288), .o (n289) );
  assign n290 = ( n277 & ~n283 ) | ( n277 & n289 ) | ( ~n283 & n289 ) ;
  buffer buf_n291( .i (n290), .o (n291) );
  assign n292 = ( n253 & n273 ) | ( n253 & n291 ) | ( n273 & n291 ) ;
  buffer buf_n293( .i (n292), .o (n293) );
  assign n296 = ( ~n253 & n273 ) | ( ~n253 & n291 ) | ( n273 & n291 ) ;
  buffer buf_n297( .i (n296), .o (n297) );
  assign n298 = ( n255 & ~n293 ) | ( n255 & n297 ) | ( ~n293 & n297 ) ;
  buffer buf_n299( .i (n298), .o (n299) );
  assign n300 = n251 & n299 ;
  buffer buf_n301( .i (n300), .o (n301) );
  assign n302 = n251 | n299 ;
  buffer buf_n303( .i (n302), .o (n303) );
  assign n304 = ~n301 & n303 ;
  buffer buf_n305( .i (n304), .o (n305) );
  assign n306 = in_78_ & in_79_ ;
  buffer buf_n307( .i (n306), .o (n307) );
  assign n308 = in_76_ | in_77_ ;
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  assign n312 = in_68_ | in_69_ ;
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  assign n316 = in_64_ | in_65_ ;
  buffer buf_n317( .i (n316), .o (n317) );
  assign n318 = in_67_ & in_66_ ;
  buffer buf_n319( .i (n318), .o (n319) );
  assign n320 = ( n313 & n317 ) | ( n313 & n319 ) | ( n317 & n319 ) ;
  buffer buf_n321( .i (n320), .o (n321) );
  assign n326 = ( ~n313 & n317 ) | ( ~n313 & n319 ) | ( n317 & n319 ) ;
  buffer buf_n327( .i (n326), .o (n327) );
  assign n328 = ( n315 & ~n321 ) | ( n315 & n327 ) | ( ~n321 & n327 ) ;
  buffer buf_n329( .i (n328), .o (n329) );
  assign n330 = in_74_ & in_75_ ;
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  assign n334 = in_70_ & in_71_ ;
  buffer buf_n335( .i (n334), .o (n335) );
  assign n336 = in_72_ | in_73_ ;
  buffer buf_n337( .i (n336), .o (n337) );
  assign n338 = ( n331 & n335 ) | ( n331 & n337 ) | ( n335 & n337 ) ;
  buffer buf_n339( .i (n338), .o (n339) );
  assign n344 = ( ~n331 & n335 ) | ( ~n331 & n337 ) | ( n335 & n337 ) ;
  buffer buf_n345( .i (n344), .o (n345) );
  assign n346 = ( n333 & ~n339 ) | ( n333 & n345 ) | ( ~n339 & n345 ) ;
  buffer buf_n347( .i (n346), .o (n347) );
  assign n348 = ( n309 & n329 ) | ( n309 & n347 ) | ( n329 & n347 ) ;
  buffer buf_n349( .i (n348), .o (n349) );
  assign n352 = ( ~n309 & n329 ) | ( ~n309 & n347 ) | ( n329 & n347 ) ;
  buffer buf_n353( .i (n352), .o (n353) );
  assign n354 = ( n311 & ~n349 ) | ( n311 & n353 ) | ( ~n349 & n353 ) ;
  buffer buf_n355( .i (n354), .o (n355) );
  assign n356 = n307 & n355 ;
  buffer buf_n357( .i (n356), .o (n357) );
  assign n358 = n307 | n355 ;
  buffer buf_n359( .i (n358), .o (n359) );
  assign n360 = ~n357 & n359 ;
  buffer buf_n361( .i (n360), .o (n361) );
  assign n362 = n305 & n361 ;
  buffer buf_n363( .i (n362), .o (n363) );
  assign n367 = n305 | n361 ;
  buffer buf_n368( .i (n367), .o (n368) );
  assign n369 = ~n363 & n368 ;
  buffer buf_n370( .i (n369), .o (n370) );
  assign n371 = n249 & n370 ;
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  assign n378 = ( n148 & n166 ) | ( n148 & n172 ) | ( n166 & n172 ) ;
  buffer buf_n379( .i (n378), .o (n379) );
  assign n384 = ( n148 & n166 ) | ( n148 & ~n172 ) | ( n166 & ~n172 ) ;
  buffer buf_n385( .i (n384), .o (n385) );
  assign n386 = ( n174 & ~n379 ) | ( n174 & n385 ) | ( ~n379 & n385 ) ;
  buffer buf_n387( .i (n386), .o (n387) );
  assign n388 = n180 & n387 ;
  buffer buf_n389( .i (n388), .o (n389) );
  assign n390 = n180 | n387 ;
  buffer buf_n391( .i (n390), .o (n391) );
  assign n392 = ~n389 & n391 ;
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  assign n394 = ( n206 & n222 ) | ( n206 & n228 ) | ( n222 & n228 ) ;
  buffer buf_n395( .i (n394), .o (n395) );
  assign n400 = ( n206 & n222 ) | ( n206 & ~n228 ) | ( n222 & ~n228 ) ;
  buffer buf_n401( .i (n400), .o (n401) );
  assign n402 = ( n230 & ~n395 ) | ( n230 & n401 ) | ( ~n395 & n401 ) ;
  buffer buf_n403( .i (n402), .o (n403) );
  assign n404 = n236 & n403 ;
  buffer buf_n405( .i (n404), .o (n405) );
  assign n406 = n236 | n403 ;
  buffer buf_n407( .i (n406), .o (n407) );
  assign n408 = ~n405 & n407 ;
  buffer buf_n409( .i (n408), .o (n409) );
  assign n410 = n393 & n409 ;
  assign n411 = n393 | n409 ;
  assign n412 = ~n410 & n411 ;
  buffer buf_n413( .i (n412), .o (n413) );
  assign n414 = n245 & n413 ;
  assign n415 = n245 | n413 ;
  assign n416 = ~n414 & n415 ;
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  assign n418 = ( n269 & n287 ) | ( n269 & n293 ) | ( n287 & n293 ) ;
  buffer buf_n419( .i (n418), .o (n419) );
  assign n424 = ( n269 & n287 ) | ( n269 & ~n293 ) | ( n287 & ~n293 ) ;
  buffer buf_n425( .i (n424), .o (n425) );
  assign n426 = ( n295 & ~n419 ) | ( n295 & n425 ) | ( ~n419 & n425 ) ;
  buffer buf_n427( .i (n426), .o (n427) );
  assign n428 = n301 & n427 ;
  buffer buf_n429( .i (n428), .o (n429) );
  assign n430 = n301 | n427 ;
  buffer buf_n431( .i (n430), .o (n431) );
  assign n432 = ~n429 & n431 ;
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  assign n434 = ( n325 & n343 ) | ( n325 & n349 ) | ( n343 & n349 ) ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n440 = ( n325 & n343 ) | ( n325 & ~n349 ) | ( n343 & ~n349 ) ;
  buffer buf_n441( .i (n440), .o (n441) );
  assign n442 = ( n351 & ~n435 ) | ( n351 & n441 ) | ( ~n435 & n441 ) ;
  buffer buf_n443( .i (n442), .o (n443) );
  assign n444 = n357 & n443 ;
  buffer buf_n445( .i (n444), .o (n445) );
  assign n446 = n357 | n443 ;
  buffer buf_n447( .i (n446), .o (n447) );
  assign n448 = ~n445 & n447 ;
  buffer buf_n449( .i (n448), .o (n449) );
  assign n450 = n433 & n449 ;
  assign n451 = n433 | n449 ;
  assign n452 = ~n450 & n451 ;
  buffer buf_n453( .i (n452), .o (n453) );
  assign n454 = n366 & n453 ;
  assign n455 = n366 | n453 ;
  assign n456 = ~n454 & n455 ;
  buffer buf_n457( .i (n456), .o (n457) );
  assign n458 = n417 & n457 ;
  assign n459 = n417 | n457 ;
  assign n460 = ~n458 & n459 ;
  buffer buf_n461( .i (n460), .o (n461) );
  assign n462 = n377 & n461 ;
  assign n463 = n377 | n461 ;
  assign n464 = ~n462 & n463 ;
  buffer buf_n465( .i (n464), .o (n465) );
  assign n466 = n249 | n370 ;
  buffer buf_n467( .i (n466), .o (n467) );
  assign n468 = ~n372 & n467 ;
  buffer buf_n469( .i (n468), .o (n469) );
  assign n470 = in_30_ & in_31_ ;
  buffer buf_n471( .i (n470), .o (n471) );
  assign n472 = in_28_ | in_29_ ;
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  assign n476 = in_26_ & in_27_ ;
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  assign n480 = in_22_ & in_23_ ;
  buffer buf_n481( .i (n480), .o (n481) );
  assign n482 = in_24_ | in_25_ ;
  buffer buf_n483( .i (n482), .o (n483) );
  assign n484 = ( n477 & n481 ) | ( n477 & n483 ) | ( n481 & n483 ) ;
  buffer buf_n485( .i (n484), .o (n485) );
  assign n490 = ( ~n477 & n481 ) | ( ~n477 & n483 ) | ( n481 & n483 ) ;
  buffer buf_n491( .i (n490), .o (n491) );
  assign n492 = ( n479 & ~n485 ) | ( n479 & n491 ) | ( ~n485 & n491 ) ;
  buffer buf_n493( .i (n492), .o (n493) );
  assign n494 = in_20_ | in_21_ ;
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  assign n498 = in_17_ | in_16_ ;
  buffer buf_n499( .i (n498), .o (n499) );
  assign n500 = in_18_ & in_19_ ;
  buffer buf_n501( .i (n500), .o (n501) );
  assign n502 = ( n495 & n499 ) | ( n495 & n501 ) | ( n499 & n501 ) ;
  buffer buf_n503( .i (n502), .o (n503) );
  assign n508 = ( ~n495 & n499 ) | ( ~n495 & n501 ) | ( n499 & n501 ) ;
  buffer buf_n509( .i (n508), .o (n509) );
  assign n510 = ( n497 & ~n503 ) | ( n497 & n509 ) | ( ~n503 & n509 ) ;
  buffer buf_n511( .i (n510), .o (n511) );
  assign n512 = ( n473 & n493 ) | ( n473 & n511 ) | ( n493 & n511 ) ;
  buffer buf_n513( .i (n512), .o (n513) );
  assign n516 = ( ~n473 & n493 ) | ( ~n473 & n511 ) | ( n493 & n511 ) ;
  buffer buf_n517( .i (n516), .o (n517) );
  assign n518 = ( n475 & ~n513 ) | ( n475 & n517 ) | ( ~n513 & n517 ) ;
  buffer buf_n519( .i (n518), .o (n519) );
  assign n520 = n471 & n519 ;
  buffer buf_n521( .i (n520), .o (n521) );
  assign n522 = n471 | n519 ;
  buffer buf_n523( .i (n522), .o (n523) );
  assign n524 = ~n521 & n523 ;
  buffer buf_n525( .i (n524), .o (n525) );
  assign n526 = in_15_ & in_14_ ;
  buffer buf_n527( .i (n526), .o (n527) );
  assign n528 = in_13_ | in_12_ ;
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  assign n532 = in_4_ | in_5_ ;
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  assign n536 = in_1_ | in_0_ ;
  buffer buf_n537( .i (n536), .o (n537) );
  assign n538 = in_3_ & in_2_ ;
  buffer buf_n539( .i (n538), .o (n539) );
  assign n540 = ( n533 & n537 ) | ( n533 & n539 ) | ( n537 & n539 ) ;
  buffer buf_n541( .i (n540), .o (n541) );
  assign n546 = ( ~n533 & n537 ) | ( ~n533 & n539 ) | ( n537 & n539 ) ;
  buffer buf_n547( .i (n546), .o (n547) );
  assign n548 = ( n535 & ~n541 ) | ( n535 & n547 ) | ( ~n541 & n547 ) ;
  buffer buf_n549( .i (n548), .o (n549) );
  assign n550 = in_10_ & in_11_ ;
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  assign n554 = in_7_ & in_6_ ;
  buffer buf_n555( .i (n554), .o (n555) );
  assign n556 = in_9_ | in_8_ ;
  buffer buf_n557( .i (n556), .o (n557) );
  assign n558 = ( n551 & n555 ) | ( n551 & n557 ) | ( n555 & n557 ) ;
  buffer buf_n559( .i (n558), .o (n559) );
  assign n564 = ( ~n551 & n555 ) | ( ~n551 & n557 ) | ( n555 & n557 ) ;
  buffer buf_n565( .i (n564), .o (n565) );
  assign n566 = ( n553 & ~n559 ) | ( n553 & n565 ) | ( ~n559 & n565 ) ;
  buffer buf_n567( .i (n566), .o (n567) );
  assign n568 = ( n529 & n549 ) | ( n529 & n567 ) | ( n549 & n567 ) ;
  buffer buf_n569( .i (n568), .o (n569) );
  assign n572 = ( ~n529 & n549 ) | ( ~n529 & n567 ) | ( n549 & n567 ) ;
  buffer buf_n573( .i (n572), .o (n573) );
  assign n574 = ( n531 & ~n569 ) | ( n531 & n573 ) | ( ~n569 & n573 ) ;
  buffer buf_n575( .i (n574), .o (n575) );
  assign n576 = n527 & n575 ;
  buffer buf_n577( .i (n576), .o (n577) );
  assign n578 = n527 | n575 ;
  buffer buf_n579( .i (n578), .o (n579) );
  assign n580 = ~n577 & n579 ;
  buffer buf_n581( .i (n580), .o (n581) );
  assign n582 = n525 & n581 ;
  buffer buf_n583( .i (n582), .o (n583) );
  assign n587 = n525 | n581 ;
  buffer buf_n588( .i (n587), .o (n588) );
  assign n589 = ~n583 & n588 ;
  buffer buf_n590( .i (n589), .o (n590) );
  assign n591 = in_47_ & in_46_ ;
  buffer buf_n592( .i (n591), .o (n592) );
  assign n593 = in_44_ | in_45_ ;
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  assign n597 = in_36_ | in_37_ ;
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  assign n601 = in_33_ | in_32_ ;
  buffer buf_n602( .i (n601), .o (n602) );
  assign n603 = in_35_ & in_34_ ;
  buffer buf_n604( .i (n603), .o (n604) );
  assign n605 = ( n598 & n602 ) | ( n598 & n604 ) | ( n602 & n604 ) ;
  buffer buf_n606( .i (n605), .o (n606) );
  assign n611 = ( ~n598 & n602 ) | ( ~n598 & n604 ) | ( n602 & n604 ) ;
  buffer buf_n612( .i (n611), .o (n612) );
  assign n613 = ( n600 & ~n606 ) | ( n600 & n612 ) | ( ~n606 & n612 ) ;
  buffer buf_n614( .i (n613), .o (n614) );
  assign n615 = in_42_ & in_43_ ;
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  assign n619 = in_38_ & in_39_ ;
  buffer buf_n620( .i (n619), .o (n620) );
  assign n621 = in_40_ | in_41_ ;
  buffer buf_n622( .i (n621), .o (n622) );
  assign n623 = ( n616 & n620 ) | ( n616 & n622 ) | ( n620 & n622 ) ;
  buffer buf_n624( .i (n623), .o (n624) );
  assign n629 = ( ~n616 & n620 ) | ( ~n616 & n622 ) | ( n620 & n622 ) ;
  buffer buf_n630( .i (n629), .o (n630) );
  assign n631 = ( n618 & ~n624 ) | ( n618 & n630 ) | ( ~n624 & n630 ) ;
  buffer buf_n632( .i (n631), .o (n632) );
  assign n633 = ( n594 & n614 ) | ( n594 & n632 ) | ( n614 & n632 ) ;
  buffer buf_n634( .i (n633), .o (n634) );
  assign n637 = ( ~n594 & n614 ) | ( ~n594 & n632 ) | ( n614 & n632 ) ;
  buffer buf_n638( .i (n637), .o (n638) );
  assign n639 = ( n596 & ~n634 ) | ( n596 & n638 ) | ( ~n634 & n638 ) ;
  buffer buf_n640( .i (n639), .o (n640) );
  assign n641 = n592 & n640 ;
  buffer buf_n642( .i (n641), .o (n642) );
  assign n643 = n592 | n640 ;
  buffer buf_n644( .i (n643), .o (n644) );
  assign n645 = ~n642 & n644 ;
  buffer buf_n646( .i (n645), .o (n646) );
  assign n647 = in_63_ & in_62_ ;
  buffer buf_n648( .i (n647), .o (n648) );
  assign n649 = in_60_ | in_61_ ;
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  assign n653 = in_58_ & in_59_ ;
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  assign n657 = in_54_ & in_55_ ;
  buffer buf_n658( .i (n657), .o (n658) );
  assign n659 = in_56_ | in_57_ ;
  buffer buf_n660( .i (n659), .o (n660) );
  assign n661 = ( n654 & n658 ) | ( n654 & n660 ) | ( n658 & n660 ) ;
  buffer buf_n662( .i (n661), .o (n662) );
  assign n667 = ( ~n654 & n658 ) | ( ~n654 & n660 ) | ( n658 & n660 ) ;
  buffer buf_n668( .i (n667), .o (n668) );
  assign n669 = ( n656 & ~n662 ) | ( n656 & n668 ) | ( ~n662 & n668 ) ;
  buffer buf_n670( .i (n669), .o (n670) );
  assign n671 = in_53_ | in_52_ ;
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  assign n675 = in_49_ | in_48_ ;
  buffer buf_n676( .i (n675), .o (n676) );
  assign n677 = in_50_ & in_51_ ;
  buffer buf_n678( .i (n677), .o (n678) );
  assign n679 = ( n672 & n676 ) | ( n672 & n678 ) | ( n676 & n678 ) ;
  buffer buf_n680( .i (n679), .o (n680) );
  assign n685 = ( ~n672 & n676 ) | ( ~n672 & n678 ) | ( n676 & n678 ) ;
  buffer buf_n686( .i (n685), .o (n686) );
  assign n687 = ( n674 & ~n680 ) | ( n674 & n686 ) | ( ~n680 & n686 ) ;
  buffer buf_n688( .i (n687), .o (n688) );
  assign n689 = ( n650 & n670 ) | ( n650 & n688 ) | ( n670 & n688 ) ;
  buffer buf_n690( .i (n689), .o (n690) );
  assign n693 = ( ~n650 & n670 ) | ( ~n650 & n688 ) | ( n670 & n688 ) ;
  buffer buf_n694( .i (n693), .o (n694) );
  assign n695 = ( n652 & ~n690 ) | ( n652 & n694 ) | ( ~n690 & n694 ) ;
  buffer buf_n696( .i (n695), .o (n696) );
  assign n697 = n648 & n696 ;
  buffer buf_n698( .i (n697), .o (n698) );
  assign n699 = n648 | n696 ;
  buffer buf_n700( .i (n699), .o (n700) );
  assign n701 = ~n698 & n700 ;
  buffer buf_n702( .i (n701), .o (n702) );
  assign n703 = n646 | n702 ;
  buffer buf_n704( .i (n703), .o (n704) );
  assign n705 = n646 & n702 ;
  buffer buf_n706( .i (n705), .o (n706) );
  assign n710 = n704 & ~n706 ;
  buffer buf_n711( .i (n710), .o (n711) );
  assign n712 = n590 & n711 ;
  buffer buf_n713( .i (n712), .o (n713) );
  assign n719 = n590 | n711 ;
  buffer buf_n720( .i (n719), .o (n720) );
  assign n721 = ~n713 & n720 ;
  buffer buf_n722( .i (n721), .o (n722) );
  assign n723 = n469 & n722 ;
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  assign n732 = ( n489 & n507 ) | ( n489 & n513 ) | ( n507 & n513 ) ;
  buffer buf_n733( .i (n732), .o (n733) );
  assign n738 = ( n489 & n507 ) | ( n489 & ~n513 ) | ( n507 & ~n513 ) ;
  buffer buf_n739( .i (n738), .o (n739) );
  assign n740 = ( n515 & ~n733 ) | ( n515 & n739 ) | ( ~n733 & n739 ) ;
  buffer buf_n741( .i (n740), .o (n741) );
  assign n742 = n521 | n741 ;
  buffer buf_n743( .i (n742), .o (n743) );
  assign n744 = n521 & n741 ;
  buffer buf_n745( .i (n744), .o (n745) );
  assign n746 = n743 & ~n745 ;
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  assign n748 = ( n545 & n563 ) | ( n545 & n569 ) | ( n563 & n569 ) ;
  buffer buf_n749( .i (n748), .o (n749) );
  assign n754 = ( n545 & n563 ) | ( n545 & ~n569 ) | ( n563 & ~n569 ) ;
  buffer buf_n755( .i (n754), .o (n755) );
  assign n756 = ( n571 & ~n749 ) | ( n571 & n755 ) | ( ~n749 & n755 ) ;
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = n577 & n757 ;
  buffer buf_n759( .i (n758), .o (n759) );
  assign n760 = n577 | n757 ;
  buffer buf_n761( .i (n760), .o (n761) );
  assign n762 = ~n759 & n761 ;
  buffer buf_n763( .i (n762), .o (n763) );
  assign n764 = n747 & n763 ;
  assign n765 = n747 | n763 ;
  assign n766 = ~n764 & n765 ;
  buffer buf_n767( .i (n766), .o (n767) );
  assign n768 = n586 & n767 ;
  assign n769 = n586 | n767 ;
  assign n770 = ~n768 & n769 ;
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  assign n772 = ( n666 & n684 ) | ( n666 & n690 ) | ( n684 & n690 ) ;
  buffer buf_n773( .i (n772), .o (n773) );
  assign n778 = ( n666 & n684 ) | ( n666 & ~n690 ) | ( n684 & ~n690 ) ;
  buffer buf_n779( .i (n778), .o (n779) );
  assign n780 = ( n692 & ~n773 ) | ( n692 & n779 ) | ( ~n773 & n779 ) ;
  buffer buf_n781( .i (n780), .o (n781) );
  assign n782 = n698 & n781 ;
  buffer buf_n783( .i (n782), .o (n783) );
  assign n784 = n698 | n781 ;
  buffer buf_n785( .i (n784), .o (n785) );
  assign n786 = ~n783 & n785 ;
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  assign n788 = ( n610 & n628 ) | ( n610 & n634 ) | ( n628 & n634 ) ;
  buffer buf_n789( .i (n788), .o (n789) );
  assign n794 = ( n610 & n628 ) | ( n610 & ~n634 ) | ( n628 & ~n634 ) ;
  buffer buf_n795( .i (n794), .o (n795) );
  assign n796 = ( n636 & ~n789 ) | ( n636 & n795 ) | ( ~n789 & n795 ) ;
  buffer buf_n797( .i (n796), .o (n797) );
  assign n798 = n642 & n797 ;
  buffer buf_n799( .i (n798), .o (n799) );
  assign n800 = n642 | n797 ;
  buffer buf_n801( .i (n800), .o (n801) );
  assign n802 = ~n799 & n801 ;
  buffer buf_n803( .i (n802), .o (n803) );
  assign n804 = n787 & n803 ;
  assign n805 = n787 | n803 ;
  assign n806 = ~n804 & n805 ;
  buffer buf_n807( .i (n806), .o (n807) );
  assign n808 = n709 & n807 ;
  assign n809 = n709 | n807 ;
  assign n810 = ~n808 & n809 ;
  buffer buf_n811( .i (n810), .o (n811) );
  assign n812 = n771 & n811 ;
  assign n813 = n771 | n811 ;
  assign n814 = ~n812 & n813 ;
  buffer buf_n815( .i (n814), .o (n815) );
  assign n816 = n718 & n815 ;
  assign n817 = n718 | n815 ;
  assign n818 = ~n816 & n817 ;
  buffer buf_n819( .i (n818), .o (n819) );
  assign n820 = ( n465 & n728 ) | ( n465 & n819 ) | ( n728 & n819 ) ;
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  assign n825 = ( n715 & n771 ) | ( n715 & n811 ) | ( n771 & n811 ) ;
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  assign n830 = ( n583 & n747 ) | ( n583 & n763 ) | ( n747 & n763 ) ;
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  assign n835 = n737 & n745 ;
  buffer buf_n836( .i (n835), .o (n836) );
  assign n841 = n737 | n745 ;
  buffer buf_n842( .i (n841), .o (n842) );
  assign n843 = ~n836 & n842 ;
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  assign n845 = n753 & n759 ;
  buffer buf_n846( .i (n845), .o (n846) );
  assign n851 = n753 | n759 ;
  buffer buf_n852( .i (n851), .o (n852) );
  assign n853 = ~n846 & n852 ;
  buffer buf_n854( .i (n853), .o (n854) );
  assign n855 = n844 & n854 ;
  assign n856 = n844 | n854 ;
  assign n857 = ~n855 & n856 ;
  buffer buf_n858( .i (n857), .o (n858) );
  assign n859 = n834 & n858 ;
  assign n860 = n834 | n858 ;
  assign n861 = ~n859 & n860 ;
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  assign n863 = n793 & n799 ;
  buffer buf_n864( .i (n863), .o (n864) );
  assign n869 = n793 | n799 ;
  buffer buf_n870( .i (n869), .o (n870) );
  assign n871 = ~n864 & n870 ;
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  assign n873 = n777 & n783 ;
  buffer buf_n874( .i (n873), .o (n874) );
  assign n879 = n777 | n783 ;
  buffer buf_n880( .i (n879), .o (n880) );
  assign n881 = ~n874 & n880 ;
  buffer buf_n882( .i (n881), .o (n882) );
  assign n883 = n872 & n882 ;
  assign n884 = n872 | n882 ;
  assign n885 = ~n883 & n884 ;
  buffer buf_n886( .i (n885), .o (n886) );
  assign n887 = ( n706 & n787 ) | ( n706 & n803 ) | ( n787 & n803 ) ;
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  assign n892 = n886 & n891 ;
  assign n893 = n886 | n891 ;
  assign n894 = ~n892 & n893 ;
  buffer buf_n895( .i (n894), .o (n895) );
  assign n896 = n862 & n895 ;
  assign n897 = n862 | n895 ;
  assign n898 = ~n896 & n897 ;
  buffer buf_n899( .i (n898), .o (n899) );
  assign n900 = n829 & n899 ;
  assign n901 = n829 | n899 ;
  assign n902 = ~n900 & n901 ;
  buffer buf_n903( .i (n902), .o (n903) );
  assign n904 = ( n374 & n417 ) | ( n374 & n457 ) | ( n417 & n457 ) ;
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  assign n909 = ( n242 & n393 ) | ( n242 & n409 ) | ( n393 & n409 ) ;
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  assign n914 = n383 & n389 ;
  buffer buf_n915( .i (n914), .o (n915) );
  assign n920 = n383 | n389 ;
  buffer buf_n921( .i (n920), .o (n921) );
  assign n922 = ~n915 & n921 ;
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  assign n924 = n399 & n405 ;
  buffer buf_n925( .i (n924), .o (n925) );
  assign n930 = n399 | n405 ;
  buffer buf_n931( .i (n930), .o (n931) );
  assign n932 = ~n925 & n931 ;
  buffer buf_n933( .i (n932), .o (n933) );
  assign n934 = n923 & n933 ;
  assign n935 = n923 | n933 ;
  assign n936 = ~n934 & n935 ;
  buffer buf_n937( .i (n936), .o (n937) );
  assign n938 = n913 & n937 ;
  assign n939 = n913 | n937 ;
  assign n940 = ~n938 & n939 ;
  buffer buf_n941( .i (n940), .o (n941) );
  assign n942 = ( n363 & n433 ) | ( n363 & n449 ) | ( n433 & n449 ) ;
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  assign n947 = n423 & n429 ;
  buffer buf_n948( .i (n947), .o (n948) );
  assign n953 = n423 | n429 ;
  buffer buf_n954( .i (n953), .o (n954) );
  assign n955 = ~n948 & n954 ;
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  assign n957 = n439 & n445 ;
  buffer buf_n958( .i (n957), .o (n958) );
  assign n963 = n439 | n445 ;
  buffer buf_n964( .i (n963), .o (n964) );
  assign n965 = ~n958 & n964 ;
  buffer buf_n966( .i (n965), .o (n966) );
  assign n967 = n956 & n966 ;
  assign n968 = n956 | n966 ;
  assign n969 = ~n967 & n968 ;
  buffer buf_n970( .i (n969), .o (n970) );
  assign n971 = n946 & n970 ;
  assign n972 = n946 | n970 ;
  assign n973 = ~n971 & n972 ;
  buffer buf_n974( .i (n973), .o (n974) );
  assign n975 = n941 & n974 ;
  assign n976 = n941 | n974 ;
  assign n977 = ~n975 & n976 ;
  buffer buf_n978( .i (n977), .o (n978) );
  assign n979 = n908 & n978 ;
  assign n980 = n908 | n978 ;
  assign n981 = ~n979 & n980 ;
  buffer buf_n982( .i (n981), .o (n982) );
  assign n983 = n903 & n982 ;
  assign n984 = n903 | n982 ;
  assign n985 = ~n983 & n984 ;
  buffer buf_n986( .i (n985), .o (n986) );
  assign n987 = n824 & n986 ;
  assign n988 = n824 | n986 ;
  assign n989 = ~n987 & n988 ;
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  assign n990 = n465 & n819 ;
  assign n991 = n465 | n819 ;
  assign n992 = ~n990 & n991 ;
  buffer buf_n993( .i (n992), .o (n993) );
  assign n994 = n731 & n993 ;
  assign n995 = n731 | n993 ;
  assign n996 = ~n994 & n995 ;
  assign n997 = ( n826 & n862 ) | ( n826 & n895 ) | ( n862 & n895 ) ;
  buffer buf_n998( .i (n997), .o (n998) );
  assign n999 = n836 & n846 ;
  assign n1000 = n836 | n846 ;
  assign n1001 = ~n999 & n1000 ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  assign n1004 = ( n831 & n844 ) | ( n831 & n854 ) | ( n844 & n854 ) ;
  buffer buf_n1005( .i (n1004), .o (n1005) );
  assign n1006 = n1003 & n1005 ;
  assign n1007 = n1003 | n1005 ;
  assign n1008 = ~n1006 & n1007 ;
  buffer buf_n1009( .i (n1008), .o (n1009) );
  assign n1013 = n864 & n874 ;
  assign n1014 = n864 | n874 ;
  assign n1015 = ~n1013 & n1014 ;
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  assign n1018 = ( n872 & n882 ) | ( n872 & n888 ) | ( n882 & n888 ) ;
  buffer buf_n1019( .i (n1018), .o (n1019) );
  assign n1020 = n1017 & n1019 ;
  assign n1021 = n1017 | n1019 ;
  assign n1022 = ~n1020 & n1021 ;
  buffer buf_n1023( .i (n1022), .o (n1023) );
  assign n1027 = n1009 & n1023 ;
  assign n1028 = n1009 | n1023 ;
  assign n1029 = ~n1027 & n1028 ;
  buffer buf_n1030( .i (n1029), .o (n1030) );
  assign n1031 = n998 & n1030 ;
  assign n1032 = n998 | n1030 ;
  assign n1033 = ~n1031 & n1032 ;
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  assign n1038 = ( n821 & n903 ) | ( n821 & n982 ) | ( n903 & n982 ) ;
  buffer buf_n1039( .i (n1038), .o (n1039) );
  assign n1040 = n915 & n925 ;
  assign n1041 = n915 | n925 ;
  assign n1042 = ~n1040 & n1041 ;
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  assign n1045 = ( n910 & n923 ) | ( n910 & n933 ) | ( n923 & n933 ) ;
  buffer buf_n1046( .i (n1045), .o (n1046) );
  assign n1047 = n1044 & n1046 ;
  assign n1048 = n1044 | n1046 ;
  assign n1049 = ~n1047 & n1048 ;
  buffer buf_n1050( .i (n1049), .o (n1050) );
  assign n1054 = n948 & n958 ;
  assign n1055 = n948 | n958 ;
  assign n1056 = ~n1054 & n1055 ;
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  assign n1059 = ( n943 & n956 ) | ( n943 & n966 ) | ( n956 & n966 ) ;
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1061 = n1058 & n1060 ;
  assign n1062 = n1058 | n1060 ;
  assign n1063 = ~n1061 & n1062 ;
  buffer buf_n1064( .i (n1063), .o (n1064) );
  assign n1068 = n1050 & n1064 ;
  assign n1069 = n1050 | n1064 ;
  assign n1070 = ~n1068 & n1069 ;
  buffer buf_n1071( .i (n1070), .o (n1071) );
  assign n1072 = ( n905 & n941 ) | ( n905 & n974 ) | ( n941 & n974 ) ;
  buffer buf_n1073( .i (n1072), .o (n1073) );
  assign n1074 = n1071 & n1073 ;
  assign n1075 = n1071 | n1073 ;
  assign n1076 = ~n1074 & n1075 ;
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  assign n1081 = ( n1037 & n1039 ) | ( n1037 & n1080 ) | ( n1039 & n1080 ) ;
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  assign n1083 = ( n998 & n1012 ) | ( n998 & n1026 ) | ( n1012 & n1026 ) ;
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  assign n1085 = ( n840 & n850 ) | ( n840 & n1005 ) | ( n850 & n1005 ) ;
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  assign n1093 = ( n868 & n878 ) | ( n868 & n1019 ) | ( n878 & n1019 ) ;
  buffer buf_n1094( .i (n1093), .o (n1094) );
  assign n1101 = n1086 & n1094 ;
  assign n1102 = n1086 | n1094 ;
  assign n1103 = ~n1101 & n1102 ;
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  assign n1108 = n1084 & n1107 ;
  assign n1109 = n1084 | n1107 ;
  assign n1110 = ~n1108 & n1109 ;
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  assign n1115 = ( n919 & n929 ) | ( n919 & n1046 ) | ( n929 & n1046 ) ;
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  assign n1123 = ( n952 & n962 ) | ( n952 & n1060 ) | ( n962 & n1060 ) ;
  buffer buf_n1124( .i (n1123), .o (n1124) );
  assign n1131 = n1116 & n1124 ;
  assign n1132 = n1116 | n1124 ;
  assign n1133 = ~n1131 & n1132 ;
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  assign n1138 = ( n1053 & n1067 ) | ( n1053 & n1073 ) | ( n1067 & n1073 ) ;
  buffer buf_n1139( .i (n1138), .o (n1139) );
  assign n1140 = n1137 & n1139 ;
  assign n1141 = n1137 | n1139 ;
  assign n1142 = ~n1140 & n1141 ;
  buffer buf_n1143( .i (n1142), .o (n1143) );
  assign n1147 = n1111 & n1143 ;
  assign n1148 = n1111 | n1143 ;
  assign n1149 = ~n1147 & n1148 ;
  buffer buf_n1150( .i (n1149), .o (n1150) );
  assign n1151 = n1082 & n1150 ;
  assign n1152 = n1082 | n1150 ;
  assign n1153 = ~n1151 & n1152 ;
  assign n1154 = n469 | n722 ;
  buffer buf_n1155( .i (n1154), .o (n1155) );
  assign n1156 = ~n724 & n1155 ;
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  assign n1157 = ( n1084 & n1092 ) | ( n1084 & n1100 ) | ( n1092 & n1100 ) ;
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  assign n1165 = ( n1082 & n1114 ) | ( n1082 & n1146 ) | ( n1114 & n1146 ) ;
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n1167 = ( n1122 & n1130 ) | ( n1122 & n1139 ) | ( n1130 & n1139 ) ;
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  assign n1175 = ( n1164 & n1166 ) | ( n1164 & n1174 ) | ( n1166 & n1174 ) ;
  assign n1176 = n1034 & n1077 ;
  assign n1177 = n1034 | n1077 ;
  assign n1178 = ~n1176 & n1177 ;
  buffer buf_n1179( .i (n1178), .o (n1179) );
  assign n1180 = n1039 & n1179 ;
  assign n1181 = n1039 | n1179 ;
  assign n1182 = ~n1180 & n1181 ;
  assign n1183 = n1158 & n1168 ;
  assign n1184 = n1158 | n1168 ;
  assign n1185 = ~n1183 & n1184 ;
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  assign n1190 = n1166 & n1189 ;
  assign n1191 = n1166 | n1189 ;
  assign n1192 = ~n1190 & n1191 ;
  assign out_3_ = n989 ;
  assign out_2_ = n996 ;
  assign out_5_ = n1153 ;
  assign out_1_ = n1156 ;
  assign out_0_ = 1'b0 ;
  assign out_7_ = n1175 ;
  assign out_4_ = n1182 ;
  assign out_6_ = n1192 ;
endmodule
