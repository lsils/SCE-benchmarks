module multi(b_4_,a_1_,a_2_,b_1_,b_7_,a_6_,a_4_,b_2_,a_7_,a_5_,b_5_,b_3_,b_6_,b_0_,a_3_,a_0_,s_1_,s_8_,s_3_,s_5_,s_9_,s_2_,s_11_,s_15_,s_4_,s_10_,s_14_,s_7_,s_13_,s_12_,s_6_,s_0_);
    wire jinkela_wire_0;
    wire jinkela_wire_1;
    wire jinkela_wire_2;
    wire jinkela_wire_3;
    wire jinkela_wire_4;
    wire jinkela_wire_5;
    wire jinkela_wire_6;
    wire jinkela_wire_7;
    wire jinkela_wire_8;
    wire jinkela_wire_9;
    wire jinkela_wire_10;
    wire jinkela_wire_11;
    wire jinkela_wire_12;
    wire jinkela_wire_13;
    wire jinkela_wire_14;
    wire jinkela_wire_15;
    wire jinkela_wire_16;
    wire jinkela_wire_17;
    wire jinkela_wire_18;
    wire jinkela_wire_19;
    wire jinkela_wire_20;
    wire jinkela_wire_21;
    wire jinkela_wire_22;
    wire jinkela_wire_23;
    wire jinkela_wire_24;
    wire jinkela_wire_25;
    wire jinkela_wire_26;
    wire jinkela_wire_27;
    wire jinkela_wire_28;
    wire jinkela_wire_29;
    wire jinkela_wire_30;
    wire jinkela_wire_31;
    wire jinkela_wire_32;
    wire jinkela_wire_33;
    wire jinkela_wire_34;
    wire jinkela_wire_35;
    wire jinkela_wire_36;
    wire jinkela_wire_37;
    wire jinkela_wire_38;
    wire jinkela_wire_39;
    wire jinkela_wire_40;
    wire jinkela_wire_41;
    wire jinkela_wire_42;
    wire jinkela_wire_43;
    wire jinkela_wire_44;
    wire jinkela_wire_45;
    wire jinkela_wire_46;
    wire jinkela_wire_47;
    wire jinkela_wire_48;
    wire jinkela_wire_49;
    wire jinkela_wire_50;
    wire jinkela_wire_51;
    wire jinkela_wire_52;
    wire jinkela_wire_53;
    wire jinkela_wire_54;
    wire jinkela_wire_55;
    wire jinkela_wire_56;
    wire jinkela_wire_57;
    wire jinkela_wire_58;
    wire jinkela_wire_59;
    wire jinkela_wire_60;
    wire jinkela_wire_61;
    wire jinkela_wire_62;
    wire jinkela_wire_63;
    wire jinkela_wire_64;
    wire jinkela_wire_65;
    wire jinkela_wire_66;
    wire jinkela_wire_67;
    wire jinkela_wire_68;
    wire jinkela_wire_69;
    wire jinkela_wire_70;
    wire jinkela_wire_71;
    wire jinkela_wire_72;
    wire jinkela_wire_73;
    wire jinkela_wire_74;
    wire jinkela_wire_75;
    wire jinkela_wire_76;
    wire jinkela_wire_77;
    wire jinkela_wire_78;
    wire jinkela_wire_79;
    wire jinkela_wire_80;
    wire jinkela_wire_81;
    wire jinkela_wire_82;
    wire jinkela_wire_83;
    wire jinkela_wire_84;
    wire jinkela_wire_85;
    wire jinkela_wire_86;
    wire jinkela_wire_87;
    wire jinkela_wire_88;
    wire jinkela_wire_89;
    wire jinkela_wire_90;
    wire jinkela_wire_91;
    wire jinkela_wire_92;
    wire jinkela_wire_93;
    wire jinkela_wire_94;
    wire jinkela_wire_95;
    wire jinkela_wire_96;
    wire jinkela_wire_97;
    wire jinkela_wire_98;
    wire jinkela_wire_99;
    wire jinkela_wire_100;
    wire jinkela_wire_101;
    wire jinkela_wire_102;
    wire jinkela_wire_103;
    wire jinkela_wire_104;
    wire jinkela_wire_105;
    wire jinkela_wire_106;
    wire jinkela_wire_107;
    wire jinkela_wire_108;
    wire jinkela_wire_109;
    wire jinkela_wire_110;
    wire jinkela_wire_111;
    wire jinkela_wire_112;
    wire jinkela_wire_113;
    wire jinkela_wire_114;
    wire jinkela_wire_115;
    wire jinkela_wire_116;
    wire jinkela_wire_117;
    wire jinkela_wire_118;
    wire jinkela_wire_119;
    wire jinkela_wire_120;
    wire jinkela_wire_121;
    wire jinkela_wire_122;
    wire jinkela_wire_123;
    wire jinkela_wire_124;
    wire jinkela_wire_125;
    wire jinkela_wire_126;
    wire jinkela_wire_127;
    wire jinkela_wire_128;
    wire jinkela_wire_129;
    wire jinkela_wire_130;
    wire jinkela_wire_131;
    wire jinkela_wire_132;
    wire jinkela_wire_133;
    wire jinkela_wire_134;
    wire jinkela_wire_135;
    wire jinkela_wire_136;
    wire jinkela_wire_137;
    wire jinkela_wire_138;
    wire jinkela_wire_139;
    wire jinkela_wire_140;
    wire jinkela_wire_141;
    wire jinkela_wire_142;
    wire jinkela_wire_143;
    wire jinkela_wire_144;
    wire jinkela_wire_145;
    wire jinkela_wire_146;
    wire jinkela_wire_147;
    wire jinkela_wire_148;
    wire jinkela_wire_149;
    wire jinkela_wire_150;
    wire jinkela_wire_151;
    wire jinkela_wire_152;
    wire jinkela_wire_153;
    wire jinkela_wire_154;
    wire jinkela_wire_155;
    wire jinkela_wire_156;
    wire jinkela_wire_157;
    wire jinkela_wire_158;
    wire jinkela_wire_159;
    wire jinkela_wire_160;
    wire jinkela_wire_161;
    wire jinkela_wire_162;
    wire jinkela_wire_163;
    wire jinkela_wire_164;
    wire jinkela_wire_165;
    wire jinkela_wire_166;
    wire jinkela_wire_167;
    wire jinkela_wire_168;
    wire jinkela_wire_169;
    wire jinkela_wire_170;
    wire jinkela_wire_171;
    wire jinkela_wire_172;
    wire jinkela_wire_173;
    wire jinkela_wire_174;
    wire jinkela_wire_175;
    wire jinkela_wire_176;
    wire jinkela_wire_177;
    wire jinkela_wire_178;
    wire jinkela_wire_179;
    wire jinkela_wire_180;
    wire jinkela_wire_181;
    wire jinkela_wire_182;
    wire jinkela_wire_183;
    wire jinkela_wire_184;
    wire jinkela_wire_185;
    wire jinkela_wire_186;
    wire jinkela_wire_187;
    wire jinkela_wire_188;
    wire jinkela_wire_189;
    wire jinkela_wire_190;
    wire jinkela_wire_191;
    wire jinkela_wire_192;
    wire jinkela_wire_193;
    wire jinkela_wire_194;
    wire jinkela_wire_195;
    wire jinkela_wire_196;
    wire jinkela_wire_197;
    wire jinkela_wire_198;
    wire jinkela_wire_199;
    wire jinkela_wire_200;
    wire jinkela_wire_201;
    wire jinkela_wire_202;
    wire jinkela_wire_203;
    wire jinkela_wire_204;
    wire jinkela_wire_205;
    wire jinkela_wire_206;
    wire jinkela_wire_207;
    wire jinkela_wire_208;
    wire jinkela_wire_209;
    wire jinkela_wire_210;
    wire jinkela_wire_211;
    wire jinkela_wire_212;
    wire jinkela_wire_213;
    wire jinkela_wire_214;
    wire jinkela_wire_215;
    wire jinkela_wire_216;
    wire jinkela_wire_217;
    wire jinkela_wire_218;
    wire jinkela_wire_219;
    wire jinkela_wire_220;
    wire jinkela_wire_221;
    wire jinkela_wire_222;
    wire jinkela_wire_223;
    wire jinkela_wire_224;
    wire jinkela_wire_225;
    wire jinkela_wire_226;
    wire jinkela_wire_227;
    wire jinkela_wire_228;
    wire jinkela_wire_229;
    wire jinkela_wire_230;
    wire jinkela_wire_231;
    wire jinkela_wire_232;
    wire jinkela_wire_233;
    wire jinkela_wire_234;
    wire jinkela_wire_235;
    wire jinkela_wire_236;
    wire jinkela_wire_237;
    wire jinkela_wire_238;
    wire jinkela_wire_239;
    wire jinkela_wire_240;
    wire jinkela_wire_241;
    wire jinkela_wire_242;
    wire jinkela_wire_243;
    wire jinkela_wire_244;
    wire jinkela_wire_245;
    wire jinkela_wire_246;
    wire jinkela_wire_247;
    wire jinkela_wire_248;
    wire jinkela_wire_249;
    wire jinkela_wire_250;
    wire jinkela_wire_251;
    wire jinkela_wire_252;
    wire jinkela_wire_253;
    wire jinkela_wire_254;
    wire jinkela_wire_255;
    wire jinkela_wire_256;
    wire jinkela_wire_257;
    wire jinkela_wire_258;
    wire jinkela_wire_259;
    wire jinkela_wire_260;
    wire jinkela_wire_261;
    wire jinkela_wire_262;
    wire jinkela_wire_263;
    wire jinkela_wire_264;
    wire jinkela_wire_265;
    wire jinkela_wire_266;
    wire jinkela_wire_267;
    wire jinkela_wire_268;
    wire jinkela_wire_269;
    wire jinkela_wire_270;
    wire jinkela_wire_271;
    wire jinkela_wire_272;
    wire jinkela_wire_273;
    wire jinkela_wire_274;
    wire jinkela_wire_275;
    wire jinkela_wire_276;
    wire jinkela_wire_277;
    wire jinkela_wire_278;
    wire jinkela_wire_279;
    wire jinkela_wire_280;
    wire jinkela_wire_281;
    wire jinkela_wire_282;
    wire jinkela_wire_283;
    wire jinkela_wire_284;
    wire jinkela_wire_285;
    wire jinkela_wire_286;
    wire jinkela_wire_287;
    wire jinkela_wire_288;
    wire jinkela_wire_289;
    wire jinkela_wire_290;
    wire jinkela_wire_291;
    wire jinkela_wire_292;
    wire jinkela_wire_293;
    wire jinkela_wire_294;
    wire jinkela_wire_295;
    wire jinkela_wire_296;
    wire jinkela_wire_297;
    wire jinkela_wire_298;
    wire jinkela_wire_299;
    wire jinkela_wire_300;
    wire jinkela_wire_301;
    wire jinkela_wire_302;
    wire jinkela_wire_303;
    wire jinkela_wire_304;
    wire jinkela_wire_305;
    wire jinkela_wire_306;
    wire jinkela_wire_307;
    wire jinkela_wire_308;
    wire jinkela_wire_309;
    wire jinkela_wire_310;
    wire jinkela_wire_311;
    wire jinkela_wire_312;
    wire jinkela_wire_313;
    wire jinkela_wire_314;
    wire jinkela_wire_315;
    wire jinkela_wire_316;
    wire jinkela_wire_317;
    wire jinkela_wire_318;
    wire jinkela_wire_319;
    wire jinkela_wire_320;
    wire jinkela_wire_321;
    wire jinkela_wire_322;
    wire jinkela_wire_323;
    wire jinkela_wire_324;
    wire jinkela_wire_325;
    wire jinkela_wire_326;
    wire jinkela_wire_327;
    wire jinkela_wire_328;
    wire jinkela_wire_329;
    wire jinkela_wire_330;
    wire jinkela_wire_331;
    wire jinkela_wire_332;
    wire jinkela_wire_333;
    wire jinkela_wire_334;
    wire jinkela_wire_335;
    wire jinkela_wire_336;
    wire jinkela_wire_337;
    wire jinkela_wire_338;
    wire jinkela_wire_339;
    wire jinkela_wire_340;
    wire jinkela_wire_341;
    wire jinkela_wire_342;
    wire jinkela_wire_343;
    wire jinkela_wire_344;
    wire jinkela_wire_345;
    wire jinkela_wire_346;
    wire jinkela_wire_347;
    wire jinkela_wire_348;
    wire jinkela_wire_349;
    wire jinkela_wire_350;
    wire jinkela_wire_351;
    wire jinkela_wire_352;
    wire jinkela_wire_353;
    wire jinkela_wire_354;
    wire jinkela_wire_355;
    wire jinkela_wire_356;
    wire jinkela_wire_357;
    wire jinkela_wire_358;
    wire jinkela_wire_359;
    wire jinkela_wire_360;
    wire jinkela_wire_361;
    wire jinkela_wire_362;
    wire jinkela_wire_363;
    wire jinkela_wire_364;
    wire jinkela_wire_365;
    wire jinkela_wire_366;
    wire jinkela_wire_367;
    wire jinkela_wire_368;
    wire jinkela_wire_369;
    wire jinkela_wire_370;
    wire jinkela_wire_371;
    wire jinkela_wire_372;
    wire jinkela_wire_373;
    wire jinkela_wire_374;
    wire jinkela_wire_375;
    wire jinkela_wire_376;
    wire jinkela_wire_377;
    wire jinkela_wire_378;
    wire jinkela_wire_379;
    wire jinkela_wire_380;
    wire jinkela_wire_381;
    wire jinkela_wire_382;
    wire jinkela_wire_383;
    wire jinkela_wire_384;
    wire jinkela_wire_385;
    wire jinkela_wire_386;
    wire jinkela_wire_387;
    wire jinkela_wire_388;
    wire jinkela_wire_389;
    wire jinkela_wire_390;
    wire jinkela_wire_391;
    wire jinkela_wire_392;
    wire jinkela_wire_393;
    wire jinkela_wire_394;
    wire jinkela_wire_395;
    wire jinkela_wire_396;
    wire jinkela_wire_397;
    wire jinkela_wire_398;
    wire jinkela_wire_399;
    wire jinkela_wire_400;
    wire jinkela_wire_401;
    wire jinkela_wire_402;
    wire jinkela_wire_403;
    wire jinkela_wire_404;
    wire jinkela_wire_405;
    wire jinkela_wire_406;
    wire jinkela_wire_407;
    wire jinkela_wire_408;
    wire jinkela_wire_409;
    wire jinkela_wire_410;
    wire jinkela_wire_411;
    wire jinkela_wire_412;
    wire jinkela_wire_413;
    wire jinkela_wire_414;
    wire jinkela_wire_415;
    wire jinkela_wire_416;
    wire jinkela_wire_417;
    wire jinkela_wire_418;
    wire jinkela_wire_419;
    wire jinkela_wire_420;
    wire jinkela_wire_421;
    wire jinkela_wire_422;
    input b_4_;
    input a_1_;
    input a_2_;
    input b_1_;
    input b_7_;
    input a_6_;
    input a_4_;
    input b_2_;
    input a_7_;
    input a_5_;
    input b_5_;
    input b_3_;
    input b_6_;
    input b_0_;
    input a_3_;
    input a_0_;
    output s_1_;
    output s_8_;
    output s_3_;
    output s_5_;
    output s_9_;
    output s_2_;
    output s_11_;
    output s_15_;
    output s_4_;
    output s_10_;
    output s_14_;
    output s_7_;
    output s_13_;
    output s_12_;
    output s_6_;
    output s_0_;

    and_bb n_642_ (
        .a(jinkela_wire_189),
        .b(jinkela_wire_304),
        .c(jinkela_wire_312)
    );

    or_bb n_643_ (
        .a(jinkela_wire_312),
        .b(jinkela_wire_361),
        .c(jinkela_wire_11)
    );

    and_ii n_644_ (
        .a(jinkela_wire_11),
        .b(jinkela_wire_359),
        .c(jinkela_wire_179)
    );

    and_bb n_645_ (
        .a(jinkela_wire_11),
        .b(jinkela_wire_359),
        .c(jinkela_wire_52)
    );

    and_ii n_646_ (
        .a(jinkela_wire_52),
        .b(jinkela_wire_179),
        .c(s_8_)
    );

    or_bb n_647_ (
        .a(jinkela_wire_179),
        .b(jinkela_wire_361),
        .c(jinkela_wire_93)
    );

    and_ii n_648_ (
        .a(jinkela_wire_320),
        .b(jinkela_wire_318),
        .c(jinkela_wire_354)
    );

    and_ii n_649_ (
        .a(jinkela_wire_12),
        .b(jinkela_wire_215),
        .c(jinkela_wire_177)
    );

    and_ii n_650_ (
        .a(jinkela_wire_396),
        .b(jinkela_wire_213),
        .c(jinkela_wire_89)
    );

    and_ii n_651_ (
        .a(jinkela_wire_137),
        .b(jinkela_wire_176),
        .c(jinkela_wire_329)
    );

    or_bi n_652_ (
        .a(jinkela_wire_324),
        .b(jinkela_wire_172),
        .c(jinkela_wire_203)
    );

    or_ii n_653_ (
        .a(b_5_),
        .b(a_4_),
        .c(jinkela_wire_199)
    );

    or_ii n_654_ (
        .a(b_4_),
        .b(a_6_),
        .c(jinkela_wire_246)
    );

    and_bi n_655_ (
        .a(jinkela_wire_28),
        .b(jinkela_wire_246),
        .c(jinkela_wire_30)
    );

    or_ii n_656_ (
        .a(b_4_),
        .b(a_5_),
        .c(jinkela_wire_217)
    );

    and_bb n_657_ (
        .a(b_3_),
        .b(a_6_),
        .c(jinkela_wire_229)
    );

    and_bi n_658_ (
        .a(jinkela_wire_217),
        .b(jinkela_wire_229),
        .c(jinkela_wire_134)
    );

    or_bb n_659_ (
        .a(jinkela_wire_134),
        .b(jinkela_wire_30),
        .c(jinkela_wire_70)
    );

    and_ii n_660_ (
        .a(jinkela_wire_70),
        .b(jinkela_wire_199),
        .c(jinkela_wire_44)
    );

    and_bb n_661_ (
        .a(jinkela_wire_70),
        .b(jinkela_wire_199),
        .c(jinkela_wire_2)
    );

    or_bb n_662_ (
        .a(jinkela_wire_2),
        .b(jinkela_wire_44),
        .c(jinkela_wire_40)
    );

    and_ii n_663_ (
        .a(jinkela_wire_40),
        .b(jinkela_wire_203),
        .c(jinkela_wire_88)
    );

    and_bb n_664_ (
        .a(jinkela_wire_40),
        .b(jinkela_wire_203),
        .c(jinkela_wire_337)
    );

    or_bb n_665_ (
        .a(jinkela_wire_337),
        .b(jinkela_wire_88),
        .c(jinkela_wire_285)
    );

    and_ii n_666_ (
        .a(jinkela_wire_285),
        .b(jinkela_wire_329),
        .c(jinkela_wire_57)
    );

    and_bb n_667_ (
        .a(jinkela_wire_285),
        .b(jinkela_wire_329),
        .c(jinkela_wire_269)
    );

    or_bb n_668_ (
        .a(jinkela_wire_269),
        .b(jinkela_wire_57),
        .c(jinkela_wire_6)
    );

    or_ii n_669_ (
        .a(b_7_),
        .b(a_2_),
        .c(jinkela_wire_22)
    );

    and_ii n_670_ (
        .a(jinkela_wire_287),
        .b(jinkela_wire_240),
        .c(jinkela_wire_349)
    );

    or_ii n_671_ (
        .a(b_6_),
        .b(a_3_),
        .c(jinkela_wire_98)
    );

    and_ii n_672_ (
        .a(jinkela_wire_98),
        .b(jinkela_wire_349),
        .c(jinkela_wire_322)
    );

    and_bb n_673_ (
        .a(jinkela_wire_98),
        .b(jinkela_wire_349),
        .c(jinkela_wire_3)
    );

    or_bb n_674_ (
        .a(jinkela_wire_3),
        .b(jinkela_wire_322),
        .c(jinkela_wire_270)
    );

    and_ii n_675_ (
        .a(jinkela_wire_270),
        .b(jinkela_wire_22),
        .c(jinkela_wire_141)
    );

    and_bb n_676_ (
        .a(jinkela_wire_270),
        .b(jinkela_wire_22),
        .c(jinkela_wire_384)
    );

    or_bb n_677_ (
        .a(jinkela_wire_384),
        .b(jinkela_wire_141),
        .c(jinkela_wire_306)
    );

    and_ii n_678_ (
        .a(jinkela_wire_306),
        .b(jinkela_wire_6),
        .c(jinkela_wire_149)
    );

    and_bb n_679_ (
        .a(jinkela_wire_306),
        .b(jinkela_wire_6),
        .c(jinkela_wire_119)
    );

    or_bb n_680_ (
        .a(jinkela_wire_119),
        .b(jinkela_wire_149),
        .c(jinkela_wire_123)
    );

    and_ii n_681_ (
        .a(jinkela_wire_123),
        .b(jinkela_wire_89),
        .c(jinkela_wire_310)
    );

    and_bb n_682_ (
        .a(jinkela_wire_123),
        .b(jinkela_wire_89),
        .c(jinkela_wire_295)
    );

    or_bb n_683_ (
        .a(jinkela_wire_295),
        .b(jinkela_wire_310),
        .c(jinkela_wire_316)
    );

    and_bi n_471_ (
        .a(jinkela_wire_347),
        .b(jinkela_wire_79),
        .c(jinkela_wire_125)
    );

    and_ii n_513_ (
        .a(jinkela_wire_303),
        .b(jinkela_wire_165),
        .c(jinkela_wire_58)
    );

    or_ii n_555_ (
        .a(b_4_),
        .b(a_3_),
        .c(jinkela_wire_390)
    );

    and_ii n_600_ (
        .a(jinkela_wire_324),
        .b(jinkela_wire_172),
        .c(jinkela_wire_358)
    );

    or_bb n_472_ (
        .a(jinkela_wire_125),
        .b(jinkela_wire_32),
        .c(jinkela_wire_162)
    );

    and_bb n_514_ (
        .a(jinkela_wire_303),
        .b(jinkela_wire_165),
        .c(jinkela_wire_185)
    );

    and_bb n_556_ (
        .a(b_3_),
        .b(a_4_),
        .c(jinkela_wire_202)
    );

    or_ii n_601_ (
        .a(a_7_),
        .b(b_1_),
        .c(jinkela_wire_220)
    );

    and_ii n_473_ (
        .a(jinkela_wire_162),
        .b(jinkela_wire_18),
        .c(jinkela_wire_144)
    );

    or_bb n_515_ (
        .a(jinkela_wire_185),
        .b(jinkela_wire_58),
        .c(jinkela_wire_170)
    );

    and_bi n_557_ (
        .a(jinkela_wire_202),
        .b(jinkela_wire_390),
        .c(jinkela_wire_133)
    );

    and_bb n_602_ (
        .a(b_2_),
        .b(a_6_),
        .c(jinkela_wire_387)
    );

    and_bb n_474_ (
        .a(jinkela_wire_162),
        .b(jinkela_wire_18),
        .c(jinkela_wire_20)
    );

    and_ii n_516_ (
        .a(jinkela_wire_170),
        .b(jinkela_wire_255),
        .c(jinkela_wire_108)
    );

    and_bi n_558_ (
        .a(jinkela_wire_390),
        .b(jinkela_wire_202),
        .c(jinkela_wire_339)
    );

    and_bi n_603_ (
        .a(jinkela_wire_220),
        .b(jinkela_wire_387),
        .c(jinkela_wire_230)
    );

    or_bb n_475_ (
        .a(jinkela_wire_20),
        .b(jinkela_wire_144),
        .c(jinkela_wire_373)
    );

    and_bb n_517_ (
        .a(jinkela_wire_170),
        .b(jinkela_wire_255),
        .c(jinkela_wire_0)
    );

    or_bb n_559_ (
        .a(jinkela_wire_339),
        .b(jinkela_wire_133),
        .c(jinkela_wire_116)
    );

    or_bb n_604_ (
        .a(jinkela_wire_230),
        .b(jinkela_wire_358),
        .c(jinkela_wire_120)
    );

    and_ii n_476_ (
        .a(jinkela_wire_373),
        .b(jinkela_wire_186),
        .c(jinkela_wire_74)
    );

    or_bb n_518_ (
        .a(jinkela_wire_0),
        .b(jinkela_wire_108),
        .c(jinkela_wire_1)
    );

    and_ii n_560_ (
        .a(jinkela_wire_116),
        .b(jinkela_wire_302),
        .c(jinkela_wire_68)
    );

    and_ii n_605_ (
        .a(jinkela_wire_120),
        .b(jinkela_wire_419),
        .c(jinkela_wire_176)
    );

    and_bb n_477_ (
        .a(jinkela_wire_373),
        .b(jinkela_wire_186),
        .c(jinkela_wire_145)
    );

    or_bb n_519_ (
        .a(jinkela_wire_1),
        .b(jinkela_wire_397),
        .c(jinkela_wire_341)
    );

    and_bb n_561_ (
        .a(jinkela_wire_116),
        .b(jinkela_wire_302),
        .c(jinkela_wire_364)
    );

    and_bb n_606_ (
        .a(jinkela_wire_120),
        .b(jinkela_wire_419),
        .c(jinkela_wire_226)
    );

    or_bb n_478_ (
        .a(jinkela_wire_145),
        .b(jinkela_wire_74),
        .c(jinkela_wire_236)
    );

    or_ii n_520_ (
        .a(jinkela_wire_1),
        .b(jinkela_wire_397),
        .c(jinkela_wire_327)
    );

    or_bb n_562_ (
        .a(jinkela_wire_364),
        .b(jinkela_wire_68),
        .c(jinkela_wire_279)
    );

    or_bb n_607_ (
        .a(jinkela_wire_226),
        .b(jinkela_wire_176),
        .c(jinkela_wire_112)
    );

    or_bb n_479_ (
        .a(jinkela_wire_236),
        .b(jinkela_wire_184),
        .c(jinkela_wire_200)
    );

    or_ii n_521_ (
        .a(jinkela_wire_327),
        .b(jinkela_wire_341),
        .c(jinkela_wire_100)
    );

    and_ii n_563_ (
        .a(jinkela_wire_279),
        .b(jinkela_wire_51),
        .c(jinkela_wire_150)
    );

    or_ii n_608_ (
        .a(b_5_),
        .b(a_3_),
        .c(jinkela_wire_401)
    );

    or_ii n_480_ (
        .a(jinkela_wire_236),
        .b(jinkela_wire_184),
        .c(jinkela_wire_8)
    );

    and_ii n_522_ (
        .a(jinkela_wire_144),
        .b(jinkela_wire_32),
        .c(jinkela_wire_153)
    );

    and_bb n_564_ (
        .a(jinkela_wire_279),
        .b(jinkela_wire_51),
        .c(jinkela_wire_294)
    );

    or_ii n_609_ (
        .a(b_4_),
        .b(a_4_),
        .c(jinkela_wire_418)
    );

    or_ii n_481_ (
        .a(jinkela_wire_8),
        .b(jinkela_wire_200),
        .c(jinkela_wire_164)
    );

    or_ii n_523_ (
        .a(b_6_),
        .b(a_0_),
        .c(jinkela_wire_323)
    );

    or_bb n_565_ (
        .a(jinkela_wire_294),
        .b(jinkela_wire_150),
        .c(jinkela_wire_406)
    );

    and_bb n_610_ (
        .a(b_3_),
        .b(a_5_),
        .c(jinkela_wire_28)
    );

    and_ii n_482_ (
        .a(jinkela_wire_164),
        .b(jinkela_wire_283),
        .c(jinkela_wire_410)
    );

    or_bb n_524_ (
        .a(jinkela_wire_323),
        .b(jinkela_wire_153),
        .c(jinkela_wire_377)
    );

    or_bb n_566_ (
        .a(jinkela_wire_406),
        .b(jinkela_wire_281),
        .c(jinkela_wire_175)
    );

    and_bi n_611_ (
        .a(jinkela_wire_28),
        .b(jinkela_wire_418),
        .c(jinkela_wire_240)
    );

    and_bb n_483_ (
        .a(jinkela_wire_164),
        .b(jinkela_wire_283),
        .c(jinkela_wire_227)
    );

    and_bb n_525_ (
        .a(jinkela_wire_323),
        .b(jinkela_wire_153),
        .c(jinkela_wire_128)
    );

    or_ii n_567_ (
        .a(jinkela_wire_406),
        .b(jinkela_wire_281),
        .c(jinkela_wire_371)
    );

    and_bi n_612_ (
        .a(jinkela_wire_418),
        .b(jinkela_wire_28),
        .c(jinkela_wire_205)
    );

    or_bb n_484_ (
        .a(jinkela_wire_227),
        .b(jinkela_wire_410),
        .c(jinkela_wire_300)
    );

    or_bi n_526_ (
        .a(jinkela_wire_128),
        .b(jinkela_wire_377),
        .c(jinkela_wire_336)
    );

    or_ii n_568_ (
        .a(jinkela_wire_371),
        .b(jinkela_wire_175),
        .c(jinkela_wire_208)
    );

    or_bb n_613_ (
        .a(jinkela_wire_205),
        .b(jinkela_wire_240),
        .c(jinkela_wire_297)
    );

    or_bb n_485_ (
        .a(jinkela_wire_300),
        .b(jinkela_wire_4),
        .c(jinkela_wire_81)
    );

    and_ii n_527_ (
        .a(jinkela_wire_336),
        .b(jinkela_wire_100),
        .c(jinkela_wire_370)
    );

    or_ii n_569_ (
        .a(b_7_),
        .b(a_0_),
        .c(jinkela_wire_271)
    );

    and_ii n_614_ (
        .a(jinkela_wire_297),
        .b(jinkela_wire_401),
        .c(jinkela_wire_287)
    );

    and_bb n_486_ (
        .a(jinkela_wire_300),
        .b(jinkela_wire_4),
        .c(jinkela_wire_207)
    );

    and_bb n_528_ (
        .a(jinkela_wire_336),
        .b(jinkela_wire_100),
        .c(jinkela_wire_131)
    );

    and_bi n_570_ (
        .a(jinkela_wire_420),
        .b(jinkela_wire_58),
        .c(jinkela_wire_66)
    );

    and_bb n_615_ (
        .a(jinkela_wire_297),
        .b(jinkela_wire_401),
        .c(jinkela_wire_206)
    );

    or_bi n_487_ (
        .a(jinkela_wire_207),
        .b(jinkela_wire_81),
        .c(jinkela_wire_325)
    );

    or_bb n_529_ (
        .a(jinkela_wire_131),
        .b(jinkela_wire_370),
        .c(jinkela_wire_130)
    );

    or_ii n_571_ (
        .a(b_6_),
        .b(a_1_),
        .c(jinkela_wire_39)
    );

    or_bb n_616_ (
        .a(jinkela_wire_206),
        .b(jinkela_wire_287),
        .c(jinkela_wire_63)
    );

    or_bb n_488_ (
        .a(jinkela_wire_325),
        .b(jinkela_wire_19),
        .c(jinkela_wire_369)
    );

    or_bb n_530_ (
        .a(jinkela_wire_130),
        .b(jinkela_wire_221),
        .c(jinkela_wire_235)
    );

    and_ii n_572_ (
        .a(jinkela_wire_39),
        .b(jinkela_wire_66),
        .c(jinkela_wire_385)
    );

    and_ii n_617_ (
        .a(jinkela_wire_63),
        .b(jinkela_wire_112),
        .c(jinkela_wire_137)
    );

    and_bb n_489_ (
        .a(jinkela_wire_325),
        .b(jinkela_wire_19),
        .c(jinkela_wire_60)
    );

    and_bb n_531_ (
        .a(jinkela_wire_130),
        .b(jinkela_wire_221),
        .c(jinkela_wire_14)
    );

    and_bb n_573_ (
        .a(jinkela_wire_39),
        .b(jinkela_wire_66),
        .c(jinkela_wire_127)
    );

    and_bb n_618_ (
        .a(jinkela_wire_63),
        .b(jinkela_wire_112),
        .c(jinkela_wire_99)
    );

    and_bi n_490_ (
        .a(jinkela_wire_369),
        .b(jinkela_wire_60),
        .c(s_5_)
    );

    or_bi n_532_ (
        .a(jinkela_wire_14),
        .b(jinkela_wire_235),
        .c(jinkela_wire_309)
    );

    or_bb n_577_ (
        .a(jinkela_wire_421),
        .b(jinkela_wire_95),
        .c(jinkela_wire_129)
    );

    or_bb n_619_ (
        .a(jinkela_wire_99),
        .b(jinkela_wire_137),
        .c(jinkela_wire_196)
    );

    and_bi n_491_ (
        .a(jinkela_wire_200),
        .b(jinkela_wire_410),
        .c(jinkela_wire_221)
    );

    or_bb n_533_ (
        .a(jinkela_wire_309),
        .b(jinkela_wire_81),
        .c(jinkela_wire_188)
    );

    and_ii n_578_ (
        .a(jinkela_wire_129),
        .b(jinkela_wire_208),
        .c(jinkela_wire_298)
    );

    and_ii n_620_ (
        .a(jinkela_wire_196),
        .b(jinkela_wire_124),
        .c(jinkela_wire_213)
    );

    and_bi n_492_ (
        .a(jinkela_wire_183),
        .b(jinkela_wire_74),
        .c(jinkela_wire_397)
    );

    or_ii n_534_ (
        .a(jinkela_wire_309),
        .b(jinkela_wire_81),
        .c(jinkela_wire_402)
    );

    and_bb n_579_ (
        .a(jinkela_wire_129),
        .b(jinkela_wire_208),
        .c(jinkela_wire_267)
    );

    and_bb n_621_ (
        .a(jinkela_wire_196),
        .b(jinkela_wire_124),
        .c(jinkela_wire_113)
    );

    and_bi n_493_ (
        .a(jinkela_wire_151),
        .b(jinkela_wire_352),
        .c(jinkela_wire_201)
    );

    or_ii n_535_ (
        .a(jinkela_wire_402),
        .b(jinkela_wire_188),
        .c(jinkela_wire_407)
    );

    or_bb n_580_ (
        .a(jinkela_wire_267),
        .b(jinkela_wire_298),
        .c(jinkela_wire_234)
    );

    or_bb n_622_ (
        .a(jinkela_wire_113),
        .b(jinkela_wire_213),
        .c(jinkela_wire_169)
    );

    or_ii n_494_ (
        .a(b_2_),
        .b(a_4_),
        .c(jinkela_wire_187)
    );

    and_ii n_536_ (
        .a(jinkela_wire_407),
        .b(jinkela_wire_369),
        .c(jinkela_wire_363)
    );

    or_bb n_581_ (
        .a(jinkela_wire_234),
        .b(jinkela_wire_132),
        .c(jinkela_wire_38)
    );

    or_ii n_623_ (
        .a(b_7_),
        .b(a_1_),
        .c(jinkela_wire_249)
    );

    or_ii n_495_ (
        .a(a_6_),
        .b(b_1_),
        .c(jinkela_wire_172)
    );

    and_bb n_537_ (
        .a(jinkela_wire_407),
        .b(jinkela_wire_369),
        .c(jinkela_wire_280)
    );

    or_ii n_582_ (
        .a(jinkela_wire_234),
        .b(jinkela_wire_132),
        .c(jinkela_wire_277)
    );

    and_ii n_624_ (
        .a(jinkela_wire_68),
        .b(jinkela_wire_133),
        .c(jinkela_wire_107)
    );

    or_bb n_496_ (
        .a(jinkela_wire_172),
        .b(jinkela_wire_331),
        .c(jinkela_wire_122)
    );

    and_ii n_538_ (
        .a(jinkela_wire_280),
        .b(jinkela_wire_363),
        .c(s_6_)
    );

    or_ii n_583_ (
        .a(jinkela_wire_277),
        .b(jinkela_wire_38),
        .c(jinkela_wire_408)
    );

    or_ii n_625_ (
        .a(b_6_),
        .b(a_2_),
        .c(jinkela_wire_315)
    );

    or_ii n_497_ (
        .a(a_5_),
        .b(b_1_),
        .c(jinkela_wire_362)
    );

    and_bi n_539_ (
        .a(jinkela_wire_188),
        .b(jinkela_wire_363),
        .c(jinkela_wire_376)
    );

    and_ii n_584_ (
        .a(jinkela_wire_408),
        .b(jinkela_wire_377),
        .c(jinkela_wire_31)
    );

    and_ii n_626_ (
        .a(jinkela_wire_315),
        .b(jinkela_wire_107),
        .c(jinkela_wire_215)
    );

    and_bb n_498_ (
        .a(b_0_),
        .b(a_6_),
        .c(jinkela_wire_282)
    );

    and_bi n_540_ (
        .a(jinkela_wire_341),
        .b(jinkela_wire_370),
        .c(jinkela_wire_132)
    );

    and_bb n_585_ (
        .a(jinkela_wire_408),
        .b(jinkela_wire_377),
        .c(jinkela_wire_97)
    );

    and_bb n_627_ (
        .a(jinkela_wire_315),
        .b(jinkela_wire_107),
        .c(jinkela_wire_102)
    );

    or_bi n_499_ (
        .a(jinkela_wire_282),
        .b(jinkela_wire_362),
        .c(jinkela_wire_192)
    );

    and_bi n_541_ (
        .a(jinkela_wire_368),
        .b(jinkela_wire_108),
        .c(jinkela_wire_281)
    );

    or_bb n_586_ (
        .a(jinkela_wire_97),
        .b(jinkela_wire_31),
        .c(jinkela_wire_244)
    );

    or_bb n_628_ (
        .a(jinkela_wire_102),
        .b(jinkela_wire_215),
        .c(jinkela_wire_152)
    );

    or_ii n_500_ (
        .a(jinkela_wire_192),
        .b(jinkela_wire_122),
        .c(jinkela_wire_374)
    );

    and_bi n_542_ (
        .a(jinkela_wire_122),
        .b(jinkela_wire_25),
        .c(jinkela_wire_109)
    );

    or_bb n_587_ (
        .a(jinkela_wire_244),
        .b(jinkela_wire_235),
        .c(jinkela_wire_48)
    );

    and_ii n_629_ (
        .a(jinkela_wire_152),
        .b(jinkela_wire_249),
        .c(jinkela_wire_12)
    );

    and_ii n_501_ (
        .a(jinkela_wire_374),
        .b(jinkela_wire_187),
        .c(jinkela_wire_25)
    );

    or_ii n_543_ (
        .a(b_2_),
        .b(a_5_),
        .c(jinkela_wire_386)
    );

    or_ii n_588_ (
        .a(jinkela_wire_244),
        .b(jinkela_wire_235),
        .c(jinkela_wire_156)
    );

    and_bb n_630_ (
        .a(jinkela_wire_152),
        .b(jinkela_wire_249),
        .c(jinkela_wire_311)
    );

    and_bb n_502_ (
        .a(jinkela_wire_374),
        .b(jinkela_wire_187),
        .c(jinkela_wire_167)
    );

    or_ii n_544_ (
        .a(b_0_),
        .b(a_7_),
        .c(jinkela_wire_21)
    );

    or_ii n_589_ (
        .a(jinkela_wire_156),
        .b(jinkela_wire_48),
        .c(jinkela_wire_59)
    );

    or_bb n_631_ (
        .a(jinkela_wire_311),
        .b(jinkela_wire_12),
        .c(jinkela_wire_103)
    );

    or_bb n_503_ (
        .a(jinkela_wire_167),
        .b(jinkela_wire_25),
        .c(jinkela_wire_340)
    );

    or_bb n_545_ (
        .a(jinkela_wire_21),
        .b(jinkela_wire_172),
        .c(jinkela_wire_350)
    );

    and_ii n_590_ (
        .a(jinkela_wire_59),
        .b(jinkela_wire_376),
        .c(jinkela_wire_256)
    );

    and_ii n_632_ (
        .a(jinkela_wire_103),
        .b(jinkela_wire_169),
        .c(jinkela_wire_396)
    );

    or_bb n_504_ (
        .a(jinkela_wire_340),
        .b(jinkela_wire_201),
        .c(jinkela_wire_368)
    );

    or_ii n_546_ (
        .a(jinkela_wire_21),
        .b(jinkela_wire_172),
        .c(jinkela_wire_212)
    );

    and_bb n_591_ (
        .a(jinkela_wire_59),
        .b(jinkela_wire_376),
        .c(jinkela_wire_49)
    );

    and_bb n_633_ (
        .a(jinkela_wire_103),
        .b(jinkela_wire_169),
        .c(jinkela_wire_332)
    );

    or_ii n_505_ (
        .a(jinkela_wire_340),
        .b(jinkela_wire_201),
        .c(jinkela_wire_389)
    );

    or_ii n_547_ (
        .a(jinkela_wire_212),
        .b(jinkela_wire_350),
        .c(jinkela_wire_422)
    );

    and_ii n_592_ (
        .a(jinkela_wire_49),
        .b(jinkela_wire_256),
        .c(s_7_)
    );

    or_bb n_634_ (
        .a(jinkela_wire_332),
        .b(jinkela_wire_396),
        .c(jinkela_wire_9)
    );

    or_ii n_506_ (
        .a(jinkela_wire_389),
        .b(jinkela_wire_368),
        .c(jinkela_wire_255)
    );

    and_ii n_548_ (
        .a(jinkela_wire_422),
        .b(jinkela_wire_386),
        .c(jinkela_wire_138)
    );

    and_bi n_593_ (
        .a(jinkela_wire_48),
        .b(jinkela_wire_256),
        .c(jinkela_wire_359)
    );

    and_ii n_635_ (
        .a(jinkela_wire_9),
        .b(jinkela_wire_266),
        .c(jinkela_wire_318)
    );

    or_ii n_507_ (
        .a(b_5_),
        .b(a_1_),
        .c(jinkela_wire_165)
    );

    and_bb n_549_ (
        .a(jinkela_wire_422),
        .b(jinkela_wire_386),
        .c(jinkela_wire_104)
    );

    and_bi n_594_ (
        .a(jinkela_wire_38),
        .b(jinkela_wire_31),
        .c(jinkela_wire_304)
    );

    and_bb n_636_ (
        .a(jinkela_wire_9),
        .b(jinkela_wire_266),
        .c(jinkela_wire_252)
    );

    or_ii n_508_ (
        .a(b_4_),
        .b(a_2_),
        .c(jinkela_wire_348)
    );

    or_bb n_550_ (
        .a(jinkela_wire_104),
        .b(jinkela_wire_138),
        .c(jinkela_wire_342)
    );

    and_ii n_595_ (
        .a(jinkela_wire_95),
        .b(jinkela_wire_385),
        .c(jinkela_wire_344)
    );

    or_bb n_637_ (
        .a(jinkela_wire_252),
        .b(jinkela_wire_318),
        .c(jinkela_wire_284)
    );

    or_ii n_509_ (
        .a(b_3_),
        .b(a_3_),
        .c(jinkela_wire_204)
    );

    or_bb n_551_ (
        .a(jinkela_wire_342),
        .b(jinkela_wire_109),
        .c(jinkela_wire_219)
    );

    and_bi n_596_ (
        .a(jinkela_wire_175),
        .b(jinkela_wire_298),
        .c(jinkela_wire_266)
    );

    and_ii n_638_ (
        .a(jinkela_wire_284),
        .b(jinkela_wire_344),
        .c(jinkela_wire_320)
    );

    or_bb n_510_ (
        .a(jinkela_wire_204),
        .b(jinkela_wire_348),
        .c(jinkela_wire_420)
    );

    or_ii n_552_ (
        .a(jinkela_wire_342),
        .b(jinkela_wire_109),
        .c(jinkela_wire_77)
    );

    and_bi n_597_ (
        .a(jinkela_wire_219),
        .b(jinkela_wire_150),
        .c(jinkela_wire_124)
    );

    and_bb n_639_ (
        .a(jinkela_wire_284),
        .b(jinkela_wire_344),
        .c(jinkela_wire_15)
    );

    or_ii n_553_ (
        .a(jinkela_wire_77),
        .b(jinkela_wire_219),
        .c(jinkela_wire_51)
    );

    and_bi n_598_ (
        .a(jinkela_wire_350),
        .b(jinkela_wire_138),
        .c(jinkela_wire_419)
    );

    or_bb n_640_ (
        .a(jinkela_wire_15),
        .b(jinkela_wire_320),
        .c(jinkela_wire_189)
    );

    or_ii n_511_ (
        .a(jinkela_wire_204),
        .b(jinkela_wire_348),
        .c(jinkela_wire_214)
    );

    or_ii n_512_ (
        .a(jinkela_wire_214),
        .b(jinkela_wire_420),
        .c(jinkela_wire_303)
    );

    or_ii n_554_ (
        .a(b_5_),
        .b(a_2_),
        .c(jinkela_wire_302)
    );

    or_ii n_599_ (
        .a(b_2_),
        .b(a_7_),
        .c(jinkela_wire_324)
    );

    and_ii n_641_ (
        .a(jinkela_wire_189),
        .b(jinkela_wire_304),
        .c(jinkela_wire_361)
    );

    and_ii n_575_ (
        .a(jinkela_wire_292),
        .b(jinkela_wire_271),
        .c(jinkela_wire_95)
    );

    and_bb n_576_ (
        .a(jinkela_wire_292),
        .b(jinkela_wire_271),
        .c(jinkela_wire_421)
    );

    or_bb n_574_ (
        .a(jinkela_wire_127),
        .b(jinkela_wire_385),
        .c(jinkela_wire_292)
    );

    or_ii n_429_ (
        .a(b_0_),
        .b(a_4_),
        .c(jinkela_wire_26)
    );

    or_bb n_430_ (
        .a(jinkela_wire_26),
        .b(jinkela_wire_37),
        .c(jinkela_wire_154)
    );

    or_ii n_431_ (
        .a(jinkela_wire_26),
        .b(jinkela_wire_37),
        .c(jinkela_wire_260)
    );

    or_ii n_432_ (
        .a(jinkela_wire_260),
        .b(jinkela_wire_154),
        .c(jinkela_wire_416)
    );

    and_ii n_433_ (
        .a(jinkela_wire_416),
        .b(jinkela_wire_382),
        .c(jinkela_wire_158)
    );

    and_bb n_434_ (
        .a(jinkela_wire_416),
        .b(jinkela_wire_382),
        .c(jinkela_wire_413)
    );

    or_bb n_435_ (
        .a(jinkela_wire_413),
        .b(jinkela_wire_158),
        .c(jinkela_wire_91)
    );

    or_bb n_436_ (
        .a(jinkela_wire_91),
        .b(jinkela_wire_356),
        .c(jinkela_wire_46)
    );

    or_ii n_437_ (
        .a(jinkela_wire_91),
        .b(jinkela_wire_356),
        .c(jinkela_wire_218)
    );

    or_ii n_438_ (
        .a(jinkela_wire_218),
        .b(jinkela_wire_46),
        .c(jinkela_wire_55)
    );

    or_ii n_439_ (
        .a(b_4_),
        .b(a_1_),
        .c(jinkela_wire_347)
    );

    or_bb n_440_ (
        .a(jinkela_wire_347),
        .b(jinkela_wire_118),
        .c(jinkela_wire_283)
    );

    or_ii n_441_ (
        .a(b_3_),
        .b(a_1_),
        .c(jinkela_wire_143)
    );

    and_bb n_442_ (
        .a(b_4_),
        .b(a_0_),
        .c(jinkela_wire_33)
    );

    and_bi n_443_ (
        .a(jinkela_wire_143),
        .b(jinkela_wire_33),
        .c(jinkela_wire_290)
    );

    or_bi n_444_ (
        .a(jinkela_wire_290),
        .b(jinkela_wire_283),
        .c(jinkela_wire_328)
    );

    and_ii n_445_ (
        .a(jinkela_wire_328),
        .b(jinkela_wire_55),
        .c(jinkela_wire_265)
    );

    and_bb n_446_ (
        .a(jinkela_wire_328),
        .b(jinkela_wire_55),
        .c(jinkela_wire_111)
    );

    or_bb n_447_ (
        .a(jinkela_wire_111),
        .b(jinkela_wire_265),
        .c(jinkela_wire_168)
    );

    or_bb n_448_ (
        .a(jinkela_wire_168),
        .b(jinkela_wire_393),
        .c(jinkela_wire_4)
    );

    and_bb n_449_ (
        .a(jinkela_wire_168),
        .b(jinkela_wire_393),
        .c(jinkela_wire_135)
    );

    or_bi n_450_ (
        .a(jinkela_wire_135),
        .b(jinkela_wire_4),
        .c(jinkela_wire_159)
    );

    or_bb n_451_ (
        .a(jinkela_wire_159),
        .b(jinkela_wire_273),
        .c(jinkela_wire_19)
    );

    and_bb n_452_ (
        .a(jinkela_wire_159),
        .b(jinkela_wire_273),
        .c(jinkela_wire_209)
    );

    and_bi n_453_ (
        .a(jinkela_wire_19),
        .b(jinkela_wire_209),
        .c(s_4_)
    );

    and_bi n_454_ (
        .a(jinkela_wire_46),
        .b(jinkela_wire_265),
        .c(jinkela_wire_184)
    );

    and_bi n_455_ (
        .a(jinkela_wire_154),
        .b(jinkela_wire_158),
        .c(jinkela_wire_248)
    );

    or_ii n_456_ (
        .a(b_2_),
        .b(a_3_),
        .c(jinkela_wire_259)
    );

    or_ii n_457_ (
        .a(a_4_),
        .b(b_1_),
        .c(jinkela_wire_245)
    );

    or_ii n_458_ (
        .a(b_0_),
        .b(a_5_),
        .c(jinkela_wire_331)
    );

    or_bb n_459_ (
        .a(jinkela_wire_331),
        .b(jinkela_wire_245),
        .c(jinkela_wire_151)
    );

    or_ii n_460_ (
        .a(jinkela_wire_331),
        .b(jinkela_wire_245),
        .c(jinkela_wire_378)
    );

    or_ii n_461_ (
        .a(jinkela_wire_378),
        .b(jinkela_wire_151),
        .c(jinkela_wire_173)
    );

    and_ii n_462_ (
        .a(jinkela_wire_173),
        .b(jinkela_wire_259),
        .c(jinkela_wire_352)
    );

    and_bb n_463_ (
        .a(jinkela_wire_173),
        .b(jinkela_wire_259),
        .c(jinkela_wire_69)
    );

    or_bb n_464_ (
        .a(jinkela_wire_69),
        .b(jinkela_wire_352),
        .c(jinkela_wire_101)
    );

    or_bb n_465_ (
        .a(jinkela_wire_101),
        .b(jinkela_wire_248),
        .c(jinkela_wire_183)
    );

    or_ii n_466_ (
        .a(jinkela_wire_101),
        .b(jinkela_wire_248),
        .c(jinkela_wire_314)
    );

    or_ii n_467_ (
        .a(jinkela_wire_314),
        .b(jinkela_wire_183),
        .c(jinkela_wire_186)
    );

    or_ii n_468_ (
        .a(b_5_),
        .b(a_0_),
        .c(jinkela_wire_18)
    );

    and_bb n_469_ (
        .a(b_3_),
        .b(a_2_),
        .c(jinkela_wire_79)
    );

    and_bi n_470_ (
        .a(jinkela_wire_79),
        .b(jinkela_wire_347),
        .c(jinkela_wire_32)
    );

    and_bi n_426_ (
        .a(jinkela_wire_405),
        .b(jinkela_wire_210),
        .c(jinkela_wire_356)
    );

    and_bi n_424_ (
        .a(jinkela_wire_273),
        .b(jinkela_wire_85),
        .c(s_3_)
    );

    and_ii n_425_ (
        .a(jinkela_wire_379),
        .b(jinkela_wire_225),
        .c(jinkela_wire_393)
    );

    and_bb n_423_ (
        .a(jinkela_wire_190),
        .b(jinkela_wire_73),
        .c(jinkela_wire_85)
    );

    or_ii n_427_ (
        .a(b_2_),
        .b(a_2_),
        .c(jinkela_wire_382)
    );

    or_ii n_428_ (
        .a(a_3_),
        .b(b_1_),
        .c(jinkela_wire_37)
    );

    and_ii n_768_ (
        .a(jinkela_wire_142),
        .b(jinkela_wire_296),
        .c(jinkela_wire_139)
    );

    and_bb n_810_ (
        .a(jinkela_wire_35),
        .b(jinkela_wire_383),
        .c(jinkela_wire_372)
    );

    and_ii n_852_ (
        .a(jinkela_wire_262),
        .b(jinkela_wire_136),
        .c(jinkela_wire_210)
    );

    and_ii n_769_ (
        .a(jinkela_wire_84),
        .b(jinkela_wire_317),
        .c(jinkela_wire_360)
    );

    or_bb n_811_ (
        .a(jinkela_wire_372),
        .b(jinkela_wire_275),
        .c(jinkela_wire_92)
    );

    and_bb n_853_ (
        .a(jinkela_wire_262),
        .b(jinkela_wire_136),
        .c(jinkela_wire_308)
    );

    and_ii n_770_ (
        .a(jinkela_wire_333),
        .b(jinkela_wire_67),
        .c(jinkela_wire_193)
    );

    and_ii n_812_ (
        .a(jinkela_wire_92),
        .b(jinkela_wire_71),
        .c(jinkela_wire_56)
    );

    or_bb n_854_ (
        .a(jinkela_wire_308),
        .b(jinkela_wire_210),
        .c(jinkela_wire_411)
    );

    or_ii n_771_ (
        .a(b_7_),
        .b(a_5_),
        .c(jinkela_wire_78)
    );

    and_bb n_813_ (
        .a(jinkela_wire_92),
        .b(jinkela_wire_71),
        .c(jinkela_wire_355)
    );

    and_ii n_855_ (
        .a(jinkela_wire_411),
        .b(jinkela_wire_166),
        .c(jinkela_wire_225)
    );

    and_bi n_772_ (
        .a(b_6_),
        .b(jinkela_wire_121),
        .c(jinkela_wire_163)
    );

    and_ii n_814_ (
        .a(jinkela_wire_355),
        .b(jinkela_wire_56),
        .c(s_13_)
    );

    and_bb n_856_ (
        .a(jinkela_wire_411),
        .b(jinkela_wire_166),
        .c(jinkela_wire_86)
    );

    and_bb n_773_ (
        .a(b_6_),
        .b(a_6_),
        .c(jinkela_wire_353)
    );

    and_ii n_815_ (
        .a(jinkela_wire_56),
        .b(jinkela_wire_275),
        .c(jinkela_wire_334)
    );

    or_bb n_857_ (
        .a(jinkela_wire_86),
        .b(jinkela_wire_225),
        .c(jinkela_wire_345)
    );

    and_bi n_774_ (
        .a(jinkela_wire_121),
        .b(jinkela_wire_353),
        .c(jinkela_wire_415)
    );

    or_bb n_816_ (
        .a(jinkela_wire_247),
        .b(jinkela_wire_353),
        .c(jinkela_wire_381)
    );

    and_ii n_858_ (
        .a(jinkela_wire_345),
        .b(jinkela_wire_118),
        .c(jinkela_wire_379)
    );

    or_bb n_775_ (
        .a(jinkela_wire_415),
        .b(jinkela_wire_163),
        .c(jinkela_wire_110)
    );

    and_ii n_817_ (
        .a(jinkela_wire_335),
        .b(jinkela_wire_36),
        .c(jinkela_wire_399)
    );

    and_bb n_859_ (
        .a(jinkela_wire_345),
        .b(jinkela_wire_118),
        .c(jinkela_wire_23)
    );

    and_ii n_776_ (
        .a(jinkela_wire_110),
        .b(jinkela_wire_78),
        .c(jinkela_wire_140)
    );

    and_ii n_818_ (
        .a(jinkela_wire_399),
        .b(jinkela_wire_381),
        .c(jinkela_wire_83)
    );

    or_bb n_860_ (
        .a(jinkela_wire_23),
        .b(jinkela_wire_379),
        .c(jinkela_wire_190)
    );

    and_bb n_777_ (
        .a(jinkela_wire_110),
        .b(jinkela_wire_78),
        .c(jinkela_wire_351)
    );

    and_bb n_819_ (
        .a(jinkela_wire_399),
        .b(jinkela_wire_381),
        .c(jinkela_wire_251)
    );

    or_bb n_861_ (
        .a(jinkela_wire_190),
        .b(jinkela_wire_73),
        .c(jinkela_wire_273)
    );

    or_bb n_778_ (
        .a(jinkela_wire_351),
        .b(jinkela_wire_140),
        .c(jinkela_wire_211)
    );

    or_bb n_820_ (
        .a(jinkela_wire_251),
        .b(jinkela_wire_83),
        .c(jinkela_wire_115)
    );

    or_bb n_779_ (
        .a(jinkela_wire_211),
        .b(jinkela_wire_105),
        .c(jinkela_wire_146)
    );

    and_ii n_821_ (
        .a(jinkela_wire_115),
        .b(jinkela_wire_334),
        .c(jinkela_wire_228)
    );

    and_bb n_780_ (
        .a(jinkela_wire_211),
        .b(jinkela_wire_105),
        .c(jinkela_wire_61)
    );

    or_ii n_822_ (
        .a(jinkela_wire_115),
        .b(jinkela_wire_334),
        .c(jinkela_wire_161)
    );

    or_bi n_781_ (
        .a(jinkela_wire_61),
        .b(jinkela_wire_146),
        .c(jinkela_wire_375)
    );

    and_bi n_823_ (
        .a(jinkela_wire_161),
        .b(jinkela_wire_228),
        .c(s_14_)
    );

    and_ii n_782_ (
        .a(jinkela_wire_375),
        .b(jinkela_wire_276),
        .c(jinkela_wire_404)
    );

    or_bb n_824_ (
        .a(jinkela_wire_83),
        .b(jinkela_wire_72),
        .c(jinkela_wire_293)
    );

    and_bb n_783_ (
        .a(jinkela_wire_375),
        .b(jinkela_wire_276),
        .c(jinkela_wire_367)
    );

    or_bb n_825_ (
        .a(jinkela_wire_293),
        .b(jinkela_wire_228),
        .c(s_15_)
    );

    or_bb n_784_ (
        .a(jinkela_wire_367),
        .b(jinkela_wire_404),
        .c(jinkela_wire_224)
    );

    and_bb n_826_ (
        .a(b_0_),
        .b(a_0_),
        .c(s_0_)
    );

    and_ii n_785_ (
        .a(jinkela_wire_224),
        .b(jinkela_wire_193),
        .c(jinkela_wire_41)
    );

    or_ii n_827_ (
        .a(b_0_),
        .b(a_1_),
        .c(jinkela_wire_278)
    );

    and_bb n_786_ (
        .a(jinkela_wire_224),
        .b(jinkela_wire_193),
        .c(jinkela_wire_232)
    );

    and_bb n_828_ (
        .a(b_1_),
        .b(a_0_),
        .c(jinkela_wire_53)
    );

    or_bb n_787_ (
        .a(jinkela_wire_232),
        .b(jinkela_wire_41),
        .c(jinkela_wire_388)
    );

    or_bi n_829_ (
        .a(jinkela_wire_278),
        .b(jinkela_wire_53),
        .c(jinkela_wire_17)
    );

    and_ii n_788_ (
        .a(jinkela_wire_388),
        .b(jinkela_wire_360),
        .c(jinkela_wire_357)
    );

    and_bi n_830_ (
        .a(jinkela_wire_278),
        .b(jinkela_wire_53),
        .c(jinkela_wire_182)
    );

    and_bb n_789_ (
        .a(jinkela_wire_388),
        .b(jinkela_wire_360),
        .c(jinkela_wire_54)
    );

    and_bi n_831_ (
        .a(jinkela_wire_17),
        .b(jinkela_wire_182),
        .c(s_1_)
    );

    or_bb n_790_ (
        .a(jinkela_wire_54),
        .b(jinkela_wire_357),
        .c(jinkela_wire_10)
    );

    or_ii n_832_ (
        .a(b_2_),
        .b(a_0_),
        .c(jinkela_wire_326)
    );

    and_ii n_791_ (
        .a(jinkela_wire_10),
        .b(jinkela_wire_139),
        .c(jinkela_wire_50)
    );

    or_ii n_833_ (
        .a(a_1_),
        .b(b_1_),
        .c(jinkela_wire_7)
    );

    and_bb n_792_ (
        .a(jinkela_wire_10),
        .b(jinkela_wire_139),
        .c(jinkela_wire_5)
    );

    and_bb n_834_ (
        .a(b_0_),
        .b(a_2_),
        .c(jinkela_wire_180)
    );

    and_ii n_793_ (
        .a(jinkela_wire_5),
        .b(jinkela_wire_50),
        .c(s_12_)
    );

    and_bi n_835_ (
        .a(jinkela_wire_180),
        .b(jinkela_wire_7),
        .c(jinkela_wire_243)
    );

    and_ii n_794_ (
        .a(jinkela_wire_50),
        .b(jinkela_wire_357),
        .c(jinkela_wire_71)
    );

    and_bi n_836_ (
        .a(jinkela_wire_7),
        .b(jinkela_wire_180),
        .c(jinkela_wire_65)
    );

    and_ii n_795_ (
        .a(jinkela_wire_41),
        .b(jinkela_wire_404),
        .c(jinkela_wire_383)
    );

    or_bb n_837_ (
        .a(jinkela_wire_65),
        .b(jinkela_wire_243),
        .c(jinkela_wire_330)
    );

    and_ii n_796_ (
        .a(jinkela_wire_140),
        .b(jinkela_wire_163),
        .c(jinkela_wire_264)
    );

    and_ii n_838_ (
        .a(jinkela_wire_330),
        .b(jinkela_wire_326),
        .c(jinkela_wire_395)
    );

    or_ii n_797_ (
        .a(b_7_),
        .b(a_7_),
        .c(jinkela_wire_247)
    );

    and_bb n_839_ (
        .a(jinkela_wire_330),
        .b(jinkela_wire_326),
        .c(jinkela_wire_286)
    );

    and_bi n_798_ (
        .a(jinkela_wire_353),
        .b(jinkela_wire_247),
        .c(jinkela_wire_72)
    );

    or_bb n_840_ (
        .a(jinkela_wire_286),
        .b(jinkela_wire_395),
        .c(jinkela_wire_94)
    );

    or_ii n_799_ (
        .a(b_6_),
        .b(a_7_),
        .c(jinkela_wire_319)
    );

    or_bb n_841_ (
        .a(jinkela_wire_94),
        .b(jinkela_wire_17),
        .c(jinkela_wire_73)
    );

    and_bb n_800_ (
        .a(b_7_),
        .b(a_6_),
        .c(jinkela_wire_45)
    );

    and_bb n_842_ (
        .a(jinkela_wire_94),
        .b(jinkela_wire_17),
        .c(jinkela_wire_233)
    );

    and_bi n_801_ (
        .a(jinkela_wire_319),
        .b(jinkela_wire_45),
        .c(jinkela_wire_238)
    );

    and_bi n_843_ (
        .a(jinkela_wire_73),
        .b(jinkela_wire_233),
        .c(s_2_)
    );

    or_bb n_802_ (
        .a(jinkela_wire_238),
        .b(jinkela_wire_72),
        .c(jinkela_wire_160)
    );

    or_ii n_844_ (
        .a(b_3_),
        .b(a_0_),
        .c(jinkela_wire_118)
    );

    and_ii n_803_ (
        .a(jinkela_wire_160),
        .b(jinkela_wire_146),
        .c(jinkela_wire_36)
    );

    and_ii n_845_ (
        .a(jinkela_wire_395),
        .b(jinkela_wire_243),
        .c(jinkela_wire_166)
    );

    and_bb n_804_ (
        .a(jinkela_wire_160),
        .b(jinkela_wire_146),
        .c(jinkela_wire_268)
    );

    or_ii n_846_ (
        .a(b_2_),
        .b(a_1_),
        .c(jinkela_wire_136)
    );

    or_bb n_805_ (
        .a(jinkela_wire_268),
        .b(jinkela_wire_36),
        .c(jinkela_wire_90)
    );

    or_ii n_847_ (
        .a(a_2_),
        .b(b_1_),
        .c(jinkela_wire_338)
    );

    and_ii n_806_ (
        .a(jinkela_wire_90),
        .b(jinkela_wire_264),
        .c(jinkela_wire_335)
    );

    or_ii n_848_ (
        .a(b_0_),
        .b(a_3_),
        .c(jinkela_wire_366)
    );

    and_bb n_807_ (
        .a(jinkela_wire_90),
        .b(jinkela_wire_264),
        .c(jinkela_wire_403)
    );

    or_bb n_849_ (
        .a(jinkela_wire_366),
        .b(jinkela_wire_338),
        .c(jinkela_wire_405)
    );

    or_bb n_808_ (
        .a(jinkela_wire_403),
        .b(jinkela_wire_335),
        .c(jinkela_wire_35)
    );

    or_ii n_850_ (
        .a(jinkela_wire_366),
        .b(jinkela_wire_338),
        .c(jinkela_wire_400)
    );

    and_ii n_809_ (
        .a(jinkela_wire_35),
        .b(jinkela_wire_383),
        .c(jinkela_wire_275)
    );

    or_ii n_851_ (
        .a(jinkela_wire_400),
        .b(jinkela_wire_405),
        .c(jinkela_wire_262)
    );

    or_bb n_726_ (
        .a(jinkela_wire_299),
        .b(jinkela_wire_237),
        .c(jinkela_wire_241)
    );

    and_ii n_684_ (
        .a(jinkela_wire_316),
        .b(jinkela_wire_177),
        .c(jinkela_wire_231)
    );

    and_ii n_727_ (
        .a(jinkela_wire_241),
        .b(jinkela_wire_417),
        .c(jinkela_wire_82)
    );

    and_bb n_685_ (
        .a(jinkela_wire_316),
        .b(jinkela_wire_177),
        .c(jinkela_wire_155)
    );

    and_bb n_728_ (
        .a(jinkela_wire_241),
        .b(jinkela_wire_417),
        .c(jinkela_wire_96)
    );

    and_ii n_686_ (
        .a(jinkela_wire_155),
        .b(jinkela_wire_231),
        .c(jinkela_wire_75)
    );

    or_bb n_729_ (
        .a(jinkela_wire_96),
        .b(jinkela_wire_82),
        .c(jinkela_wire_258)
    );

    and_bi n_687_ (
        .a(jinkela_wire_75),
        .b(jinkela_wire_354),
        .c(jinkela_wire_222)
    );

    and_bi n_688_ (
        .a(jinkela_wire_354),
        .b(jinkela_wire_75),
        .c(jinkela_wire_13)
    );

    and_ii n_730_ (
        .a(jinkela_wire_222),
        .b(jinkela_wire_93),
        .c(jinkela_wire_223)
    );

    and_ii n_689_ (
        .a(jinkela_wire_13),
        .b(jinkela_wire_222),
        .c(jinkela_wire_34)
    );

    or_bb n_731_ (
        .a(jinkela_wire_223),
        .b(jinkela_wire_13),
        .c(jinkela_wire_64)
    );

    or_bb n_690_ (
        .a(jinkela_wire_34),
        .b(jinkela_wire_93),
        .c(jinkela_wire_254)
    );

    and_ii n_732_ (
        .a(jinkela_wire_64),
        .b(jinkela_wire_258),
        .c(jinkela_wire_148)
    );

    and_bb n_691_ (
        .a(jinkela_wire_34),
        .b(jinkela_wire_93),
        .c(jinkela_wire_394)
    );

    and_bb n_733_ (
        .a(jinkela_wire_64),
        .b(jinkela_wire_258),
        .c(jinkela_wire_216)
    );

    and_bi n_692_ (
        .a(jinkela_wire_254),
        .b(jinkela_wire_394),
        .c(s_9_)
    );

    and_ii n_734_ (
        .a(jinkela_wire_216),
        .b(jinkela_wire_148),
        .c(s_10_)
    );

    and_ii n_693_ (
        .a(jinkela_wire_231),
        .b(jinkela_wire_310),
        .c(jinkela_wire_417)
    );

    and_ii n_735_ (
        .a(jinkela_wire_148),
        .b(jinkela_wire_82),
        .c(jinkela_wire_47)
    );

    and_ii n_694_ (
        .a(jinkela_wire_141),
        .b(jinkela_wire_322),
        .c(jinkela_wire_147)
    );

    and_ii n_736_ (
        .a(jinkela_wire_237),
        .b(jinkela_wire_157),
        .c(jinkela_wire_80)
    );

    and_ii n_695_ (
        .a(jinkela_wire_149),
        .b(jinkela_wire_57),
        .c(jinkela_wire_29)
    );

    and_ii n_737_ (
        .a(jinkela_wire_414),
        .b(jinkela_wire_346),
        .c(jinkela_wire_197)
    );

    and_ii n_696_ (
        .a(jinkela_wire_88),
        .b(jinkela_wire_358),
        .c(jinkela_wire_126)
    );

    and_ii n_738_ (
        .a(jinkela_wire_27),
        .b(jinkela_wire_181),
        .c(jinkela_wire_263)
    );

    and_bb n_766_ (
        .a(jinkela_wire_392),
        .b(jinkela_wire_47),
        .c(jinkela_wire_272)
    );

    or_ii n_697_ (
        .a(b_5_),
        .b(a_5_),
        .c(jinkela_wire_305)
    );

    or_ii n_739_ (
        .a(b_5_),
        .b(a_7_),
        .c(jinkela_wire_105)
    );

    or_ii n_698_ (
        .a(b_4_),
        .b(a_7_),
        .c(jinkela_wire_106)
    );

    or_bb n_740_ (
        .a(jinkela_wire_105),
        .b(jinkela_wire_246),
        .c(jinkela_wire_121)
    );

    and_bi n_699_ (
        .a(jinkela_wire_229),
        .b(jinkela_wire_106),
        .c(jinkela_wire_250)
    );

    and_bb n_741_ (
        .a(b_5_),
        .b(a_6_),
        .c(jinkela_wire_365)
    );

    and_bb n_700_ (
        .a(b_3_),
        .b(a_7_),
        .c(jinkela_wire_42)
    );

    and_bi n_742_ (
        .a(jinkela_wire_106),
        .b(jinkela_wire_365),
        .c(jinkela_wire_398)
    );

    and_bi n_701_ (
        .a(jinkela_wire_246),
        .b(jinkela_wire_42),
        .c(jinkela_wire_194)
    );

    or_bi n_743_ (
        .a(jinkela_wire_398),
        .b(jinkela_wire_121),
        .c(jinkela_wire_114)
    );

    and_ii n_767_ (
        .a(jinkela_wire_272),
        .b(jinkela_wire_142),
        .c(s_11_)
    );

    or_bb n_702_ (
        .a(jinkela_wire_194),
        .b(jinkela_wire_250),
        .c(jinkela_wire_313)
    );

    or_ii n_744_ (
        .a(b_7_),
        .b(a_4_),
        .c(jinkela_wire_178)
    );

    and_ii n_703_ (
        .a(jinkela_wire_313),
        .b(jinkela_wire_305),
        .c(jinkela_wire_291)
    );

    and_ii n_745_ (
        .a(jinkela_wire_291),
        .b(jinkela_wire_250),
        .c(jinkela_wire_171)
    );

    and_bb n_704_ (
        .a(jinkela_wire_313),
        .b(jinkela_wire_305),
        .c(jinkela_wire_195)
    );

    or_ii n_746_ (
        .a(b_6_),
        .b(a_5_),
        .c(jinkela_wire_412)
    );

    or_bb n_705_ (
        .a(jinkela_wire_195),
        .b(jinkela_wire_291),
        .c(jinkela_wire_261)
    );

    and_ii n_747_ (
        .a(jinkela_wire_412),
        .b(jinkela_wire_171),
        .c(jinkela_wire_67)
    );

    and_ii n_706_ (
        .a(jinkela_wire_261),
        .b(jinkela_wire_126),
        .c(jinkela_wire_181)
    );

    and_bb n_748_ (
        .a(jinkela_wire_412),
        .b(jinkela_wire_171),
        .c(jinkela_wire_16)
    );

    and_bb n_707_ (
        .a(jinkela_wire_261),
        .b(jinkela_wire_126),
        .c(jinkela_wire_174)
    );

    or_bb n_749_ (
        .a(jinkela_wire_16),
        .b(jinkela_wire_67),
        .c(jinkela_wire_257)
    );

    or_bb n_708_ (
        .a(jinkela_wire_174),
        .b(jinkela_wire_181),
        .c(jinkela_wire_274)
    );

    and_ii n_750_ (
        .a(jinkela_wire_257),
        .b(jinkela_wire_178),
        .c(jinkela_wire_333)
    );

    or_ii n_709_ (
        .a(b_7_),
        .b(a_3_),
        .c(jinkela_wire_289)
    );

    and_bb n_751_ (
        .a(jinkela_wire_257),
        .b(jinkela_wire_178),
        .c(jinkela_wire_62)
    );

    and_ii n_710_ (
        .a(jinkela_wire_44),
        .b(jinkela_wire_30),
        .c(jinkela_wire_239)
    );

    or_bb n_752_ (
        .a(jinkela_wire_62),
        .b(jinkela_wire_333),
        .c(jinkela_wire_24)
    );

    or_ii n_711_ (
        .a(b_6_),
        .b(a_4_),
        .c(jinkela_wire_343)
    );

    or_bb n_753_ (
        .a(jinkela_wire_24),
        .b(jinkela_wire_114),
        .c(jinkela_wire_276)
    );

    and_ii n_712_ (
        .a(jinkela_wire_343),
        .b(jinkela_wire_239),
        .c(jinkela_wire_346)
    );

    and_bb n_754_ (
        .a(jinkela_wire_24),
        .b(jinkela_wire_114),
        .c(jinkela_wire_117)
    );

    and_bb n_713_ (
        .a(jinkela_wire_343),
        .b(jinkela_wire_239),
        .c(jinkela_wire_380)
    );

    or_bi n_755_ (
        .a(jinkela_wire_117),
        .b(jinkela_wire_276),
        .c(jinkela_wire_301)
    );

    or_bb n_714_ (
        .a(jinkela_wire_380),
        .b(jinkela_wire_346),
        .c(jinkela_wire_87)
    );

    and_ii n_756_ (
        .a(jinkela_wire_301),
        .b(jinkela_wire_263),
        .c(jinkela_wire_317)
    );

    and_ii n_715_ (
        .a(jinkela_wire_87),
        .b(jinkela_wire_289),
        .c(jinkela_wire_414)
    );

    and_bb n_757_ (
        .a(jinkela_wire_301),
        .b(jinkela_wire_263),
        .c(jinkela_wire_198)
    );

    and_bb n_716_ (
        .a(jinkela_wire_87),
        .b(jinkela_wire_289),
        .c(jinkela_wire_391)
    );

    or_bb n_758_ (
        .a(jinkela_wire_198),
        .b(jinkela_wire_317),
        .c(jinkela_wire_307)
    );

    or_bb n_717_ (
        .a(jinkela_wire_391),
        .b(jinkela_wire_414),
        .c(jinkela_wire_409)
    );

    and_ii n_759_ (
        .a(jinkela_wire_307),
        .b(jinkela_wire_197),
        .c(jinkela_wire_84)
    );

    and_ii n_718_ (
        .a(jinkela_wire_409),
        .b(jinkela_wire_274),
        .c(jinkela_wire_27)
    );

    and_bb n_760_ (
        .a(jinkela_wire_307),
        .b(jinkela_wire_197),
        .c(jinkela_wire_288)
    );

    and_bb n_719_ (
        .a(jinkela_wire_409),
        .b(jinkela_wire_274),
        .c(jinkela_wire_43)
    );

    or_bb n_761_ (
        .a(jinkela_wire_288),
        .b(jinkela_wire_84),
        .c(jinkela_wire_76)
    );

    or_bb n_720_ (
        .a(jinkela_wire_43),
        .b(jinkela_wire_27),
        .c(jinkela_wire_191)
    );

    and_ii n_762_ (
        .a(jinkela_wire_76),
        .b(jinkela_wire_80),
        .c(jinkela_wire_296)
    );

    and_ii n_721_ (
        .a(jinkela_wire_191),
        .b(jinkela_wire_29),
        .c(jinkela_wire_157)
    );

    and_bb n_763_ (
        .a(jinkela_wire_76),
        .b(jinkela_wire_80),
        .c(jinkela_wire_253)
    );

    and_bb n_722_ (
        .a(jinkela_wire_191),
        .b(jinkela_wire_29),
        .c(jinkela_wire_242)
    );

    or_bb n_764_ (
        .a(jinkela_wire_253),
        .b(jinkela_wire_296),
        .c(jinkela_wire_392)
    );

    or_bb n_723_ (
        .a(jinkela_wire_242),
        .b(jinkela_wire_157),
        .c(jinkela_wire_321)
    );

    and_ii n_765_ (
        .a(jinkela_wire_392),
        .b(jinkela_wire_47),
        .c(jinkela_wire_142)
    );

    and_ii n_724_ (
        .a(jinkela_wire_321),
        .b(jinkela_wire_147),
        .c(jinkela_wire_237)
    );

    and_bb n_725_ (
        .a(jinkela_wire_321),
        .b(jinkela_wire_147),
        .c(jinkela_wire_299)
    );

endmodule
