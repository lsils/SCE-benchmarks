module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 );
  input G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 ;
  output G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 ;
  wire n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 ;
  buffer buf_n160( .i (G115), .o (n160) );
  buffer buf_n213( .i (G124), .o (n213) );
  buffer buf_n275( .i (G137), .o (n275) );
  buffer buf_n320( .i (G32), .o (n320) );
  buffer buf_n159( .i (G106), .o (n159) );
  buffer buf_n323( .i (G64), .o (n323) );
  buffer buf_n324( .i (G76), .o (n324) );
  buffer buf_n322( .i (G53), .o (n322) );
  buffer buf_n331( .i (G96), .o (n331) );
  buffer buf_n321( .i (G43), .o (n321) );
  buffer buf_n330( .i (G86), .o (n330) );
  buffer buf_n300( .i (G141), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n305( .i (G142), .o (n305) );
  assign n332 = n301 | n305 ;
  buffer buf_n286( .i (G139), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n294( .i (G140), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  assign n333 = n290 | n295 ;
  assign n334 = n332 | n333 ;
  buffer buf_n206( .i (G121), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  assign n335 = G2 | n208 ;
  assign n336 = G11 | n335 ;
  buffer buf_n161( .i (n160), .o (n161) );
  assign n337 = ~G74 & n161 ;
  assign n338 = G7 | n207 ;
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n180( .i (G119), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  assign n340 = n185 | n339 ;
  buffer buf_n310( .i (G147), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  assign n341 = n315 | n339 ;
  assign n342 = n322 & ~n331 ;
  assign n343 = n321 | n330 ;
  assign n344 = n342 & ~n343 ;
  buffer buf_n345( .i (n344), .o (n345) );
  assign n346 = ~n159 & n320 ;
  assign n347 = n323 | n324 ;
  assign n348 = n346 & ~n347 ;
  buffer buf_n349( .i (n348), .o (n349) );
  assign n350 = n345 | n349 ;
  buffer buf_n351( .i (n350), .o (n351) );
  assign n352 = n310 & ~n349 ;
  assign n353 = n180 & ~n345 ;
  assign n354 = n352 | n353 ;
  buffer buf_n355( .i (n354), .o (n355) );
  assign n356 = G145 | G146 ;
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  assign n372 = G109 & ~n360 ;
  assign n373 = G79 & ~n360 ;
  assign n374 = n372 | n373 ;
  assign n375 = G89 & ~n360 ;
  buffer buf_n376( .i (n359), .o (n376) );
  assign n377 = G99 & ~n376 ;
  assign n378 = n375 | n377 ;
  assign n379 = n374 | n378 ;
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  assign n396 = G108 | n370 ;
  assign n397 = G98 & ~n370 ;
  assign n398 = n396 & ~n397 ;
  assign n399 = G88 & ~n370 ;
  buffer buf_n400( .i (n369), .o (n400) );
  assign n401 = G78 & ~n400 ;
  assign n402 = n399 | n401 ;
  assign n403 = n398 & ~n402 ;
  buffer buf_n404( .i (n403), .o (n404) );
  assign n407 = G80 | n376 ;
  assign n408 = G90 & ~n376 ;
  assign n409 = n407 & ~n408 ;
  assign n410 = G100 & ~n376 ;
  buffer buf_n411( .i (n359), .o (n411) );
  assign n412 = G110 & ~n411 ;
  assign n413 = n410 | n412 ;
  assign n414 = n409 & ~n413 ;
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n162( .i (G117), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  assign n427 = ~G36 & n169 ;
  buffer buf_n191( .i (G120), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  assign n428 = ~G68 & n168 ;
  assign n429 = n198 | n428 ;
  assign n430 = n427 & ~n429 ;
  assign n431 = n162 | n191 ;
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  assign n445 = G46 & ~n437 ;
  assign n446 = G57 & ~n437 ;
  assign n447 = n445 | n446 ;
  assign n448 = n430 & ~n447 ;
  buffer buf_n449( .i (n448), .o (n449) );
  assign n451 = ~G37 & n168 ;
  assign n452 = ~G69 & n167 ;
  assign n453 = n197 | n452 ;
  assign n454 = n451 & ~n453 ;
  assign n455 = G47 & ~n436 ;
  assign n456 = G58 & ~n436 ;
  assign n457 = n455 | n456 ;
  assign n458 = n454 & ~n457 ;
  buffer buf_n459( .i (n458), .o (n459) );
  assign n469 = ~G38 & n168 ;
  assign n470 = ~G70 & n167 ;
  assign n471 = n197 | n470 ;
  assign n472 = n469 & ~n471 ;
  assign n473 = G48 & ~n436 ;
  buffer buf_n474( .i (n435), .o (n474) );
  assign n475 = G59 & ~n474 ;
  assign n476 = n473 | n475 ;
  assign n477 = n472 & ~n476 ;
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n209( .i (G122), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  assign n488 = ~G31 & n167 ;
  assign n489 = ~G63 & n166 ;
  assign n490 = n196 | n489 ;
  assign n491 = n488 & ~n490 ;
  assign n492 = G42 & ~n435 ;
  assign n493 = G52 & ~n435 ;
  assign n494 = n492 | n493 ;
  assign n495 = n491 & ~n494 ;
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  assign n509 = n210 | n508 ;
  assign n510 = G116 | n206 ;
  assign n511 = n355 | n510 ;
  buffer buf_n512( .i (n511), .o (n512) );
  assign n513 = G28 | n512 ;
  assign n514 = G1 & ~G3 ;
  assign n515 = n512 | n514 ;
  buffer buf_n516( .i (n166), .o (n516) );
  assign n517 = G39 | n516 ;
  assign n518 = ~G71 & n166 ;
  assign n519 = n196 | n518 ;
  assign n520 = n517 & ~n519 ;
  buffer buf_n521( .i (n434), .o (n521) );
  assign n522 = G49 & ~n521 ;
  assign n523 = G60 & ~n521 ;
  assign n524 = n522 | n523 ;
  assign n525 = n520 | n524 ;
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  assign n537 = G56 & ~n440 ;
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  assign n538 = G35 | n171 ;
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  assign n539 = ~G67 & n170 ;
  assign n540 = n200 | n539 ;
  assign n541 = n538 & ~n540 ;
  assign n542 = n537 & ~n541 ;
  buffer buf_n543( .i (n542), .o (n543) );
  assign n545 = ~G34 & n169 ;
  buffer buf_n546( .i (n516), .o (n546) );
  assign n547 = ~G66 & n546 ;
  assign n548 = n198 | n547 ;
  assign n549 = n545 & ~n548 ;
  assign n550 = G45 & ~n437 ;
  buffer buf_n551( .i (n474), .o (n551) );
  assign n552 = G55 & ~n551 ;
  assign n553 = n550 | n552 ;
  assign n554 = n549 & ~n553 ;
  buffer buf_n555( .i (n554), .o (n555) );
  assign n562 = ~G33 & n169 ;
  assign n563 = ~G65 & n546 ;
  assign n564 = n198 | n563 ;
  assign n565 = n562 & ~n564 ;
  assign n566 = G44 & ~n551 ;
  assign n567 = G54 & ~n551 ;
  assign n568 = n566 | n567 ;
  assign n569 = n565 & ~n568 ;
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n211( .i (G123), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  assign n574 = ~G40 & n516 ;
  buffer buf_n575( .i (n165), .o (n575) );
  assign n576 = ~G72 & n575 ;
  assign n577 = n196 | n576 ;
  assign n578 = n574 & ~n577 ;
  assign n579 = G50 & ~n521 ;
  assign n580 = G61 & ~n521 ;
  assign n581 = n579 | n580 ;
  assign n582 = n578 & ~n581 ;
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  assign n596 = n212 | n593 ;
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  assign n597 = n212 & ~n487 ;
  assign n598 = n596 & ~n597 ;
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  assign n600 = n212 | n536 ;
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  assign n601 = ~n212 & n468 ;
  assign n602 = n600 & ~n601 ;
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n177( .i (G118), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  assign n604 = n179 & ~n209 ;
  assign n605 = n595 | n604 ;
  buffer buf_n606( .i (n211), .o (n606) );
  assign n607 = ~n506 & n606 ;
  assign n608 = n177 | n211 ;
  assign n609 = n593 & ~n608 ;
  assign n610 = n607 | n609 ;
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n309( .i (G143), .o (n309) );
  buffer buf_n371( .i (n370), .o (n371) );
  assign n612 = G77 & ~n371 ;
  assign n613 = G97 & ~n371 ;
  assign n614 = n612 & ~n613 ;
  assign n615 = G107 & ~n371 ;
  assign n616 = G87 & ~n371 ;
  assign n617 = n615 | n616 ;
  assign n618 = n614 & ~n617 ;
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  assign n627 = n309 | n626 ;
  assign n628 = n309 & ~n626 ;
  assign n629 = n627 & ~n628 ;
  assign n630 = G144 | n629 ;
  buffer buf_n158( .i (G10), .o (n158) );
  inverter inv_n972( .i (n158), .o (n972) );
  buffer buf_n263( .i (G135), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n316( .i (G23), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  assign n631 = ~G19 & n318 ;
  buffer buf_n632( .i (n400), .o (n632) );
  assign n633 = G75 & ~n632 ;
  assign n634 = G85 & ~n632 ;
  assign n635 = n633 & ~n634 ;
  assign n636 = G95 & ~n632 ;
  assign n637 = G105 & ~n632 ;
  assign n638 = n636 | n637 ;
  assign n639 = n635 & ~n638 ;
  buffer buf_n640( .i (n639), .o (n640) );
  assign n642 = n318 & ~n640 ;
  assign n643 = n631 & ~n642 ;
  assign n644 = n264 & ~n643 ;
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n214( .i (G125), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n186( .i (G12), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  assign n648 = ~G13 & n188 ;
  assign n649 = n188 & ~n498 ;
  assign n650 = n648 & ~n649 ;
  assign n651 = n220 & ~n650 ;
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n242( .i (G130), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  assign n655 = ~G15 & n188 ;
  buffer buf_n656( .i (n187), .o (n656) );
  assign n657 = n460 & ~n656 ;
  assign n658 = n655 & ~n657 ;
  assign n659 = n246 & ~n658 ;
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  assign n663 = n654 | n662 ;
  assign n664 = n647 | n663 ;
  buffer buf_n237( .i (G129), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  assign n665 = ~G5 & n656 ;
  assign n666 = ~n479 & n656 ;
  assign n667 = n665 & ~n666 ;
  assign n668 = n241 & ~n667 ;
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  assign n671 = ~G21 & n318 ;
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n672( .i (n317), .o (n672) );
  assign n673 = ~n426 & n672 ;
  assign n674 = n671 & ~n673 ;
  assign n675 = n299 & ~n674 ;
  buffer buf_n676( .i (n675), .o (n676) );
  assign n677 = n670 | n676 ;
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  assign n678 = ~G27 & n317 ;
  assign n679 = n317 & ~n404 ;
  assign n680 = n678 & ~n679 ;
  assign n681 = n308 & ~n680 ;
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  assign n684 = n645 | n683 ;
  assign n685 = n677 | n684 ;
  buffer buf_n229( .i (G128), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  assign n686 = ~G14 & n656 ;
  buffer buf_n687( .i (n187), .o (n687) );
  assign n688 = n528 & ~n687 ;
  assign n689 = n686 & ~n688 ;
  assign n690 = n236 & ~n689 ;
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n221( .i (G126), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  assign n693 = ~G4 & n687 ;
  assign n694 = ~n585 & n687 ;
  assign n695 = n693 & ~n694 ;
  assign n696 = n228 & ~n695 ;
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  assign n699 = n692 | n698 ;
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n700( .i (n316), .o (n700) );
  assign n701 = ~G26 & n700 ;
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  assign n702 = ~n390 & n700 ;
  assign n703 = n701 & ~n702 ;
  assign n704 = n304 & ~n703 ;
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  assign n707 = n676 | n706 ;
  assign n708 = n699 | n707 ;
  assign n709 = n685 | n708 ;
  assign n710 = n664 | n709 ;
  buffer buf_n265( .i (G136), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n319( .i (n318), .o (n319) );
  assign n711 = ~G24 & n319 ;
  buffer buf_n712( .i (n400), .o (n712) );
  assign n713 = G93 & ~n712 ;
  assign n714 = G103 & ~n712 ;
  assign n715 = n713 & ~n714 ;
  assign n716 = G113 & ~n712 ;
  assign n717 = G83 & ~n712 ;
  assign n718 = n716 | n717 ;
  assign n719 = n715 & ~n718 ;
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  assign n722 = n319 & ~n721 ;
  assign n723 = n711 & ~n722 ;
  buffer buf_n724( .i (n723), .o (n724) );
  assign n725 = n274 | n724 ;
  assign n726 = n274 & ~n724 ;
  assign n727 = n725 & ~n726 ;
  buffer buf_n247( .i (G131), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n189( .i (n188), .o (n189) );
  assign n728 = ~G16 & n189 ;
  buffer buf_n450( .i (n449), .o (n450) );
  assign n729 = n189 & ~n450 ;
  assign n730 = n728 & ~n729 ;
  buffer buf_n731( .i (n730), .o (n731) );
  assign n732 = n252 | n731 ;
  assign n733 = n252 & ~n731 ;
  assign n734 = n732 & ~n733 ;
  buffer buf_n276( .i (G138), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  assign n735 = ~G20 & n672 ;
  buffer buf_n736( .i (n400), .o (n736) );
  assign n737 = G82 & ~n736 ;
  assign n738 = G102 & ~n736 ;
  assign n739 = n737 & ~n738 ;
  assign n740 = G112 & ~n736 ;
  assign n741 = G92 & ~n736 ;
  assign n742 = n740 | n741 ;
  assign n743 = n739 & ~n742 ;
  buffer buf_n744( .i (n743), .o (n744) );
  assign n747 = n672 & ~n744 ;
  assign n748 = n735 & ~n747 ;
  buffer buf_n749( .i (n748), .o (n749) );
  assign n750 = n285 | n749 ;
  assign n751 = n285 & ~n749 ;
  assign n752 = n750 & ~n751 ;
  assign n753 = n734 | n752 ;
  assign n754 = n727 | n753 ;
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  assign n755 = ~G25 & n700 ;
  buffer buf_n756( .i (n369), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = G81 & ~n757 ;
  assign n759 = G101 & ~n757 ;
  assign n760 = n758 & ~n759 ;
  assign n761 = G111 & ~n757 ;
  assign n762 = G91 & ~n757 ;
  assign n763 = n761 | n762 ;
  assign n764 = n760 & ~n763 ;
  assign n765 = n700 & ~n764 ;
  assign n766 = n755 & ~n765 ;
  assign n767 = n293 & ~n766 ;
  buffer buf_n768( .i (n767), .o (n768) );
  assign n769 = n660 | n768 ;
  buffer buf_n261( .i (G134), .o (n261) );
  assign n770 = ~G18 & n687 ;
  buffer buf_n771( .i (n187), .o (n771) );
  assign n772 = ~n570 & n771 ;
  assign n773 = n770 & ~n772 ;
  assign n774 = n261 & ~n773 ;
  buffer buf_n775( .i (n774), .o (n775) );
  assign n776 = n697 | n775 ;
  assign n777 = n769 | n776 ;
  buffer buf_n255( .i (G133), .o (n255) );
  assign n778 = ~G6 & n771 ;
  assign n779 = ~n555 & n771 ;
  assign n780 = n778 & ~n779 ;
  assign n781 = n255 & ~n780 ;
  buffer buf_n782( .i (n781), .o (n782) );
  assign n783 = n319 & ~n620 ;
  assign n784 = ~G22 & n672 ;
  assign n785 = G9 | n784 ;
  assign n786 = n783 | n785 ;
  assign n787 = n782 | n786 ;
  assign n788 = n682 | n782 ;
  assign n789 = n787 | n788 ;
  assign n790 = n777 | n789 ;
  assign n791 = n669 | n705 ;
  assign n792 = n652 | n691 ;
  assign n793 = n791 | n792 ;
  assign n794 = n768 | n775 ;
  buffer buf_n253( .i (G132), .o (n253) );
  buffer buf_n190( .i (n189), .o (n190) );
  assign n795 = ~G17 & n190 ;
  assign n796 = n190 & ~n543 ;
  assign n797 = n795 & ~n796 ;
  assign n798 = n253 & ~n797 ;
  assign n799 = n794 | n798 ;
  assign n800 = n793 | n799 ;
  assign n801 = n790 | n800 ;
  assign n802 = n754 | n801 ;
  assign n803 = n710 | n802 ;
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  assign n805 = ~G41 & n176 ;
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  assign n806 = ~G73 & n175 ;
  assign n807 = n205 | n806 ;
  assign n808 = n805 & ~n807 ;
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  assign n809 = G51 & ~n444 ;
  assign n810 = G62 & ~n444 ;
  assign n811 = n809 | n810 ;
  assign n812 = n808 & ~n811 ;
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  assign n816 = n209 & ~n815 ;
  assign n817 = n210 | n816 ;
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  assign n818 = n406 | n620 ;
  assign n819 = n406 & ~n620 ;
  assign n820 = n818 & ~n819 ;
  buffer buf_n821( .i (n820), .o (n821) );
  assign n822 = n395 | n821 ;
  assign n823 = ~n395 & n821 ;
  assign n824 = n822 & ~n823 ;
  assign n825 = G29 | n824 ;
  buffer buf_n826( .i (n825), .o (n826) );
  inverter inv_n973( .i (n826), .o (n973) );
  assign n827 = n211 & ~n813 ;
  assign n828 = n606 | n827 ;
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n325( .i (G8), .o (n325) );
  assign n830 = G127 | n415 ;
  buffer buf_n831( .i (n830), .o (n831) );
  assign n832 = G30 | n380 ;
  buffer buf_n833( .i (n832), .o (n833) );
  assign n834 = n831 | n833 ;
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  assign n840 = ~n325 & n837 ;
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  assign n851 = ~n260 & n850 ;
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  assign n852 = n325 | n837 ;
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  assign n862 = n561 | n861 ;
  buffer buf_n254( .i (n253), .o (n254) );
  assign n863 = ~n254 & n848 ;
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  assign n864 = n237 & n839 ;
  assign n865 = n294 & ~n839 ;
  assign n866 = n864 & ~n865 ;
  assign n867 = n479 & ~n866 ;
  buffer buf_n868( .i (n867), .o (n868) );
  assign n869 = ~n229 & n836 ;
  assign n870 = n286 & ~n836 ;
  assign n871 = n869 | n870 ;
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  assign n875 = ~n528 & n874 ;
  assign n876 = ~n221 & n836 ;
  buffer buf_n877( .i (n835), .o (n877) );
  assign n878 = n276 & ~n877 ;
  assign n879 = n876 | n878 ;
  buffer buf_n880( .i (n879), .o (n880) );
  assign n881 = n583 | n880 ;
  assign n882 = ~n214 & n837 ;
  buffer buf_n883( .i (n877), .o (n883) );
  assign n884 = n265 & ~n883 ;
  assign n885 = n882 | n884 ;
  assign n886 = ~n496 & n885 ;
  assign n887 = n881 & n886 ;
  assign n888 = n583 & n880 ;
  assign n889 = n526 & n872 ;
  assign n890 = n888 | n889 ;
  assign n891 = n887 | n890 ;
  assign n892 = ~n875 & n891 ;
  assign n893 = n868 | n892 ;
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  assign n894 = n328 & ~n459 ;
  assign n895 = n242 & n841 ;
  assign n896 = n300 & ~n853 ;
  assign n897 = n895 & ~n896 ;
  assign n898 = n894 & ~n897 ;
  buffer buf_n899( .i (n898), .o (n899) );
  assign n901 = n868 | n899 ;
  assign n902 = n893 & ~n901 ;
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n329( .i (n328), .o (n329) );
  assign n903 = n329 & ~n449 ;
  assign n904 = n247 & n842 ;
  assign n905 = n305 & ~n854 ;
  assign n906 = n904 & ~n905 ;
  assign n907 = n903 & ~n906 ;
  buffer buf_n908( .i (n907), .o (n908) );
  assign n910 = n900 | n908 ;
  assign n911 = n902 | n910 ;
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n544( .i (n543), .o (n544) );
  assign n912 = n544 & ~n858 ;
  assign n913 = n909 | n912 ;
  assign n914 = n911 & ~n913 ;
  assign n915 = n863 | n914 ;
  assign n916 = n862 & n915 ;
  assign n917 = n851 | n916 ;
  assign n918 = n831 & ~n833 ;
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  assign n931 = n270 | n720 ;
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  assign n935 = n930 & ~n934 ;
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  assign n936 = n284 | n746 ;
  assign n937 = n929 & ~n936 ;
  buffer buf_n938( .i (n937), .o (n938) );
  assign n942 = n935 & ~n938 ;
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n641( .i (n640), .o (n641) );
  assign n944 = n263 | n641 ;
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  assign n948 = n262 & ~n573 ;
  assign n949 = n945 & ~n948 ;
  assign n950 = n930 & ~n949 ;
  assign n951 = n938 | n950 ;
  assign n952 = n263 & ~n641 ;
  assign n953 = n932 & ~n952 ;
  assign n954 = n929 & ~n953 ;
  buffer buf_n955( .i (n954), .o (n955) );
  assign n957 = n262 | n573 ;
  assign n958 = n929 & ~n957 ;
  buffer buf_n959( .i (n958), .o (n959) );
  assign n960 = n955 | n959 ;
  assign n961 = n951 | n960 ;
  assign n962 = n943 & ~n961 ;
  assign n963 = n917 & n962 ;
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  assign n964 = n947 & ~n959 ;
  assign n965 = n956 & ~n964 ;
  assign n966 = n943 & ~n965 ;
  assign n967 = n941 | n966 ;
  assign n968 = ~n963 & ~n967 ;
  assign n969 = n158 & ~n355 ;
  assign n970 = n826 & n969 ;
  inverter inv_n971( .i (n970), .o (n971) );
  assign G2531 = n160 ;
  assign G2532 = n160 ;
  assign G2533 = n160 ;
  assign G2534 = n213 ;
  assign G2535 = n213 ;
  assign G2536 = n275 ;
  assign G2537 = n275 ;
  assign G2538 = n275 ;
  assign G2539 = n320 ;
  assign G2540 = n159 ;
  assign G2541 = n323 ;
  assign G2542 = n324 ;
  assign G2543 = n322 ;
  assign G2544 = n331 ;
  assign G2545 = n321 ;
  assign G2546 = n330 ;
  assign G2547 = n334 ;
  assign G2548 = n336 ;
  assign G2549 = n161 ;
  assign G2550 = n337 ;
  assign G2551 = n339 ;
  assign G2552 = n340 ;
  assign G2553 = n341 ;
  assign G2554 = n351 ;
  assign G2555 = n351 ;
  assign G2556 = n355 ;
  assign G2557 = n380 ;
  assign G2558 = n404 ;
  assign G2559 = n415 ;
  assign G2560 = n449 ;
  assign G2561 = n459 ;
  assign G2562 = n478 ;
  assign G2563 = n509 ;
  assign G2564 = n513 ;
  assign G2565 = n515 ;
  assign G2566 = n526 ;
  assign G2567 = n478 ;
  assign G2568 = n459 ;
  assign G2569 = n449 ;
  assign G2570 = n543 ;
  assign G2571 = n555 ;
  assign G2572 = n570 ;
  assign G2573 = n599 ;
  assign G2574 = n599 ;
  assign G2575 = n603 ;
  assign G2576 = n603 ;
  assign G2577 = n605 ;
  assign G2578 = n611 ;
  assign G2579 = n611 ;
  assign G2580 = n630 ;
  assign G2581 = n972 ;
  assign G2582 = 1'b0 ;
  assign G2583 = 1'b0 ;
  assign G2584 = n804 ;
  assign G2585 = n804 ;
  assign G2586 = n817 ;
  assign G2587 = n973 ;
  assign G2588 = n829 ;
  assign G2589 = n829 ;
  assign G2590 = 1'b0 ;
  assign G2591 = n968 ;
  assign G2592 = 1'b0 ;
  assign G2593 = n971 ;
  assign G2594 = n971 ;
endmodule
