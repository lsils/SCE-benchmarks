module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n2 , n3 , n4 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n66 , n67 , n68 , n69 , n70 , n71 , n73 , n74 , n75 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n150 , n151 , n152 , n153 , n154 , n156 , n157 , n158 , n162 , n163 , n164 , n165 , n167 , n168 , n169 , n170 , n171 , n172 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n182 , n183 , n184 , n185 , n186 , n187 , n189 , n190 , n191 , n192 , n193 , n195 , n196 , n197 , n198 , n199 , n201 , n202 , n203 , n204 , n205 , n206 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 ;
  buffer buf_n40( .i (x4), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n97( .i (x11), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  assign n209 = n46 | n103 ;
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n120( .i (x13), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n150( .i (x16), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  assign n212 = n121 & n151 ;
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n109( .i (x12), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n139( .i (x15), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  assign n219 = n116 & n146 ;
  assign n220 = ( n210 & ~n218 ) | ( n210 & n219 ) | ( ~n218 & n219 ) ;
  assign n221 = ~n211 & n220 ;
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n131( .i (x14), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  assign n224 = n103 | n137 ;
  assign n225 = n115 & ~n216 ;
  assign n226 = ( n116 & ~n224 ) | ( n116 & n225 ) | ( ~n224 & n225 ) ;
  assign n227 = ~n111 & n133 ;
  buffer buf_n228( .i (n227), .o (n228) );
  assign n229 = n44 | n228 ;
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  assign n234 = n226 | n232 ;
  assign n235 = ( n129 & ~n148 ) | ( n129 & n234 ) | ( ~n148 & n234 ) ;
  buffer buf_n152( .i (n151), .o (n152) );
  assign n236 = n99 | n152 ;
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  assign n239 = ~n114 & n238 ;
  assign n240 = ( ~n126 & n145 ) | ( ~n126 & n239 ) | ( n145 & n239 ) ;
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  assign n244 = n235 | n243 ;
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n18( .i (x2), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n167( .i (x21), .o (n167) );
  buffer buf_n182( .i (x23), .o (n182) );
  assign n246 = ~n167 & n182 ;
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n174( .i (x22), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  assign n253 = n18 | n174 ;
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n189( .i (x24), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n201( .i (x26), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  assign n258 = n190 & n202 ;
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  assign n261 = ( n178 & n256 ) | ( n178 & n260 ) | ( n256 & n260 ) ;
  buffer buf_n262( .i (n261), .o (n262) );
  assign n265 = n251 & ~n262 ;
  buffer buf_n266( .i (n265), .o (n266) );
  assign n268 = n26 & n266 ;
  buffer buf_n162( .i (x20), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  assign n269 = x18 | x19 ;
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n156( .i (x17), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  assign n275 = n133 & ~n158 ;
  assign n276 = ( ~n165 & n272 ) | ( ~n165 & n275 ) | ( n272 & n275 ) ;
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n273( .i (n272), .o (n273) );
  assign n278 = n101 & ~n273 ;
  assign n279 = n277 & n278 ;
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  assign n284 = n268 & n282 ;
  buffer buf_n285( .i (n284), .o (n285) );
  assign n286 = n222 | n285 ;
  assign n287 = ( n223 & ~n245 ) | ( n223 & n286 ) | ( ~n245 & n286 ) ;
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n233( .i (n232), .o (n233) );
  assign n289 = n142 & n213 ;
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  assign n293 = n280 & n292 ;
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n257( .i (n256), .o (n257) );
  assign n294 = n206 & ~n257 ;
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = n252 & n295 ;
  assign n297 = n293 & n296 ;
  assign n298 = ~n99 & n152 ;
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  assign n301 = ~n144 & n300 ;
  buffer buf_n302( .i (n301), .o (n302) );
  assign n303 = ~n231 & n302 ;
  buffer buf_n304( .i (n303), .o (n304) );
  assign n305 = ( ~n233 & n297 ) | ( ~n233 & n304 ) | ( n297 & n304 ) ;
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n104( .i (n103), .o (n104) );
  assign n310 = ~n123 & n142 ;
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  assign n314 = n104 & ~n313 ;
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n27( .i (n26), .o (n27) );
  assign n318 = ~n116 & n146 ;
  buffer buf_n319( .i (n318), .o (n319) );
  assign n320 = ~n27 & n319 ;
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n274( .i (n273), .o (n274) );
  assign n322 = ~n274 & n277 ;
  assign n323 = n291 & n322 ;
  buffer buf_n324( .i (n323), .o (n324) );
  assign n326 = n214 & n228 ;
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n195( .i (x25), .o (n195) );
  assign n330 = ( n18 & n195 ) | ( n18 & n201 ) | ( n195 & n201 ) ;
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n183( .i (n182), .o (n183) );
  assign n335 = n183 | n190 ;
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  assign n338 = n167 & n174 ;
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  assign n343 = ( n333 & ~n337 ) | ( n333 & n341 ) | ( ~n337 & n341 ) ;
  assign n344 = ~n334 & n343 ;
  assign n345 = n327 | n344 ;
  buffer buf_n346( .i (n345), .o (n346) );
  assign n347 = ( n324 & n329 ) | ( n324 & n346 ) | ( n329 & n346 ) ;
  buffer buf_n348( .i (n347), .o (n348) );
  assign n349 = n316 & ~n348 ;
  assign n350 = ( n317 & n321 ) | ( n317 & n349 ) | ( n321 & n349 ) ;
  buffer buf_n29( .i (x3), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  assign n351 = n35 & ~n115 ;
  assign n352 = ( n36 & n292 ) | ( n36 & n351 ) | ( n292 & n351 ) ;
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  assign n356 = n122 | n152 ;
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  assign n360 = n144 & n358 ;
  assign n361 = ( n137 & n359 ) | ( n137 & ~n360 ) | ( n359 & ~n360 ) ;
  assign n362 = n121 & n132 ;
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  assign n366 = ~n102 & n365 ;
  assign n367 = n140 & ~n151 ;
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  assign n372 = ( ~n103 & n366 ) | ( ~n103 & n371 ) | ( n366 & n371 ) ;
  assign n373 = n361 & ~n372 ;
  assign n374 = n140 & n151 ;
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  assign n377 = n135 & n376 ;
  buffer buf_n378( .i (n377), .o (n378) );
  assign n379 = n115 & ~n378 ;
  assign n380 = ~n47 & n379 ;
  assign n381 = ( ~n48 & n373 ) | ( ~n48 & n380 ) | ( n373 & n380 ) ;
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  assign n383 = ~n143 & n154 ;
  assign n384 = ~n22 & n135 ;
  assign n385 = ( n23 & n383 ) | ( n23 & ~n384 ) | ( n383 & ~n384 ) ;
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  assign n389 = n106 | n388 ;
  assign n390 = ( ~n354 & n382 ) | ( ~n354 & n389 ) | ( n382 & n389 ) ;
  assign n391 = n355 & n390 ;
  assign n392 = ~n350 & n391 ;
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  assign n394 = ~n20 & n169 ;
  assign n395 = ( n170 & n259 ) | ( n170 & n394 ) | ( n259 & n394 ) ;
  assign n396 = ~n178 & n395 ;
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  assign n397 = ( n185 & n192 ) | ( n185 & n198 ) | ( n192 & n198 ) ;
  assign n398 = n192 | n204 ;
  assign n399 = n397 & n398 ;
  assign n400 = n396 & ~n399 ;
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n403 = n196 & n202 ;
  buffer buf_n404( .i (n403), .o (n404) );
  assign n407 = n169 | n191 ;
  assign n408 = ( n170 & n404 ) | ( n170 & n407 ) | ( n404 & n407 ) ;
  assign n409 = n186 | n408 ;
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  assign n412 = n182 & n189 ;
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n199( .i (n198), .o (n199) );
  assign n420 = n18 | n201 ;
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  assign n424 = n199 & n423 ;
  assign n425 = n337 & n341 ;
  assign n426 = ( n342 & n424 ) | ( n342 & n425 ) | ( n424 & n425 ) ;
  assign n427 = ( n410 & n417 ) | ( n410 & n426 ) | ( n417 & n426 ) ;
  assign n428 = n411 & ~n427 ;
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  assign n429 = ~n189 & n195 ;
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  assign n434 = n19 & n202 ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n436 = n185 & ~n435 ;
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n193( .i (n192), .o (n193) );
  assign n438 = n20 & n197 ;
  buffer buf_n439( .i (n438), .o (n439) );
  assign n441 = ( n193 & n260 ) | ( n193 & ~n439 ) | ( n260 & ~n439 ) ;
  assign n442 = ( n433 & ~n437 ) | ( n433 & n441 ) | ( ~n437 & n441 ) ;
  assign n443 = n180 | n442 ;
  assign n444 = n401 | n443 ;
  assign n445 = ( n402 & ~n428 ) | ( n402 & n444 ) | ( ~n428 & n444 ) ;
  assign n446 = n174 | n182 ;
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = ( ~n169 & n254 ) | ( ~n169 & n339 ) | ( n254 & n339 ) ;
  assign n450 = n430 & ~n447 ;
  assign n451 = ( n448 & n449 ) | ( n448 & n450 ) | ( n449 & n450 ) ;
  assign n452 = ~n203 & n331 ;
  assign n453 = ~n247 & n331 ;
  assign n454 = ( n204 & n452 ) | ( n204 & ~n453 ) | ( n452 & ~n453 ) ;
  assign n455 = n451 | n454 ;
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  assign n458 = ~n171 & n205 ;
  assign n459 = ( ~n172 & n433 ) | ( ~n172 & n458 ) | ( n433 & n458 ) ;
  assign n460 = n189 & ~n195 ;
  buffer buf_n461( .i (n460), .o (n461) );
  assign n465 = n203 | n461 ;
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  assign n468 = n19 & ~n190 ;
  buffer buf_n469( .i (n468), .o (n469) );
  assign n472 = n185 & ~n469 ;
  assign n473 = ( n171 & n466 ) | ( n171 & ~n472 ) | ( n466 & ~n472 ) ;
  assign n474 = ~n467 & n473 ;
  assign n475 = ( ~n456 & n459 ) | ( ~n456 & n474 ) | ( n459 & n474 ) ;
  assign n476 = n197 | n421 ;
  assign n477 = ~n336 & n476 ;
  assign n478 = ( ~n20 & n203 ) | ( ~n20 & n413 ) | ( n203 & n413 ) ;
  assign n479 = ( n198 & n435 ) | ( n198 & n478 ) | ( n435 & n478 ) ;
  assign n480 = n477 | n479 ;
  buffer buf_n481( .i (n480), .o (n481) );
  assign n482 = ~n170 & n177 ;
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  assign n485 = ~n481 & n484 ;
  assign n486 = n475 | n485 ;
  buffer buf_n487( .i (n486), .o (n487) );
  assign n489 = n445 & ~n487 ;
  assign n490 = n283 & ~n489 ;
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n77( .i (x9), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  assign n492 = n178 | n470 ;
  assign n493 = ( n467 & n471 ) | ( n467 & n492 ) | ( n471 & n492 ) ;
  assign n494 = n83 & n493 ;
  buffer buf_n495( .i (n177), .o (n495) );
  assign n496 = ( ~n199 & n205 ) | ( ~n199 & n495 ) | ( n205 & n495 ) ;
  assign n497 = n334 | n496 ;
  assign n498 = ~n172 & n250 ;
  assign n499 = ( n172 & ~n250 ) | ( n172 & n433 ) | ( ~n250 & n433 ) ;
  assign n500 = ( n497 & n498 ) | ( n497 & ~n499 ) | ( n498 & ~n499 ) ;
  assign n501 = ( n252 & ~n494 ) | ( n252 & n500 ) | ( ~n494 & n500 ) ;
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n440( .i (n439), .o (n440) );
  assign n512 = ~n437 & n440 ;
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n66( .i (x7), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  assign n514 = n69 & n123 ;
  buffer buf_n515( .i (n514), .o (n515) );
  assign n516 = n483 & n515 ;
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  assign n517 = ~n186 & n193 ;
  assign n518 = ( n406 & n464 ) | ( n406 & n517 ) | ( n464 & n517 ) ;
  assign n519 = n516 & ~n518 ;
  assign n520 = ~n513 & n519 ;
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n50( .i (x5), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  assign n504 = n52 & ~n79 ;
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n187( .i (n186), .o (n187) );
  assign n508 = ~n179 & n187 ;
  assign n509 = ( n56 & n507 ) | ( n56 & ~n508 ) | ( n507 & ~n508 ) ;
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  assign n523 = n511 | n521 ;
  assign n524 = ( n503 & n522 ) | ( n503 & n523 ) | ( n522 & n523 ) ;
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n525( .i (n168), .o (n525) );
  assign n526 = n52 & n525 ;
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  assign n529 = n463 & n527 ;
  assign n530 = ( n515 & n528 ) | ( n515 & ~n529 ) | ( n528 & ~n529 ) ;
  assign n531 = n172 & n416 ;
  assign n532 = n530 & ~n531 ;
  assign n533 = ~n457 & n532 ;
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  assign n537 = n524 | n536 ;
  assign n538 = n491 & n537 ;
  assign n539 = x27 | x28 ;
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n88( .i (x10), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  assign n543 = n68 & n90 ;
  assign n544 = n542 & n543 ;
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  assign n553 = ~n238 & n311 ;
  assign n554 = n507 & n553 ;
  assign n555 = ( n123 & n363 ) | ( n123 & n375 ) | ( n363 & n375 ) ;
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  assign n559 = n52 & ~n99 ;
  assign n560 = ( n53 & n368 ) | ( n53 & n559 ) | ( n368 & n559 ) ;
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n562( .i (n150), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  assign n564 = n141 | n563 ;
  buffer buf_n565( .i (n564), .o (n565) );
  assign n568 = n69 & ~n100 ;
  assign n569 = ( n70 & ~n565 ) | ( n70 & n568 ) | ( ~n565 & n568 ) ;
  buffer buf_n58( .i (x6), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  assign n570 = n62 & ~n237 ;
  assign n571 = ( ~n561 & n569 ) | ( ~n561 & n570 ) | ( n569 & n570 ) ;
  assign n572 = n556 & ~n561 ;
  assign n573 = ~n571 & n572 ;
  assign n574 = ( n554 & n558 ) | ( n554 & ~n573 ) | ( n558 & ~n573 ) ;
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  assign n575 = ~n47 & n95 ;
  assign n576 = n69 & n142 ;
  assign n577 = ( n299 & ~n357 ) | ( n299 & n576 ) | ( ~n357 & n576 ) ;
  assign n578 = n98 & ~n121 ;
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  assign n581 = ( n237 & n505 ) | ( n237 & n580 ) | ( n505 & n580 ) ;
  buffer buf_n73( .i (x8), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  assign n582 = n75 & ~n141 ;
  assign n583 = n579 & ~n582 ;
  buffer buf_n584( .i (n583), .o (n584) );
  assign n585 = ( n577 & n581 ) | ( n577 & ~n584 ) | ( n581 & ~n584 ) ;
  assign n586 = ~n45 & n114 ;
  assign n587 = ( ~n230 & n585 ) | ( ~n230 & n586 ) | ( n585 & n586 ) ;
  assign n588 = n95 & n587 ;
  assign n589 = ( n574 & n575 ) | ( n574 & n588 ) | ( n575 & n588 ) ;
  buffer buf_n590( .i (n589), .o (n590) );
  assign n591 = n550 | n590 ;
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n594( .i (n171), .o (n594) );
  assign n595 = n23 & ~n594 ;
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  assign n598 = n187 & n433 ;
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  assign n601 = n295 & n599 ;
  assign n602 = ( n597 & n600 ) | ( n597 & n601 ) | ( n600 & n601 ) ;
  assign n603 = n267 | n602 ;
  assign n604 = n488 | n603 ;
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  assign n605 = n101 | n505 ;
  assign n606 = ~n290 & n605 ;
  buffer buf_n71( .i (n70), .o (n71) );
  assign n607 = n71 | n566 ;
  assign n608 = ( ~n567 & n606 ) | ( ~n567 & n607 ) | ( n606 & n607 ) ;
  assign n609 = ~n55 & n114 ;
  assign n610 = n54 | n70 ;
  buffer buf_n611( .i (n113), .o (n611) );
  assign n612 = ~n610 & n611 ;
  assign n613 = ( n378 & n609 ) | ( n378 & n612 ) | ( n609 & n612 ) ;
  buffer buf_n614( .i (n611), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  assign n616 = ( ~n608 & n613 ) | ( ~n608 & n615 ) | ( n613 & n615 ) ;
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  assign n619 = n590 & ~n618 ;
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  assign n620 = n64 & n291 ;
  assign n621 = n280 & n620 ;
  buffer buf_n622( .i (n621), .o (n622) );
  assign n623 = n617 & ~n622 ;
  assign n624 = n590 & ~n623 ;
  assign n625 = ( n604 & n619 ) | ( n604 & n624 ) | ( n619 & n624 ) ;
  assign n626 = n552 | n625 ;
  assign n627 = ( n538 & n593 ) | ( n538 & n626 ) | ( n593 & n626 ) ;
  buffer buf_n107( .i (n106), .o (n107) );
  assign n628 = n136 & n311 ;
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  assign n633 = n86 & ~n106 ;
  assign n634 = ( n107 & n632 ) | ( n107 & ~n633 ) | ( n632 & ~n633 ) ;
  assign n635 = ~n187 & n483 ;
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  assign n638 = n324 & n637 ;
  assign n639 = ~n81 & n193 ;
  buffer buf_n640( .i (n639), .o (n640) );
  assign n641 = n481 & ~n640 ;
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  assign n644 = n638 & ~n643 ;
  assign n645 = n228 & n376 ;
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  assign n646 = n4 & ~n42 ;
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  assign n649 = ~n645 & n648 ;
  buffer buf_n650( .i (n649), .o (n650) );
  assign n651 = ( n104 & n629 ) | ( n104 & ~n650 ) | ( n629 & ~n650 ) ;
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  assign n654 = n118 | n652 ;
  assign n655 = ( ~n644 & n653 ) | ( ~n644 & n654 ) | ( n653 & n654 ) ;
  assign n656 = n634 & ~n655 ;
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  assign n659 = n38 & ~n319 ;
  assign n660 = n348 & ~n659 ;
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  assign n661 = ( ~n264 & n266 ) | ( ~n264 & n419 ) | ( n266 & n419 ) ;
  assign n662 = n325 & n661 ;
  assign n663 = n37 | n117 ;
  assign n664 = ( n106 & n315 ) | ( n106 & n663 ) | ( n315 & n663 ) ;
  assign n665 = ~n662 & n664 ;
  assign n666 = ~n660 & n665 ;
  buffer buf_n6( .i (x1), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  assign n667 = n16 & n382 ;
  buffer buf_n668( .i (n667), .o (n668) );
  assign n669 = ~n666 & n668 ;
  buffer buf_n670( .i (n669), .o (n670) );
  assign n671 = n245 | n491 ;
  buffer buf_n672( .i (n671), .o (n672) );
  assign y0 = n288 ;
  assign y1 = n309 ;
  assign y2 = n393 ;
  assign y3 = n627 ;
  assign y4 = n658 ;
  assign y5 = n670 ;
  assign y6 = n672 ;
endmodule
