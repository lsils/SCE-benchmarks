module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 ;
  assign n129 = x101 & x115 ;
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  assign n139 = x44 | x94 ;
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  assign n147 = x28 | x39 ;
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  assign n151 = x11 | x87 ;
  buffer buf_n152( .i (n151), .o (n152) );
  assign n153 = x49 & x64 ;
  buffer buf_n154( .i (n153), .o (n154) );
  assign n155 = ( n148 & n152 ) | ( n148 & n154 ) | ( n152 & n154 ) ;
  buffer buf_n156( .i (n155), .o (n156) );
  assign n161 = ( ~n148 & n152 ) | ( ~n148 & n154 ) | ( n152 & n154 ) ;
  buffer buf_n162( .i (n161), .o (n162) );
  assign n163 = ( n150 & ~n156 ) | ( n150 & n162 ) | ( ~n156 & n162 ) ;
  buffer buf_n164( .i (n163), .o (n164) );
  assign n165 = x53 & x93 ;
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = x7 & x89 ;
  buffer buf_n170( .i (n169), .o (n170) );
  assign n171 = x41 | x111 ;
  buffer buf_n172( .i (n171), .o (n172) );
  assign n173 = ( n166 & n170 ) | ( n166 & n172 ) | ( n170 & n172 ) ;
  buffer buf_n174( .i (n173), .o (n174) );
  assign n179 = ( ~n166 & n170 ) | ( ~n166 & n172 ) | ( n170 & n172 ) ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = ( n168 & ~n174 ) | ( n168 & n180 ) | ( ~n174 & n180 ) ;
  buffer buf_n182( .i (n181), .o (n182) );
  assign n183 = ( n144 & n164 ) | ( n144 & n182 ) | ( n164 & n182 ) ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n187 = ( ~n144 & n164 ) | ( ~n144 & n182 ) | ( n164 & n182 ) ;
  buffer buf_n188( .i (n187), .o (n188) );
  assign n189 = ( n146 & ~n184 ) | ( n146 & n188 ) | ( ~n184 & n188 ) ;
  buffer buf_n190( .i (n189), .o (n190) );
  assign n191 = n138 & n190 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = n138 | n190 ;
  buffer buf_n194( .i (n193), .o (n194) );
  assign n195 = ~n192 & n194 ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n197 = x59 & x124 ;
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  assign n207 = x3 | x27 ;
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n215 = x8 | x18 ;
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  assign n219 = x102 | x112 ;
  buffer buf_n220( .i (n219), .o (n220) );
  assign n221 = x114 & x119 ;
  buffer buf_n222( .i (n221), .o (n222) );
  assign n223 = ( ~n216 & n220 ) | ( ~n216 & n222 ) | ( n220 & n222 ) ;
  buffer buf_n224( .i (n223), .o (n224) );
  assign n225 = ( n216 & n220 ) | ( n216 & n222 ) | ( n220 & n222 ) ;
  buffer buf_n226( .i (n225), .o (n226) );
  assign n231 = ( n218 & n224 ) | ( n218 & ~n226 ) | ( n224 & ~n226 ) ;
  buffer buf_n232( .i (n231), .o (n232) );
  assign n233 = x5 & x80 ;
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  assign n237 = x29 & x69 ;
  buffer buf_n238( .i (n237), .o (n238) );
  assign n239 = x19 | x42 ;
  buffer buf_n240( .i (n239), .o (n240) );
  assign n241 = ( n234 & n238 ) | ( n234 & n240 ) | ( n238 & n240 ) ;
  buffer buf_n242( .i (n241), .o (n242) );
  assign n247 = ( ~n234 & n238 ) | ( ~n234 & n240 ) | ( n238 & n240 ) ;
  buffer buf_n248( .i (n247), .o (n248) );
  assign n249 = ( n236 & ~n242 ) | ( n236 & n248 ) | ( ~n242 & n248 ) ;
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = ( n212 & n232 ) | ( n212 & n250 ) | ( n232 & n250 ) ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n255 = ( ~n212 & n232 ) | ( ~n212 & n250 ) | ( n232 & n250 ) ;
  buffer buf_n256( .i (n255), .o (n256) );
  assign n257 = ( n214 & ~n252 ) | ( n214 & n256 ) | ( ~n252 & n256 ) ;
  buffer buf_n258( .i (n257), .o (n258) );
  assign n259 = n206 & n258 ;
  buffer buf_n260( .i (n259), .o (n260) );
  assign n261 = n206 | n258 ;
  buffer buf_n262( .i (n261), .o (n262) );
  assign n263 = ~n260 & n262 ;
  buffer buf_n264( .i (n263), .o (n264) );
  assign n265 = n196 & n264 ;
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  assign n270 = n196 | n264 ;
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  assign n273 = ~n267 & n272 ;
  buffer buf_n274( .i (n273), .o (n274) );
  assign n275 = x26 & x108 ;
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  assign n285 = x73 | x96 ;
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  assign n293 = x36 | x82 ;
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  assign n297 = x48 | x76 ;
  buffer buf_n298( .i (n297), .o (n298) );
  assign n299 = x58 & x66 ;
  buffer buf_n300( .i (n299), .o (n300) );
  assign n301 = ( n294 & n298 ) | ( n294 & n300 ) | ( n298 & n300 ) ;
  buffer buf_n302( .i (n301), .o (n302) );
  assign n307 = ( ~n294 & n298 ) | ( ~n294 & n300 ) | ( n298 & n300 ) ;
  buffer buf_n308( .i (n307), .o (n308) );
  assign n309 = ( n296 & ~n302 ) | ( n296 & n308 ) | ( ~n302 & n308 ) ;
  buffer buf_n310( .i (n309), .o (n310) );
  assign n311 = x75 & x117 ;
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  assign n315 = x62 & x67 ;
  buffer buf_n316( .i (n315), .o (n316) );
  assign n317 = x14 | x50 ;
  buffer buf_n318( .i (n317), .o (n318) );
  assign n319 = ( n312 & n316 ) | ( n312 & n318 ) | ( n316 & n318 ) ;
  buffer buf_n320( .i (n319), .o (n320) );
  assign n325 = ( ~n312 & n316 ) | ( ~n312 & n318 ) | ( n316 & n318 ) ;
  buffer buf_n326( .i (n325), .o (n326) );
  assign n327 = ( n314 & ~n320 ) | ( n314 & n326 ) | ( ~n320 & n326 ) ;
  buffer buf_n328( .i (n327), .o (n328) );
  assign n329 = ( n290 & n310 ) | ( n290 & n328 ) | ( n310 & n328 ) ;
  buffer buf_n330( .i (n329), .o (n330) );
  assign n333 = ( ~n290 & n310 ) | ( ~n290 & n328 ) | ( n310 & n328 ) ;
  buffer buf_n334( .i (n333), .o (n334) );
  assign n335 = ( n292 & ~n330 ) | ( n292 & n334 ) | ( ~n330 & n334 ) ;
  buffer buf_n336( .i (n335), .o (n336) );
  assign n337 = n284 & n336 ;
  buffer buf_n338( .i (n337), .o (n338) );
  assign n339 = n284 | n336 ;
  buffer buf_n340( .i (n339), .o (n340) );
  assign n341 = ~n338 & n340 ;
  buffer buf_n342( .i (n341), .o (n342) );
  assign n343 = x23 & x55 ;
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  assign n353 = x33 | x90 ;
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  assign n361 = x60 | x110 ;
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  assign n365 = x43 | x68 ;
  buffer buf_n366( .i (n365), .o (n366) );
  assign n367 = x30 & x126 ;
  buffer buf_n368( .i (n367), .o (n368) );
  assign n369 = ( n362 & n366 ) | ( n362 & n368 ) | ( n366 & n368 ) ;
  buffer buf_n370( .i (n369), .o (n370) );
  assign n375 = ( ~n362 & n366 ) | ( ~n362 & n368 ) | ( n366 & n368 ) ;
  buffer buf_n376( .i (n375), .o (n376) );
  assign n377 = ( n364 & ~n370 ) | ( n364 & n376 ) | ( ~n370 & n376 ) ;
  buffer buf_n378( .i (n377), .o (n378) );
  assign n379 = x63 & x71 ;
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  assign n383 = x16 & x121 ;
  buffer buf_n384( .i (n383), .o (n384) );
  assign n385 = x38 | x77 ;
  buffer buf_n386( .i (n385), .o (n386) );
  assign n387 = ( n380 & n384 ) | ( n380 & n386 ) | ( n384 & n386 ) ;
  buffer buf_n388( .i (n387), .o (n388) );
  assign n393 = ( ~n380 & n384 ) | ( ~n380 & n386 ) | ( n384 & n386 ) ;
  buffer buf_n394( .i (n393), .o (n394) );
  assign n395 = ( n382 & ~n388 ) | ( n382 & n394 ) | ( ~n388 & n394 ) ;
  buffer buf_n396( .i (n395), .o (n396) );
  assign n397 = ( n358 & n378 ) | ( n358 & n396 ) | ( n378 & n396 ) ;
  buffer buf_n398( .i (n397), .o (n398) );
  assign n401 = ( ~n358 & n378 ) | ( ~n358 & n396 ) | ( n378 & n396 ) ;
  buffer buf_n402( .i (n401), .o (n402) );
  assign n403 = ( n360 & ~n398 ) | ( n360 & n402 ) | ( ~n398 & n402 ) ;
  buffer buf_n404( .i (n403), .o (n404) );
  assign n405 = n352 & n404 ;
  buffer buf_n406( .i (n405), .o (n406) );
  assign n407 = n352 | n404 ;
  buffer buf_n408( .i (n407), .o (n408) );
  assign n409 = ~n406 & n408 ;
  buffer buf_n410( .i (n409), .o (n410) );
  assign n411 = n342 & n410 ;
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  assign n416 = n342 | n410 ;
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  assign n419 = ~n413 & n418 ;
  buffer buf_n420( .i (n419), .o (n420) );
  assign n421 = n274 & n420 ;
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  assign n427 = ( n160 & n178 ) | ( n160 & n184 ) | ( n178 & n184 ) ;
  buffer buf_n428( .i (n427), .o (n428) );
  assign n433 = ( n160 & n178 ) | ( n160 & ~n184 ) | ( n178 & ~n184 ) ;
  buffer buf_n434( .i (n433), .o (n434) );
  assign n435 = ( n186 & ~n428 ) | ( n186 & n434 ) | ( ~n428 & n434 ) ;
  buffer buf_n436( .i (n435), .o (n436) );
  assign n437 = n192 & n436 ;
  buffer buf_n438( .i (n437), .o (n438) );
  assign n439 = n192 | n436 ;
  buffer buf_n440( .i (n439), .o (n440) );
  assign n441 = ~n438 & n440 ;
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  assign n443 = ( n230 & n246 ) | ( n230 & n252 ) | ( n246 & n252 ) ;
  buffer buf_n444( .i (n443), .o (n444) );
  assign n449 = ( n230 & n246 ) | ( n230 & ~n252 ) | ( n246 & ~n252 ) ;
  buffer buf_n450( .i (n449), .o (n450) );
  assign n451 = ( n254 & ~n444 ) | ( n254 & n450 ) | ( ~n444 & n450 ) ;
  buffer buf_n452( .i (n451), .o (n452) );
  assign n453 = n260 & n452 ;
  buffer buf_n454( .i (n453), .o (n454) );
  assign n455 = n260 | n452 ;
  buffer buf_n456( .i (n455), .o (n456) );
  assign n457 = ~n454 & n456 ;
  buffer buf_n458( .i (n457), .o (n458) );
  assign n459 = n442 & n458 ;
  assign n460 = n442 | n458 ;
  assign n461 = ~n459 & n460 ;
  buffer buf_n462( .i (n461), .o (n462) );
  assign n463 = n269 & n462 ;
  assign n464 = n269 | n462 ;
  assign n465 = ~n463 & n464 ;
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  assign n467 = ( n306 & n324 ) | ( n306 & n330 ) | ( n324 & n330 ) ;
  buffer buf_n468( .i (n467), .o (n468) );
  assign n473 = ( n306 & n324 ) | ( n306 & ~n330 ) | ( n324 & ~n330 ) ;
  buffer buf_n474( .i (n473), .o (n474) );
  assign n475 = ( n332 & ~n468 ) | ( n332 & n474 ) | ( ~n468 & n474 ) ;
  buffer buf_n476( .i (n475), .o (n476) );
  assign n477 = n338 & n476 ;
  buffer buf_n478( .i (n477), .o (n478) );
  assign n479 = n338 | n476 ;
  buffer buf_n480( .i (n479), .o (n480) );
  assign n481 = ~n478 & n480 ;
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  assign n483 = ( n374 & n392 ) | ( n374 & n398 ) | ( n392 & n398 ) ;
  buffer buf_n484( .i (n483), .o (n484) );
  assign n489 = ( n374 & n392 ) | ( n374 & ~n398 ) | ( n392 & ~n398 ) ;
  buffer buf_n490( .i (n489), .o (n490) );
  assign n491 = ( n400 & ~n484 ) | ( n400 & n490 ) | ( ~n484 & n490 ) ;
  buffer buf_n492( .i (n491), .o (n492) );
  assign n493 = n406 & n492 ;
  buffer buf_n494( .i (n493), .o (n494) );
  assign n495 = n406 | n492 ;
  buffer buf_n496( .i (n495), .o (n496) );
  assign n497 = ~n494 & n496 ;
  buffer buf_n498( .i (n497), .o (n498) );
  assign n499 = n482 & n498 ;
  assign n500 = n482 | n498 ;
  assign n501 = ~n499 & n500 ;
  buffer buf_n502( .i (n501), .o (n502) );
  assign n503 = n415 & n502 ;
  assign n504 = n415 | n502 ;
  assign n505 = ~n503 & n504 ;
  buffer buf_n506( .i (n505), .o (n506) );
  assign n507 = n466 & n506 ;
  assign n508 = n466 | n506 ;
  assign n509 = ~n507 & n508 ;
  buffer buf_n510( .i (n509), .o (n510) );
  assign n511 = n426 & n510 ;
  assign n512 = n426 | n510 ;
  assign n513 = ~n511 & n512 ;
  buffer buf_n514( .i (n513), .o (n514) );
  assign n515 = n274 | n420 ;
  buffer buf_n516( .i (n515), .o (n516) );
  assign n517 = ~n422 & n516 ;
  buffer buf_n518( .i (n517), .o (n518) );
  assign n519 = x13 & x56 ;
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  assign n529 = x20 | x24 ;
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  assign n537 = x118 & x120 ;
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  assign n541 = x103 & x123 ;
  buffer buf_n542( .i (n541), .o (n542) );
  assign n543 = x51 | x79 ;
  buffer buf_n544( .i (n543), .o (n544) );
  assign n545 = ( n538 & n542 ) | ( n538 & n544 ) | ( n542 & n544 ) ;
  buffer buf_n546( .i (n545), .o (n546) );
  assign n551 = ( ~n538 & n542 ) | ( ~n538 & n544 ) | ( n542 & n544 ) ;
  buffer buf_n552( .i (n551), .o (n552) );
  assign n553 = ( n540 & ~n546 ) | ( n540 & n552 ) | ( ~n546 & n552 ) ;
  buffer buf_n554( .i (n553), .o (n554) );
  assign n555 = x35 | x107 ;
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  assign n559 = x37 | x40 ;
  buffer buf_n560( .i (n559), .o (n560) );
  assign n561 = x0 & x127 ;
  buffer buf_n562( .i (n561), .o (n562) );
  assign n563 = ( n556 & n560 ) | ( n556 & n562 ) | ( n560 & n562 ) ;
  buffer buf_n564( .i (n563), .o (n564) );
  assign n569 = ( ~n556 & n560 ) | ( ~n556 & n562 ) | ( n560 & n562 ) ;
  buffer buf_n570( .i (n569), .o (n570) );
  assign n571 = ( n558 & ~n564 ) | ( n558 & n570 ) | ( ~n564 & n570 ) ;
  buffer buf_n572( .i (n571), .o (n572) );
  assign n573 = ( n534 & n554 ) | ( n534 & n572 ) | ( n554 & n572 ) ;
  buffer buf_n574( .i (n573), .o (n574) );
  assign n577 = ( ~n534 & n554 ) | ( ~n534 & n572 ) | ( n554 & n572 ) ;
  buffer buf_n578( .i (n577), .o (n578) );
  assign n579 = ( n536 & ~n574 ) | ( n536 & n578 ) | ( ~n574 & n578 ) ;
  buffer buf_n580( .i (n579), .o (n580) );
  assign n581 = n528 & n580 ;
  buffer buf_n582( .i (n581), .o (n582) );
  assign n583 = n528 | n580 ;
  buffer buf_n584( .i (n583), .o (n584) );
  assign n585 = ~n582 & n584 ;
  buffer buf_n586( .i (n585), .o (n586) );
  assign n587 = x97 & x116 ;
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  assign n597 = x4 | x86 ;
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  assign n605 = x72 | x100 ;
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  assign n609 = x1 | x10 ;
  buffer buf_n610( .i (n609), .o (n610) );
  assign n611 = x9 & x61 ;
  buffer buf_n612( .i (n611), .o (n612) );
  assign n613 = ( n606 & n610 ) | ( n606 & n612 ) | ( n610 & n612 ) ;
  buffer buf_n614( .i (n613), .o (n614) );
  assign n619 = ( ~n606 & n610 ) | ( ~n606 & n612 ) | ( n610 & n612 ) ;
  buffer buf_n620( .i (n619), .o (n620) );
  assign n621 = ( n608 & ~n614 ) | ( n608 & n620 ) | ( ~n614 & n620 ) ;
  buffer buf_n622( .i (n621), .o (n622) );
  assign n623 = x21 & x113 ;
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  assign n627 = x2 & x70 ;
  buffer buf_n628( .i (n627), .o (n628) );
  assign n629 = x22 | x122 ;
  buffer buf_n630( .i (n629), .o (n630) );
  assign n631 = ( n624 & n628 ) | ( n624 & n630 ) | ( n628 & n630 ) ;
  buffer buf_n632( .i (n631), .o (n632) );
  assign n637 = ( ~n624 & n628 ) | ( ~n624 & n630 ) | ( n628 & n630 ) ;
  buffer buf_n638( .i (n637), .o (n638) );
  assign n639 = ( n626 & ~n632 ) | ( n626 & n638 ) | ( ~n632 & n638 ) ;
  buffer buf_n640( .i (n639), .o (n640) );
  assign n641 = ( n602 & n622 ) | ( n602 & n640 ) | ( n622 & n640 ) ;
  buffer buf_n642( .i (n641), .o (n642) );
  assign n645 = ( ~n602 & n622 ) | ( ~n602 & n640 ) | ( n622 & n640 ) ;
  buffer buf_n646( .i (n645), .o (n646) );
  assign n647 = ( n604 & ~n642 ) | ( n604 & n646 ) | ( ~n642 & n646 ) ;
  buffer buf_n648( .i (n647), .o (n648) );
  assign n649 = n596 & n648 ;
  buffer buf_n650( .i (n649), .o (n650) );
  assign n651 = n596 | n648 ;
  buffer buf_n652( .i (n651), .o (n652) );
  assign n653 = ~n650 & n652 ;
  buffer buf_n654( .i (n653), .o (n654) );
  assign n655 = n586 & n654 ;
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  assign n660 = n586 | n654 ;
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  assign n663 = ~n657 & n662 ;
  buffer buf_n664( .i (n663), .o (n664) );
  assign n665 = x34 & x78 ;
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  assign n675 = x31 | x74 ;
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  assign n683 = x57 | x81 ;
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  assign n687 = x52 | x88 ;
  buffer buf_n688( .i (n687), .o (n688) );
  assign n689 = x15 & x91 ;
  buffer buf_n690( .i (n689), .o (n690) );
  assign n691 = ( n684 & n688 ) | ( n684 & n690 ) | ( n688 & n690 ) ;
  buffer buf_n692( .i (n691), .o (n692) );
  assign n697 = ( ~n684 & n688 ) | ( ~n684 & n690 ) | ( n688 & n690 ) ;
  buffer buf_n698( .i (n697), .o (n698) );
  assign n699 = ( n686 & ~n692 ) | ( n686 & n698 ) | ( ~n692 & n698 ) ;
  buffer buf_n700( .i (n699), .o (n700) );
  assign n701 = x46 & x104 ;
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  assign n705 = x17 & x84 ;
  buffer buf_n706( .i (n705), .o (n706) );
  assign n707 = x47 | x92 ;
  buffer buf_n708( .i (n707), .o (n708) );
  assign n709 = ( n702 & n706 ) | ( n702 & n708 ) | ( n706 & n708 ) ;
  buffer buf_n710( .i (n709), .o (n710) );
  assign n715 = ( ~n702 & n706 ) | ( ~n702 & n708 ) | ( n706 & n708 ) ;
  buffer buf_n716( .i (n715), .o (n716) );
  assign n717 = ( n704 & ~n710 ) | ( n704 & n716 ) | ( ~n710 & n716 ) ;
  buffer buf_n718( .i (n717), .o (n718) );
  assign n719 = ( n680 & n700 ) | ( n680 & n718 ) | ( n700 & n718 ) ;
  buffer buf_n720( .i (n719), .o (n720) );
  assign n723 = ( ~n680 & n700 ) | ( ~n680 & n718 ) | ( n700 & n718 ) ;
  buffer buf_n724( .i (n723), .o (n724) );
  assign n725 = ( n682 & ~n720 ) | ( n682 & n724 ) | ( ~n720 & n724 ) ;
  buffer buf_n726( .i (n725), .o (n726) );
  assign n727 = n674 & n726 ;
  buffer buf_n728( .i (n727), .o (n728) );
  assign n729 = n674 | n726 ;
  buffer buf_n730( .i (n729), .o (n730) );
  assign n731 = ~n728 & n730 ;
  buffer buf_n732( .i (n731), .o (n732) );
  assign n733 = x85 & x125 ;
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  assign n743 = x25 | x54 ;
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  assign n751 = x45 & x109 ;
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  assign n755 = x6 & x98 ;
  buffer buf_n756( .i (n755), .o (n756) );
  assign n757 = x12 | x32 ;
  buffer buf_n758( .i (n757), .o (n758) );
  assign n759 = ( n752 & n756 ) | ( n752 & n758 ) | ( n756 & n758 ) ;
  buffer buf_n760( .i (n759), .o (n760) );
  assign n765 = ( ~n752 & n756 ) | ( ~n752 & n758 ) | ( n756 & n758 ) ;
  buffer buf_n766( .i (n765), .o (n766) );
  assign n767 = ( n754 & ~n760 ) | ( n754 & n766 ) | ( ~n760 & n766 ) ;
  buffer buf_n768( .i (n767), .o (n768) );
  assign n769 = x65 | x105 ;
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  assign n773 = x83 | x95 ;
  buffer buf_n774( .i (n773), .o (n774) );
  assign n775 = x99 & x106 ;
  buffer buf_n776( .i (n775), .o (n776) );
  assign n777 = ( n770 & n774 ) | ( n770 & n776 ) | ( n774 & n776 ) ;
  buffer buf_n778( .i (n777), .o (n778) );
  assign n783 = ( ~n770 & n774 ) | ( ~n770 & n776 ) | ( n774 & n776 ) ;
  buffer buf_n784( .i (n783), .o (n784) );
  assign n785 = ( n772 & ~n778 ) | ( n772 & n784 ) | ( ~n778 & n784 ) ;
  buffer buf_n786( .i (n785), .o (n786) );
  assign n787 = ( n748 & n768 ) | ( n748 & n786 ) | ( n768 & n786 ) ;
  buffer buf_n788( .i (n787), .o (n788) );
  assign n791 = ( ~n748 & n768 ) | ( ~n748 & n786 ) | ( n768 & n786 ) ;
  buffer buf_n792( .i (n791), .o (n792) );
  assign n793 = ( n750 & ~n788 ) | ( n750 & n792 ) | ( ~n788 & n792 ) ;
  buffer buf_n794( .i (n793), .o (n794) );
  assign n795 = n742 & n794 ;
  buffer buf_n796( .i (n795), .o (n796) );
  assign n797 = n742 | n794 ;
  buffer buf_n798( .i (n797), .o (n798) );
  assign n799 = ~n796 & n798 ;
  buffer buf_n800( .i (n799), .o (n800) );
  assign n801 = n732 | n800 ;
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  assign n804 = n732 & n800 ;
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  assign n809 = n803 & ~n806 ;
  buffer buf_n810( .i (n809), .o (n810) );
  assign n811 = n664 & n810 ;
  buffer buf_n812( .i (n811), .o (n812) );
  assign n817 = n664 | n810 ;
  buffer buf_n818( .i (n817), .o (n818) );
  assign n819 = ~n812 & n818 ;
  buffer buf_n820( .i (n819), .o (n820) );
  assign n821 = n518 & n820 ;
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  assign n829 = ( n550 & n568 ) | ( n550 & n574 ) | ( n568 & n574 ) ;
  buffer buf_n830( .i (n829), .o (n830) );
  assign n835 = ( n550 & n568 ) | ( n550 & ~n574 ) | ( n568 & ~n574 ) ;
  buffer buf_n836( .i (n835), .o (n836) );
  assign n837 = ( n576 & ~n830 ) | ( n576 & n836 ) | ( ~n830 & n836 ) ;
  buffer buf_n838( .i (n837), .o (n838) );
  assign n839 = n582 | n838 ;
  buffer buf_n840( .i (n839), .o (n840) );
  assign n841 = n582 & n838 ;
  buffer buf_n842( .i (n841), .o (n842) );
  assign n843 = n840 & ~n842 ;
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  assign n845 = ( n618 & n636 ) | ( n618 & n642 ) | ( n636 & n642 ) ;
  buffer buf_n846( .i (n845), .o (n846) );
  assign n851 = ( n618 & n636 ) | ( n618 & ~n642 ) | ( n636 & ~n642 ) ;
  buffer buf_n852( .i (n851), .o (n852) );
  assign n853 = ( n644 & ~n846 ) | ( n644 & n852 ) | ( ~n846 & n852 ) ;
  buffer buf_n854( .i (n853), .o (n854) );
  assign n855 = n650 & n854 ;
  buffer buf_n856( .i (n855), .o (n856) );
  assign n857 = n650 | n854 ;
  buffer buf_n858( .i (n857), .o (n858) );
  assign n859 = ~n856 & n858 ;
  buffer buf_n860( .i (n859), .o (n860) );
  assign n861 = n844 & n860 ;
  assign n862 = n844 | n860 ;
  assign n863 = ~n861 & n862 ;
  buffer buf_n864( .i (n863), .o (n864) );
  assign n865 = n659 & n864 ;
  assign n866 = n659 | n864 ;
  assign n867 = ~n865 & n866 ;
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  assign n869 = ( n764 & n782 ) | ( n764 & n788 ) | ( n782 & n788 ) ;
  buffer buf_n870( .i (n869), .o (n870) );
  assign n875 = ( n764 & n782 ) | ( n764 & ~n788 ) | ( n782 & ~n788 ) ;
  buffer buf_n876( .i (n875), .o (n876) );
  assign n877 = ( n790 & ~n870 ) | ( n790 & n876 ) | ( ~n870 & n876 ) ;
  buffer buf_n878( .i (n877), .o (n878) );
  assign n879 = n796 & n878 ;
  buffer buf_n880( .i (n879), .o (n880) );
  assign n881 = n796 | n878 ;
  buffer buf_n882( .i (n881), .o (n882) );
  assign n883 = ~n880 & n882 ;
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  assign n885 = ( n696 & n714 ) | ( n696 & n720 ) | ( n714 & n720 ) ;
  buffer buf_n886( .i (n885), .o (n886) );
  assign n891 = ( n696 & n714 ) | ( n696 & ~n720 ) | ( n714 & ~n720 ) ;
  buffer buf_n892( .i (n891), .o (n892) );
  assign n893 = ( n722 & ~n886 ) | ( n722 & n892 ) | ( ~n886 & n892 ) ;
  buffer buf_n894( .i (n893), .o (n894) );
  assign n895 = n728 & n894 ;
  buffer buf_n896( .i (n895), .o (n896) );
  assign n897 = n728 | n894 ;
  buffer buf_n898( .i (n897), .o (n898) );
  assign n899 = ~n896 & n898 ;
  buffer buf_n900( .i (n899), .o (n900) );
  assign n901 = n884 & n900 ;
  assign n902 = n884 | n900 ;
  assign n903 = ~n901 & n902 ;
  buffer buf_n904( .i (n903), .o (n904) );
  assign n905 = n808 & n904 ;
  assign n906 = n808 | n904 ;
  assign n907 = ~n905 & n906 ;
  buffer buf_n908( .i (n907), .o (n908) );
  assign n909 = n868 & n908 ;
  assign n910 = n868 | n908 ;
  assign n911 = ~n909 & n910 ;
  buffer buf_n912( .i (n911), .o (n912) );
  assign n913 = n816 & n912 ;
  assign n914 = n816 | n912 ;
  assign n915 = ~n913 & n914 ;
  buffer buf_n916( .i (n915), .o (n916) );
  assign n917 = ( n514 & n825 ) | ( n514 & n916 ) | ( n825 & n916 ) ;
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  assign n922 = ( n813 & n868 ) | ( n813 & n908 ) | ( n868 & n908 ) ;
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  assign n927 = ( n656 & n844 ) | ( n656 & n860 ) | ( n844 & n860 ) ;
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  assign n932 = n834 & n842 ;
  buffer buf_n933( .i (n932), .o (n933) );
  assign n938 = n834 | n842 ;
  buffer buf_n939( .i (n938), .o (n939) );
  assign n940 = ~n933 & n939 ;
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  assign n942 = n850 & n856 ;
  buffer buf_n943( .i (n942), .o (n943) );
  assign n948 = n850 | n856 ;
  buffer buf_n949( .i (n948), .o (n949) );
  assign n950 = ~n943 & n949 ;
  buffer buf_n951( .i (n950), .o (n951) );
  assign n952 = n941 & n951 ;
  assign n953 = n941 | n951 ;
  assign n954 = ~n952 & n953 ;
  buffer buf_n955( .i (n954), .o (n955) );
  assign n956 = n931 & n955 ;
  assign n957 = n931 | n955 ;
  assign n958 = ~n956 & n957 ;
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  assign n960 = n890 & n896 ;
  buffer buf_n961( .i (n960), .o (n961) );
  assign n966 = n890 | n896 ;
  buffer buf_n967( .i (n966), .o (n967) );
  assign n968 = ~n961 & n967 ;
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  assign n970 = n874 & n880 ;
  buffer buf_n971( .i (n970), .o (n971) );
  assign n976 = n874 | n880 ;
  buffer buf_n977( .i (n976), .o (n977) );
  assign n978 = ~n971 & n977 ;
  buffer buf_n979( .i (n978), .o (n979) );
  assign n980 = n969 & n979 ;
  assign n981 = n969 | n979 ;
  assign n982 = ~n980 & n981 ;
  buffer buf_n983( .i (n982), .o (n983) );
  assign n984 = ( n805 & n884 ) | ( n805 & n900 ) | ( n884 & n900 ) ;
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  assign n989 = n983 & n988 ;
  assign n990 = n983 | n988 ;
  assign n991 = ~n989 & n990 ;
  buffer buf_n992( .i (n991), .o (n992) );
  assign n993 = n959 & n992 ;
  assign n994 = n959 | n992 ;
  assign n995 = ~n993 & n994 ;
  buffer buf_n996( .i (n995), .o (n996) );
  assign n997 = n926 & n996 ;
  assign n998 = n926 | n996 ;
  assign n999 = ~n997 & n998 ;
  buffer buf_n1000( .i (n999), .o (n1000) );
  assign n1001 = ( n423 & n466 ) | ( n423 & n506 ) | ( n466 & n506 ) ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  assign n1006 = ( n266 & n442 ) | ( n266 & n458 ) | ( n442 & n458 ) ;
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  assign n1011 = n432 & n438 ;
  buffer buf_n1012( .i (n1011), .o (n1012) );
  assign n1017 = n432 | n438 ;
  buffer buf_n1018( .i (n1017), .o (n1018) );
  assign n1019 = ~n1012 & n1018 ;
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  assign n1021 = n448 & n454 ;
  buffer buf_n1022( .i (n1021), .o (n1022) );
  assign n1027 = n448 | n454 ;
  buffer buf_n1028( .i (n1027), .o (n1028) );
  assign n1029 = ~n1022 & n1028 ;
  buffer buf_n1030( .i (n1029), .o (n1030) );
  assign n1031 = n1020 & n1030 ;
  assign n1032 = n1020 | n1030 ;
  assign n1033 = ~n1031 & n1032 ;
  buffer buf_n1034( .i (n1033), .o (n1034) );
  assign n1035 = n1010 & n1034 ;
  assign n1036 = n1010 | n1034 ;
  assign n1037 = ~n1035 & n1036 ;
  buffer buf_n1038( .i (n1037), .o (n1038) );
  assign n1039 = ( n412 & n482 ) | ( n412 & n498 ) | ( n482 & n498 ) ;
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  assign n1044 = n472 & n478 ;
  buffer buf_n1045( .i (n1044), .o (n1045) );
  assign n1050 = n472 | n478 ;
  buffer buf_n1051( .i (n1050), .o (n1051) );
  assign n1052 = ~n1045 & n1051 ;
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  assign n1054 = n488 & n494 ;
  buffer buf_n1055( .i (n1054), .o (n1055) );
  assign n1060 = n488 | n494 ;
  buffer buf_n1061( .i (n1060), .o (n1061) );
  assign n1062 = ~n1055 & n1061 ;
  buffer buf_n1063( .i (n1062), .o (n1063) );
  assign n1064 = n1053 & n1063 ;
  assign n1065 = n1053 | n1063 ;
  assign n1066 = ~n1064 & n1065 ;
  buffer buf_n1067( .i (n1066), .o (n1067) );
  assign n1068 = n1043 & n1067 ;
  assign n1069 = n1043 | n1067 ;
  assign n1070 = ~n1068 & n1069 ;
  buffer buf_n1071( .i (n1070), .o (n1071) );
  assign n1072 = n1038 & n1071 ;
  assign n1073 = n1038 | n1071 ;
  assign n1074 = ~n1072 & n1073 ;
  buffer buf_n1075( .i (n1074), .o (n1075) );
  assign n1076 = n1005 & n1075 ;
  assign n1077 = n1005 | n1075 ;
  assign n1078 = ~n1076 & n1077 ;
  buffer buf_n1079( .i (n1078), .o (n1079) );
  assign n1080 = n1000 & n1079 ;
  assign n1081 = n1000 | n1079 ;
  assign n1082 = ~n1080 & n1081 ;
  buffer buf_n1083( .i (n1082), .o (n1083) );
  assign n1084 = n921 & n1083 ;
  assign n1085 = n921 | n1083 ;
  assign n1086 = ~n1084 & n1085 ;
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  assign n1090 = n514 & n916 ;
  assign n1091 = n514 | n916 ;
  assign n1092 = ~n1090 & n1091 ;
  buffer buf_n1093( .i (n1092), .o (n1093) );
  assign n1094 = n828 & n1093 ;
  assign n1095 = n828 | n1093 ;
  assign n1096 = ~n1094 & n1095 ;
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  assign n1102 = ( n923 & n959 ) | ( n923 & n992 ) | ( n959 & n992 ) ;
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  assign n1105 = n935 & n945 ;
  assign n1106 = n935 | n945 ;
  assign n1107 = ~n1105 & n1106 ;
  buffer buf_n1108( .i (n1107), .o (n1108) );
  assign n1109 = ( n928 & n941 ) | ( n928 & n951 ) | ( n941 & n951 ) ;
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  assign n1112 = n1108 & n1111 ;
  assign n1113 = n1108 | n1111 ;
  assign n1114 = ~n1112 & n1113 ;
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  assign n1118 = n963 & n973 ;
  assign n1119 = n963 | n973 ;
  assign n1120 = ~n1118 & n1119 ;
  buffer buf_n1121( .i (n1120), .o (n1121) );
  assign n1122 = ( n969 & n979 ) | ( n969 & n985 ) | ( n979 & n985 ) ;
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  assign n1125 = n1121 & n1124 ;
  assign n1126 = n1121 | n1124 ;
  assign n1127 = ~n1125 & n1126 ;
  buffer buf_n1128( .i (n1127), .o (n1128) );
  assign n1131 = n1115 & n1128 ;
  assign n1132 = n1115 | n1128 ;
  assign n1133 = ~n1131 & n1132 ;
  buffer buf_n1134( .i (n1133), .o (n1134) );
  assign n1135 = n1104 & n1134 ;
  assign n1136 = n1104 | n1134 ;
  assign n1137 = ~n1135 & n1136 ;
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  assign n1141 = ( n918 & n1000 ) | ( n918 & n1079 ) | ( n1000 & n1079 ) ;
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  assign n1145 = n1014 & n1024 ;
  assign n1146 = n1014 | n1024 ;
  assign n1147 = ~n1145 & n1146 ;
  buffer buf_n1148( .i (n1147), .o (n1148) );
  assign n1149 = ( n1007 & n1020 ) | ( n1007 & n1030 ) | ( n1020 & n1030 ) ;
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  assign n1152 = n1148 & n1151 ;
  assign n1153 = n1148 | n1151 ;
  assign n1154 = ~n1152 & n1153 ;
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  assign n1158 = n1047 & n1057 ;
  assign n1159 = n1047 | n1057 ;
  assign n1160 = ~n1158 & n1159 ;
  buffer buf_n1161( .i (n1160), .o (n1161) );
  assign n1162 = ( n1040 & n1053 ) | ( n1040 & n1063 ) | ( n1053 & n1063 ) ;
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  assign n1165 = n1161 & n1164 ;
  assign n1166 = n1161 | n1164 ;
  assign n1167 = ~n1165 & n1166 ;
  buffer buf_n1168( .i (n1167), .o (n1168) );
  assign n1171 = n1155 & n1168 ;
  assign n1172 = n1155 | n1168 ;
  assign n1173 = ~n1171 & n1172 ;
  buffer buf_n1174( .i (n1173), .o (n1174) );
  assign n1175 = ( n1002 & n1038 ) | ( n1002 & n1071 ) | ( n1038 & n1071 ) ;
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  assign n1178 = n1174 & n1177 ;
  assign n1179 = n1174 | n1177 ;
  assign n1180 = ~n1178 & n1179 ;
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  assign n1184 = ( n1140 & n1142 ) | ( n1140 & n1183 ) | ( n1142 & n1183 ) ;
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n1187 = ( n1103 & n1117 ) | ( n1103 & n1130 ) | ( n1117 & n1130 ) ;
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  assign n1189 = ( n937 & n947 ) | ( n937 & n1110 ) | ( n947 & n1110 ) ;
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  assign n1197 = ( n965 & n975 ) | ( n965 & n1123 ) | ( n975 & n1123 ) ;
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  assign n1205 = n1193 & n1201 ;
  assign n1206 = n1193 | n1201 ;
  assign n1207 = ~n1205 & n1206 ;
  buffer buf_n1208( .i (n1207), .o (n1208) );
  assign n1209 = n1188 & n1208 ;
  assign n1210 = n1188 | n1208 ;
  assign n1211 = ~n1209 & n1210 ;
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  assign n1216 = ( n1016 & n1026 ) | ( n1016 & n1150 ) | ( n1026 & n1150 ) ;
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  assign n1224 = ( n1049 & n1059 ) | ( n1049 & n1163 ) | ( n1059 & n1163 ) ;
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  assign n1232 = n1220 & n1228 ;
  assign n1233 = n1220 | n1228 ;
  assign n1234 = ~n1232 & n1233 ;
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  assign n1236 = ( n1157 & n1170 ) | ( n1157 & n1176 ) | ( n1170 & n1176 ) ;
  buffer buf_n1237( .i (n1236), .o (n1237) );
  assign n1238 = n1235 & n1237 ;
  assign n1239 = n1235 | n1237 ;
  assign n1240 = ~n1238 & n1239 ;
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  assign n1245 = n1213 & n1242 ;
  assign n1246 = n1213 | n1242 ;
  assign n1247 = ~n1245 & n1246 ;
  buffer buf_n1248( .i (n1247), .o (n1248) );
  assign n1249 = n1186 & n1248 ;
  assign n1250 = n1186 | n1248 ;
  assign n1251 = ~n1249 & n1250 ;
  buffer buf_n1252( .i (n1251), .o (n1252) );
  assign n1253 = n518 | n820 ;
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  assign n1256 = ~n823 & n1255 ;
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  assign n1268 = ( n1188 & n1196 ) | ( n1188 & n1204 ) | ( n1196 & n1204 ) ;
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  assign n1276 = ( n1185 & n1215 ) | ( n1185 & n1244 ) | ( n1215 & n1244 ) ;
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  assign n1278 = ( n1223 & n1231 ) | ( n1223 & n1237 ) | ( n1231 & n1237 ) ;
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  assign n1286 = ( n1275 & n1277 ) | ( n1275 & n1285 ) | ( n1277 & n1285 ) ;
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  assign n1288 = n1139 & n1182 ;
  assign n1289 = n1139 | n1182 ;
  assign n1290 = ~n1288 & n1289 ;
  buffer buf_n1291( .i (n1290), .o (n1291) );
  assign n1292 = n1144 & n1291 ;
  assign n1293 = n1144 | n1291 ;
  assign n1294 = ~n1292 & n1293 ;
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  assign n1297 = n1272 & n1282 ;
  assign n1298 = n1272 | n1282 ;
  assign n1299 = ~n1297 & n1298 ;
  buffer buf_n1300( .i (n1299), .o (n1300) );
  assign n1301 = n1277 & n1300 ;
  assign n1302 = n1277 | n1300 ;
  assign n1303 = ~n1301 & n1302 ;
  assign y0 = n1089 ;
  assign y1 = n1101 ;
  assign y2 = n1252 ;
  assign y3 = n1267 ;
  assign y4 = 1'b0 ;
  assign y5 = n1287 ;
  assign y6 = n1296 ;
  assign y7 = n1303 ;
endmodule
