module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n19 , n20 , n21 , n22 , n23 , n25 , n26 , n27 , n28 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n38 , n39 , n40 , n41 , n42 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n68 , n70 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n104 , n105 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n135 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n148 , n149 , n150 , n151 , n152 , n153 , n155 , n156 , n157 , n158 , n159 , n160 , n162 , n163 , n164 , n165 , n166 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n206 , n207 , n208 , n209 , n210 , n211 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n283 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n296 , n298 , n300 , n302 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n323 , n324 , n325 , n326 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n341 , n342 , n343 , n344 , n345 , n347 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 ;
  buffer buf_n236( .i (x28), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n246( .i (x29), .o (n246) );
  buffer buf_n257( .i (x30), .o (n257) );
  assign n361 = ~n246 & n257 ;
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  assign n373 = ~n240 & n364 ;
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n168( .i (x21), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n148( .i (x18), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n155( .i (x19), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  assign n379 = ~n149 & n156 ;
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  assign n385 = n173 & n382 ;
  assign n386 = n374 & n385 ;
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n81( .i (x10), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n206( .i (x25), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  assign n389 = n84 & n209 ;
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n198( .i (x24), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n213( .i (x26), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  assign n397 = n203 | n218 ;
  buffer buf_n398( .i (n397), .o (n398) );
  assign n400 = n392 | n398 ;
  assign n401 = n387 & n400 ;
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  assign n406 = n202 & n364 ;
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n162( .i (x20), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  assign n411 = n163 & n169 ;
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  assign n415 = n148 & n155 ;
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  assign n421 = n413 & n418 ;
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  assign n426 = n148 | n155 ;
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  assign n430 = n413 & ~n429 ;
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  assign n435 = n423 | n432 ;
  buffer buf_n436( .i (n435), .o (n436) );
  assign n437 = n410 & n436 ;
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  assign n439 = n148 & ~n155 ;
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  assign n444 = ~n162 & n168 ;
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  assign n451 = n441 & n446 ;
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  assign n458 = n378 & n457 ;
  assign n459 = n438 | n458 ;
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  assign n461 = n14 & ~n404 ;
  assign n462 = ( n405 & n460 ) | ( n405 & ~n461 ) | ( n460 & ~n461 ) ;
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  assign n467 = ~n13 & n438 ;
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n219( .i (n218), .o (n219) );
  assign n474 = n219 | n391 ;
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  assign n477 = n388 & n476 ;
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  assign n486 = ~n9 & n423 ;
  assign n487 = n409 & n486 ;
  buffer buf_n399( .i (n398), .o (n399) );
  assign n488 = n387 & n399 ;
  assign n489 = n487 | n488 ;
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  assign n498 = n5 & n363 ;
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n241( .i (n240), .o (n241) );
  assign n505 = ~n241 & n452 ;
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  assign n508 = n171 & n239 ;
  assign n509 = n381 & n508 ;
  buffer buf_n510( .i (n509), .o (n510) );
  assign n515 = n422 | n510 ;
  buffer buf_n516( .i (n515), .o (n516) );
  assign n518 = n507 | n516 ;
  buffer buf_n519( .i (n518), .o (n519) );
  assign n520 = n409 & n502 ;
  assign n521 = n436 & n520 ;
  assign n522 = ( n504 & n519 ) | ( n504 & n521 ) | ( n519 & n521 ) ;
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n44( .i (x5), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  assign n530 = n46 | n238 ;
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n258( .i (n257), .o (n258) );
  assign n536 = n247 & ~n258 ;
  buffer buf_n537( .i (n536), .o (n537) );
  assign n545 = n5 & n537 ;
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  assign n548 = ~n533 & n547 ;
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n177( .i (x22), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  assign n551 = n162 & ~n168 ;
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  assign n555 = n381 & n554 ;
  buffer buf_n556( .i (n555), .o (n556) );
  assign n559 = n183 & n556 ;
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n30( .i (x3), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  assign n563 = n163 | n169 ;
  buffer buf_n564( .i (n563), .o (n564) );
  assign n567 = n428 | n564 ;
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  assign n572 = n36 | n569 ;
  buffer buf_n573( .i (n572), .o (n573) );
  assign n574 = ~n560 & n573 ;
  assign n575 = n550 & ~n574 ;
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n123( .i (x15), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  assign n577 = n127 | n531 ;
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n442( .i (n441), .o (n442) );
  assign n579 = n413 & n442 ;
  buffer buf_n580( .i (n579), .o (n580) );
  assign n582 = ~n578 & n580 ;
  assign n583 = n431 & n500 ;
  assign n584 = ( n501 & n582 ) | ( n501 & n583 ) | ( n582 & n583 ) ;
  buffer buf_n585( .i (n584), .o (n585) );
  assign n586 = n182 | n390 ;
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  assign n590 = ~n159 & n217 ;
  assign n591 = n414 & n590 ;
  buffer buf_n592( .i (n591), .o (n592) );
  assign n596 = n587 | n592 ;
  buffer buf_n597( .i (n596), .o (n597) );
  assign n598 = n585 & n597 ;
  assign n599 = n500 & ~n578 ;
  buffer buf_n600( .i (n599), .o (n600) );
  assign n601 = n180 & n412 ;
  buffer buf_n602( .i (n601), .o (n602) );
  assign n606 = n382 & n602 ;
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  assign n612 = n600 & n608 ;
  buffer buf_n613( .i (n612), .o (n613) );
  assign n622 = n598 | n613 ;
  assign n623 = n576 | n622 ;
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  assign n627 = n5 & ~n260 ;
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  assign n632 = n416 & n552 ;
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n226( .i (x27), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  assign n640 = n34 & ~n250 ;
  assign n641 = n231 & n640 ;
  assign n642 = n635 & n641 ;
  buffer buf_n643( .i (n642), .o (n643) );
  assign n647 = n631 & n643 ;
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n189( .i (x23), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  assign n652 = n191 & ~n238 ;
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  assign n656 = n547 & n655 ;
  assign n657 = ~n428 & n553 ;
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  assign n665 = n656 & n660 ;
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  assign n670 = n648 | n667 ;
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n25( .i (x2), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  assign n672 = n27 & ~n32 ;
  buffer buf_n673( .i (n672), .o (n673) );
  assign n674 = n236 & ~n246 ;
  buffer buf_n675( .i (n674), .o (n675) );
  assign n681 = n259 & n675 ;
  buffer buf_n682( .i (n681), .o (n682) );
  assign n689 = n673 & n682 ;
  buffer buf_n690( .i (n689), .o (n690) );
  assign n696 = n7 & ~n568 ;
  assign n697 = n690 & n696 ;
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  assign n703 = n671 | n702 ;
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n534( .i (n533), .o (n534) );
  assign n709 = n9 & ~n534 ;
  assign n710 = n248 & n259 ;
  buffer buf_n711( .i (n710), .o (n711) );
  assign n717 = ~n230 & n711 ;
  assign n718 = n634 & n717 ;
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  assign n721 = n709 & n720 ;
  buffer buf_n722( .i (n721), .o (n722) );
  assign n723 = ~n673 & n682 ;
  buffer buf_n724( .i (n723), .o (n724) );
  assign n729 = n6 & ~n34 ;
  assign n730 = n658 & n729 ;
  assign n731 = n724 & n730 ;
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  assign n736 = n722 | n734 ;
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  assign n740 = n704 | n739 ;
  assign n741 = n626 | n740 ;
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n538( .i (n537), .o (n538) );
  assign n743 = n240 & n538 ;
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  assign n748 = n7 & n182 ;
  assign n749 = n556 & n748 ;
  buffer buf_n38( .i (x4), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  assign n750 = n42 | n230 ;
  assign n751 = n7 | n750 ;
  assign n752 = n635 & ~n751 ;
  assign n753 = ( n745 & n749 ) | ( n745 & n752 ) | ( n749 & n752 ) ;
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = n440 & n552 ;
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  assign n762 = n417 & ~n564 ;
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  assign n768 = n761 | n764 ;
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n242( .i (n241), .o (n242) );
  assign n772 = n8 & n242 ;
  assign n773 = n367 & n772 ;
  buffer buf_n774( .i (n773), .o (n774) );
  assign n777 = n222 & n774 ;
  assign n778 = n771 & n777 ;
  buffer buf_n779( .i (n778), .o (n779) );
  assign n780 = n757 | n779 ;
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  assign n786 = n546 & n763 ;
  buffer buf_n787( .i (n786), .o (n787) );
  assign n790 = n587 & n787 ;
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  assign n794 = ~n238 & n248 ;
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  assign n802 = n628 & n796 ;
  buffer buf_n803( .i (n802), .o (n803) );
  assign n805 = n220 & n803 ;
  assign n806 = n769 & n805 ;
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  assign n809 = n793 | n808 ;
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  assign n813 = n782 | n812 ;
  buffer buf_n814( .i (n813), .o (n814) );
  assign n815 = n742 | n814 ;
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  assign n816 = n585 | n789 ;
  buffer buf_n817( .i (n816), .o (n817) );
  assign n818 = n396 & n817 ;
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n92( .i (x11), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  assign n825 = n217 & n759 ;
  buffer buf_n826( .i (n825), .o (n826) );
  assign n827 = n98 & n826 ;
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  assign n833 = n219 & n764 ;
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  assign n838 = ~n102 & n836 ;
  assign n839 = ( n776 & n831 ) | ( n776 & n838 ) | ( n831 & n838 ) ;
  assign n840 = n757 | n839 ;
  assign n841 = n98 & ~n183 ;
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  assign n845 = n597 & ~n843 ;
  buffer buf_n846( .i (n845), .o (n846) );
  assign n847 = n817 & n846 ;
  assign n848 = n549 & ~n573 ;
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  assign n851 = n613 | n734 ;
  assign n852 = n850 | n851 ;
  assign n853 = n847 | n852 ;
  assign n854 = n840 | n853 ;
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  assign n859 = ~n171 & n380 ;
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n19( .i (x1), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n164( .i (n163), .o (n164) );
  assign n864 = n21 & ~n164 ;
  buffer buf_n865( .i (n864), .o (n865) );
  assign n867 = n538 & n865 ;
  assign n868 = n860 & n867 ;
  buffer buf_n869( .i (n868), .o (n869) );
  assign n870 = n196 & n869 ;
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n261( .i (n260), .o (n261) );
  assign n873 = n261 & n795 ;
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n137( .i (x17), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  assign n879 = ~n140 & n216 ;
  assign n880 = n759 & n879 ;
  buffer buf_n881( .i (n880), .o (n881) );
  assign n887 = n874 & n881 ;
  buffer buf_n888( .i (n887), .o (n888) );
  assign n899 = n744 & n826 ;
  buffer buf_n900( .i (n899), .o (n900) );
  assign n911 = n888 | n900 ;
  buffer buf_n912( .i (n911), .o (n912) );
  assign n915 = n872 | n912 ;
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  assign n918 = n519 & n544 ;
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n746( .i (n745), .o (n746) );
  assign n920 = ~n571 & n746 ;
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n747( .i (n746), .o (n747) );
  assign n923 = n747 & n835 ;
  assign n924 = n921 | n923 ;
  buffer buf_n443( .i (n442), .o (n443) );
  assign n925 = n173 & n443 ;
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n210( .i (n209), .o (n210) );
  assign n930 = n181 | n210 ;
  buffer buf_n931( .i (n930), .o (n931) );
  assign n935 = n797 & n931 ;
  assign n936 = n926 & n935 ;
  buffer buf_n937( .i (n936), .o (n937) );
  assign n939 = n542 & ~n842 ;
  assign n940 = n937 & n939 ;
  buffer buf_n941( .i (n940), .o (n941) );
  assign n944 = n924 | n941 ;
  assign n945 = n919 | n944 ;
  assign n946 = n917 | n945 ;
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n243( .i (n242), .o (n243) );
  assign n950 = n243 & n719 ;
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n712( .i (n711), .o (n712) );
  assign n955 = n182 & n712 ;
  assign n956 = n556 & n955 ;
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  assign n960 = n952 | n959 ;
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  assign n963 = ~n240 & n538 ;
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  assign n969 = n142 & n218 ;
  assign n970 = n761 & n969 ;
  buffer buf_n971( .i (n970), .o (n971) );
  assign n972 = n966 & n971 ;
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n72( .i (x9), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  assign n977 = ~n427 & n445 ;
  buffer buf_n978( .i (n977), .o (n978) );
  assign n982 = n178 & ~n237 ;
  assign n983 = n362 & n982 ;
  buffer buf_n984( .i (n983), .o (n984) );
  assign n989 = n978 & n984 ;
  buffer buf_n990( .i (n989), .o (n990) );
  assign n993 = ~n78 & n990 ;
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  assign n999 = n975 | n998 ;
  assign n1000 = n962 | n999 ;
  assign n1001 = n422 & n540 ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  assign n1004 = n659 & n744 ;
  buffer buf_n1005( .i (n1004), .o (n1005) );
  assign n1006 = n1002 | n1005 ;
  buffer buf_n1007( .i (n1006), .o (n1007) );
  assign n1011 = n659 & n874 ;
  buffer buf_n1012( .i (n1011), .o (n1012) );
  assign n1014 = n231 & n365 ;
  assign n1015 = n635 & n1014 ;
  buffer buf_n1016( .i (n1015), .o (n1016) );
  assign n1021 = n1012 | n1016 ;
  buffer buf_n1022( .i (n1021), .o (n1022) );
  assign n1025 = n1007 | n1022 ;
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  assign n1028 = ~n230 & n633 ;
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  assign n1034 = n248 | n259 ;
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  assign n1037 = n241 & ~n1036 ;
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  assign n1042 = n1031 & n1039 ;
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  assign n1047 = ~n570 & n875 ;
  assign n1048 = ( n834 & n876 ) | ( n834 & n1047 ) | ( n876 & n1047 ) ;
  buffer buf_n1049( .i (n1048), .o (n1049) );
  assign n1053 = n1043 | n1049 ;
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n184( .i (n183), .o (n184) );
  assign n1056 = n184 & n869 ;
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n932( .i (n931), .o (n932) );
  assign n1060 = n714 & n932 ;
  assign n1061 = n766 & n1060 ;
  buffer buf_n1062( .i (n1061), .o (n1062) );
  assign n1064 = n1058 | n1062 ;
  buffer buf_n1065( .i (n1064), .o (n1065) );
  assign n1066 = n1054 | n1065 ;
  assign n1067 = n1027 | n1066 ;
  assign n1068 = n1000 | n1067 ;
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n349( .i (x44), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  assign n1070 = n181 & n978 ;
  buffer buf_n1071( .i (n1070), .o (n1071) );
  assign n1075 = n75 | n239 ;
  buffer buf_n1076( .i (n537), .o (n1076) );
  assign n1077 = ~n1075 & n1076 ;
  buffer buf_n1078( .i (n1077), .o (n1078) );
  assign n1080 = n1071 & n1078 ;
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n304( .i (x38), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n328( .i (x41), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  assign n1084 = n307 | n331 ;
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n315( .i (x39), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n341( .i (x42), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  assign n1086 = n318 | n344 ;
  buffer buf_n1087( .i (n1086), .o (n1087) );
  assign n1088 = n1085 | n1087 ;
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n323( .i (x40), .o (n323) );
  buffer buf_n347( .i (x43), .o (n347) );
  assign n1093 = n323 | n347 ;
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  assign n1100 = n1089 | n1099 ;
  buffer buf_n1101( .i (n1100), .o (n1101) );
  assign n1102 = n1082 & ~n1101 ;
  buffer buf_n1103( .i (n1102), .o (n1103) );
  assign n1107 = n360 & n1103 ;
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n866( .i (n865), .o (n866) );
  assign n1110 = n180 | n192 ;
  buffer buf_n1111( .i (n1110), .o (n1111) );
  assign n1112 = n866 & n1111 ;
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  assign n1116 = n388 & n1115 ;
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n211( .i (n210), .o (n211) );
  assign n1120 = n211 & n796 ;
  buffer buf_n1121( .i (n1120), .o (n1121) );
  assign n1122 = n581 & n1121 ;
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  assign n1125 = n100 & ~n265 ;
  assign n1126 = n1123 & n1125 ;
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  assign n1129 = n1118 | n1128 ;
  assign n1130 = n1108 | n1129 ;
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n1132( .i (n237), .o (n1132) );
  assign n1133 = n215 & ~n1132 ;
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n1135( .i (n1134), .o (n1135) );
  assign n1138 = n443 & ~n1135 ;
  assign n1139 = n252 & ~n1138 ;
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  assign n1142 = n594 & n1141 ;
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  assign n1145 = n432 & n541 ;
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  assign n1149 = n180 & n260 ;
  buffer buf_n1150( .i (n1149), .o (n1150) );
  assign n1155 = n796 & n1150 ;
  assign n1156 = n980 & n1155 ;
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  assign n1161 = n1148 | n1160 ;
  assign n1162 = n1144 | n1161 ;
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  assign n1163 = n512 & n542 ;
  assign n1164 = ( n543 & n609 ) | ( n543 & n1163 ) | ( n609 & n1163 ) ;
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  assign n1168 = n1162 | n1167 ;
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  assign n1169 = n1079 & n1089 ;
  assign n1170 = n1073 & n1169 ;
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n270( .i (x31), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n285( .i (x33), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  assign n1173 = n275 | n290 ;
  assign n1174 = n321 & ~n1173 ;
  assign n1175 = n79 & n1174 ;
  assign n1176 = n992 & n1175 ;
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  assign n1181 = n1172 | n1178 ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  assign n1184 = n1168 | n1183 ;
  assign n1185 = n1131 | n1184 ;
  assign n1186 = n1069 | n1185 ;
  assign n1187 = n949 | n1186 ;
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  assign n1188 = n263 & n1136 ;
  assign n1189 = n765 & n1188 ;
  assign n1190 = n957 | n1189 ;
  buffer buf_n1191( .i (n1190), .o (n1191) );
  assign n1192 = n801 & n1191 ;
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n976( .i (n975), .o (n976) );
  assign n1196 = ~n323 & n347 ;
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  assign n1203 = ~n1089 & n1202 ;
  buffer buf_n1204( .i (n1203), .o (n1204) );
  assign n1207 = ~n355 & n1078 ;
  assign n1208 = n1072 & n1207 ;
  buffer buf_n1209( .i (n1208), .o (n1209) );
  assign n1213 = n1204 & n1209 ;
  buffer buf_n1214( .i (n1213), .o (n1214) );
  assign n1218 = n834 & n1039 ;
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  assign n1221 = n1214 | n1220 ;
  buffer buf_n1222( .i (n1221), .o (n1222) );
  assign n1225 = n976 | n1222 ;
  assign n1226 = n1195 | n1225 ;
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1228( .i (n229), .o (n1228) );
  assign n1229 = n633 & n1228 ;
  buffer buf_n1230( .i (n1229), .o (n1230) );
  assign n1233 = n35 | n1036 ;
  assign n1234 = n1230 & ~n1233 ;
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  assign n1239 = n1143 | n1238 ;
  buffer buf_n1240( .i (n1239), .o (n1240) );
  assign n1241 = n1046 | n1240 ;
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n938( .i (n937), .o (n938) );
  assign n1242 = ~n844 & n938 ;
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  assign n1244 = n101 & n1123 ;
  assign n1245 = n878 & n1244 ;
  buffer buf_n1246( .i (n1245), .o (n1246) );
  assign n1247 = n1243 | n1246 ;
  assign n1248 = n1027 | n1247 ;
  assign n1249 = n1241 | n1248 ;
  buffer buf_n447( .i (n446), .o (n447) );
  assign n1250 = n381 & n447 ;
  assign n1251 = n1111 & n1250 ;
  assign n1252 = n964 & n1251 ;
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n253( .i (n252), .o (n253) );
  assign n1256 = n252 & n510 ;
  assign n1257 = ( n253 & n607 ) | ( n253 & n1256 ) | ( n607 & n1256 ) ;
  assign n1258 = n1253 | n1257 ;
  buffer buf_n1259( .i (n1258), .o (n1259) );
  assign n1262 = n745 | n875 ;
  assign n1263 = ~n571 & n1262 ;
  buffer buf_n1264( .i (n1263), .o (n1264) );
  assign n1265 = n1259 | n1264 ;
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  assign n1269 = n971 & n1039 ;
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n433( .i (n432), .o (n433) );
  assign n1273 = n433 | n507 ;
  assign n1274 = n255 & n1273 ;
  assign n1275 = n1270 | n1274 ;
  buffer buf_n1276( .i (n1275), .o (n1276) );
  assign n1278 = n1118 | n1276 ;
  buffer buf_n1279( .i (n1278), .o (n1279) );
  assign n1280 = n1268 | n1279 ;
  assign n1281 = n1249 | n1280 ;
  assign n1282 = n1227 | n1281 ;
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  assign n1284 = n1240 | n1277 ;
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  assign n1285 = n261 & n418 ;
  buffer buf_n1286( .i (n1285), .o (n1286) );
  assign n1289 = n449 & n1286 ;
  buffer buf_n1290( .i (n1289), .o (n1290) );
  assign n1293 = n475 & n1290 ;
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  assign n1296 = n242 & ~n263 ;
  assign n1297 = n220 & n1296 ;
  assign n1298 = n766 & n1297 ;
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  assign n1301 = n1295 | n1300 ;
  buffer buf_n1302( .i (n1301), .o (n1302) );
  assign n1303 = n917 | n1302 ;
  assign n1304 = n1284 | n1303 ;
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  assign n1307 = n253 & n423 ;
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  assign n1310 = n938 | n1309 ;
  buffer buf_n1311( .i (n1310), .o (n1311) );
  assign n1312 = n1266 | n1311 ;
  buffer buf_n1313( .i (n1312), .o (n1313) );
  assign n1314 = n1106 | n1313 ;
  buffer buf_n1315( .i (n1314), .o (n1315) );
  assign n1316 = n1069 | n1315 ;
  assign n1317 = n1306 | n1316 ;
  assign n1318 = n181 & n364 ;
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  assign n1320 = n382 & ~n566 ;
  assign n1321 = n1319 & n1320 ;
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  assign n1325 = n425 & n716 ;
  assign n1326 = n1324 | n1325 ;
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n165( .i (n164), .o (n165) );
  assign n1328 = ~n165 & n192 ;
  buffer buf_n1329( .i (n363), .o (n1329) );
  assign n1330 = n1328 & n1329 ;
  buffer buf_n1331( .i (n1330), .o (n1331) );
  assign n1332 = n861 & n1331 ;
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  assign n1335 = n871 | n1334 ;
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  assign n1337 = n764 & n1151 ;
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  assign n1342 = n1336 | n1341 ;
  assign n1343 = n1327 | n1342 ;
  assign n1344 = n1157 | n1235 ;
  assign n1345 = n951 | n1344 ;
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  assign n1347 = ~n1085 & n1087 ;
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  assign n1352 = n1083 & n1351 ;
  assign n1353 = n1346 | n1352 ;
  buffer buf_n1354( .i (n1353), .o (n1354) );
  assign n1355 = n1343 | n1354 ;
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  assign n1358 = n374 & n1029 ;
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n767( .i (n766), .o (n767) );
  assign n1363 = n1134 & n1329 ;
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  assign n1368 = n767 & n1367 ;
  buffer buf_n1369( .i (n1368), .o (n1369) );
  assign n1370 = n1362 | n1369 ;
  buffer buf_n1371( .i (n1370), .o (n1371) );
  assign n1372 = n172 | n429 ;
  buffer buf_n1373( .i (n1372), .o (n1373) );
  assign n1374 = n374 & ~n1373 ;
  assign n1375 = ~n194 & n658 ;
  buffer buf_n1376( .i (n1375), .o (n1376) );
  assign n1379 = n1374 & ~n1376 ;
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  assign n1385 = n1371 | n1384 ;
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  assign n1387 = n861 & n986 ;
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n557( .i (n556), .o (n557) );
  assign n1392 = n653 & n1329 ;
  buffer buf_n1393( .i (n1392), .o (n1393) );
  assign n1395 = n1364 | n1393 ;
  assign n1396 = n557 & n1395 ;
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  assign n1400 = n1058 | n1398 ;
  assign n1401 = n1391 | n1400 ;
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  assign n1405 = n1386 | n1404 ;
  assign n1406 = n1357 | n1405 ;
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  assign n1407 = n1062 | n1299 ;
  assign n1408 = n1271 | n1407 ;
  assign n1409 = n1179 | n1408 ;
  buffer buf_n115( .i (x14), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  assign n1410 = n229 | n239 ;
  assign n1411 = n1035 | n1410 ;
  buffer buf_n1412( .i (n1411), .o (n1412) );
  assign n1413 = n121 & ~n1412 ;
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n107( .i (x13), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  assign n1416 = n111 & n172 ;
  assign n1417 = ~n120 & n1416 ;
  assign n1418 = ~n1412 & n1417 ;
  buffer buf_n1419( .i (n1418), .o (n1419) );
  assign n1422 = n1414 | n1419 ;
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  assign n1426 = n761 & n1364 ;
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  assign n1430 = n367 & n765 ;
  buffer buf_n1431( .i (n1430), .o (n1431) );
  assign n1433 = n394 & n1431 ;
  assign n1434 = n1429 | n1433 ;
  buffer buf_n1435( .i (n1434), .o (n1435) );
  assign n1436 = n1425 | n1435 ;
  assign n1437 = n1409 | n1436 ;
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  assign n1440 = n241 & n1150 ;
  buffer buf_n1441( .i (n1440), .o (n1441) );
  assign n1442 = n557 & n1441 ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  assign n1445 = ~n693 & n1443 ;
  buffer buf_n1446( .i (n1445), .o (n1446) );
  assign n1448 = n761 & n1151 ;
  buffer buf_n1449( .i (n1448), .o (n1449) );
  assign n1452 = n194 & n262 ;
  buffer buf_n1453( .i (n760), .o (n1453) );
  assign n1454 = n1452 & n1453 ;
  buffer buf_n1455( .i (n1454), .o (n1455) );
  assign n1459 = n1449 | n1455 ;
  buffer buf_n1460( .i (n1459), .o (n1460) );
  assign n1461 = n1294 | n1460 ;
  assign n1462 = n1446 | n1461 ;
  assign n1463 = n914 | n1462 ;
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  assign n1466 = n1131 | n1465 ;
  assign n1467 = n1439 | n1466 ;
  assign n1468 = n1406 | n1467 ;
  buffer buf_n513( .i (n512), .o (n513) );
  assign n1469 = n513 & n716 ;
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  assign n1472 = n1238 | n1300 ;
  assign n1473 = n1471 | n1472 ;
  assign n1474 = n1128 | n1179 ;
  assign n1475 = n1473 | n1474 ;
  buffer buf_n1476( .i (n380), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  assign n1478 = n866 & n1477 ;
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n174( .i (n173), .o (n174) );
  assign n1481 = n174 & n195 ;
  assign n1482 = n375 & n1481 ;
  assign n1483 = n1480 & n1482 ;
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  assign n1486 = n1446 | n1485 ;
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  assign n1488 = n223 & n1292 ;
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  assign n1491 = n1487 | n1490 ;
  assign n1492 = n1475 | n1491 ;
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  assign n1495 = ~n313 & n1082 ;
  buffer buf_n1496( .i (n1495), .o (n1496) );
  assign n1497 = n339 & n1496 ;
  assign n1498 = n1065 | n1497 ;
  assign n1499 = n917 | n1498 ;
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  assign n1502 = n326 | n344 ;
  assign n1503 = ~n319 & n1502 ;
  assign n1504 = n1085 | n1503 ;
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  assign n1507 = n1081 & n1506 ;
  buffer buf_n1508( .i (n1507), .o (n1508) );
  assign n1511 = ~n1092 & n1508 ;
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  assign n1512 = n79 & n991 ;
  buffer buf_n1513( .i (n1512), .o (n1513) );
  assign n1516 = n294 & n1513 ;
  buffer buf_n1517( .i (n1516), .o (n1517) );
  assign n1518 = n1511 | n1517 ;
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  assign n1520 = n268 & n1143 ;
  assign n1521 = n954 | n1520 ;
  assign n1522 = n1519 | n1521 ;
  buffer buf_n1523( .i (n1522), .o (n1523) );
  assign n1524 = n317 & ~n343 ;
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  assign n1533 = n1496 & n1532 ;
  buffer buf_n1074( .i (n1073), .o (n1074) );
  assign n1534 = n609 | n1074 ;
  assign n1535 = n878 & n1534 ;
  assign n1536 = n1271 | n1535 ;
  assign n1537 = n1533 | n1536 ;
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  assign n1540 = n1523 | n1539 ;
  assign n1541 = n1501 | n1540 ;
  assign n1542 = n1494 | n1541 ;
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  assign n1543 = n1063 | n1148 ;
  assign n1544 = n1009 | n1543 ;
  assign n1545 = n1119 | n1544 ;
  buffer buf_n1059( .i (n1058), .o (n1059) );
  assign n1546 = n593 & n966 ;
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  assign n1550 = n1059 | n1548 ;
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n1551( .i (n1132), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  assign n1553 = ~n42 & n1552 ;
  buffer buf_n1554( .i (n1553), .o (n1554) );
  assign n1555 = n540 & ~n1554 ;
  buffer buf_n1556( .i (n1555), .o (n1556) );
  assign n1557 = n244 & n1556 ;
  assign n1558 = n1032 & n1557 ;
  buffer buf_n1559( .i (n1558), .o (n1559) );
  assign n1561 = n1127 | n1559 ;
  assign n1562 = n1550 | n1561 ;
  buffer buf_n1563( .i (n1562), .o (n1563) );
  assign n1565 = n1545 | n1563 ;
  assign n1566 = n947 | n1565 ;
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n981( .i (n980), .o (n981) );
  assign n1568 = n195 & n540 ;
  assign n1569 = n981 & n1568 ;
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n296( .i (x34), .o (n296) );
  buffer buf_n298( .i (x35), .o (n298) );
  assign n1573 = n296 | n298 ;
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n300( .i (x36), .o (n300) );
  buffer buf_n302( .i (x37), .o (n302) );
  assign n1585 = ~n300 & n302 ;
  buffer buf_n1586( .i (n1585), .o (n1586) );
  assign n1587 = n1574 | n1586 ;
  buffer buf_n283( .i (x32), .o (n283) );
  assign n1588 = n270 | n283 ;
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  assign n1591 = n287 & ~n1589 ;
  assign n1592 = ( n1587 & n1590 ) | ( n1587 & ~n1591 ) | ( n1590 & ~n1591 ) ;
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  assign n1600 = n1572 & n1599 ;
  assign n1601 = n1166 | n1600 ;
  assign n1602 = n962 | n1601 ;
  buffer buf_n1013( .i (n1012), .o (n1013) );
  assign n1603 = n1013 | n1323 ;
  assign n1604 = n1423 | n1603 ;
  buffer buf_n1605( .i (n1604), .o (n1605) );
  assign n1607 = n980 & n1331 ;
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  assign n1610 = n407 & n659 ;
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  assign n1613 = n1609 | n1612 ;
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  assign n1620 = n146 & n1428 ;
  buffer buf_n1621( .i (n1620), .o (n1621) );
  assign n1622 = n1614 | n1621 ;
  assign n1623 = n1605 | n1622 ;
  buffer buf_n1624( .i (n1623), .o (n1624) );
  assign n1627 = n1602 | n1624 ;
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n987( .i (n986), .o (n987) );
  assign n1628 = n987 & n1479 ;
  buffer buf_n1629( .i (n1628), .o (n1629) );
  assign n1630 = n1146 | n1629 ;
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  assign n1632 = n966 & n1232 ;
  buffer buf_n1633( .i (n1632), .o (n1633) );
  assign n1634 = n981 & n1441 ;
  buffer buf_n1635( .i (n1634), .o (n1635) );
  buffer buf_n1636( .i (n1635), .o (n1636) );
  assign n1637 = n1633 | n1636 ;
  assign n1638 = n1631 | n1637 ;
  buffer buf_n1639( .i (n1638), .o (n1639) );
  assign n1640 = n1055 | n1639 ;
  buffer buf_n47( .i (n46), .o (n47) );
  assign n1641 = n47 & ~n1551 ;
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  assign n1646 = n719 & n1644 ;
  buffer buf_n1647( .i (n1646), .o (n1647) );
  assign n1650 = ~n570 & n965 ;
  assign n1651 = n35 | n1642 ;
  assign n1652 = n569 | n1651 ;
  buffer buf_n1653( .i (n1652), .o (n1653) );
  assign n1657 = n1650 & n1653 ;
  assign n1658 = n1647 | n1657 ;
  buffer buf_n1659( .i (n1658), .o (n1659) );
  assign n1662 = n1369 | n1659 ;
  buffer buf_n1663( .i (n1662), .o (n1663) );
  assign n1666 = n499 | n539 ;
  buffer buf_n1667( .i (n1666), .o (n1667) );
  assign n1670 = n506 & n1667 ;
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  assign n1674 = n457 & n1041 ;
  assign n1675 = n1673 | n1674 ;
  assign n1676 = n975 | n1675 ;
  assign n1677 = n1663 | n1676 ;
  assign n1678 = n1640 | n1677 ;
  assign n1679 = n1627 | n1678 ;
  assign n1680 = n698 | n732 ;
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n58( .i (x6), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n661( .i (n660), .o (n661) );
  assign n1683 = n66 & n661 ;
  assign n1684 = n727 & n1683 ;
  assign n1685 = n1681 | n1684 ;
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  assign n1689 = n694 & n1444 ;
  assign n1690 = n541 & n1644 ;
  assign n1691 = n560 & n1690 ;
  buffer buf_n1692( .i (n1691), .o (n1692) );
  assign n1695 = n648 | n1692 ;
  assign n1696 = n1689 | n1695 ;
  assign n1697 = n1686 | n1696 ;
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  assign n1699 = n1019 | n1206 ;
  assign n1700 = ( n1020 & n1212 ) | ( n1020 & n1699 ) | ( n1212 & n1699 ) ;
  buffer buf_n1701( .i (n1700), .o (n1701) );
  assign n1702 = n1698 | n1701 ;
  buffer buf_n1703( .i (n1702), .o (n1703) );
  assign n1704 = n1679 | n1703 ;
  assign n1705 = n1567 | n1704 ;
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  assign n1706 = n223 & n1147 ;
  buffer buf_n1707( .i (n1706), .o (n1707) );
  assign n1708 = n1045 | n1707 ;
  assign n1709 = n651 | n1708 ;
  assign n1710 = n1688 | n1709 ;
  assign n1711 = n1665 | n1710 ;
  assign n1712 = n994 | n1359 ;
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n1716( .i (n539), .o (n1716) );
  assign n1717 = n204 & n1716 ;
  buffer buf_n1718( .i (n1717), .o (n1718) );
  assign n1719 = n661 & n1718 ;
  buffer buf_n1720( .i (n1719), .o (n1720) );
  assign n1721 = n1451 | n1720 ;
  buffer buf_n1722( .i (n658), .o (n1722) );
  assign n1723 = n1319 & n1722 ;
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  assign n1735 = n1721 | n1727 ;
  assign n1736 = n1715 | n1735 ;
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  assign n1739 = n1444 | n1692 ;
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  assign n1743 = n1109 | n1742 ;
  assign n1744 = n1738 | n1743 ;
  assign n1745 = n1711 | n1744 ;
  buffer buf_n1746( .i (n634), .o (n1746) );
  assign n1747 = n964 & n1746 ;
  buffer buf_n1748( .i (n1747), .o (n1748) );
  assign n1751 = n1338 | n1748 ;
  assign n1752 = n1397 | n1751 ;
  assign n1753 = n1171 | n1752 ;
  assign n1754 = n1346 | n1753 ;
  assign n1755 = n916 | n1754 ;
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  assign n1759 = n1438 | n1564 ;
  assign n1760 = n1758 | n1759 ;
  assign n1761 = n1745 | n1760 ;
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  assign n1762 = n1217 | n1279 ;
  assign n1763 = n1523 | n1762 ;
  assign n1764 = n1626 | n1763 ;
  assign n1765 = n1191 | n1299 ;
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  buffer buf_n1584( .i (n1583), .o (n1584) );
  assign n1768 = n300 | n302 ;
  buffer buf_n1769( .i (n1768), .o (n1769) );
  assign n1770 = n1574 | n1769 ;
  buffer buf_n1771( .i (n1770), .o (n1771) );
  assign n1772 = n283 | n285 ;
  buffer buf_n1773( .i (n1772), .o (n1773) );
  assign n1784 = n272 | n1773 ;
  buffer buf_n1785( .i (n1784), .o (n1785) );
  assign n1786 = n1771 & ~n1785 ;
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  assign n1792 = n1571 & n1791 ;
  buffer buf_n1793( .i (n1792), .o (n1793) );
  assign n1794 = ~n1584 & n1793 ;
  assign n1795 = n1767 | n1794 ;
  buffer buf_n1394( .i (n1393), .o (n1394) );
  assign n1796 = n557 & n1394 ;
  assign n1797 = n1005 | n1796 ;
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  assign n1802 = n455 & n686 ;
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  assign n1805 = n1063 | n1804 ;
  assign n1806 = n1800 | n1805 ;
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  assign n1807 = n1018 | n1750 ;
  buffer buf_n1808( .i (n1807), .o (n1808) );
  assign n1809 = n975 | n1808 ;
  assign n1810 = n1806 | n1809 ;
  assign n1811 = n1795 | n1810 ;
  assign n1812 = n1313 | n1464 ;
  assign n1813 = n1811 | n1812 ;
  assign n1814 = ~n360 & n1103 ;
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n450( .i (n449), .o (n450) );
  assign n1815 = n184 & n450 ;
  assign n1816 = n1288 & n1815 ;
  assign n1817 = n1635 | n1816 ;
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n595( .i (n594), .o (n595) );
  assign n1819 = n101 & n877 ;
  assign n1820 = n595 & n1819 ;
  assign n1821 = n1818 | n1820 ;
  assign n1822 = n1814 | n1821 ;
  buffer buf_n1823( .i (n1822), .o (n1823) );
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1825( .i (n1824), .o (n1825) );
  assign n1826 = n1813 | n1825 ;
  assign n1827 = n1764 | n1826 ;
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  assign n1828 = n378 & n639 ;
  assign n1829 = n1451 | n1803 ;
  assign n1830 = n1828 | n1829 ;
  assign n1831 = n942 | n1830 ;
  assign n1832 = n1606 | n1831 ;
  assign n1833 = n1195 | n1832 ;
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  assign n1836 = n1380 | n1629 ;
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  assign n1839 = n377 & n884 ;
  assign n1840 = n973 | n1839 ;
  assign n1841 = n1837 | n1840 ;
  buffer buf_n1842( .i (n1841), .o (n1842) );
  assign n1843 = n1402 | n1842 ;
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  assign n1845 = n1264 | n1633 ;
  buffer buf_n1846( .i (n1845), .o (n1846) );
  assign n1847 = n1793 | n1846 ;
  assign n1848 = n1010 | n1847 ;
  assign n1849 = n433 & n1718 ;
  assign n1850 = n1612 | n1849 ;
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  assign n1854 = n443 & ~n566 ;
  buffer buf_n1855( .i (n1854), .o (n1855) );
  assign n1857 = n211 & n262 ;
  buffer buf_n1858( .i (n1857), .o (n1858) );
  assign n1860 = n1855 & n1858 ;
  buffer buf_n1861( .i (n1860), .o (n1861) );
  assign n1862 = n90 & n1861 ;
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n224( .i (n223), .o (n224) );
  assign n1865 = ~n224 & n1148 ;
  assign n1866 = n1864 | n1865 ;
  assign n1867 = n1853 | n1866 ;
  assign n1868 = n1848 | n1867 ;
  assign n1869 = n1844 | n1868 ;
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  assign n1870 = n589 & n1431 ;
  buffer buf_n1871( .i (n1870), .o (n1871) );
  buffer buf_n1872( .i (n1871), .o (n1872) );
  assign n1873 = n1485 | n1673 ;
  assign n1874 = n1872 | n1873 ;
  assign n1875 = n1017 | n1236 ;
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  assign n1878 = n1165 | n1336 ;
  assign n1879 = n1877 | n1878 ;
  assign n1880 = n1874 | n1879 ;
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  assign n1883 = n1869 | n1882 ;
  assign n1884 = n1835 | n1883 ;
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1885( .i (n974), .o (n1885) );
  assign n1886 = n1272 | n1885 ;
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n1888( .i (n1887), .o (n1888) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  assign n1889 = n727 | n877 ;
  assign n1890 = n562 & n1889 ;
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  assign n1894 = n1052 | n1371 ;
  assign n1895 = n1893 | n1894 ;
  assign n1896 = n1888 | n1895 ;
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  assign n1897 = ~n281 & n1572 ;
  assign n1898 = n1783 & n1897 ;
  assign n1899 = n1801 | n1898 ;
  assign n1900 = n1388 | n1427 ;
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  assign n1904 = n1322 | n1333 ;
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1907( .i (n1906), .o (n1907) );
  assign n1908 = n1903 | n1907 ;
  buffer buf_n1909( .i (n1908), .o (n1909) );
  assign n1910 = n1899 | n1909 ;
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  assign n1911 = n922 | n1458 ;
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1549( .i (n1548), .o (n1549) );
  assign n1914 = n1045 | n1549 ;
  assign n1915 = n1729 | n1914 ;
  assign n1916 = n1913 | n1915 ;
  assign n1917 = n1910 | n1916 ;
  assign n1918 = n1896 | n1917 ;
  assign n1919 = ~n296 & n298 ;
  assign n1920 = ~n271 & n1919 ;
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  assign n1928 = n1570 & n1927 ;
  assign n1929 = n1381 | n1928 ;
  buffer buf_n1003( .i (n1002), .o (n1003) );
  assign n1930 = n1003 | n1013 ;
  assign n1931 = n1720 | n1930 ;
  assign n1932 = n1929 | n1931 ;
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n1934( .i (n1933), .o (n1934) );
  buffer buf_n943( .i (n942), .o (n943) );
  assign n1935 = n943 | n1639 ;
  assign n1936 = n1934 | n1935 ;
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  assign n1938 = n1224 | n1881 ;
  assign n1939 = n1937 | n1938 ;
  assign n1940 = n1918 | n1939 ;
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n434( .i (n433), .o (n434) );
  assign n1941 = ~n85 & n210 ;
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  assign n1949 = n715 | n1944 ;
  assign n1950 = n434 & n1949 ;
  assign n1951 = n211 | n218 ;
  buffer buf_n1952( .i (n1951), .o (n1952) );
  assign n1953 = n450 & n1952 ;
  assign n1954 = n1288 & n1953 ;
  buffer buf_n1955( .i (n1954), .o (n1955) );
  assign n1956 = n1950 | n1955 ;
  buffer buf_n1957( .i (n1956), .o (n1957) );
  assign n1958 = n1447 | n1957 ;
  assign n1959 = n1180 | n1958 ;
  assign n1960 = n1887 | n1959 ;
  assign n1961 = n1757 | n1960 ;
  assign n1962 = n1703 | n1961 ;
  assign n1963 = n387 & n1944 ;
  assign n1964 = n1861 | n1963 ;
  buffer buf_n1965( .i (n1964), .o (n1965) );
  assign n1966 = n1659 | n1965 ;
  assign n1967 = n1766 | n1966 ;
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  assign n1968 = n1031 & n1556 ;
  assign n1969 = n1671 | n1968 ;
  assign n1970 = n1713 | n1969 ;
  buffer buf_n1971( .i (n1970), .o (n1971) );
  assign n1975 = n1261 | n1971 ;
  assign n1976 = n1967 | n1975 ;
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  assign n1979 = n1460 | n1901 ;
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  assign n1982 = n454 & n680 ;
  buffer buf_n1983( .i (n1982), .o (n1983) );
  buffer buf_n1984( .i (n1983), .o (n1984) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  assign n1985 = n798 & n1952 ;
  buffer buf_n1986( .i (n1985), .o (n1986) );
  assign n1987 = n928 & n1986 ;
  assign n1988 = n1984 | n1987 ;
  assign n1989 = n1058 | n1484 ;
  assign n1990 = n1988 | n1989 ;
  assign n1991 = n1980 | n1990 ;
  assign n1992 = n1079 & ~n1202 ;
  buffer buf_n1993( .i (n1992), .o (n1993) );
  assign n1994 = n1074 & n1993 ;
  buffer buf_n1995( .i (n1994), .o (n1995) );
  assign n1996 = n1818 | n1995 ;
  buffer buf_n1859( .i (n1858), .o (n1859) );
  assign n1997 = n766 & n1859 ;
  assign n1998 = n1609 | n1997 ;
  assign n1999 = n1043 | n1998 ;
  buffer buf_n1415( .i (n1414), .o (n1415) );
  assign n2000 = n1308 | n1415 ;
  assign n2001 = ~n453 & n1373 ;
  buffer buf_n2002( .i (n2001), .o (n2002) );
  assign n2003 = n876 & ~n2002 ;
  buffer buf_n2004( .i (n2003), .o (n2004) );
  assign n2005 = n2000 | n2004 ;
  assign n2006 = n1999 | n2005 ;
  assign n2007 = n1996 | n2006 ;
  assign n2008 = n1991 | n2007 ;
  buffer buf_n2009( .i (n2008), .o (n2009) );
  assign n2010 = n1771 | n1785 ;
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n2012( .i (n2011), .o (n2012) );
  buffer buf_n2013( .i (n2012), .o (n2013) );
  buffer buf_n2014( .i (n2013), .o (n2014) );
  buffer buf_n2015( .i (n2014), .o (n2015) );
  assign n2016 = n1571 & n2015 ;
  assign n2017 = n1631 | n2016 ;
  assign n2018 = n293 & n992 ;
  buffer buf_n2019( .i (n2018), .o (n2019) );
  buffer buf_n2020( .i (n2019), .o (n2020) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n2021 = n186 & n800 ;
  assign n2022 = n929 & n2021 ;
  assign n2023 = n2020 | n2022 ;
  assign n2024 = n2017 | n2023 ;
  assign n2025 = n1933 | n2024 ;
  buffer buf_n160( .i (n159), .o (n160) );
  assign n2026 = ~n160 & n414 ;
  buffer buf_n2027( .i (n2026), .o (n2027) );
  assign n2028 = n366 & n1942 ;
  assign n2029 = n2027 & n2028 ;
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  assign n2031 = n600 | n1645 ;
  assign n2032 = n2030 & n2031 ;
  buffer buf_n2033( .i (n2032), .o (n2033) );
  assign n2034 = n1611 | n1724 ;
  buffer buf_n2035( .i (n2034), .o (n2035) );
  assign n2044 = n1905 | n2035 ;
  assign n2045 = n2033 | n2044 ;
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  assign n2048 = n2025 | n2047 ;
  assign n2049 = n2009 | n2048 ;
  assign n2050 = n1978 | n2049 ;
  assign n2051 = n1962 | n2050 ;
  assign n2052 = n1549 | n1707 ;
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  buffer buf_n2055( .i (n2054), .o (n2055) );
  buffer buf_n2056( .i (n2055), .o (n2056) );
  buffer buf_n2057( .i (n2056), .o (n2057) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  assign n2058 = n934 & n1431 ;
  assign n2059 = n1421 | n2058 ;
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  assign n2064 = n1386 | n2063 ;
  assign n2065 = n1619 | n2064 ;
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  assign n2066 = n371 & n664 ;
  buffer buf_n187( .i (n186), .o (n187) );
  assign n2067 = n187 | n223 ;
  buffer buf_n2068( .i (n2067), .o (n2068) );
  assign n2069 = n2066 & n2068 ;
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  assign n2070 = n424 | n1856 ;
  assign n2071 = n1154 & n2070 ;
  buffer buf_n2072( .i (n2071), .o (n2072) );
  assign n2073 = n1399 | n2072 ;
  assign n2074 = n1907 | n2073 ;
  assign n2075 = n2069 | n2074 ;
  buffer buf_n2076( .i (n2075), .o (n2076) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  assign n2077 = n1948 & n1957 ;
  assign n2078 = n1981 | n2077 ;
  assign n2079 = n1965 | n2033 ;
  buffer buf_n2080( .i (n2079), .o (n2080) );
  buffer buf_n2081( .i (n2080), .o (n2081) );
  assign n2082 = n2078 | n2081 ;
  assign n2083 = n2076 | n2082 ;
  buffer buf_n2084( .i (n2083), .o (n2084) );
  assign n2085 = n2065 | n2084 ;
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n988( .i (n987), .o (n988) );
  assign n2086 = n558 & n988 ;
  assign n2087 = n1360 | n2086 ;
  buffer buf_n2088( .i (n2087), .o (n2088) );
  assign n2089 = n1382 | n2088 ;
  buffer buf_n2090( .i (n2089), .o (n2090) );
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  assign n2096 = n1560 | n1660 ;
  buffer buf_n2097( .i (n2096), .o (n2097) );
  assign n2098 = n1698 | n2097 ;
  buffer buf_n2099( .i (n2098), .o (n2099) );
  buffer buf_n2100( .i (n2099), .o (n2100) );
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n517( .i (n516), .o (n517) );
  assign n2102 = n517 & n716 ;
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  assign n2105 = n1255 | n1803 ;
  assign n2106 = n1727 | n2105 ;
  assign n2107 = n2104 | n2106 ;
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n68( .i (x7), .o (n68) );
  buffer buf_n135( .i (x16), .o (n135) );
  assign n2108 = n68 & ~n135 ;
  buffer buf_n70( .i (x8), .o (n70) );
  assign n2109 = n70 & n135 ;
  assign n2110 = n2108 | n2109 ;
  buffer buf_n2111( .i (n2110), .o (n2111) );
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  assign n2119 = n1041 & n2118 ;
  assign n2120 = n611 & n2119 ;
  assign n2121 = n1246 | n2120 ;
  assign n2122 = n2107 | n2121 ;
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  assign n2125 = n53 & ~n2030 ;
  assign n2126 = n375 & n581 ;
  assign n2127 = ( n376 & n608 ) | ( n376 & n2126 ) | ( n608 & n2126 ) ;
  buffer buf_n2128( .i (n2127), .o (n2128) );
  assign n2129 = n2125 & n2128 ;
  buffer buf_n2130( .i (n2129), .o (n2130) );
  assign n2131 = n1957 | n2130 ;
  assign n2132 = n243 & n581 ;
  buffer buf_n2133( .i (n2132), .o (n2133) );
  assign n2135 = n2117 & n2133 ;
  buffer buf_n2136( .i (n2135), .o (n2136) );
  assign n2137 = n1571 | n1720 ;
  assign n2138 = n2136 | n2137 ;
  assign n2139 = n222 & n369 ;
  assign n2140 = n663 & n2139 ;
  assign n2141 = n2072 | n2140 ;
  assign n2142 = n2138 | n2141 ;
  assign n2143 = n2131 | n2142 ;
  buffer buf_n2144( .i (n2143), .o (n2144) );
  assign n2145 = n1823 | n2081 ;
  assign n2146 = n2144 | n2145 ;
  assign n2147 = n2124 | n2146 ;
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  assign n2149 = n808 & ~n886 ;
  buffer buf_n2150( .i (n2149), .o (n2150) );
  assign n2151 = n524 | n2150 ;
  buffer buf_n2152( .i (n2151), .o (n2152) );
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  assign n2155 = n742 | n2154 ;
  buffer buf_n804( .i (n803), .o (n804) );
  assign n2156 = n804 & n883 ;
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n2158( .i (n2157), .o (n2158) );
  assign n2159 = n754 | n791 ;
  buffer buf_n2160( .i (n2159), .o (n2160) );
  assign n2161 = n2158 | n2160 ;
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n2163( .i (n2162), .o (n2163) );
  buffer buf_n2164( .i (n2163), .o (n2164) );
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n2166( .i (n2165), .o (n2166) );
  buffer buf_n2167( .i (n2166), .o (n2167) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  assign n2168 = n121 | n1412 ;
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n104( .i (x12), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  assign n2172 = n105 | n108 ;
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n2175( .i (n2174), .o (n2175) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  buffer buf_n2177( .i (n2176), .o (n2177) );
  assign n2178 = n175 & ~n2177 ;
  assign n2179 = ~n2169 & n2178 ;
  buffer buf_n2180( .i (n2179), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  buffer buf_n2182( .i (n2181), .o (n2182) );
  buffer buf_n2183( .i (n2182), .o (n2183) );
  buffer buf_n2184( .i (n2183), .o (n2184) );
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  buffer buf_n2187( .i (n2186), .o (n2187) );
  buffer buf_n2188( .i (n2187), .o (n2188) );
  assign n2189 = n650 | n1020 ;
  buffer buf_n535( .i (n534), .o (n535) );
  assign n2190 = n535 & n720 ;
  buffer buf_n2191( .i (n2190), .o (n2191) );
  buffer buf_n2192( .i (n2191), .o (n2192) );
  buffer buf_n2193( .i (n2192), .o (n2193) );
  assign n2194 = n1560 | n2193 ;
  assign n2195 = n2189 | n2194 ;
  buffer buf_n2196( .i (n2195), .o (n2196) );
  buffer buf_n2197( .i (n2196), .o (n2197) );
  buffer buf_n2198( .i (n2197), .o (n2198) );
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  assign n2200 = n688 & n1033 ;
  assign n2201 = n735 | n2200 ;
  buffer buf_n2202( .i (n2201), .o (n2202) );
  buffer buf_n2203( .i (n2202), .o (n2203) );
  assign n2204 = n561 | n1032 ;
  assign n2205 = n1041 & n2204 ;
  buffer buf_n2206( .i (n2205), .o (n2206) );
  buffer buf_n2207( .i (n2206), .o (n2207) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  assign n2208 = n1510 | n1891 ;
  assign n2209 = n2207 | n2208 ;
  assign n2210 = n2203 | n2209 ;
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  assign n2211 = n513 & n1669 ;
  assign n2212 = n2004 | n2211 ;
  assign n2213 = n266 & n928 ;
  assign n2214 = ~n99 & n1121 ;
  buffer buf_n2215( .i (n2214), .o (n2215) );
  buffer buf_n2216( .i (n2215), .o (n2216) );
  assign n2217 = n2213 & n2216 ;
  assign n2218 = n2212 | n2217 ;
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  assign n2221 = n781 | n2220 ;
  assign n2222 = n2210 | n2221 ;
  buffer buf_n2223( .i (n2222), .o (n2223) );
  buffer buf_n2224( .i (n1038), .o (n2224) );
  assign n2225 = ~n2002 & n2224 ;
  buffer buf_n2226( .i (n2225), .o (n2226) );
  assign n2228 = n799 & n927 ;
  assign n2229 = ~n98 & n219 ;
  assign n2230 = ( n264 & n1152 ) | ( n264 & n2229 ) | ( n1152 & n2229 ) ;
  buffer buf_n2231( .i (n2230), .o (n2231) );
  assign n2232 = n2228 & n2231 ;
  assign n2233 = n2226 | n2232 ;
  assign n2234 = n701 | n2233 ;
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  assign n2235 = n402 | n722 ;
  assign n2236 = n1515 | n2235 ;
  assign n2237 = n2234 | n2236 ;
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  assign n2240 = n1109 | n1538 ;
  assign n2241 = n2239 | n2240 ;
  assign n2242 = n1227 | n2241 ;
  assign n2243 = n2223 | n2242 ;
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n2244( .i (n965), .o (n2244) );
  assign n2245 = n605 & n2244 ;
  assign n2246 = n1146 | n2245 ;
  assign n2247 = n807 | n2246 ;
  assign n2248 = n2160 | n2247 ;
  buffer buf_n2249( .i (n2248), .o (n2249) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n28( .i (n27), .o (n28) );
  assign n2250 = n28 | n33 ;
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  assign n2255 = n571 | n2254 ;
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  assign n2257 = ~n234 & n368 ;
  assign n2258 = n638 & n2257 ;
  assign n2259 = ( n370 & ~n2256 ) | ( n370 & n2258 ) | ( ~n2256 & n2258 ) ;
  assign n2260 = n1682 | n2259 ;
  assign n2261 = n523 | n2260 ;
  assign n2262 = n2249 | n2261 ;
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  assign n2263 = n184 | n1137 ;
  buffer buf_n2264( .i (n2263), .o (n2264) );
  buffer buf_n2265( .i (n2264), .o (n2265) );
  assign n2266 = n1432 & n2265 ;
  assign n2267 = ~n66 & n661 ;
  assign n2268 = n727 & n2267 ;
  buffer buf_n2269( .i (n2268), .o (n2269) );
  assign n2270 = n2266 | n2269 ;
  assign n2271 = n779 | n2270 ;
  assign n2272 = n624 | n2271 ;
  assign n2273 = n2262 | n2272 ;
  buffer buf_n2274( .i (n2273), .o (n2274) );
  buffer buf_n2275( .i (n2274), .o (n2275) );
  buffer buf_n345( .i (n344), .o (n345) );
  assign n2276 = n319 & n345 ;
  assign n2277 = ~n1085 & n2276 ;
  buffer buf_n2278( .i (n2277), .o (n2278) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  buffer buf_n2280( .i (n2279), .o (n2280) );
  buffer buf_n2281( .i (n2280), .o (n2281) );
  assign n2282 = n1083 & n2281 ;
  assign n2283 = n1127 | n2282 ;
  assign n2284 = n919 | n2283 ;
  buffer buf_n2285( .i (n2284), .o (n2285) );
  assign n2286 = n1389 | n1609 ;
  buffer buf_n2287( .i (n2286), .o (n2287) );
  assign n2288 = n1876 | n2287 ;
  assign n2289 = n942 | n2288 ;
  buffer buf_n1838( .i (n1837), .o (n1838) );
  assign n2290 = n1435 | n1838 ;
  assign n2291 = n2289 | n2290 ;
  assign n2292 = n2285 | n2291 ;
  buffer buf_n2293( .i (n2292), .o (n2293) );
  buffer buf_n1972( .i (n1971), .o (n1972) );
  buffer buf_n1973( .i (n1972), .o (n1973) );
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  assign n2294 = n1649 | n1906 ;
  buffer buf_n2295( .i (n2294), .o (n2295) );
  assign n2296 = n1853 | n2295 ;
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  assign n2297 = n669 | n1549 ;
  assign n2298 = n1487 | n2297 ;
  assign n2299 = n2296 | n2298 ;
  assign n2300 = n1974 | n2299 ;
  assign n2301 = n2293 | n2300 ;
  assign n2302 = n2275 | n2301 ;
  assign n2303 = n1519 | n2249 ;
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  assign n2307 = n1219 | n2134 ;
  assign n2308 = ~n2136 & n2307 ;
  buffer buf_n2170( .i (n2169), .o (n2170) );
  buffer buf_n2171( .i (n2170), .o (n2171) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  assign n2309 = n113 | n174 ;
  buffer buf_n2310( .i (n2309), .o (n2310) );
  assign n2311 = n175 & n2177 ;
  assign n2312 = ( n1856 & n2310 ) | ( n1856 & ~n2311 ) | ( n2310 & ~n2311 ) ;
  assign n2313 = n1378 | n2312 ;
  assign n2314 = ~n2171 & n2313 ;
  assign n2315 = n1270 | n1547 ;
  assign n2316 = n2314 | n2315 ;
  assign n2317 = n2308 | n2316 ;
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  assign n2320 = n133 & n2128 ;
  buffer buf_n2321( .i (n2320), .o (n2321) );
  assign n2323 = ~n56 & n2321 ;
  buffer buf_n2324( .i (n2323), .o (n2324) );
  assign n2325 = n2285 | n2324 ;
  assign n2326 = n2319 | n2325 ;
  buffer buf_n1124( .i (n1123), .o (n1124) );
  assign n2327 = ~n102 & n1124 ;
  assign n2328 = n1238 | n2327 ;
  buffer buf_n2329( .i (n2328), .o (n2329) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  assign n2330 = n968 & n1033 ;
  buffer buf_n2331( .i (n2330), .o (n2331) );
  buffer buf_n2227( .i (n2226), .o (n2227) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n2332( .i (n179), .o (n2332) );
  buffer buf_n2333( .i (n2332), .o (n2333) );
  assign n2334 = n166 & n2333 ;
  buffer buf_n2335( .i (n2334), .o (n2335) );
  assign n2336 = n383 & n2335 ;
  buffer buf_n2337( .i (n2336), .o (n2337) );
  assign n2338 = n2224 & n2337 ;
  buffer buf_n2339( .i (n2338), .o (n2339) );
  assign n2340 = ~n2118 & n2339 ;
  assign n2341 = n2227 | n2340 ;
  assign n2342 = n2331 | n2341 ;
  assign n2343 = n2329 | n2342 ;
  assign n2344 = n403 | n576 ;
  buffer buf_n2345( .i (n2344), .o (n2345) );
  assign n2346 = n671 | n2206 ;
  assign n2347 = n2345 | n2346 ;
  assign n2348 = n2343 | n2347 ;
  buffer buf_n2349( .i (n2348), .o (n2349) );
  assign n2350 = n2326 | n2349 ;
  assign n2351 = n2306 | n2350 ;
  assign n2352 = n2238 | n2318 ;
  assign n2353 = n1212 | n1740 ;
  assign n2354 = n671 | n1026 ;
  assign n2355 = n2353 | n2354 ;
  assign n2356 = n1756 | n2355 ;
  assign n2357 = n2352 | n2356 ;
  assign n2358 = n2274 | n2357 ;
  assign n2359 = n1977 | n2144 ;
  buffer buf_n2322( .i (n2321), .o (n2322) );
  assign n2360 = n2046 | n2322 ;
  buffer buf_n728( .i (n727), .o (n728) );
  assign n2361 = n663 & n728 ;
  buffer buf_n2362( .i (n2361), .o (n2362) );
  assign n2363 = n175 & n220 ;
  assign n2364 = n1288 & n2363 ;
  buffer buf_n2365( .i (n2364), .o (n2365) );
  assign n2366 = n2339 | n2365 ;
  assign n2367 = n922 | n2366 ;
  assign n2368 = n2362 | n2367 ;
  assign n2369 = n1842 | n2368 ;
  assign n2370 = n2360 | n2369 ;
  assign n2371 = n2009 | n2370 ;
  assign n2372 = n2359 | n2371 ;
  assign n2373 = n2358 | n2372 ;
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n695( .i (n694), .o (n695) );
  assign n2374 = n664 & n695 ;
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  assign n2375 = n767 & n934 ;
  assign n2376 = n544 & n2375 ;
  assign n2377 = n646 | n2376 ;
  assign n2378 = n2374 | n2377 ;
  buffer buf_n2379( .i (n2378), .o (n2379) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  assign n2380 = n728 | n968 ;
  assign n2381 = ~n1656 & n2380 ;
  buffer buf_n2382( .i (n2381), .o (n2382) );
  assign n2383 = n460 | n2382 ;
  assign n2384 = n2379 | n2383 ;
  buffer buf_n832( .i (n831), .o (n832) );
  assign n2385 = n687 | n967 ;
  buffer buf_n2386( .i (n2385), .o (n2386) );
  buffer buf_n2387( .i (n2386), .o (n2387) );
  buffer buf_n837( .i (n836), .o (n837) );
  assign n2388 = n837 & n2386 ;
  assign n2389 = ( n832 & n2387 ) | ( n832 & n2388 ) | ( n2387 & n2388 ) ;
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  assign n2390 = ~n153 & n602 ;
  assign n2391 = ( ~n578 & n580 ) | ( ~n578 & n2390 ) | ( n580 & n2390 ) ;
  buffer buf_n2392( .i (n2391), .o (n2392) );
  buffer buf_n2393( .i (n2392), .o (n2393) );
  buffer buf_n2394( .i (n2393), .o (n2394) );
  buffer buf_n2395( .i (n2394), .o (n2395) );
  buffer buf_n514( .i (n513), .o (n514) );
  assign n2396 = n221 | n933 ;
  assign n2397 = n434 & n2396 ;
  assign n2398 = n514 | n2397 ;
  assign n2399 = n2395 | n2398 ;
  assign n2400 = n372 & n2399 ;
  assign n2401 = n2389 | n2400 ;
  assign n2402 = ~n16 & n2401 ;
  assign n2403 = ( ~n17 & n2384 ) | ( ~n17 & n2402 ) | ( n2384 & n2402 ) ;
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  assign n2404 = n542 & n863 ;
  assign n2405 = n388 | n2404 ;
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  assign n2406 = n23 | n166 ;
  assign n2407 = n1111 & ~n2406 ;
  buffer buf_n2408( .i (n2407), .o (n2408) );
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  buffer buf_n2411( .i (n2410), .o (n2411) );
  assign n2412 = n2405 & n2411 ;
  assign n2413 = ~n6 & n554 ;
  assign n2414 = n429 | n653 ;
  assign n2415 = n2413 & n2414 ;
  assign n2416 = ~n1230 & n2415 ;
  buffer buf_n2417( .i (n2416), .o (n2417) );
  buffer buf_n2418( .i (n2417), .o (n2418) );
  buffer buf_n384( .i (n383), .o (n384) );
  assign n2419 = n183 & ~n1643 ;
  assign n2420 = n384 & ~n2419 ;
  assign n2421 = n1140 & ~n2420 ;
  assign n2422 = n2418 & n2421 ;
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  assign n2423 = n420 & ~n1554 ;
  buffer buf_n2424( .i (n2423), .o (n2424) );
  buffer buf_n2425( .i (n2424), .o (n2425) );
  assign n2426 = n266 | n2425 ;
  assign n2427 = ~n535 & n2424 ;
  assign n2428 = n266 & n2427 ;
  assign n2429 = ( n2422 & ~n2426 ) | ( n2422 & n2428 ) | ( ~n2426 & n2428 ) ;
  assign n2430 = n2412 | n2429 ;
  buffer buf_n2431( .i (n2430), .o (n2431) );
  buffer buf_n2432( .i (n2431), .o (n2432) );
  buffer buf_n2433( .i (n2432), .o (n2433) );
  buffer buf_n2434( .i (n2433), .o (n2434) );
  assign n2435 = n2403 | n2434 ;
  buffer buf_n2436( .i (n2435), .o (n2436) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  assign n2437 = n1024 | n1166 ;
  assign n2438 = ~n1447 & n1740 ;
  assign n2439 = n2437 | n2438 ;
  buffer buf_n2440( .i (n2439), .o (n2440) );
  buffer buf_n2441( .i (n2440), .o (n2441) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  assign n2443 = n1567 | n2442 ;
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  assign n2444 = n1694 | n2130 ;
  assign n2445 = n1661 | n2444 ;
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n2448( .i (n2447), .o (n2448) );
  buffer buf_n2449( .i (n2448), .o (n2449) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n2036( .i (n2035), .o (n2036) );
  buffer buf_n2037( .i (n2036), .o (n2037) );
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  assign y0 = n466 ;
  assign y1 = n473 ;
  assign y2 = 1'b0 ;
  assign y3 = n485 ;
  assign y4 = n497 ;
  assign y5 = n529 ;
  assign y6 = n815 ;
  assign y7 = n824 ;
  assign y8 = n858 ;
  assign y9 = n708 ;
  assign y10 = n1187 ;
  assign y11 = n1283 ;
  assign y12 = n1317 ;
  assign y13 = n1468 ;
  assign y14 = n1542 ;
  assign y15 = n1705 ;
  assign y16 = n1761 ;
  assign y17 = n1827 ;
  assign y18 = n1884 ;
  assign y19 = n1940 ;
  assign y20 = n898 ;
  assign y21 = n910 ;
  assign y22 = n2051 ;
  assign y23 = n2057 ;
  assign y24 = n1734 ;
  assign y25 = n2085 ;
  assign y26 = n2095 ;
  assign y27 = n2101 ;
  assign y28 = n2148 ;
  assign y29 = n2155 ;
  assign y30 = n2167 ;
  assign y31 = n785 ;
  assign y32 = n2188 ;
  assign y33 = n2199 ;
  assign y34 = n2243 ;
  assign y35 = n2302 ;
  assign y36 = n2351 ;
  assign y37 = n2373 ;
  assign y38 = n2436 ;
  assign y39 = n2443 ;
  assign y40 = n2449 ;
  assign y41 = n621 ;
  assign y42 = 1'b0 ;
  assign y43 = n2043 ;
  assign y44 = n1734 ;
endmodule
