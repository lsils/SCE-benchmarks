module top( G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G6 , G7 , G8 , G9 , G3519 , G3520 , G3521 , G3522 , G3523 , G3524 , G3525 , G3526 , G3527 , G3528 , G3529 , G3530 , G3531 , G3532 , G3533 , G3534 , G3535 , G3536 , G3537 , G3538 , G3539 , G3540 );
  input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G6 , G7 , G8 , G9 ;
  output G3519 , G3520 , G3521 , G3522 , G3523 , G3524 , G3525 , G3526 , G3527 , G3528 , G3529 , G3530 , G3531 , G3532 , G3533 , G3534 , G3535 , G3536 , G3537 , G3538 , G3539 , G3540 ;
  wire n686 , n688 , n692 , n743 , n745 , n795 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n816 , n820 , n822 , n830 , n835 , n837 , n838 , n839 , n840 , n841 , n884 , n885 , n886 , n888 , n889 , n890 , n892 , n893 , n894 , n896 , n897 , n898 , n900 , n901 , n902 , n904 , n905 , n906 , n908 , n909 , n910 , n956 , n957 , n959 , n960 , n962 , n963 , n964 , n966 , n967 , n968 , n970 , n971 , n972 , n974 , n975 , n976 , n978 , n979 , n980 , n1025 , n1031 , n1032 , n1037 , n1039 , n1040 , n1041 , n1045 , n1047 , n1048 , n1049 , n1050 , n1053 , n1055 , n1056 , n1059 , n1060 , n1061 , n1062 , n1065 , n1068 , n1080 , n1082 , n1089 , n1095 , n1099 , n1101 , n1103 , n1105 , n1108 , n1109 , n1111 , n1112 , n1113 , n1114 , n1115 , n1118 , n1120 , n1121 , n1123 , n1128 , n1129 , n1132 , n1134 , n1135 , n1136 , n1137 , n1138 , n1140 , n1149 , n1150 , n1151 , n1152 , n1156 , n1159 , n1161 , n1164 , n1166 , n1167 , n1168 , n1169 , n1170 , n1173 , n1175 , n1176 , n1178 , n1179 , n1181 , n1183 , n1185 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1194 , n1195 , n1198 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1212 , n1214 , n1215 , n1217 , n1218 , n1220 , n1232 , n1234 , n1235 , n1236 , n1237 , n1238 , n1241 , n1242 , n1244 , n1247 , n1249 , n1250 , n1254 , n1255 , n1256 , n1257 , n1258 , n1261 , n1263 , n1264 , n1266 , n1267 , n1270 , n1272 , n1274 , n1282 , n1283 , n1285 , n1286 , n1287 , n1288 , n1289 , n1292 , n1293 , n1294 , n1296 , n1297 , n1298 , n1299 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1308 , n1309 , n1310 , n1312 , n1313 , n1315 , n1318 , n1322 , n1325 , n1328 , n1332 , n1333 , n1334 , n1335 , n1336 , n1341 , n1342 , n1344 , n1345 , n1346 , n1350 , n1351 , n1354 , n1359 , n1361 , n1363 , n1365 , n1366 , n1367 , n1368 , n1369 , n1371 , n1374 , n1377 , n1378 , n1381 , n1382 , n1384 , n1386 , n1388 , n1389 , n1390 , n1391 , n1392 , n1396 , n1398 , n1400 , n1401 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1411 , n1413 , n1414 , n1420 , n1421 , n1423 , n1427 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1439 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1452 , n1454 , n1455 , n1463 , n1464 , n1466 , n1472 , n1474 , n1504 , n1505 , n1506 , n1507 , n1511 , n1513 , n1515 , n1516 , n1517 , n1520 , n1521 , n1522 , n1526 , n1534 , n1562 , n1604 , n1620 , n1624 , n1625 , n1626 , n1629 , n1634 , n1635 , n1636 , n1638 , n1639 , n1671 , n1700 , n1717 , n1725 , n1726 , n1753 , n1769 , n1770 , n1791 , n1792 , n1806 , n1810 , n1812 , n1814 , n1820 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1830 , n1833 , n1835 , n1838 , n1839 , n1840 , n1844 , n1852 , n1853 , n1859 , n1868 , n1869 , n1870 , n1871 , n1874 , n1879 , n1881 , n1885 , n1886 , n1888 , n1889 , n1890 , n1891 , n1893 , n1894 , n1895 , n1896 , n1898 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1913 , n1915 , n1919 , n1920 , n1921 , n1922 , n1952 , n1957 , n1958 , n1959 , n1969 , n1971 , n1972 , n1973 , n1975 , n1976 , n1977 , n1981 , n1982 , n1983 , n1984 , n1985 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1997 , n1998 , n1999 , n2002 , n2003 , n2006 , n2007 , n2010 , n2011 , n2012 , n2013 , n2014 , n2019 , n2031 , n2032 , n2033 , n2035 , n2037 , n2038 , n2041 , n2042 , n2043 , n2044 , n2053 , n2054 , n2056 , n2060 , n2062 , n2063 , n2065 , n2067 , n2068 , n2069 , n2070 , n2090 , n2094 , n2098 , n2099 , n2100 , n2111 , n2119 , n2126 , n2131 , n2132 , n2133 , n2138 , n2145 , n2146 , n2147 , n2151 , n2155 , n2156 , n2158 , n2164 , n2177 , n2178 , n2180 , n2182 , n2192 , n2197 , n2198 , n2199 , n2201 , n2202 , n2203 , n2204 , n2206 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2243 , n2272 , n2289 , n2290 , n2325 , n2330 , n2332 , n2337 , n2339 , n2340 , n2341 , n2343 , n2344 , n2349 , n2354 , n2355 , n2356 , n2362 , n2369 , n2371 , n2373 , n2375 , n2377 , n2379 , n2382 , n2384 , n2385 , n2386 , n2387 , n2398 , n2401 , n2405 , n2406 , n2407 , n2418 , n2419 , n2420 , n2422 , n2423 , n2424 , n2427 , n2428 , n2429 , n2432 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2452 , n2453 , n2456 , n2457 , n2458 , n2460 , n2462 , n2463 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2476 , n2492 , n2510 , n2513 , n2514 , n2515 , n2516 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2528 , n2529 , n2530 , n2534 , n2536 , n2537 , n2538 , n2541 , n2542 , n2543 , n2546 , n2549 , n2550 , n2553 , n2558 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2570 , n2577 , n2580 , n2602 , n2605 , n2607 , n2608 , n2609 , n2610 , n2612 , n2613 , n2614 , n2618 , n2619 , n2620 , n2622 , n2627 , n2628 , n2631 , n2632 , n2633 , n2634 , n2636 , n2637 , n2638 , n2639 , n2641 , n2645 , n2646 , n2649 , n2650 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2662 , n2674 , n2675 , n2677 , n2678 , n2679 , n2698 , n2700 , n2702 , n2704 , n2709 , n2710 , n2718 , n2722 , n2723 , n2724 , n2726 , n2727 , n2728 , n2730 , n2735 , n2737 , n2738 , n2739 , n2741 , n2743 , n2744 , n2747 , n2750 , n2751 , n2754 , n2755 , n2757 , n2759 , n2760 , n2761 , n2762 , n2763 , n2765 , n2766 , n2770 , n2771 , n2773 , n2774 , n2775 , n2776 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2788 , n2807 , n2808 , n2820 , n2825 , n2826 , n2827 , n2836 , n2837 , n2839 , n2844 , n2848 , n2849 , n2851 , n2852 , n2861 , n2862 , n2863 , n2864 , n2867 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2877 , n2878 , n2879 , n2881 , n2882 , n2884 , n2885 , n2886 , n2887 , n2891 , n2910 , n2914 , n2915 , n2918 , n2919 , n2920 , n2921 , n2922 , n2925 , n2926 , n2927 , n2934 , n2935 , n2948 , n2949 , n2950 , n2953 , n2954 , n2955 , n2956 , n2957 , n2959 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2970 , n2973 , n2974 , n2975 , n2976 , n2977 , n2980 , n2981 , n2983 , n2984 , n2985 , n2987 , n2988 , n2991 , n2995 , n3010 , n3011 , n3015 , n3028 , n3030 , n3032 , n3034 , n3041 , n3045 , n3046 , n3054 , n3057 , n3058 , n3063 , n3065 , n3067 , n3069 , n3076 , n3078 , n3080 , n3081 , n3082 , n3085 , n3086 , n3087 , n3091 , n3093 , n3097 , n3099 , n3100 , n3101 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 ;
  buffer buf_n661( .i (G8), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n672( .i (G9), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  assign n686 = n662 | n673 ;
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n79( .i (G10), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n648( .i (G7), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  assign n688 = n80 | n649 ;
  buffer buf_n689( .i (n688), .o (n689) );
  assign n692 = n687 | n689 ;
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n92( .i (G11), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n104( .i (G12), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n118( .i (G13), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  assign n743 = n106 | n120 ;
  buffer buf_n744( .i (n743), .o (n744) );
  assign n745 = n96 & n744 ;
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n51( .i (G1), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n330( .i (G3), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  assign n795 = n56 | n335 ;
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n352( .i (G32), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  assign n797 = n355 & ~n675 ;
  buffer buf_n346( .i (G31), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  assign n798 = n349 & ~n664 ;
  assign n799 = n797 | n798 ;
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n381( .i (G36), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  assign n800 = ~n121 & n384 ;
  buffer buf_n131( .i (G14), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n389( .i (G37), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  assign n801 = ~n134 & n392 ;
  assign n802 = n800 | n801 ;
  assign n803 = n799 | n802 ;
  buffer buf_n364( .i (G34), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  assign n804 = ~n95 & n367 ;
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n373( .i (G35), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  assign n805 = ~n107 & n376 ;
  assign n806 = n804 | n805 ;
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n358( .i (G33), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  assign n807 = ~n82 & n361 ;
  buffer buf_n340( .i (G30), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  assign n808 = n343 & ~n651 ;
  assign n809 = n807 | n808 ;
  assign n810 = n806 | n809 ;
  assign n811 = n803 | n810 ;
  assign n812 = n796 & n811 ;
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n185( .i (G2), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n816 = ~n52 & n186 ;
  buffer buf_n817( .i (n816), .o (n817) );
  assign n820 = ~n333 & n817 ;
  buffer buf_n821( .i (n820), .o (n821) );
  assign n822 = ~n651 & n687 ;
  buffer buf_n823( .i (n822), .o (n823) );
  assign n830 = n821 & n823 ;
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  assign n835 = n192 | n796 ;
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  assign n837 = n380 | n388 ;
  assign n838 = n372 & n837 ;
  assign n839 = ~n836 & n838 ;
  assign n840 = n834 | n839 ;
  assign n841 = n815 | n840 ;
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  assign n884 = n382 | n390 ;
  assign n885 = n382 & n390 ;
  assign n886 = n884 & ~n885 ;
  buffer buf_n887( .i (n886), .o (n887) );
  assign n888 = n365 & ~n374 ;
  assign n889 = ~n365 & n374 ;
  assign n890 = n888 | n889 ;
  buffer buf_n891( .i (n890), .o (n891) );
  assign n892 = n887 | n891 ;
  assign n893 = n887 & n891 ;
  assign n894 = n892 & ~n893 ;
  buffer buf_n895( .i (n894), .o (n895) );
  assign n896 = n341 & ~n347 ;
  assign n897 = ~n341 & n347 ;
  assign n898 = n896 | n897 ;
  buffer buf_n899( .i (n898), .o (n899) );
  assign n900 = n353 | n359 ;
  assign n901 = n353 & n359 ;
  assign n902 = n900 & ~n901 ;
  buffer buf_n903( .i (n902), .o (n903) );
  assign n904 = n899 | n903 ;
  assign n905 = n899 & n903 ;
  assign n906 = n904 & ~n905 ;
  buffer buf_n907( .i (n906), .o (n907) );
  assign n908 = n895 | n907 ;
  assign n909 = n895 & n907 ;
  assign n910 = n908 & ~n909 ;
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  assign n956 = n663 & n674 ;
  assign n957 = n687 & ~n956 ;
  buffer buf_n958( .i (n957), .o (n958) );
  assign n959 = n81 & n650 ;
  assign n960 = n689 & ~n959 ;
  buffer buf_n961( .i (n960), .o (n961) );
  assign n962 = ~n958 & n961 ;
  assign n963 = n958 & ~n961 ;
  assign n964 = n962 | n963 ;
  buffer buf_n965( .i (n964), .o (n965) );
  assign n966 = ~n94 & n120 ;
  assign n967 = n94 & ~n120 ;
  assign n968 = n966 | n967 ;
  buffer buf_n969( .i (n968), .o (n969) );
  assign n970 = n106 | n133 ;
  assign n971 = n106 & n133 ;
  assign n972 = n970 & ~n971 ;
  buffer buf_n973( .i (n972), .o (n973) );
  assign n974 = n969 & ~n973 ;
  assign n975 = ~n969 & n973 ;
  assign n976 = n974 | n975 ;
  buffer buf_n977( .i (n976), .o (n977) );
  assign n978 = n965 & n977 ;
  assign n979 = n965 | n977 ;
  assign n980 = ~n978 & n979 ;
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  assign n1025 = n333 & n817 ;
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  assign n1031 = n657 | n1030 ;
  assign n1032 = ~n53 & n332 ;
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  assign n1037 = n53 & n187 ;
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n418( .i (G4), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  assign n1039 = n53 & n332 ;
  assign n1040 = n421 & n1039 ;
  assign n1041 = n1038 | n1040 ;
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  assign n1045 = n1036 | n1043 ;
  buffer buf_n1046( .i (n1045), .o (n1046) );
  assign n1047 = n657 & n1046 ;
  assign n1048 = n1031 & ~n1047 ;
  buffer buf_n1044( .i (n1043), .o (n1044) );
  assign n1049 = n651 | n687 ;
  assign n1050 = n334 & n1049 ;
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n218( .i (G21), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  assign n1053 = n333 | n421 ;
  buffer buf_n1054( .i (n1053), .o (n1054) );
  assign n1055 = n223 & ~n1054 ;
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  assign n1056 = ~n332 & n420 ;
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  assign n1059 = ~n666 & n1058 ;
  assign n1060 = n1055 | n1059 ;
  assign n1061 = n1052 | n1060 ;
  assign n1062 = n1044 & n1061 ;
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  assign n1065 = n1048 | n1064 ;
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n261( .i (G25), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n264( .i (G26), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  assign n1068 = n262 | n265 ;
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n572( .i (G5), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n636( .i (G6), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  assign n1080 = n573 | n637 ;
  buffer buf_n1081( .i (n52), .o (n1081) );
  assign n1082 = n1080 & ~n1081 ;
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n396( .i (G38), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n574( .i (n573), .o (n574) );
  assign n1089 = n420 & n574 ;
  buffer buf_n1090( .i (n1089), .o (n1090) );
  assign n1095 = n1038 & ~n1090 ;
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  assign n1099 = n403 & ~n1097 ;
  buffer buf_n1100( .i (n1099), .o (n1100) );
  assign n1101 = n1088 & n1100 ;
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  assign n1103 = n345 & ~n1084 ;
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n318( .i (G28), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n569( .i (G49), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  assign n1105 = n420 | n571 ;
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  assign n1108 = n323 & ~n1107 ;
  assign n1109 = n82 & ~n421 ;
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n324( .i (G29), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n422( .i (n421), .o (n422) );
  assign n1111 = n328 & n422 ;
  assign n1112 = n1110 | n1111 ;
  assign n1113 = n1108 | n1112 ;
  assign n1114 = n1104 | n1113 ;
  assign n1115 = ~n1098 & n1114 ;
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  assign n1118 = n1102 | n1117 ;
  buffer buf_n1119( .i (n1118), .o (n1119) );
  assign n1120 = n1079 & ~n1119 ;
  assign n1121 = n1067 | n1120 ;
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n241( .i (G23), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (G24), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  assign n1123 = n249 | n258 ;
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  assign n1128 = ~n1119 & n1127 ;
  assign n1129 = n1067 & n1128 ;
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n1132 = n1122 & ~n1130 ;
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  assign n1134 = n670 & n1046 ;
  assign n1135 = n670 | n1030 ;
  assign n1136 = ~n1134 & n1135 ;
  assign n1137 = n335 & n958 ;
  buffer buf_n676( .i (n675), .o (n676) );
  assign n1138 = ~n676 & n1057 ;
  buffer buf_n230( .i (G22), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n1139( .i (n331), .o (n1139) );
  assign n1140 = n232 & ~n1139 ;
  buffer buf_n1141( .i (n1140), .o (n1141) );
  assign n1149 = ~n422 & n1141 ;
  assign n1150 = n1138 | n1149 ;
  assign n1151 = n1137 | n1150 ;
  assign n1152 = n1043 & n1151 ;
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  assign n1156 = n1136 | n1155 ;
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  assign n1159 = n351 & ~n1084 ;
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n329( .i (n328), .o (n329) );
  assign n1161 = n329 & ~n1107 ;
  buffer buf_n1162( .i (n419), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  assign n1164 = n95 | n1163 ;
  buffer buf_n1165( .i (n1164), .o (n1165) );
  assign n1166 = ~n344 & n422 ;
  assign n1167 = n1165 & ~n1166 ;
  assign n1168 = n1161 | n1167 ;
  assign n1169 = n1160 | n1168 ;
  assign n1170 = ~n1098 & n1169 ;
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  assign n1173 = n1102 | n1172 ;
  buffer buf_n1174( .i (n1173), .o (n1174) );
  assign n1175 = n1079 & ~n1174 ;
  assign n1176 = n1158 | n1175 ;
  buffer buf_n1177( .i (n1176), .o (n1177) );
  assign n1178 = n1127 & ~n1174 ;
  assign n1179 = n1158 & n1178 ;
  buffer buf_n1180( .i (n1179), .o (n1180) );
  assign n1181 = n1177 & ~n1180 ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  assign n1183 = n1133 & n1182 ;
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  assign n1185 = n337 & n1043 ;
  buffer buf_n1186( .i (n1185), .o (n1186) );
  assign n1187 = n1046 & ~n1186 ;
  assign n1188 = n89 & ~n1187 ;
  assign n1189 = ~n86 & n1028 ;
  assign n1190 = n666 | n1054 ;
  buffer buf_n97( .i (n96), .o (n97) );
  assign n1191 = ~n97 & n1058 ;
  assign n1192 = n1190 & ~n1191 ;
  buffer buf_n1193( .i (n1042), .o (n1193) );
  assign n1194 = ~n1192 & n1193 ;
  assign n1195 = n1189 | n1194 ;
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  assign n1198 = n1188 | n1197 ;
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  assign n1201 = n363 & ~n1084 ;
  assign n1202 = n350 & ~n1106 ;
  assign n1203 = n121 | n1163 ;
  assign n1204 = ~n355 & n1163 ;
  assign n1205 = n1203 & ~n1204 ;
  assign n1206 = n1202 | n1205 ;
  assign n1207 = n1201 | n1206 ;
  assign n1208 = ~n1097 & n1207 ;
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  assign n1212 = n1102 | n1211 ;
  buffer buf_n1213( .i (n1212), .o (n1213) );
  assign n1214 = n1079 & ~n1213 ;
  assign n1215 = n1200 | n1214 ;
  buffer buf_n1216( .i (n1215), .o (n1216) );
  assign n1217 = n1127 & ~n1213 ;
  assign n1218 = n1200 & n1217 ;
  buffer buf_n1219( .i (n1218), .o (n1219) );
  assign n1220 = n1216 & ~n1219 ;
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  assign n1232 = n1030 | n1186 ;
  buffer buf_n1233( .i (n1232), .o (n1233) );
  assign n1234 = ~n683 & n1233 ;
  assign n1235 = n653 & ~n1054 ;
  assign n1236 = n84 & n1058 ;
  assign n1237 = n1235 | n1236 ;
  assign n1238 = n1193 & n1237 ;
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  assign n1241 = n681 & ~n1046 ;
  assign n1242 = n1240 | n1241 ;
  buffer buf_n1243( .i (n1242), .o (n1243) );
  assign n1244 = n1234 | n1243 ;
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n1246( .i (n1083), .o (n1246) );
  assign n1247 = n357 & ~n1246 ;
  buffer buf_n1248( .i (n1247), .o (n1248) );
  assign n1249 = n345 & ~n1107 ;
  assign n1250 = n107 | n1163 ;
  buffer buf_n1251( .i (n1250), .o (n1251) );
  buffer buf_n1252( .i (n1162), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  assign n1254 = ~n350 & n1253 ;
  assign n1255 = n1251 & ~n1254 ;
  assign n1256 = n1249 | n1255 ;
  assign n1257 = n1248 | n1256 ;
  assign n1258 = ~n1098 & n1257 ;
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  assign n1261 = n1102 | n1260 ;
  buffer buf_n1262( .i (n1261), .o (n1262) );
  assign n1263 = n1079 & ~n1262 ;
  assign n1264 = n1245 | n1263 ;
  buffer buf_n1265( .i (n1264), .o (n1265) );
  assign n1266 = n1127 & ~n1262 ;
  assign n1267 = n1245 & n1266 ;
  buffer buf_n1268( .i (n1267), .o (n1268) );
  assign n1270 = n1265 & ~n1268 ;
  buffer buf_n1271( .i (n1270), .o (n1271) );
  assign n1272 = n1221 & n1271 ;
  buffer buf_n1273( .i (n1272), .o (n1273) );
  assign n1274 = n1184 & n1273 ;
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  assign n1282 = n96 | n744 ;
  assign n1283 = n335 & n1282 ;
  buffer buf_n1284( .i (n1283), .o (n1284) );
  assign n1285 = n677 | n1054 ;
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  assign n1286 = ~n109 & n1058 ;
  assign n1287 = n1285 & ~n1286 ;
  assign n1288 = ~n1284 & n1287 ;
  assign n1289 = n1044 & ~n1288 ;
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n423( .i (n422), .o (n423) );
  assign n1292 = ~n56 & n423 ;
  assign n1293 = n1027 | n1292 ;
  assign n1294 = n1193 | n1293 ;
  buffer buf_n1295( .i (n1294), .o (n1295) );
  assign n1296 = n101 & ~n1295 ;
  assign n1297 = ~n101 & n1030 ;
  assign n1298 = n1296 | n1297 ;
  assign n1299 = n1291 | n1298 ;
  buffer buf_n1300( .i (n1299), .o (n1300) );
  assign n1301 = n357 & ~n1107 ;
  buffer buf_n135( .i (n134), .o (n135) );
  assign n1302 = n135 | n1253 ;
  assign n1303 = ~n362 & n1253 ;
  assign n1304 = n1302 & ~n1303 ;
  assign n1305 = n1301 | n1304 ;
  buffer buf_n638( .i (n637), .o (n638) );
  assign n1306 = n638 | n1081 ;
  buffer buf_n1307( .i (n1306), .o (n1307) );
  assign n1308 = n400 | n1307 ;
  assign n1309 = ~n368 & n1307 ;
  assign n1310 = n1308 & ~n1309 ;
  buffer buf_n1311( .i (n1310), .o (n1311) );
  assign n1312 = n1305 | n1311 ;
  assign n1313 = ~n1098 & n1312 ;
  buffer buf_n1314( .i (n1313), .o (n1314) );
  assign n1315 = n1124 & ~n1314 ;
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  assign n1318 = n1300 & n1317 ;
  buffer buf_n1319( .i (n1318), .o (n1319) );
  assign n1322 = n1076 & ~n1314 ;
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  assign n1325 = n1300 | n1324 ;
  buffer buf_n1326( .i (n1325), .o (n1326) );
  assign n1328 = ~n1319 & n1326 ;
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n1331( .i (n1029), .o (n1331) );
  assign n1332 = n113 | n1331 ;
  assign n1333 = n113 & n1295 ;
  assign n1334 = n1332 & ~n1333 ;
  assign n1335 = n107 & n121 ;
  assign n1336 = n744 & ~n1335 ;
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  assign n1341 = n1186 & n1340 ;
  assign n1342 = ~n334 & n1038 ;
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n122( .i (n121), .o (n122) );
  assign n1344 = n122 & n1253 ;
  assign n1345 = n1110 | n1344 ;
  assign n1346 = n1343 & n1345 ;
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  assign n1350 = n1341 | n1349 ;
  assign n1351 = n1334 | n1350 ;
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  assign n1354 = n576 | n1307 ;
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  assign n1359 = n1100 & ~n1358 ;
  buffer buf_n1360( .i (n1359), .o (n1360) );
  assign n1361 = n379 & n1355 ;
  buffer buf_n1362( .i (n1106), .o (n1362) );
  assign n1363 = n363 & ~n1362 ;
  buffer buf_n404( .i (G39), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n1364( .i (n1252), .o (n1364) );
  assign n1365 = n408 | n1364 ;
  assign n1366 = ~n368 & n1364 ;
  assign n1367 = n1365 & ~n1366 ;
  assign n1368 = n1363 | n1367 ;
  assign n1369 = n1361 | n1368 ;
  buffer buf_n1370( .i (n1097), .o (n1370) );
  assign n1371 = n1369 & ~n1370 ;
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  assign n1374 = n1360 | n1373 ;
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1126), .o (n1376) );
  assign n1377 = ~n1375 & n1376 ;
  assign n1378 = n1353 & n1377 ;
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1380( .i (n1078), .o (n1380) );
  assign n1381 = ~n1375 & n1380 ;
  assign n1382 = n1353 | n1381 ;
  buffer buf_n1383( .i (n1382), .o (n1383) );
  assign n1384 = ~n1379 & n1383 ;
  buffer buf_n1385( .i (n1384), .o (n1385) );
  assign n1386 = n1330 & n1385 ;
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  assign n1388 = ~n129 & n1233 ;
  assign n1389 = n127 & ~n1295 ;
  assign n1390 = n135 & n1364 ;
  assign n1391 = n1165 & ~n1390 ;
  assign n1392 = n1343 & ~n1391 ;
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  assign n1396 = n1389 | n1395 ;
  buffer buf_n1397( .i (n1396), .o (n1397) );
  assign n1398 = n1388 | n1397 ;
  buffer buf_n1399( .i (n1398), .o (n1399) );
  assign n1400 = n387 & n1355 ;
  assign n1401 = n377 & n1364 ;
  buffer buf_n438( .i (G40), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n1402( .i (n1252), .o (n1402) );
  assign n1403 = n442 & ~n1402 ;
  assign n1404 = n1401 | n1403 ;
  assign n1405 = n369 & ~n1362 ;
  assign n1406 = n1404 | n1405 ;
  assign n1407 = n1400 | n1406 ;
  assign n1408 = ~n1370 & n1407 ;
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  assign n1411 = n1360 | n1410 ;
  buffer buf_n1412( .i (n1411), .o (n1412) );
  assign n1413 = n1376 & ~n1412 ;
  assign n1414 = n1399 & n1413 ;
  buffer buf_n1415( .i (n1414), .o (n1415) );
  assign n1420 = n1380 & ~n1412 ;
  assign n1421 = n1399 | n1420 ;
  buffer buf_n1422( .i (n1421), .o (n1422) );
  assign n1423 = ~n1415 & n1422 ;
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  assign n1427 = n1387 & n1426 ;
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  assign n1429 = ~n1186 & n1295 ;
  assign n1430 = n141 & ~n1429 ;
  assign n1431 = ~n137 & n1027 ;
  assign n1432 = n408 & n1402 ;
  assign n1433 = n1251 & ~n1432 ;
  assign n1434 = n1343 & ~n1433 ;
  assign n1435 = n1431 | n1434 ;
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  assign n1439 = n1430 | n1438 ;
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  assign n1442 = n395 & n1355 ;
  assign n1443 = n385 & n1402 ;
  buffer buf_n449( .i (G41), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  assign n1444 = n453 & ~n1402 ;
  assign n1445 = n1443 | n1444 ;
  assign n1446 = n378 & ~n1362 ;
  assign n1447 = n1445 | n1446 ;
  assign n1448 = n1442 | n1447 ;
  assign n1449 = ~n1370 & n1448 ;
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  assign n1452 = n1360 | n1451 ;
  buffer buf_n1453( .i (n1452), .o (n1453) );
  assign n1454 = n1376 & ~n1453 ;
  assign n1455 = n1441 & n1454 ;
  buffer buf_n1456( .i (n1455), .o (n1456) );
  assign n1463 = n1380 & ~n1453 ;
  assign n1464 = n1441 | n1463 ;
  buffer buf_n1465( .i (n1464), .o (n1465) );
  assign n1466 = ~n1456 & n1465 ;
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  assign n1472 = n1428 & n1471 ;
  buffer buf_n1473( .i (n1472), .o (n1473) );
  assign n1474 = n1277 & n1473 ;
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n1488( .i (n1487), .o (n1488) );
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  assign n1504 = n1428 & n1462 ;
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  assign n1505 = n1387 & n1419 ;
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  assign n1506 = n1327 & n1379 ;
  assign n1507 = n1321 | n1506 ;
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  assign n1511 = n1505 | n1510 ;
  buffer buf_n1512( .i (n1511), .o (n1512) );
  assign n1513 = n1504 | n1512 ;
  buffer buf_n1514( .i (n1513), .o (n1514) );
  assign n1515 = n1278 & n1514 ;
  buffer buf_n1269( .i (n1268), .o (n1269) );
  assign n1516 = n1219 & n1265 ;
  assign n1517 = n1269 | n1516 ;
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  assign n1520 = n1184 & n1519 ;
  buffer buf_n1131( .i (n1130), .o (n1131) );
  assign n1521 = n1122 & n1180 ;
  assign n1522 = n1131 | n1521 ;
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  assign n1526 = n1520 | n1525 ;
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  assign n1534 = n1515 | n1530 ;
  buffer buf_n1535( .i (n1534), .o (n1535) );
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n1556( .i (n1555), .o (n1556) );
  buffer buf_n1557( .i (n1556), .o (n1557) );
  buffer buf_n1558( .i (n1557), .o (n1558) );
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n269( .i (G27), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n522( .i (G48), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  assign n1562 = n276 & n529 ;
  buffer buf_n1563( .i (n1562), .o (n1563) );
  assign n1604 = ~n836 & n1563 ;
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  assign n1620 = n1399 & n1608 ;
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  assign n1624 = n1424 | n1623 ;
  assign n1625 = n1424 & n1623 ;
  assign n1626 = n1624 & ~n1625 ;
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n494( .i (G47), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  assign n1629 = n1440 & n1607 ;
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n1633( .i (n1632), .o (n1633) );
  assign n1634 = n1467 | n1633 ;
  assign n1635 = n1467 & n1633 ;
  assign n1636 = n1634 & ~n1635 ;
  buffer buf_n1637( .i (n1636), .o (n1637) );
  assign n1638 = n515 & n1637 ;
  assign n1639 = ~n1628 & n1638 ;
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  buffer buf_n1658( .i (n1657), .o (n1658) );
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  assign n1671 = n581 & ~n836 ;
  buffer buf_n1672( .i (n1671), .o (n1672) );
  assign n1700 = n829 & ~n1672 ;
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  assign n1717 = n1514 & ~n1619 ;
  buffer buf_n1718( .i (n1717), .o (n1718) );
  assign n1725 = ~n78 & n1718 ;
  assign n1726 = n1716 | n1725 ;
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1057), .o (n1752) );
  assign n1753 = ~n190 & n1752 ;
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  assign n1769 = n1637 & n1768 ;
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  assign n1770 = ~n647 & n1672 ;
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  assign n1791 = ~n243 & n1139 ;
  assign n1792 = n817 & ~n1791 ;
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n263( .i (n262), .o (n263) );
  assign n1806 = n263 & n1139 ;
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  assign n1810 = n252 & n1139 ;
  buffer buf_n1811( .i (n1810), .o (n1811) );
  assign n1812 = n268 & ~n1811 ;
  buffer buf_n1813( .i (n1812), .o (n1813) );
  assign n1814 = n1809 & n1813 ;
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n470( .i (G43), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  assign n1820 = n412 | n478 ;
  buffer buf_n1821( .i (n1820), .o (n1821) );
  assign n1822 = ~n1817 & n1821 ;
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  assign n1823 = ~n339 & n458 ;
  assign n1824 = n428 & ~n1823 ;
  assign n1825 = ~n1822 & n1824 ;
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  assign n1826 = n253 | n1069 ;
  assign n1827 = n334 & n1826 ;
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  assign n1830 = n445 & n1829 ;
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n481( .i (G44), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  assign n1833 = n268 | n1811 ;
  buffer buf_n1834( .i (n1833), .o (n1834) );
  assign n1835 = n1809 | n1834 ;
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  assign n1838 = n490 & n1837 ;
  assign n1839 = n1832 | n1838 ;
  assign n1840 = ~n1809 & n1813 ;
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n491( .i (G45), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  assign n1844 = n450 | n492 ;
  buffer buf_n1845( .i (n1844), .o (n1845) );
  buffer buf_n1846( .i (n1845), .o (n1846) );
  buffer buf_n1847( .i (n1846), .o (n1847) );
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  assign n1852 = ~n1842 & n1851 ;
  assign n1853 = n1809 & ~n1834 ;
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n460( .i (G42), .o (n460) );
  buffer buf_n493( .i (G46), .o (n493) );
  assign n1859 = n460 | n493 ;
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  assign n1868 = ~n1855 & n1867 ;
  assign n1869 = n1852 | n1868 ;
  assign n1870 = n1839 | n1869 ;
  assign n1871 = n1825 & ~n1870 ;
  buffer buf_n1872( .i (n1871), .o (n1872) );
  buffer buf_n1873( .i (n1872), .o (n1873) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  assign n1874 = n338 & n1841 ;
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n1876( .i (n1875), .o (n1876) );
  assign n1879 = n103 | n1876 ;
  buffer buf_n1880( .i (n1879), .o (n1880) );
  assign n1881 = n127 | n1816 ;
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  assign n1885 = n1880 & n1884 ;
  assign n1886 = n681 | n1816 ;
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  assign n1888 = n658 | n1843 ;
  assign n1889 = n1887 & n1888 ;
  buffer buf_n1856( .i (n1855), .o (n1856) );
  assign n1890 = n89 | n1856 ;
  assign n1891 = ~n670 & n1837 ;
  buffer buf_n1892( .i (n1891), .o (n1892) );
  assign n1893 = n1890 & ~n1892 ;
  assign n1894 = n1889 & n1893 ;
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  assign n1895 = n239 & ~n1855 ;
  assign n1896 = n428 | n1895 ;
  buffer buf_n1897( .i (n1896), .o (n1897) );
  assign n1898 = ~n111 & n1829 ;
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  assign n1903 = n1897 | n1902 ;
  assign n1904 = n1894 & ~n1903 ;
  assign n1905 = n1885 & n1904 ;
  assign n1906 = n1873 | n1905 ;
  assign n1907 = ~n1804 & n1906 ;
  assign n1908 = n1775 & ~n1907 ;
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  assign n1913 = ~n1769 & n1912 ;
  buffer buf_n1914( .i (n1913), .o (n1914) );
  assign n1915 = n515 & ~n1637 ;
  buffer buf_n1916( .i (n1915), .o (n1916) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  assign n1919 = ~n515 & n1637 ;
  assign n1920 = n1780 | n1919 ;
  assign n1921 = n1916 | n1920 ;
  assign n1922 = ~n1914 & n1921 ;
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  buffer buf_n1930( .i (n1929), .o (n1930) );
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n1934( .i (n1933), .o (n1934) );
  buffer buf_n1935( .i (n1934), .o (n1935) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  assign n1952 = n1199 & n1607 ;
  buffer buf_n1953( .i (n1952), .o (n1953) );
  buffer buf_n1954( .i (n1953), .o (n1954) );
  buffer buf_n1955( .i (n1954), .o (n1955) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  assign n1957 = n1221 | n1956 ;
  assign n1958 = n1221 & n1956 ;
  assign n1959 = n1957 & ~n1958 ;
  buffer buf_n1960( .i (n1959), .o (n1960) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  assign n1969 = ~n204 & n437 ;
  buffer buf_n1970( .i (n1969), .o (n1970) );
  assign n1971 = n1960 & n1970 ;
  buffer buf_n205( .i (G20), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n1972 = n214 & n1837 ;
  assign n1973 = ~n668 & n1829 ;
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n175( .i (G19), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  assign n1975 = n183 & ~n1841 ;
  assign n1976 = n1974 | n1975 ;
  assign n1977 = n1972 | n1976 ;
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  assign n1981 = n660 | n1877 ;
  buffer buf_n165( .i (G18), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  assign n1982 = n174 & ~n1855 ;
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  assign n1983 = ~n226 & n680 ;
  assign n1984 = n1816 | n1983 ;
  assign n1985 = ~n1982 & n1984 ;
  buffer buf_n1986( .i (n1985), .o (n1986) );
  assign n1987 = ~n1897 & n1986 ;
  assign n1988 = n1981 & n1987 ;
  assign n1989 = ~n1980 & n1988 ;
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  assign n1990 = n447 & n1837 ;
  assign n1991 = n1900 | n1990 ;
  assign n1992 = n458 & ~n1842 ;
  assign n1993 = n99 & ~n411 ;
  buffer buf_n1994( .i (n1993), .o (n1994) );
  buffer buf_n1996( .i (n1815), .o (n1996) );
  assign n1997 = n1994 | n1996 ;
  assign n1998 = ~n1992 & n1997 ;
  assign n1999 = ~n1991 & n1998 ;
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n2001( .i (n2000), .o (n2001) );
  buffer buf_n130( .i (n129), .o (n130) );
  assign n2002 = n130 | n1877 ;
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  assign n2003 = n138 & ~n467 ;
  buffer buf_n2004( .i (n2003), .o (n2004) );
  buffer buf_n2005( .i (n1854), .o (n2005) );
  assign n2006 = n2004 | n2005 ;
  assign n2007 = n428 & n2006 ;
  buffer buf_n2008( .i (n2007), .o (n2008) );
  buffer buf_n2009( .i (n2008), .o (n2009) );
  assign n2010 = n2002 & n2009 ;
  assign n2011 = n2001 & n2010 ;
  assign n2012 = n1989 | n2011 ;
  assign n2013 = ~n1804 & n2012 ;
  assign n2014 = n1775 & ~n2013 ;
  buffer buf_n2015( .i (n2014), .o (n2015) );
  buffer buf_n2016( .i (n2015), .o (n2016) );
  buffer buf_n2017( .i (n2016), .o (n2017) );
  buffer buf_n2018( .i (n2017), .o (n2018) );
  assign n2019 = ~n1971 & n2018 ;
  buffer buf_n2020( .i (n2019), .o (n2020) );
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2028( .i (n2027), .o (n2028) );
  buffer buf_n2029( .i (n2028), .o (n2029) );
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  assign n2031 = n1409 | n1450 ;
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  assign n2032 = n260 | n1314 ;
  assign n2033 = n2031 | n2032 ;
  buffer buf_n2034( .i (n2033), .o (n2034) );
  assign n2035 = n1375 | n2034 ;
  buffer buf_n2036( .i (n2035), .o (n2036) );
  assign n2037 = n1412 & n1453 ;
  assign n2038 = n260 & n1314 ;
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  assign n2041 = n1375 & n2040 ;
  assign n2042 = n2037 & n2041 ;
  assign n2043 = n2036 & ~n2042 ;
  assign n2044 = n1610 | n2043 ;
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  assign n2053 = n1473 & n1618 ;
  assign n2054 = n2052 & ~n2053 ;
  buffer buf_n2055( .i (n2054), .o (n2055) );
  assign n2056 = n521 & ~n2055 ;
  buffer buf_n2057( .i (n2056), .o (n2057) );
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1966( .i (n1965), .o (n1966) );
  assign n2060 = ~n1718 & n1966 ;
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1719( .i (n1718), .o (n1719) );
  assign n2062 = ~n1231 & n1719 ;
  assign n2063 = n2061 | n2062 ;
  buffer buf_n2064( .i (n2063), .o (n2064) );
  assign n2065 = n2059 | n2064 ;
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  assign n2067 = n2059 & n2064 ;
  assign n2068 = n1790 | n2067 ;
  assign n2069 = n2066 & ~n2068 ;
  assign n2070 = n2030 | n2069 ;
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n2073( .i (n2072), .o (n2073) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n2075( .i (n2074), .o (n2075) );
  buffer buf_n2076( .i (n2075), .o (n2076) );
  buffer buf_n2077( .i (n2076), .o (n2077) );
  buffer buf_n2078( .i (n2077), .o (n2078) );
  buffer buf_n2079( .i (n2078), .o (n2079) );
  buffer buf_n2080( .i (n2079), .o (n2080) );
  buffer buf_n2081( .i (n2080), .o (n2081) );
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2089( .i (n2088), .o (n2089) );
  assign n2090 = n521 & n2055 ;
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  assign n2094 = n1245 & n1608 ;
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  assign n2098 = n1271 & ~n2097 ;
  assign n2099 = ~n1271 & n2097 ;
  assign n2100 = n2098 | n2099 ;
  buffer buf_n2101( .i (n2100), .o (n2101) );
  assign n2111 = n1960 & n2101 ;
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  assign n2119 = n278 & ~n836 ;
  buffer buf_n2120( .i (n2119), .o (n2120) );
  buffer buf_n2121( .i (n2120), .o (n2121) );
  buffer buf_n2122( .i (n2121), .o (n2122) );
  assign n2126 = n1157 & n2122 ;
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  buffer buf_n2129( .i (n2128), .o (n2129) );
  buffer buf_n2130( .i (n2129), .o (n2130) );
  assign n2131 = n1182 | n2130 ;
  assign n2132 = n1182 & n2130 ;
  assign n2133 = n2131 & ~n2132 ;
  buffer buf_n2134( .i (n2133), .o (n2134) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  assign n2138 = n2112 & n2136 ;
  buffer buf_n2139( .i (n2138), .o (n2139) );
  assign n2145 = n1278 & n2139 ;
  assign n2146 = n1278 | n2139 ;
  assign n2147 = ~n2145 & n2146 ;
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n2150( .i (n2149), .o (n2150) );
  assign n2151 = n2092 & ~n2150 ;
  buffer buf_n2152( .i (n2151), .o (n2152) );
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  assign n2155 = n1281 | n1719 ;
  assign n2156 = ~n1533 & n2155 ;
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n2137( .i (n2136), .o (n2137) );
  assign n2158 = n1268 & ~n1610 ;
  buffer buf_n2159( .i (n2158), .o (n2159) );
  buffer buf_n2160( .i (n2159), .o (n2160) );
  buffer buf_n2161( .i (n2160), .o (n2161) );
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n2163( .i (n2162), .o (n2163) );
  assign n2164 = n1219 & ~n1610 ;
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n2166( .i (n2165), .o (n2166) );
  buffer buf_n2167( .i (n2166), .o (n2167) );
  buffer buf_n2168( .i (n2167), .o (n2168) );
  assign n2177 = n2101 & ~n2168 ;
  assign n2178 = n2163 | n2177 ;
  buffer buf_n2179( .i (n2178), .o (n2179) );
  assign n2180 = n2137 & n2179 ;
  buffer buf_n2181( .i (n2180), .o (n2181) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  assign n2182 = n1180 & ~n2125 ;
  buffer buf_n2183( .i (n2182), .o (n2183) );
  buffer buf_n2184( .i (n2183), .o (n2184) );
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  buffer buf_n2187( .i (n2186), .o (n2187) );
  buffer buf_n2188( .i (n2187), .o (n2188) );
  buffer buf_n2189( .i (n2188), .o (n2189) );
  buffer buf_n2190( .i (n2189), .o (n2190) );
  buffer buf_n2191( .i (n2190), .o (n2191) );
  assign n2192 = n2181 | n2191 ;
  buffer buf_n2193( .i (n2192), .o (n2193) );
  buffer buf_n2194( .i (n2193), .o (n2194) );
  buffer buf_n2195( .i (n2194), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  assign n2197 = n2157 & n2196 ;
  assign n2198 = n2157 | n2196 ;
  assign n2199 = ~n2197 & n2198 ;
  buffer buf_n2200( .i (n2199), .o (n2200) );
  assign n2201 = n2154 & n2200 ;
  assign n2202 = n2154 | n2200 ;
  assign n2203 = ~n2201 & n2202 ;
  assign n2204 = n56 | n190 ;
  buffer buf_n2205( .i (n2204), .o (n2205) );
  assign n2206 = n796 & n2205 ;
  buffer buf_n2207( .i (n2206), .o (n2207) );
  buffer buf_n2208( .i (n2207), .o (n2208) );
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n2211( .i (n2210), .o (n2211) );
  buffer buf_n2212( .i (n2211), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  buffer buf_n2214( .i (n2213), .o (n2214) );
  buffer buf_n2215( .i (n2214), .o (n2215) );
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n2221( .i (n2220), .o (n2221) );
  buffer buf_n2222( .i (n2221), .o (n2222) );
  buffer buf_n2223( .i (n2222), .o (n2223) );
  buffer buf_n2224( .i (n2223), .o (n2224) );
  buffer buf_n2225( .i (n2224), .o (n2225) );
  buffer buf_n2226( .i (n2225), .o (n2226) );
  buffer buf_n2227( .i (n2226), .o (n2227) );
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  buffer buf_n2231( .i (n2230), .o (n2231) );
  buffer buf_n2232( .i (n2231), .o (n2232) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  assign n2235 = ~n2203 & n2234 ;
  assign n2236 = n653 & ~n677 ;
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  assign n2237 = n691 | n958 ;
  assign n2238 = ~n2236 & n2237 ;
  assign n2239 = n2205 | n2238 ;
  assign n2240 = ~n136 & n821 ;
  assign n2241 = ~n1337 & n2240 ;
  buffer buf_n2242( .i (n2241), .o (n2242) );
  assign n2243 = n2239 & ~n2242 ;
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  buffer buf_n2250( .i (n2249), .o (n2250) );
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  buffer buf_n2265( .i (n2264), .o (n2265) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  buffer buf_n2269( .i (n2268), .o (n2269) );
  buffer buf_n2270( .i (n2269), .o (n2270) );
  buffer buf_n2271( .i (n2270), .o (n2271) );
  assign n2272 = ~n2235 & n2271 ;
  buffer buf_n2273( .i (n2272), .o (n2273) );
  buffer buf_n2274( .i (n2273), .o (n2274) );
  buffer buf_n2275( .i (n2274), .o (n2275) );
  buffer buf_n2276( .i (n2275), .o (n2276) );
  buffer buf_n2277( .i (n2276), .o (n2277) );
  buffer buf_n2278( .i (n2277), .o (n2278) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  buffer buf_n2280( .i (n2279), .o (n2280) );
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  assign n2289 = ~n1033 & n1307 ;
  assign n2290 = ~n819 & n2289 ;
  buffer buf_n2291( .i (n2290), .o (n2291) );
  buffer buf_n2292( .i (n2291), .o (n2292) );
  buffer buf_n2293( .i (n2292), .o (n2293) );
  buffer buf_n2294( .i (n2293), .o (n2294) );
  buffer buf_n2295( .i (n2294), .o (n2295) );
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n2297( .i (n2296), .o (n2297) );
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  buffer buf_n2307( .i (n2306), .o (n2307) );
  buffer buf_n2308( .i (n2307), .o (n2308) );
  buffer buf_n2309( .i (n2308), .o (n2309) );
  buffer buf_n2310( .i (n2309), .o (n2310) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1917( .i (n1916), .o (n1917) );
  buffer buf_n1918( .i (n1917), .o (n1918) );
  buffer buf_n2324( .i (n1609), .o (n2324) );
  assign n2325 = n1456 & ~n2324 ;
  buffer buf_n2326( .i (n2325), .o (n2326) );
  buffer buf_n2327( .i (n2326), .o (n2327) );
  buffer buf_n2328( .i (n2327), .o (n2328) );
  buffer buf_n2329( .i (n2328), .o (n2329) );
  assign n2330 = n1627 | n2329 ;
  buffer buf_n2331( .i (n2330), .o (n2331) );
  assign n2332 = n1424 & n2326 ;
  buffer buf_n2333( .i (n2332), .o (n2333) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n2335( .i (n2334), .o (n2335) );
  buffer buf_n2336( .i (n2335), .o (n2336) );
  assign n2337 = n2331 & ~n2336 ;
  buffer buf_n2338( .i (n2337), .o (n2338) );
  assign n2339 = n1918 | n2338 ;
  assign n2340 = n1918 & n2338 ;
  assign n2341 = n2339 & ~n2340 ;
  buffer buf_n2342( .i (n2341), .o (n2342) );
  assign n2343 = n1719 & n2342 ;
  assign n2344 = n1690 | n2343 ;
  buffer buf_n2345( .i (n2344), .o (n2345) );
  buffer buf_n2346( .i (n2345), .o (n2346) );
  buffer buf_n2347( .i (n2346), .o (n2347) );
  buffer buf_n2348( .i (n2347), .o (n2348) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  assign n2349 = n1352 & n1607 ;
  buffer buf_n2350( .i (n2349), .o (n2350) );
  buffer buf_n2351( .i (n2350), .o (n2351) );
  buffer buf_n2352( .i (n2351), .o (n2352) );
  buffer buf_n2353( .i (n2352), .o (n2353) );
  assign n2354 = n1385 | n2353 ;
  assign n2355 = n1385 & n2353 ;
  assign n2356 = n2354 & ~n2355 ;
  buffer buf_n2357( .i (n2356), .o (n2357) );
  buffer buf_n2358( .i (n2357), .o (n2358) );
  buffer buf_n2359( .i (n2358), .o (n2359) );
  buffer buf_n2360( .i (n2359), .o (n2360) );
  buffer buf_n2361( .i (n2360), .o (n2361) );
  assign n2362 = n1415 & ~n2324 ;
  buffer buf_n2363( .i (n2362), .o (n2363) );
  buffer buf_n2364( .i (n2363), .o (n2364) );
  buffer buf_n2365( .i (n2364), .o (n2365) );
  buffer buf_n2366( .i (n2365), .o (n2366) );
  buffer buf_n2367( .i (n2366), .o (n2367) );
  buffer buf_n2368( .i (n2367), .o (n2368) );
  assign n2369 = n2331 & ~n2368 ;
  buffer buf_n2370( .i (n2369), .o (n2370) );
  assign n2371 = n2361 | n2370 ;
  buffer buf_n2372( .i (n2371), .o (n2372) );
  assign n2373 = n2361 & n2370 ;
  buffer buf_n2374( .i (n2373), .o (n2374) );
  assign n2375 = n2372 & ~n2374 ;
  buffer buf_n2376( .i (n2375), .o (n2376) );
  assign n2377 = ~n1645 & n2376 ;
  buffer buf_n2378( .i (n2377), .o (n2378) );
  assign n2379 = n1645 & ~n2376 ;
  buffer buf_n2380( .i (n2379), .o (n2380) );
  assign n2382 = n2378 | n2380 ;
  buffer buf_n2383( .i (n2382), .o (n2383) );
  assign n2384 = n1724 & ~n2383 ;
  assign n2385 = n2348 | n2384 ;
  assign n2386 = ~n2319 & n2385 ;
  buffer buf_n2381( .i (n2380), .o (n2381) );
  assign n2387 = n1379 & ~n2324 ;
  buffer buf_n2388( .i (n2387), .o (n2388) );
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2391( .i (n2390), .o (n2391) );
  buffer buf_n2392( .i (n2391), .o (n2392) );
  buffer buf_n2393( .i (n2392), .o (n2393) );
  buffer buf_n2394( .i (n2393), .o (n2394) );
  buffer buf_n2395( .i (n2394), .o (n2395) );
  buffer buf_n2396( .i (n2395), .o (n2396) );
  buffer buf_n2397( .i (n2396), .o (n2397) );
  assign n2398 = n2372 & ~n2397 ;
  buffer buf_n2399( .i (n2398), .o (n2399) );
  buffer buf_n2400( .i (n1606), .o (n2400) );
  assign n2401 = n1300 & n2400 ;
  buffer buf_n2402( .i (n2401), .o (n2402) );
  buffer buf_n2403( .i (n2402), .o (n2403) );
  buffer buf_n2404( .i (n2403), .o (n2404) );
  assign n2405 = n1329 | n2404 ;
  assign n2406 = n1329 & n2404 ;
  assign n2407 = n2405 & ~n2406 ;
  buffer buf_n2408( .i (n2407), .o (n2408) );
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  buffer buf_n2411( .i (n2410), .o (n2411) );
  buffer buf_n2412( .i (n2411), .o (n2412) );
  buffer buf_n2413( .i (n2412), .o (n2413) );
  buffer buf_n2414( .i (n2413), .o (n2414) );
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n2416( .i (n2415), .o (n2416) );
  buffer buf_n2417( .i (n2416), .o (n2417) );
  assign n2418 = n2399 & ~n2417 ;
  assign n2419 = ~n2399 & n2417 ;
  assign n2420 = n2418 | n2419 ;
  buffer buf_n2421( .i (n2420), .o (n2421) );
  assign n2422 = n2381 & ~n2421 ;
  assign n2423 = ~n2381 & n2421 ;
  assign n2424 = n2422 | n2423 ;
  buffer buf_n2425( .i (n2424), .o (n2425) );
  buffer buf_n2426( .i (n2425), .o (n2426) );
  assign n2427 = ~n2386 & n2426 ;
  assign n2428 = n1767 & n2408 ;
  assign n2429 = ~n182 & n655 ;
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  assign n2432 = n1856 | n2431 ;
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n2433( .i (n1836), .o (n2433) );
  assign n2434 = n227 & n2433 ;
  assign n2435 = n214 & ~n1842 ;
  assign n2436 = n2434 | n2435 ;
  assign n2437 = n2432 & ~n2436 ;
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n240( .i (n239), .o (n240) );
  assign n2438 = n89 & ~n240 ;
  assign n2439 = n1818 | n2438 ;
  assign n2440 = n2437 & n2439 ;
  assign n2441 = ~n679 & n1829 ;
  buffer buf_n2442( .i (n2441), .o (n2442) );
  buffer buf_n2443( .i (n2442), .o (n2443) );
  buffer buf_n2444( .i (n2443), .o (n2444) );
  buffer buf_n671( .i (n670), .o (n671) );
  assign n2445 = n671 | n1875 ;
  assign n2446 = ~n2444 & n2445 ;
  assign n2447 = ~n430 & n2446 ;
  assign n2448 = n2440 & n2447 ;
  assign n2449 = n1821 & ~n1856 ;
  assign n2450 = n112 & ~n446 ;
  buffer buf_n2451( .i (n2450), .o (n2451) );
  assign n2452 = n1817 | n2451 ;
  assign n2453 = ~n2449 & n2452 ;
  buffer buf_n2454( .i (n2453), .o (n2454) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n2455( .i (n1841), .o (n2455) );
  assign n2456 = n469 & ~n2455 ;
  assign n2457 = n458 & n2433 ;
  assign n2458 = n2456 | n2457 ;
  buffer buf_n2459( .i (n2458), .o (n2459) );
  assign n2460 = n141 | n1875 ;
  buffer buf_n2461( .i (n1828), .o (n2461) );
  assign n2462 = ~n125 & n2461 ;
  assign n2463 = n426 & ~n2462 ;
  buffer buf_n2464( .i (n2463), .o (n2464) );
  buffer buf_n2465( .i (n2464), .o (n2465) );
  assign n2466 = n2460 & n2465 ;
  assign n2467 = ~n2459 & n2466 ;
  assign n2468 = n2454 & n2467 ;
  assign n2469 = n2448 | n2468 ;
  assign n2470 = ~n1803 & n2469 ;
  assign n2471 = n1774 & ~n2470 ;
  buffer buf_n2472( .i (n2471), .o (n2472) );
  buffer buf_n2473( .i (n2472), .o (n2473) );
  buffer buf_n2474( .i (n2473), .o (n2474) );
  buffer buf_n2475( .i (n2474), .o (n2475) );
  assign n2476 = ~n2428 & n2475 ;
  buffer buf_n2477( .i (n2476), .o (n2477) );
  buffer buf_n2478( .i (n2477), .o (n2478) );
  buffer buf_n2479( .i (n2478), .o (n2479) );
  buffer buf_n2480( .i (n2479), .o (n2480) );
  buffer buf_n2481( .i (n2480), .o (n2481) );
  buffer buf_n2482( .i (n2481), .o (n2482) );
  buffer buf_n2483( .i (n2482), .o (n2483) );
  buffer buf_n2484( .i (n2483), .o (n2484) );
  buffer buf_n2485( .i (n2484), .o (n2485) );
  buffer buf_n2486( .i (n2485), .o (n2486) );
  buffer buf_n2487( .i (n2486), .o (n2487) );
  buffer buf_n2488( .i (n2487), .o (n2488) );
  buffer buf_n2489( .i (n2488), .o (n2489) );
  buffer buf_n2490( .i (n2489), .o (n2490) );
  buffer buf_n2491( .i (n2490), .o (n2491) );
  assign n2492 = n2427 | n2491 ;
  buffer buf_n2493( .i (n2492), .o (n2493) );
  buffer buf_n2494( .i (n2493), .o (n2494) );
  buffer buf_n2495( .i (n2494), .o (n2495) );
  buffer buf_n2496( .i (n2495), .o (n2496) );
  buffer buf_n2497( .i (n2496), .o (n2497) );
  buffer buf_n2498( .i (n2497), .o (n2498) );
  buffer buf_n2499( .i (n2498), .o (n2499) );
  buffer buf_n2500( .i (n2499), .o (n2500) );
  buffer buf_n2501( .i (n2500), .o (n2501) );
  buffer buf_n2502( .i (n2501), .o (n2502) );
  buffer buf_n2503( .i (n2502), .o (n2503) );
  buffer buf_n2504( .i (n2503), .o (n2504) );
  buffer buf_n2505( .i (n2504), .o (n2505) );
  buffer buf_n2506( .i (n2505), .o (n2506) );
  buffer buf_n2507( .i (n2506), .o (n2507) );
  buffer buf_n2508( .i (n2507), .o (n2508) );
  buffer buf_n2509( .i (n1718), .o (n2509) );
  assign n2510 = n2342 | n2509 ;
  buffer buf_n2511( .i (n2510), .o (n2511) );
  buffer buf_n2512( .i (n2511), .o (n2512) );
  assign n2513 = ~n2345 & n2512 ;
  assign n2514 = n2312 & ~n2342 ;
  assign n2515 = n1627 & n1768 ;
  buffer buf_n1805( .i (n1804), .o (n1805) );
  assign n2516 = n411 & n2461 ;
  buffer buf_n2517( .i (n2516), .o (n2517) );
  buffer buf_n2518( .i (n2517), .o (n2518) );
  assign n2519 = n490 & ~n2455 ;
  assign n2520 = n2518 | n2519 ;
  assign n2521 = n1851 & ~n2005 ;
  buffer buf_n479( .i (n478), .o (n479) );
  assign n2522 = n479 & n2433 ;
  assign n2523 = n2521 | n2522 ;
  assign n2524 = n2520 | n2523 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n2525 = n448 & ~n1875 ;
  assign n2526 = n1996 | n2004 ;
  buffer buf_n2527( .i (n427), .o (n2527) );
  assign n2528 = n2526 & n2527 ;
  assign n2529 = ~n2525 & n2528 ;
  assign n2530 = ~n2524 & n2529 ;
  buffer buf_n2531( .i (n2530), .o (n2531) );
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n2532), .o (n2533) );
  assign n2534 = ~n657 & n2433 ;
  buffer buf_n2535( .i (n2534), .o (n2535) );
  assign n2536 = n240 & ~n1843 ;
  assign n2537 = n2535 | n2536 ;
  assign n2538 = n113 | n1996 ;
  buffer buf_n2539( .i (n2538), .o (n2539) );
  buffer buf_n2540( .i (n2005), .o (n2540) );
  assign n2541 = n682 | n2540 ;
  assign n2542 = n2539 & n2541 ;
  assign n2543 = ~n2537 & n2542 ;
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  assign n2546 = n91 | n1877 ;
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2548( .i (n669), .o (n2548) );
  assign n2549 = n1996 | n2548 ;
  assign n2550 = ~n2527 & n2549 ;
  buffer buf_n2551( .i (n2550), .o (n2551) );
  buffer buf_n2552( .i (n2551), .o (n2552) );
  assign n2553 = ~n99 & n2461 ;
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2555( .i (n2554), .o (n2555) );
  buffer buf_n2556( .i (n2555), .o (n2556) );
  buffer buf_n2557( .i (n2556), .o (n2557) );
  buffer buf_n228( .i (n227), .o (n228) );
  assign n2558 = n228 & ~n2540 ;
  buffer buf_n2559( .i (n2558), .o (n2559) );
  assign n2560 = n2557 | n2559 ;
  assign n2561 = n2552 & ~n2560 ;
  assign n2562 = n2547 & n2561 ;
  assign n2563 = n2545 & n2562 ;
  assign n2564 = n2533 | n2563 ;
  assign n2565 = ~n1805 & n2564 ;
  assign n2566 = n1776 & ~n2565 ;
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n2568( .i (n2567), .o (n2568) );
  buffer buf_n2569( .i (n2568), .o (n2569) );
  assign n2570 = ~n2515 & n2569 ;
  buffer buf_n2571( .i (n2570), .o (n2571) );
  buffer buf_n2572( .i (n2571), .o (n2572) );
  buffer buf_n2573( .i (n2572), .o (n2573) );
  buffer buf_n2574( .i (n2573), .o (n2574) );
  buffer buf_n2575( .i (n2574), .o (n2575) );
  buffer buf_n2576( .i (n2575), .o (n2576) );
  assign n2577 = n2514 | n2576 ;
  buffer buf_n2578( .i (n2577), .o (n2578) );
  buffer buf_n2579( .i (n2578), .o (n2579) );
  assign n2580 = n2513 | n2579 ;
  buffer buf_n2581( .i (n2580), .o (n2581) );
  buffer buf_n2582( .i (n2581), .o (n2582) );
  buffer buf_n2583( .i (n2582), .o (n2583) );
  buffer buf_n2584( .i (n2583), .o (n2584) );
  buffer buf_n2585( .i (n2584), .o (n2585) );
  buffer buf_n2586( .i (n2585), .o (n2586) );
  buffer buf_n2587( .i (n2586), .o (n2587) );
  buffer buf_n2588( .i (n2587), .o (n2588) );
  buffer buf_n2589( .i (n2588), .o (n2589) );
  buffer buf_n2590( .i (n2589), .o (n2590) );
  buffer buf_n2591( .i (n2590), .o (n2591) );
  buffer buf_n2592( .i (n2591), .o (n2592) );
  buffer buf_n2593( .i (n2592), .o (n2593) );
  buffer buf_n2594( .i (n2593), .o (n2594) );
  buffer buf_n2595( .i (n2594), .o (n2595) );
  buffer buf_n2596( .i (n2595), .o (n2596) );
  buffer buf_n2597( .i (n2596), .o (n2597) );
  buffer buf_n2598( .i (n2597), .o (n2598) );
  buffer buf_n2599( .i (n2598), .o (n2599) );
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  assign n2602 = ~n1691 & n2511 ;
  buffer buf_n2603( .i (n2602), .o (n2603) );
  buffer buf_n2604( .i (n2603), .o (n2604) );
  assign n2605 = ~n2383 & n2604 ;
  buffer buf_n2606( .i (n2605), .o (n2606) );
  assign n2607 = n1768 & n2357 ;
  assign n2608 = n228 & ~n1843 ;
  assign n2609 = n2005 | n2548 ;
  assign n2610 = n100 & n656 ;
  buffer buf_n2611( .i (n1815), .o (n2611) );
  assign n2612 = n2610 | n2611 ;
  assign n2613 = n2609 & n2612 ;
  assign n2614 = ~n2608 & n2613 ;
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  buffer buf_n2617( .i (n2616), .o (n2617) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  assign n2618 = n685 | n1878 ;
  buffer buf_n215( .i (n214), .o (n215) );
  assign n2619 = n215 & ~n2540 ;
  assign n2620 = n429 | n2619 ;
  buffer buf_n2621( .i (n2620), .o (n2621) );
  assign n2622 = ~n86 & n2461 ;
  buffer buf_n2623( .i (n2622), .o (n2623) );
  buffer buf_n2624( .i (n2623), .o (n2624) );
  buffer buf_n2626( .i (n1836), .o (n2626) );
  assign n2627 = n239 & n2626 ;
  assign n2628 = n2624 | n2627 ;
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  assign n2631 = n2621 | n2630 ;
  assign n2632 = n2618 & ~n2631 ;
  assign n2633 = n2617 & n2632 ;
  assign n2634 = n469 & n2626 ;
  buffer buf_n2635( .i (n2634), .o (n2635) );
  assign n2636 = n447 | n490 ;
  assign n2637 = ~n2540 & n2636 ;
  assign n2638 = n2635 | n2637 ;
  buffer buf_n480( .i (n479), .o (n480) );
  assign n2639 = n480 & ~n1843 ;
  buffer buf_n2640( .i (n1828), .o (n2640) );
  assign n2641 = ~n138 & n2640 ;
  buffer buf_n2642( .i (n2641), .o (n2642) );
  buffer buf_n2643( .i (n2642), .o (n2643) );
  buffer buf_n2644( .i (n2643), .o (n2644) );
  assign n2645 = n2639 | n2644 ;
  assign n2646 = n2638 | n2645 ;
  buffer buf_n2647( .i (n2646), .o (n2647) );
  buffer buf_n2648( .i (n2647), .o (n2648) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  assign n2649 = n417 & ~n1878 ;
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n459( .i (n458), .o (n459) );
  assign n2650 = n128 & ~n459 ;
  buffer buf_n2651( .i (n2650), .o (n2651) );
  assign n2652 = n1819 | n2651 ;
  assign n2653 = n431 & n2652 ;
  assign n2654 = ~n2649 & n2653 ;
  assign n2655 = ~n2648 & n2654 ;
  assign n2656 = n2633 | n2655 ;
  assign n2657 = ~n1805 & n2656 ;
  assign n2658 = n1776 & ~n2657 ;
  buffer buf_n2659( .i (n2658), .o (n2659) );
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2660), .o (n2661) );
  assign n2662 = ~n2607 & n2661 ;
  buffer buf_n2663( .i (n2662), .o (n2663) );
  buffer buf_n2664( .i (n2663), .o (n2664) );
  buffer buf_n2665( .i (n2664), .o (n2665) );
  buffer buf_n2666( .i (n2665), .o (n2666) );
  buffer buf_n2667( .i (n2666), .o (n2667) );
  buffer buf_n2668( .i (n2667), .o (n2668) );
  buffer buf_n2669( .i (n2668), .o (n2669) );
  buffer buf_n2670( .i (n2669), .o (n2670) );
  buffer buf_n2671( .i (n2670), .o (n2671) );
  buffer buf_n2672( .i (n2671), .o (n2672) );
  buffer buf_n2673( .i (n2672), .o (n2673) );
  assign n2674 = n1691 | n2511 ;
  assign n2675 = ~n2315 & n2674 ;
  buffer buf_n2676( .i (n2675), .o (n2676) );
  assign n2677 = n2383 & ~n2676 ;
  assign n2678 = n2673 | n2677 ;
  assign n2679 = n2606 | n2678 ;
  buffer buf_n2680( .i (n2679), .o (n2680) );
  buffer buf_n2681( .i (n2680), .o (n2681) );
  buffer buf_n2682( .i (n2681), .o (n2682) );
  buffer buf_n2683( .i (n2682), .o (n2683) );
  buffer buf_n2684( .i (n2683), .o (n2684) );
  buffer buf_n2685( .i (n2684), .o (n2685) );
  buffer buf_n2686( .i (n2685), .o (n2686) );
  buffer buf_n2687( .i (n2686), .o (n2687) );
  buffer buf_n2688( .i (n2687), .o (n2688) );
  buffer buf_n2689( .i (n2688), .o (n2689) );
  buffer buf_n2690( .i (n2689), .o (n2690) );
  buffer buf_n2691( .i (n2690), .o (n2691) );
  buffer buf_n2692( .i (n2691), .o (n2692) );
  buffer buf_n2693( .i (n2692), .o (n2693) );
  buffer buf_n2694( .i (n2693), .o (n2694) );
  buffer buf_n2695( .i (n2694), .o (n2695) );
  buffer buf_n2696( .i (n2695), .o (n2696) );
  buffer buf_n2697( .i (n2696), .o (n2697) );
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n2143( .i (n2142), .o (n2143) );
  buffer buf_n2144( .i (n2143), .o (n2144) );
  assign n2698 = n2092 & n2144 ;
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  assign n2700 = n2091 & n2118 ;
  buffer buf_n2701( .i (n2700), .o (n2701) );
  assign n2702 = n2137 | n2179 ;
  buffer buf_n2703( .i (n2702), .o (n2703) );
  assign n2704 = ~n2181 & n2703 ;
  buffer buf_n2705( .i (n2704), .o (n2705) );
  buffer buf_n2706( .i (n2705), .o (n2706) );
  buffer buf_n2707( .i (n2706), .o (n2707) );
  buffer buf_n2708( .i (n2707), .o (n2708) );
  assign n2709 = ~n2701 & n2708 ;
  assign n2710 = n2699 | n2709 ;
  buffer buf_n2711( .i (n2710), .o (n2711) );
  buffer buf_n2712( .i (n2711), .o (n2712) );
  buffer buf_n2713( .i (n2712), .o (n2713) );
  buffer buf_n2714( .i (n2713), .o (n2714) );
  buffer buf_n2715( .i (n2714), .o (n2715) );
  buffer buf_n2716( .i (n2715), .o (n2716) );
  buffer buf_n2717( .i (n2716), .o (n2717) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n2321( .i (n2320), .o (n2321) );
  buffer buf_n2322( .i (n2321), .o (n2322) );
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  buffer buf_n2171( .i (n2170), .o (n2171) );
  buffer buf_n2172( .i (n2171), .o (n2172) );
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n2175( .i (n2174), .o (n2175) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  assign n2718 = n2061 | n2176 ;
  buffer buf_n2719( .i (n2718), .o (n2719) );
  buffer buf_n2720( .i (n2719), .o (n2720) );
  buffer buf_n2721( .i (n2720), .o (n2721) );
  buffer buf_n2102( .i (n2101), .o (n2102) );
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n1967( .i (n1966), .o (n1967) );
  buffer buf_n1968( .i (n1967), .o (n1968) );
  assign n2722 = n1968 & n2091 ;
  assign n2723 = n2110 | n2722 ;
  assign n2724 = ~n2701 & n2723 ;
  buffer buf_n2725( .i (n2724), .o (n2725) );
  assign n2726 = n2721 | n2725 ;
  assign n2727 = n2721 & n2725 ;
  assign n2728 = n2726 & ~n2727 ;
  buffer buf_n2729( .i (n2728), .o (n2729) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  assign n2730 = n2093 & ~n2157 ;
  buffer buf_n2731( .i (n2730), .o (n2731) );
  buffer buf_n2732( .i (n2731), .o (n2732) );
  buffer buf_n2733( .i (n2732), .o (n2733) );
  buffer buf_n2734( .i (n2733), .o (n2734) );
  assign n2735 = n2729 | n2734 ;
  buffer buf_n2736( .i (n2735), .o (n2736) );
  assign n2737 = n1699 | n2736 ;
  assign n2738 = ~n2323 & n2737 ;
  assign n2739 = n2717 & ~n2738 ;
  buffer buf_n2740( .i (n2739), .o (n2740) );
  assign n2741 = ~n1699 & n2736 ;
  buffer buf_n2742( .i (n2741), .o (n2742) );
  assign n2743 = ~n2717 & n2742 ;
  assign n2744 = n1970 & n2134 ;
  buffer buf_n2745( .i (n1854), .o (n2745) );
  buffer buf_n2746( .i (n2745), .o (n2746) );
  assign n2747 = n2451 | n2746 ;
  buffer buf_n2748( .i (n2747), .o (n2748) );
  buffer buf_n2749( .i (n2748), .o (n2749) );
  assign n2750 = n1880 & n2749 ;
  assign n2751 = ~n140 & n2626 ;
  buffer buf_n2752( .i (n2751), .o (n2752) );
  buffer buf_n2753( .i (n2752), .o (n2753) );
  buffer buf_n2625( .i (n2624), .o (n2625) );
  assign n2754 = n1887 & ~n2625 ;
  assign n2755 = ~n2753 & n2754 ;
  buffer buf_n2756( .i (n2455), .o (n2756) );
  assign n2757 = n414 & ~n2756 ;
  buffer buf_n2758( .i (n2757), .o (n2758) );
  assign n2759 = n429 & n1882 ;
  assign n2760 = ~n2758 & n2759 ;
  assign n2761 = n2755 & n2760 ;
  assign n2762 = n2750 & n2761 ;
  buffer buf_n143( .i (G16), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  assign n2763 = n153 & ~n2746 ;
  buffer buf_n2764( .i (n2763), .o (n2764) );
  buffer buf_n154( .i (G17), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  assign n2765 = n164 & ~n2756 ;
  assign n2766 = n237 & n2640 ;
  buffer buf_n2767( .i (n2766), .o (n2767) );
  buffer buf_n2768( .i (n2767), .o (n2768) );
  buffer buf_n2769( .i (n2768), .o (n2769) );
  assign n2770 = n2765 | n2769 ;
  assign n2771 = n2764 | n2770 ;
  buffer buf_n2772( .i (n2771), .o (n2772) );
  buffer buf_n229( .i (n228), .o (n229) );
  assign n2773 = n229 & ~n1876 ;
  assign n2774 = n174 & n2626 ;
  assign n2775 = n2430 | n2611 ;
  assign n2776 = ~n2774 & n2775 ;
  buffer buf_n2777( .i (n2776), .o (n2777) );
  assign n2778 = ~n2773 & n2777 ;
  assign n2779 = ~n2621 & n2778 ;
  assign n2780 = ~n2772 & n2779 ;
  assign n2781 = n2762 | n2780 ;
  assign n2782 = ~n1804 & n2781 ;
  assign n2783 = n1775 & ~n2782 ;
  buffer buf_n2784( .i (n2783), .o (n2784) );
  buffer buf_n2785( .i (n2784), .o (n2785) );
  buffer buf_n2786( .i (n2785), .o (n2786) );
  buffer buf_n2787( .i (n2786), .o (n2787) );
  assign n2788 = ~n2744 & n2787 ;
  buffer buf_n2789( .i (n2788), .o (n2789) );
  buffer buf_n2790( .i (n2789), .o (n2790) );
  buffer buf_n2791( .i (n2790), .o (n2791) );
  buffer buf_n2792( .i (n2791), .o (n2792) );
  buffer buf_n2793( .i (n2792), .o (n2793) );
  buffer buf_n2794( .i (n2793), .o (n2794) );
  buffer buf_n2795( .i (n2794), .o (n2795) );
  buffer buf_n2796( .i (n2795), .o (n2796) );
  buffer buf_n2797( .i (n2796), .o (n2797) );
  buffer buf_n2798( .i (n2797), .o (n2798) );
  buffer buf_n2799( .i (n2798), .o (n2799) );
  buffer buf_n2800( .i (n2799), .o (n2800) );
  buffer buf_n2801( .i (n2800), .o (n2801) );
  buffer buf_n2802( .i (n2801), .o (n2802) );
  buffer buf_n2803( .i (n2802), .o (n2803) );
  buffer buf_n2804( .i (n2803), .o (n2804) );
  buffer buf_n2805( .i (n2804), .o (n2805) );
  buffer buf_n2806( .i (n2805), .o (n2806) );
  assign n2807 = n2743 | n2806 ;
  assign n2808 = n2740 | n2807 ;
  buffer buf_n2809( .i (n2808), .o (n2809) );
  buffer buf_n2810( .i (n2809), .o (n2810) );
  buffer buf_n2811( .i (n2810), .o (n2811) );
  buffer buf_n2812( .i (n2811), .o (n2812) );
  buffer buf_n2813( .i (n2812), .o (n2813) );
  buffer buf_n2814( .i (n2813), .o (n2814) );
  buffer buf_n2815( .i (n2814), .o (n2815) );
  buffer buf_n2816( .i (n2815), .o (n2816) );
  buffer buf_n2817( .i (n2816), .o (n2817) );
  buffer buf_n2818( .i (n2817), .o (n2818) );
  buffer buf_n2819( .i (n2818), .o (n2819) );
  assign n2820 = n1066 & n2122 ;
  buffer buf_n2821( .i (n2820), .o (n2821) );
  buffer buf_n2822( .i (n2821), .o (n2822) );
  buffer buf_n2823( .i (n2822), .o (n2823) );
  buffer buf_n2824( .i (n2823), .o (n2824) );
  assign n2825 = n1133 | n2824 ;
  assign n2826 = n1133 & n2824 ;
  assign n2827 = n2825 & ~n2826 ;
  buffer buf_n2828( .i (n2827), .o (n2828) );
  assign n2836 = n1970 & n2828 ;
  assign n2837 = n173 | n238 ;
  buffer buf_n2838( .i (n2837), .o (n2838) );
  assign n2839 = ~n1817 & n2838 ;
  buffer buf_n2840( .i (n2839), .o (n2840) );
  buffer buf_n2841( .i (n2840), .o (n2841) );
  buffer buf_n2842( .i (n2841), .o (n2842) );
  buffer buf_n2843( .i (n2842), .o (n2843) );
  assign n2844 = n153 & ~n2756 ;
  buffer buf_n2845( .i (n2844), .o (n2845) );
  buffer buf_n2846( .i (n2845), .o (n2846) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n2847( .i (n1876), .o (n2847) );
  assign n2848 = n217 & ~n2847 ;
  assign n2849 = n2846 | n2848 ;
  buffer buf_n2850( .i (n1836), .o (n2850) );
  assign n2851 = n163 & n2850 ;
  buffer buf_n142( .i (G15), .o (n142) );
  assign n2852 = n142 | n175 ;
  buffer buf_n2853( .i (n2852), .o (n2853) );
  buffer buf_n2854( .i (n2853), .o (n2854) );
  buffer buf_n2855( .i (n2854), .o (n2855) );
  buffer buf_n2856( .i (n2855), .o (n2856) );
  buffer buf_n2857( .i (n2856), .o (n2857) );
  buffer buf_n2858( .i (n2857), .o (n2858) );
  buffer buf_n2859( .i (n2858), .o (n2859) );
  buffer buf_n2860( .i (n2859), .o (n2860) );
  assign n2861 = ~n2745 & n2860 ;
  assign n2862 = n2851 | n2861 ;
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  assign n2863 = n225 & n2640 ;
  assign n2864 = n1094 & ~n2863 ;
  buffer buf_n2865( .i (n2864), .o (n2865) );
  buffer buf_n2866( .i (n2865), .o (n2866) );
  assign n2867 = ~n2862 & n2866 ;
  buffer buf_n2868( .i (n2867), .o (n2868) );
  buffer buf_n2869( .i (n2868), .o (n2869) );
  assign n2870 = ~n2849 & n2869 ;
  assign n2871 = ~n2843 & n2870 ;
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  assign n2872 = n586 & n2547 ;
  assign n2873 = n141 | n2756 ;
  assign n2874 = ~n2444 & n2873 ;
  assign n2875 = ~n127 & n2850 ;
  buffer buf_n2876( .i (n2875), .o (n2876) );
  assign n2877 = n2539 & ~n2876 ;
  assign n2878 = n2874 & n2877 ;
  buffer buf_n1995( .i (n1994), .o (n1995) );
  assign n2879 = n1995 | n2746 ;
  buffer buf_n2880( .i (n2879), .o (n2880) );
  assign n2881 = n2551 & n2880 ;
  assign n2882 = n2878 & n2881 ;
  buffer buf_n2883( .i (n2882), .o (n2883) );
  assign n2884 = n2872 & n2883 ;
  assign n2885 = n2871 | n2884 ;
  assign n2886 = ~n1805 & n2885 ;
  assign n2887 = n1776 & ~n2886 ;
  buffer buf_n2888( .i (n2887), .o (n2888) );
  buffer buf_n2889( .i (n2888), .o (n2889) );
  buffer buf_n2890( .i (n2889), .o (n2890) );
  assign n2891 = ~n2836 & n2890 ;
  buffer buf_n2892( .i (n2891), .o (n2892) );
  buffer buf_n2893( .i (n2892), .o (n2893) );
  buffer buf_n2894( .i (n2893), .o (n2894) );
  buffer buf_n2895( .i (n2894), .o (n2895) );
  buffer buf_n2896( .i (n2895), .o (n2896) );
  buffer buf_n2897( .i (n2896), .o (n2897) );
  buffer buf_n2898( .i (n2897), .o (n2898) );
  buffer buf_n2899( .i (n2898), .o (n2899) );
  buffer buf_n2900( .i (n2899), .o (n2900) );
  buffer buf_n2901( .i (n2900), .o (n2901) );
  buffer buf_n2902( .i (n2901), .o (n2902) );
  buffer buf_n2903( .i (n2902), .o (n2903) );
  buffer buf_n2904( .i (n2903), .o (n2904) );
  buffer buf_n2905( .i (n2904), .o (n2905) );
  buffer buf_n2906( .i (n2905), .o (n2906) );
  buffer buf_n2907( .i (n2906), .o (n2907) );
  buffer buf_n2908( .i (n2907), .o (n2908) );
  buffer buf_n2909( .i (n2908), .o (n2909) );
  assign n2910 = n2729 & n2734 ;
  buffer buf_n2911( .i (n2910), .o (n2911) );
  assign n2914 = ~n2711 & n2732 ;
  assign n2915 = n1696 | n2914 ;
  buffer buf_n2916( .i (n2915), .o (n2916) );
  buffer buf_n2917( .i (n2916), .o (n2917) );
  assign n2918 = n2911 | n2917 ;
  assign n2919 = ~n2323 & n2918 ;
  buffer buf_n2829( .i (n2828), .o (n2829) );
  buffer buf_n2830( .i (n2829), .o (n2830) );
  buffer buf_n2831( .i (n2830), .o (n2831) );
  buffer buf_n2832( .i (n2831), .o (n2832) );
  buffer buf_n2833( .i (n2832), .o (n2833) );
  buffer buf_n2834( .i (n2833), .o (n2834) );
  buffer buf_n2835( .i (n2834), .o (n2835) );
  assign n2920 = n2193 & ~n2835 ;
  assign n2921 = ~n2193 & n2835 ;
  assign n2922 = n2920 | n2921 ;
  buffer buf_n2923( .i (n2922), .o (n2923) );
  buffer buf_n2924( .i (n2923), .o (n2924) );
  assign n2925 = n2699 & ~n2924 ;
  assign n2926 = ~n2699 & n2924 ;
  assign n2927 = n2925 | n2926 ;
  buffer buf_n2928( .i (n2927), .o (n2928) );
  buffer buf_n2929( .i (n2928), .o (n2929) );
  buffer buf_n2930( .i (n2929), .o (n2930) );
  buffer buf_n2931( .i (n2930), .o (n2931) );
  buffer buf_n2932( .i (n2931), .o (n2932) );
  buffer buf_n2933( .i (n2932), .o (n2933) );
  assign n2934 = ~n2919 & n2933 ;
  assign n2935 = n2909 | n2934 ;
  buffer buf_n2936( .i (n2935), .o (n2936) );
  buffer buf_n2937( .i (n2936), .o (n2937) );
  buffer buf_n2938( .i (n2937), .o (n2938) );
  buffer buf_n2939( .i (n2938), .o (n2939) );
  buffer buf_n2940( .i (n2939), .o (n2940) );
  buffer buf_n2941( .i (n2940), .o (n2941) );
  buffer buf_n2942( .i (n2941), .o (n2942) );
  buffer buf_n2943( .i (n2942), .o (n2943) );
  buffer buf_n2944( .i (n2943), .o (n2944) );
  buffer buf_n2945( .i (n2944), .o (n2945) );
  buffer buf_n2946( .i (n2945), .o (n2946) );
  buffer buf_n2947( .i (n2946), .o (n2947) );
  buffer buf_n2912( .i (n2911), .o (n2912) );
  buffer buf_n2913( .i (n2912), .o (n2913) );
  assign n2948 = n2742 & ~n2913 ;
  assign n2949 = n1970 & n2101 ;
  assign n2950 = n413 & n2850 ;
  buffer buf_n2951( .i (n2950), .o (n2951) );
  buffer buf_n2952( .i (n2455), .o (n2952) );
  assign n2953 = n448 & ~n2952 ;
  assign n2954 = n2951 | n2953 ;
  assign n2955 = n87 & n139 ;
  assign n2956 = n2611 | n2955 ;
  assign n2957 = ~n2555 & n2956 ;
  buffer buf_n2958( .i (n2957), .o (n2958) );
  assign n2959 = ~n2954 & n2958 ;
  buffer buf_n2960( .i (n2959), .o (n2960) );
  buffer buf_n2961( .i (n2960), .o (n2961) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  assign n2962 = n117 | n1878 ;
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  assign n2963 = n1858 | n2651 ;
  assign n2964 = n431 & n2963 ;
  assign n2965 = n2962 & n2964 ;
  assign n2966 = n2961 & n2965 ;
  assign n2967 = n164 & ~n2746 ;
  buffer buf_n2968( .i (n2967), .o (n2968) );
  buffer buf_n2969( .i (n2968), .o (n2969) );
  buffer buf_n184( .i (n183), .o (n184) );
  assign n2970 = n184 & n2850 ;
  buffer buf_n2971( .i (n2970), .o (n2971) );
  buffer buf_n2972( .i (n2971), .o (n2972) );
  assign n2973 = n2559 | n2972 ;
  assign n2974 = n2969 | n2973 ;
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  assign n2975 = n2838 & ~n2952 ;
  assign n2976 = n1148 | n2975 ;
  assign n2977 = ~n655 & n2640 ;
  buffer buf_n2978( .i (n2977), .o (n2978) );
  buffer buf_n2979( .i (n2978), .o (n2979) );
  assign n2980 = n214 & ~n2611 ;
  assign n2981 = n2979 | n2980 ;
  buffer buf_n2982( .i (n2981), .o (n2982) );
  assign n2983 = n2976 | n2982 ;
  assign n2984 = n2552 & ~n2983 ;
  assign n2985 = ~n2974 & n2984 ;
  buffer buf_n2986( .i (n2985), .o (n2986) );
  assign n2987 = n2966 | n2986 ;
  assign n2988 = ~n1805 & n2987 ;
  buffer buf_n2989( .i (n1774), .o (n2989) );
  buffer buf_n2990( .i (n2989), .o (n2990) );
  assign n2991 = ~n2988 & n2990 ;
  buffer buf_n2992( .i (n2991), .o (n2992) );
  buffer buf_n2993( .i (n2992), .o (n2993) );
  buffer buf_n2994( .i (n2993), .o (n2994) );
  assign n2995 = ~n2949 & n2994 ;
  buffer buf_n2996( .i (n2995), .o (n2996) );
  buffer buf_n2997( .i (n2996), .o (n2997) );
  buffer buf_n2998( .i (n2997), .o (n2998) );
  buffer buf_n2999( .i (n2998), .o (n2999) );
  buffer buf_n3000( .i (n2999), .o (n3000) );
  buffer buf_n3001( .i (n3000), .o (n3001) );
  buffer buf_n3002( .i (n3001), .o (n3002) );
  buffer buf_n3003( .i (n3002), .o (n3003) );
  buffer buf_n3004( .i (n3003), .o (n3004) );
  buffer buf_n3005( .i (n3004), .o (n3005) );
  buffer buf_n3006( .i (n3005), .o (n3006) );
  buffer buf_n3007( .i (n3006), .o (n3007) );
  buffer buf_n3008( .i (n3007), .o (n3008) );
  buffer buf_n3009( .i (n3008), .o (n3009) );
  assign n3010 = n2320 & ~n2729 ;
  assign n3011 = n3009 | n3010 ;
  buffer buf_n3012( .i (n3011), .o (n3012) );
  buffer buf_n3013( .i (n3012), .o (n3013) );
  buffer buf_n3014( .i (n3013), .o (n3014) );
  assign n3015 = n2948 | n3014 ;
  buffer buf_n3016( .i (n3015), .o (n3016) );
  buffer buf_n3017( .i (n3016), .o (n3017) );
  buffer buf_n3018( .i (n3017), .o (n3018) );
  buffer buf_n3019( .i (n3018), .o (n3019) );
  buffer buf_n3020( .i (n3019), .o (n3020) );
  buffer buf_n3021( .i (n3020), .o (n3021) );
  buffer buf_n3022( .i (n3021), .o (n3022) );
  buffer buf_n3023( .i (n3022), .o (n3023) );
  buffer buf_n3024( .i (n3023), .o (n3024) );
  buffer buf_n3025( .i (n3024), .o (n3025) );
  buffer buf_n3026( .i (n3025), .o (n3026) );
  buffer buf_n3027( .i (n3026), .o (n3027) );
  assign n3028 = n2809 | n2937 ;
  buffer buf_n3029( .i (n3028), .o (n3029) );
  assign n3030 = n2078 | n3016 ;
  buffer buf_n3031( .i (n3030), .o (n3031) );
  assign n3032 = n2493 | n2682 ;
  buffer buf_n3033( .i (n3032), .o (n3033) );
  assign n3034 = n1931 & ~n2581 ;
  buffer buf_n3035( .i (n3034), .o (n3035) );
  buffer buf_n3036( .i (n3035), .o (n3036) );
  buffer buf_n3037( .i (n3036), .o (n3037) );
  buffer buf_n3038( .i (n3037), .o (n3038) );
  buffer buf_n3039( .i (n3038), .o (n3039) );
  buffer buf_n3040( .i (n3039), .o (n3040) );
  assign n3041 = ~n3033 & n3040 ;
  buffer buf_n3042( .i (n3041), .o (n3042) );
  buffer buf_n3043( .i (n3042), .o (n3043) );
  buffer buf_n3044( .i (n3043), .o (n3044) );
  assign n3045 = ~n3031 & n3044 ;
  assign n3046 = ~n3029 & n3045 ;
  buffer buf_n3047( .i (n3046), .o (n3047) );
  buffer buf_n3048( .i (n3047), .o (n3048) );
  buffer buf_n3049( .i (n3048), .o (n3049) );
  buffer buf_n3050( .i (n3049), .o (n3050) );
  buffer buf_n3051( .i (n3050), .o (n3051) );
  buffer buf_n3052( .i (n3051), .o (n3052) );
  buffer buf_n3053( .i (n3052), .o (n3053) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  assign n3054 = n568 & ~n3029 ;
  buffer buf_n3055( .i (n3054), .o (n3055) );
  buffer buf_n3056( .i (n3055), .o (n3056) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  assign n3057 = n317 & ~n3047 ;
  assign n3058 = ~n3056 & n3057 ;
  buffer buf_n3059( .i (n3058), .o (n3059) );
  buffer buf_n3060( .i (n3059), .o (n3060) );
  buffer buf_n3061( .i (n3060), .o (n3061) );
  buffer buf_n3062( .i (n3061), .o (n3062) );
  assign n3063 = n2078 & n3016 ;
  buffer buf_n3064( .i (n3063), .o (n3064) );
  assign n3065 = n3031 & ~n3064 ;
  buffer buf_n3066( .i (n3065), .o (n3066) );
  assign n3067 = ~n1931 & n2581 ;
  buffer buf_n3068( .i (n3067), .o (n3068) );
  assign n3069 = n3035 | n3068 ;
  buffer buf_n3070( .i (n3069), .o (n3070) );
  buffer buf_n3071( .i (n3070), .o (n3071) );
  buffer buf_n3072( .i (n3071), .o (n3072) );
  buffer buf_n3073( .i (n3072), .o (n3073) );
  buffer buf_n3074( .i (n3073), .o (n3074) );
  buffer buf_n3075( .i (n3074), .o (n3075) );
  assign n3076 = n2493 & n2682 ;
  buffer buf_n3077( .i (n3076), .o (n3077) );
  assign n3078 = n3033 & ~n3077 ;
  buffer buf_n3079( .i (n3078), .o (n3079) );
  assign n3080 = n3075 | n3079 ;
  assign n3081 = n3075 & n3079 ;
  assign n3082 = n3080 & ~n3081 ;
  buffer buf_n3083( .i (n3082), .o (n3083) );
  buffer buf_n3084( .i (n3083), .o (n3084) );
  assign n3085 = n3066 & n3084 ;
  assign n3086 = n3066 | n3084 ;
  assign n3087 = ~n3085 & n3086 ;
  buffer buf_n3088( .i (n3087), .o (n3088) );
  buffer buf_n3089( .i (n3088), .o (n3089) );
  buffer buf_n3090( .i (n3089), .o (n3090) );
  buffer buf_n587( .i (G50), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  assign n3091 = n2809 & n2937 ;
  buffer buf_n3092( .i (n3091), .o (n3092) );
  assign n3093 = n3029 & ~n3092 ;
  buffer buf_n3094( .i (n3093), .o (n3094) );
  assign n3097 = n635 & n3094 ;
  buffer buf_n3098( .i (n3097), .o (n3098) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  assign n3099 = n635 | n3094 ;
  assign n3100 = ~n1603 & n3099 ;
  assign n3101 = ~n3098 & n3100 ;
  buffer buf_n3102( .i (n3101), .o (n3102) );
  assign n3103 = n3090 & n3102 ;
  assign n3104 = n3090 | n3102 ;
  assign n3105 = ~n3103 & n3104 ;
  buffer buf_n3095( .i (n3094), .o (n3095) );
  buffer buf_n3096( .i (n3095), .o (n3096) );
  assign n3106 = n3088 | n3096 ;
  assign n3107 = n3088 & n3096 ;
  assign n3108 = n3106 & ~n3107 ;
  buffer buf_n3109( .i (n3108), .o (n3109) );
  buffer buf_n3110( .i (n3109), .o (n3110) );
  assign G3519 = ~n742 ;
  assign G3520 = ~n794 ;
  assign G3521 = ~n883 ;
  assign G3522 = n955 ;
  assign G3523 = n1024 ;
  assign G3524 = n1503 ;
  assign G3525 = n1561 ;
  assign G3526 = n1670 ;
  assign G3527 = n1751 ;
  assign G3528 = ~n1951 ;
  assign G3529 = n2089 ;
  assign G3530 = ~n2288 ;
  assign G3531 = n2508 ;
  assign G3532 = n2601 ;
  assign G3533 = n2697 ;
  assign G3534 = n2819 ;
  assign G3535 = n2947 ;
  assign G3536 = n3027 ;
  assign G3537 = ~n3053 ;
  assign G3538 = ~n3062 ;
  assign G3539 = ~n3105 ;
  assign G3540 = n3110 ;
endmodule
