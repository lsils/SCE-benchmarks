module top( N1 , N100 , N103 , N106 , N109 , N110 , N111 , N112 , N113 , N114 , N115 , N118 , N12 , N121 , N124 , N127 , N130 , N133 , N134 , N135 , N138 , N141 , N144 , N147 , N15 , N150 , N151 , N152 , N153 , N154 , N155 , N156 , N157 , N158 , N159 , N160 , N161 , N162 , N163 , N164 , N165 , N166 , N167 , N168 , N169 , N170 , N171 , N172 , N173 , N174 , N175 , N176 , N177 , N178 , N179 , N18 , N180 , N181 , N182 , N183 , N184 , N185 , N186 , N187 , N188 , N189 , N190 , N191 , N192 , N193 , N194 , N195 , N196 , N197 , N198 , N199 , N200 , N201 , N202 , N203 , N204 , N205 , N206 , N207 , N208 , N209 , N210 , N211 , N212 , N213 , N214 , N215 , N216 , N217 , N218 , N219 , N220 , N221 , N222 , N223 , N224 , N225 , N226 , N227 , N228 , N229 , N23 , N230 , N231 , N232 , N233 , N234 , N235 , N236 , N237 , N238 , N239 , N240 , N241_I , N242 , N245 , N248 , N251 , N254 , N257 , N26 , N260 , N263 , N267 , N271 , N274 , N277 , N280 , N283 , N286 , N289 , N29 , N293 , N296 , N299 , N303 , N307 , N310 , N313 , N316 , N319 , N32 , N322 , N325 , N328 , N331 , N334 , N337 , N340 , N343 , N346 , N349 , N35 , N352 , N355 , N358 , N361 , N364 , N367 , N38 , N382 , N41 , N44 , N47 , N5 , N50 , N53 , N54 , N55 , N56 , N57 , N58 , N59 , N60 , N61 , N62 , N63 , N64 , N65 , N66 , N69 , N70 , N73 , N74 , N75 , N76 , N77 , N78 , N79 , N80 , N81 , N82 , N83 , N84 , N85 , N86 , N87 , N88 , N89 , N9 , N94 , N97 , N10025 , N10101 , N10102 , N10103 , N10104 , N10109 , N10110 , N10111 , N10112 , N10350 , N10351 , N10352 , N10353 , N10574 , N10575 , N10576 , N10628 , N10632 , N10641 , N10704 , N10706 , N10711 , N10712 , N10713 , N10714 , N10715 , N10716 , N10717 , N10718 , N10729 , N10759 , N10760 , N10761 , N10762 , N10763 , N10827 , N10837 , N10838 , N10839 , N10840 , N10868 , N10869 , N10870 , N10871 , N10905 , N10906 , N10907 , N10908 , N1110 , N1111 , N1112 , N1113 , N1114 , N11333 , N11334 , N11340 , N11342 , N1489 , N1490 , N1781 , N241_O , N387 , N388 , N478 , N482 , N484 , N486 , N489 , N492 , N501 , N505 , N507 , N509 , N511 , N513 , N515 , N517 , N519 , N535 , N537 , N539 , N541 , N543 , N545 , N547 , N549 , N551 , N553 , N556 , N559 , N561 , N563 , N565 , N567 , N569 , N571 , N573 , N582 , N643 , N707 , N813 , N881 , N882 , N883 , N884 , N885 , N889 , N945 );
  input N1 , N100 , N103 , N106 , N109 , N110 , N111 , N112 , N113 , N114 , N115 , N118 , N12 , N121 , N124 , N127 , N130 , N133 , N134 , N135 , N138 , N141 , N144 , N147 , N15 , N150 , N151 , N152 , N153 , N154 , N155 , N156 , N157 , N158 , N159 , N160 , N161 , N162 , N163 , N164 , N165 , N166 , N167 , N168 , N169 , N170 , N171 , N172 , N173 , N174 , N175 , N176 , N177 , N178 , N179 , N18 , N180 , N181 , N182 , N183 , N184 , N185 , N186 , N187 , N188 , N189 , N190 , N191 , N192 , N193 , N194 , N195 , N196 , N197 , N198 , N199 , N200 , N201 , N202 , N203 , N204 , N205 , N206 , N207 , N208 , N209 , N210 , N211 , N212 , N213 , N214 , N215 , N216 , N217 , N218 , N219 , N220 , N221 , N222 , N223 , N224 , N225 , N226 , N227 , N228 , N229 , N23 , N230 , N231 , N232 , N233 , N234 , N235 , N236 , N237 , N238 , N239 , N240 , N241_I , N242 , N245 , N248 , N251 , N254 , N257 , N26 , N260 , N263 , N267 , N271 , N274 , N277 , N280 , N283 , N286 , N289 , N29 , N293 , N296 , N299 , N303 , N307 , N310 , N313 , N316 , N319 , N32 , N322 , N325 , N328 , N331 , N334 , N337 , N340 , N343 , N346 , N349 , N35 , N352 , N355 , N358 , N361 , N364 , N367 , N38 , N382 , N41 , N44 , N47 , N5 , N50 , N53 , N54 , N55 , N56 , N57 , N58 , N59 , N60 , N61 , N62 , N63 , N64 , N65 , N66 , N69 , N70 , N73 , N74 , N75 , N76 , N77 , N78 , N79 , N80 , N81 , N82 , N83 , N84 , N85 , N86 , N87 , N88 , N89 , N9 , N94 , N97 ;
  output N10025 , N10101 , N10102 , N10103 , N10104 , N10109 , N10110 , N10111 , N10112 , N10350 , N10351 , N10352 , N10353 , N10574 , N10575 , N10576 , N10628 , N10632 , N10641 , N10704 , N10706 , N10711 , N10712 , N10713 , N10714 , N10715 , N10716 , N10717 , N10718 , N10729 , N10759 , N10760 , N10761 , N10762 , N10763 , N10827 , N10837 , N10838 , N10839 , N10840 , N10868 , N10869 , N10870 , N10871 , N10905 , N10906 , N10907 , N10908 , N1110 , N1111 , N1112 , N1113 , N1114 , N11333 , N11334 , N11340 , N11342 , N1489 , N1490 , N1781 , N241_O , N387 , N388 , N478 , N482 , N484 , N486 , N489 , N492 , N501 , N505 , N507 , N509 , N511 , N513 , N515 , N517 , N519 , N535 , N537 , N539 , N541 , N543 , N545 , N547 , N549 , N551 , N553 , N556 , N559 , N561 , N563 , N565 , N567 , N569 , N571 , N573 , N582 , N643 , N707 , N813 , N881 , N882 , N883 , N884 , N885 , N889 , N945 ;
  wire n3608 , n3610 , n3616 , n3617 , n3625 , n3629 , n3631 , n3633 , n3687 , n3748 , n3807 , n3808 , n3865 , n3867 , n3872 , n3876 , n3878 , n3885 , n3889 , n3891 , n3895 , n3899 , n3901 , n3912 , n3914 , n3915 , n3954 , n3958 , n3960 , n3967 , n3973 , n3978 , n3980 , n3984 , n3986 , n3988 , n4036 , n4038 , n4040 , n4077 , n4078 , n4113 , n4123 , n4165 , n4208 , n4211 , n4212 , n4213 , n4217 , n4219 , n4256 , n4292 , n4296 , n4298 , n4305 , n4311 , n4315 , n4317 , n4321 , n4326 , n4330 , n4332 , n4367 , n4370 , n4401 , n4403 , n4429 , n4463 , n4465 , n4494 , n4528 , n4531 , n4556 , n4558 , n4560 , n4576 , n4589 , n4591 , n4593 , n4595 , n4606 , n4617 , n4619 , n4621 , n4623 , n4630 , n4636 , n4638 , n4640 , n4642 , n4648 , n4650 , n4652 , n4654 , n4691 , n4693 , n4695 , n4723 , n4724 , n4750 , n4751 , n4774 , n4792 , n4794 , n4827 , n4864 , n4891 , n4924 , n4956 , n4958 , n4961 , n4962 , n4978 , n4980 , n4982 , n4984 , n5013 , n5042 , n5044 , n5046 , n5048 , n5056 , n5063 , n5065 , n5067 , n5069 , n5073 , n5077 , n5079 , n5081 , n5083 , n5108 , n5110 , n5132 , n5133 , n5151 , n5177 , n5203 , n5227 , n5246 , n5247 , n5264 , n5266 , n5268 , n5270 , n5296 , n5298 , n5300 , n5302 , n5306 , n5308 , n5329 , n5332 , n5336 , n5338 , n5340 , n5342 , n5344 , n5354 , n5365 , n5389 , n5391 , n5393 , n5395 , n5401 , n5409 , n5435 , n5437 , n5450 , n5452 , n5454 , n5456 , n5470 , n5483 , n5494 , n5506 , n5508 , n5510 , n5512 , n5521 , n5529 , n5531 , n5533 , n5535 , n5541 , n5547 , n5549 , n5551 , n5553 , n5556 , n5559 , n5561 , n5563 , n5565 , n5585 , n5586 , n5604 , n5605 , n5618 , n5619 , n5630 , n5632 , n5634 , n5636 , n5650 , n5663 , n5665 , n5667 , n5669 , n5680 , n5689 , n5691 , n5693 , n5695 , n5700 , n5702 , n5704 , n5706 , n5711 , n5713 , n5715 , n5719 , n5721 , n5722 , n5727 , n5730 , n5732 , n5733 , n5735 , n5737 , n5742 , n5746 , n5748 , n5750 , n5760 , n5763 , n5765 , n5766 , n5768 , n5771 , n5791 , n5809 , n5825 , n5827 , n5848 , n5867 , n5869 , n5880 , n5881 , n5885 , n5887 , n5888 , n5910 , n5912 , n5926 , n5927 , n5929 , n5930 , n5939 , n5944 , n5945 , n5947 , n5948 , n5954 , n5955 , n5962 , n5963 , n5965 , n5966 , n5974 , n6015 , n6017 , n6061 , n6109 , n6145 , n6179 , n6181 , n6182 , n6191 , n6193 , n6194 , n6197 , n6199 , n6200 , n6227 , n6228 , n6229 , n6232 , n6234 , n6236 , n6242 , n6244 , n6245 , n6248 , n6250 , n6252 , n6257 , n6259 , n6260 , n6262 , n6264 , n6266 , n6267 , n6268 , n6270 , n6272 , n6273 , n6275 , n6276 , n6277 , n6278 , n6280 , n6282 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6299 , n6301 , n6303 , n6304 , n6306 , n6307 , n6308 , n6309 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6322 , n6324 , n6326 , n6327 , n6328 , n6334 , n6336 , n6337 , n6338 , n6341 , n6343 , n6345 , n6347 , n6349 , n6350 , n6353 , n6355 , n6357 , n6359 , n6360 , n6361 , n6362 , n6364 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6378 , n6380 , n6382 , n6383 , n6385 , n6391 , n6392 , n6393 , n6394 , n6397 , n6399 , n6401 , n6404 , n6405 , n6406 , n6409 , n6411 , n6413 , n6414 , n6417 , n6419 , n6420 , n6423 , n6425 , n6427 , n6430 , n6432 , n6435 , n6436 , n6437 , n6439 , n6440 , n6441 , n6443 , n6445 , n6447 , n6448 , n6449 , n6454 , n6455 , n6456 , n6458 , n6461 , n6465 , n6466 , n6467 , n6471 , n6475 , n6476 , n6477 , n6478 , n6482 , n6484 , n6486 , n6488 , n6489 , n6490 , n6493 , n6495 , n6497 , n6499 , n6500 , n6503 , n6505 , n6506 , n6509 , n6510 , n6511 , n6514 , n6516 , n6518 , n6519 , n6522 , n6523 , n6526 , n6528 , n6530 , n6531 , n6533 , n6536 , n6538 , n6539 , n6541 , n6548 , n6549 , n6551 , n6552 , n6553 , n6556 , n6563 , n6608 , n6609 , n6610 , n6613 , n6614 , n6617 , n6619 , n6620 , n6621 , n6624 , n6626 , n6628 , n6629 , n6631 , n6635 , n6636 , n6638 , n6641 , n6642 , n6643 , n6648 , n6650 , n6652 , n6653 , n6655 , n6656 , n6661 , n6663 , n6665 , n6666 , n6668 , n6671 , n6673 , n6674 , n6676 , n6678 , n6679 , n6680 , n6685 , n6687 , n6689 , n6696 , n6698 , n6703 , n6711 , n6712 , n6713 , n6715 , n6716 , n6719 , n6721 , n6729 , n6730 , n6731 , n6732 , n6735 , n6739 , n6741 , n6743 , n6744 , n6745 , n6748 , n6752 , n6754 , n6755 , n6757 , n6759 , n6762 , n6763 , n6765 , n6767 , n6768 , n6771 , n6775 , n6777 , n6778 , n6779 , n6780 , n6784 , n6790 , n6792 , n6793 , n6795 , n6798 , n6800 , n6801 , n6803 , n6815 , n6816 , n6818 , n6819 , n6822 , n6834 , n6835 , n6836 , n6837 , n6840 , n6844 , n6846 , n6853 , n6854 , n6855 , n6858 , n6862 , n6864 , n6867 , n6869 , n6870 , n6872 , n6873 , n6876 , n6880 , n6882 , n6884 , n6886 , n6887 , n6888 , n6890 , n6891 , n6892 , n6894 , n6897 , n6898 , n6899 , n6902 , n6907 , n6909 , n6910 , n6913 , n6917 , n6921 , n6924 , n6925 , n6926 , n6928 , n6941 , n6942 , n6943 , n6945 , n6946 , n6949 , n6950 , n6958 , n6959 , n6960 , n6963 , n6976 , n6977 , n7014 , n7025 , n7027 , n7028 , n7030 , n7031 , n7032 , n7076 , n7078 , n7079 , n7080 , n7125 , n7127 , n7128 , n7130 , n7131 , n7132 , n7182 , n7184 , n7185 , n7186 , n7237 , n7248 , n7249 , n7251 , n7252 , n7253 , n7289 , n7291 , n7292 , n7294 , n7295 , n7296 , n7330 , n7332 , n7333 , n7334 , n7369 , n7370 , n7371 , n7409 , n7410 , n7411 , n7415 , n7416 , n7417 , n7419 , n7422 , n7424 , n7426 , n7427 , n7428 , n7430 , n7431 , n7432 , n7434 , n7435 , n7436 , n7438 , n7439 , n7440 , n7442 , n7443 , n7444 , n7446 , n7447 , n7448 , n7453 , n7455 , n7460 , n7461 , n7462 , n7464 , n7465 , n7466 , n7468 , n7469 , n7470 , n7472 , n7474 , n7475 , n7476 , n7480 , n7485 , n7486 , n7487 , n7489 , n7490 , n7491 , n7494 , n7495 , n7496 , n7497 , n7499 , n7501 , n7502 , n7503 , n7505 , n7506 , n7507 , n7509 , n7510 , n7511 , n7516 , n7517 , n7518 , n7523 , n7524 , n7525 , n7527 , n7531 , n7533 , n7535 , n7536 , n7537 , n7539 , n7540 , n7541 , n7543 , n7544 , n7545 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7554 , n7555 , n7556 , n7558 , n7559 , n7560 , n7565 , n7567 , n7569 , n7571 , n7572 , n7573 , n7578 , n7579 , n7580 , n7582 , n7583 , n7584 , n7586 , n7587 , n7588 , n7590 , n7591 , n7592 , n7594 , n7595 , n7596 , n7597 , n7598 , n7644 , n7646 , n7647 , n7649 , n7650 , n7651 , n7653 , n7654 , n7655 , n7657 , n7658 , n7659 , n7661 , n7662 , n7663 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7676 , n7677 , n7678 , n7680 , n7681 , n7682 , n7686 , n7687 , n7689 , n7690 , n7691 , n7694 , n7695 , n7696 , n7698 , n7699 , n7700 , n7702 , n7703 , n7704 , n7708 , n7709 , n7710 , n7712 , n7713 , n7714 , n7716 , n7717 , n7718 , n7720 , n7721 , n7722 , n7724 , n7725 , n7726 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7736 , n7737 , n7738 , n7740 , n7741 , n7742 , n7744 , n7745 , n7746 , n7750 , n7751 , n7752 , n7754 , n7755 , n7756 , n7759 , n7760 , n7761 , n7763 , n7764 , n7765 , n7767 , n7768 , n7769 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7781 , n7782 , n7783 , n7785 , n7786 , n7787 , n7792 , n7793 , n7794 , n7796 , n7797 , n7798 , n7800 , n7801 , n7802 , n7804 , n7805 , n7806 , n7808 , n7809 , n7810 , n7812 , n7813 , n7814 , n7816 , n7817 , n7818 , n7819 , n7820 , n7867 , n7872 , n7873 , n7874 , n7876 , n7877 , n7878 , n7880 , n7881 , n7882 , n7884 , n7885 , n7886 , n7890 , n7895 , n7896 , n7897 , n7899 , n7900 , n7901 , n7905 , n7906 , n7907 , n7912 , n7913 , n7914 , n7916 , n7917 , n7918 , n7920 , n7921 , n7922 , n7924 , n7925 , n7926 , n7928 , n7929 , n7930 , n7934 , n7936 , n7938 , n7939 , n7940 , n7942 , n7943 , n7944 , n7949 , n7950 , n7951 , n7952 , n7953 , n7955 , n7957 , n7958 , n7959 , n7964 , n7965 , n7966 , n7968 , n7969 , n7970 , n7972 , n7973 , n7974 , n7976 , n7977 , n7978 , n7980 , n7981 , n7982 , n7984 , n7985 , n7986 , n7988 , n7989 , n7990 , n7995 , n7996 , n7997 , n7998 , n8000 , n8002 , n8004 , n8006 , n8007 , n8008 , n8013 , n8014 , n8015 , n8017 , n8018 , n8019 , n8021 , n8022 , n8023 , n8025 , n8026 , n8027 , n8029 , n8030 , n8031 , n8033 , n8034 , n8035 , n8037 , n8038 , n8039 , n8044 , n8045 , n8046 , n8047 , n8048 , n8094 , n8096 , n8098 , n8119 , n8121 , n8123 , n8133 , n8167 , n8192 , n8194 , n8195 , n8197 , n8198 , n8199 , n8220 , n8222 , n8223 , n8224 , n8246 , n8247 , n8249 , n8250 , n8251 , n8274 , n8276 , n8277 , n8278 , n8296 , n8297 , n8329 , n8330 , n8332 , n8333 , n8334 , n8346 , n8348 , n8349 , n8350 , n8363 , n8364 , n8366 , n8367 , n8368 , n8382 , n8384 , n8385 , n8386 , n8393 , n8394 , n8395 , n8460 , n8461 , n8462 , n8527 , n8528 , n8529 , n8530 , n8595 , n8596 , n8597 , n8662 , n8663 , n8681 , n8682 , n8683 , n8726 , n8760 , n8761 , n8762 , n8782 , n8783 , n8785 , n8786 , n8787 , n8807 , n8842 , n8843 , n8845 , n8846 , n8847 , n8867 , n8902 , n8903 , n8904 , n8922 , n8924 , n8926 , n8928 , n8961 , n8962 , n8963 , n8965 , n8966 , n8967 , n8969 , n8971 , n8975 , n8976 , n8977 , n8978 , n8986 , n8987 , n9022 , n9035 , n9036 , n9038 , n9039 , n9040 , n9073 , n9098 , n9099 , n9101 , n9102 , n9103 , n9132 , n9134 , n9135 , n9136 , n9166 , n9192 , n9193 , n9194 , n9223 , n9249 , n9250 , n9252 , n9253 , n9254 , n9283 , n9284 , n9286 , n9287 , n9288 , n9317 , n9318 , n9319 , n9348 , n9413 , n9414 , n9478 , n9480 , n9487 , n9488 , n9489 , n9491 , n9493 , n9495 , n9496 , n9497 , n9499 , n9500 , n9501 , n9507 , n9508 , n9509 , n9514 , n9515 , n9516 , n9532 , n9533 , n9535 , n9537 , n9538 , n9539 , n9542 , n9544 , n9545 , n9550 , n9551 , n9552 , n9570 , n9571 , n9573 , n9574 , n9599 , n9600 , n9601 , n9604 , n9606 , n9609 , n9610 , n9612 , n9614 , n9615 , n9616 , n9618 , n9619 , n9620 , n9622 , n9623 , n9624 , n9651 , n9652 , n9653 , n9655 , n9656 , n9657 , n9664 , n9665 , n9667 , n9668 , n9669 , n9671 , n9672 , n9673 , n9675 , n9676 , n9677 , n9700 , n9701 , n9703 , n9704 , n9705 , n9721 , n9722 , n9724 , n9725 , n9726 , n9728 , n9729 , n9730 , n9732 , n9734 , n9741 , n9742 , n9743 , n9745 , n9753 , n9755 , n9757 , n9758 , n9759 , n9761 , n9762 , n9763 , n9769 , n9770 , n9771 , n9776 , n9777 , n9778 , n9805 , n9806 , n9808 , n9810 , n9811 , n9812 , n9815 , n9817 , n9818 , n9823 , n9824 , n9825 , n9854 , n9855 , n9857 , n9858 , n9859 , n9864 , n9865 , n9866 , n9868 , n9870 , n9872 , n9873 , n9875 , n9876 , n9877 , n9879 , n9880 , n9881 , n9883 , n9884 , n9885 , n9901 , n9902 , n9903 , n9905 , n9906 , n9907 , n9909 , n9910 , n9914 , n9916 , n9917 , n9918 , n9920 , n9921 , n9922 , n9937 , n9938 , n9940 , n9942 , n9944 , n9945 , n9946 , n9948 , n9949 , n9950 , n9955 , n9956 , n9957 , n9963 , n9964 , n9965 , n9967 , n9969 , n9973 , n9974 , n9979 , n9980 , n9981 , n9987 , n9988 , n9989 , n9992 , n9993 , n9995 , n9996 , n10014 , n10015 , n10016 , n10020 , n10021 , n10022 , n10048 , n10049 , n10053 , n10057 , n10058 , n10059 , n10061 , n10062 , n10068 , n10069 , n10070 , n10073 , n10074 , n10075 , n10077 , n10079 , n10080 , n10081 , n10084 , n10087 , n10088 , n10090 , n10091 , n10093 , n10094 , n10095 , n10097 , n10098 , n10099 , n10100 , n10101 , n10103 , n10104 , n10106 , n10111 , n10113 , n10118 , n10125 , n10127 , n10129 , n10130 , n10131 , n10135 , n10136 , n10137 , n10139 , n10141 , n10142 , n10143 , n10146 , n10148 , n10152 , n10153 , n10154 , n10158 , n10159 , n10160 , n10165 , n10166 , n10167 , n10169 , n10171 , n10172 , n10173 , n10174 , n10176 , n10177 , n10178 , n10193 , n10194 , n10195 , n10197 , n10198 , n10199 , n10232 , n10296 ;
  buffer buf_n3312( .i (N367), .o (n3312) );
  buffer buf_n3313( .i (n3312), .o (n3313) );
  buffer buf_n3314( .i (n3313), .o (n3314) );
  buffer buf_n3315( .i (n3314), .o (n3315) );
  buffer buf_n3316( .i (n3315), .o (n3316) );
  buffer buf_n3317( .i (n3316), .o (n3317) );
  buffer buf_n3318( .i (n3317), .o (n3318) );
  buffer buf_n3319( .i (n3318), .o (n3319) );
  buffer buf_n3320( .i (n3319), .o (n3320) );
  buffer buf_n3321( .i (n3320), .o (n3321) );
  buffer buf_n2050( .i (N310), .o (n2050) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  buffer buf_n2055( .i (n2054), .o (n2055) );
  buffer buf_n586( .i (N18), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n3447( .i (N41), .o (n3447) );
  buffer buf_n3448( .i (n3447), .o (n3448) );
  buffer buf_n3449( .i (n3448), .o (n3449) );
  buffer buf_n3450( .i (n3449), .o (n3450) );
  assign n3608 = ~n589 & n3450 ;
  buffer buf_n3609( .i (n3608), .o (n3609) );
  assign n3610 = ~n2055 & n3609 ;
  buffer buf_n3611( .i (n3610), .o (n3611) );
  assign n3616 = n589 | n3450 ;
  assign n3617 = n2054 & ~n3616 ;
  buffer buf_n3618( .i (n3617), .o (n3618) );
  buffer buf_n3619( .i (n3618), .o (n3619) );
  assign n3625 = n3611 | n3619 ;
  buffer buf_n3626( .i (n3625), .o (n3626) );
  assign n3629 = n3321 & ~n3626 ;
  buffer buf_n3630( .i (n3629), .o (n3630) );
  assign n3631 = ~n3321 & n3626 ;
  buffer buf_n3632( .i (n3631), .o (n3632) );
  assign n3633 = n3630 | n3632 ;
  buffer buf_n3634( .i (n3633), .o (n3634) );
  buffer buf_n3635( .i (n3634), .o (n3635) );
  buffer buf_n3636( .i (n3635), .o (n3636) );
  buffer buf_n3637( .i (n3636), .o (n3637) );
  buffer buf_n3638( .i (n3637), .o (n3638) );
  buffer buf_n3639( .i (n3638), .o (n3639) );
  buffer buf_n3640( .i (n3639), .o (n3640) );
  buffer buf_n3641( .i (n3640), .o (n3641) );
  buffer buf_n3642( .i (n3641), .o (n3642) );
  buffer buf_n3643( .i (n3642), .o (n3643) );
  buffer buf_n3644( .i (n3643), .o (n3644) );
  buffer buf_n3645( .i (n3644), .o (n3645) );
  buffer buf_n3646( .i (n3645), .o (n3646) );
  buffer buf_n3647( .i (n3646), .o (n3647) );
  buffer buf_n3648( .i (n3647), .o (n3648) );
  buffer buf_n3649( .i (n3648), .o (n3649) );
  buffer buf_n3650( .i (n3649), .o (n3650) );
  buffer buf_n3651( .i (n3650), .o (n3651) );
  buffer buf_n3652( .i (n3651), .o (n3652) );
  buffer buf_n3653( .i (n3652), .o (n3653) );
  buffer buf_n3654( .i (n3653), .o (n3654) );
  buffer buf_n3655( .i (n3654), .o (n3655) );
  buffer buf_n3656( .i (n3655), .o (n3656) );
  buffer buf_n3657( .i (n3656), .o (n3657) );
  buffer buf_n3658( .i (n3657), .o (n3658) );
  buffer buf_n3659( .i (n3658), .o (n3659) );
  buffer buf_n3660( .i (n3659), .o (n3660) );
  buffer buf_n3661( .i (n3660), .o (n3661) );
  buffer buf_n3662( .i (n3661), .o (n3662) );
  buffer buf_n3663( .i (n3662), .o (n3663) );
  buffer buf_n3664( .i (n3663), .o (n3664) );
  buffer buf_n3665( .i (n3664), .o (n3665) );
  buffer buf_n3666( .i (n3665), .o (n3666) );
  buffer buf_n3667( .i (n3666), .o (n3667) );
  buffer buf_n3668( .i (n3667), .o (n3668) );
  buffer buf_n3669( .i (n3668), .o (n3669) );
  buffer buf_n3670( .i (n3669), .o (n3670) );
  buffer buf_n3671( .i (n3670), .o (n3671) );
  buffer buf_n3672( .i (n3671), .o (n3672) );
  buffer buf_n3673( .i (n3672), .o (n3673) );
  buffer buf_n3674( .i (n3673), .o (n3674) );
  buffer buf_n3675( .i (n3674), .o (n3675) );
  buffer buf_n3676( .i (n3675), .o (n3676) );
  buffer buf_n3677( .i (n3676), .o (n3677) );
  buffer buf_n3678( .i (n3677), .o (n3678) );
  buffer buf_n3679( .i (n3678), .o (n3679) );
  buffer buf_n3680( .i (n3679), .o (n3680) );
  buffer buf_n3681( .i (n3680), .o (n3681) );
  buffer buf_n3682( .i (n3681), .o (n3682) );
  buffer buf_n3683( .i (n3682), .o (n3683) );
  buffer buf_n3684( .i (n3683), .o (n3684) );
  buffer buf_n3685( .i (n3684), .o (n3685) );
  buffer buf_n3686( .i (n3685), .o (n3686) );
  buffer buf_n3337( .i (N38), .o (n3337) );
  buffer buf_n3338( .i (n3337), .o (n3338) );
  buffer buf_n3339( .i (n3338), .o (n3339) );
  buffer buf_n3340( .i (n3339), .o (n3340) );
  buffer buf_n1253( .i (N267), .o (n1253) );
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n3393( .i (N382), .o (n3393) );
  buffer buf_n3394( .i (n3393), .o (n3394) );
  assign n3687 = n1254 & n3394 ;
  buffer buf_n3688( .i (n3687), .o (n3688) );
  assign n3748 = ~n3340 & n3688 ;
  buffer buf_n3749( .i (n3748), .o (n3749) );
  buffer buf_n3750( .i (n3749), .o (n3750) );
  buffer buf_n3751( .i (n3750), .o (n3751) );
  buffer buf_n3752( .i (n3751), .o (n3752) );
  buffer buf_n3753( .i (n3752), .o (n3753) );
  buffer buf_n3754( .i (n3753), .o (n3754) );
  buffer buf_n3755( .i (n3754), .o (n3755) );
  buffer buf_n3756( .i (n3755), .o (n3756) );
  buffer buf_n3757( .i (n3756), .o (n3757) );
  buffer buf_n3758( .i (n3757), .o (n3758) );
  buffer buf_n3759( .i (n3758), .o (n3759) );
  buffer buf_n3760( .i (n3759), .o (n3760) );
  buffer buf_n3761( .i (n3760), .o (n3761) );
  buffer buf_n3762( .i (n3761), .o (n3762) );
  buffer buf_n3763( .i (n3762), .o (n3763) );
  buffer buf_n3764( .i (n3763), .o (n3764) );
  buffer buf_n3765( .i (n3764), .o (n3765) );
  buffer buf_n3766( .i (n3765), .o (n3766) );
  buffer buf_n3767( .i (n3766), .o (n3767) );
  buffer buf_n3768( .i (n3767), .o (n3768) );
  buffer buf_n3769( .i (n3768), .o (n3769) );
  buffer buf_n3770( .i (n3769), .o (n3770) );
  buffer buf_n3771( .i (n3770), .o (n3771) );
  buffer buf_n3772( .i (n3771), .o (n3772) );
  buffer buf_n3773( .i (n3772), .o (n3773) );
  buffer buf_n3774( .i (n3773), .o (n3774) );
  buffer buf_n3775( .i (n3774), .o (n3775) );
  buffer buf_n3776( .i (n3775), .o (n3776) );
  buffer buf_n3777( .i (n3776), .o (n3777) );
  buffer buf_n3778( .i (n3777), .o (n3778) );
  buffer buf_n3779( .i (n3778), .o (n3779) );
  buffer buf_n3780( .i (n3779), .o (n3780) );
  buffer buf_n3781( .i (n3780), .o (n3781) );
  buffer buf_n3782( .i (n3781), .o (n3782) );
  buffer buf_n3783( .i (n3782), .o (n3783) );
  buffer buf_n3784( .i (n3783), .o (n3784) );
  buffer buf_n3785( .i (n3784), .o (n3785) );
  buffer buf_n3786( .i (n3785), .o (n3786) );
  buffer buf_n3787( .i (n3786), .o (n3787) );
  buffer buf_n3788( .i (n3787), .o (n3788) );
  buffer buf_n3789( .i (n3788), .o (n3789) );
  buffer buf_n3790( .i (n3789), .o (n3790) );
  buffer buf_n3791( .i (n3790), .o (n3791) );
  buffer buf_n3792( .i (n3791), .o (n3792) );
  buffer buf_n3793( .i (n3792), .o (n3793) );
  buffer buf_n3794( .i (n3793), .o (n3794) );
  buffer buf_n3795( .i (n3794), .o (n3795) );
  buffer buf_n3796( .i (n3795), .o (n3796) );
  buffer buf_n3797( .i (n3796), .o (n3797) );
  buffer buf_n3798( .i (n3797), .o (n3798) );
  buffer buf_n3799( .i (n3798), .o (n3799) );
  buffer buf_n3800( .i (n3799), .o (n3800) );
  buffer buf_n3801( .i (n3800), .o (n3801) );
  buffer buf_n3802( .i (n3801), .o (n3802) );
  buffer buf_n3803( .i (n3802), .o (n3803) );
  buffer buf_n3804( .i (n3803), .o (n3804) );
  buffer buf_n3805( .i (n3804), .o (n3805) );
  buffer buf_n3806( .i (n3805), .o (n3806) );
  buffer buf_n3341( .i (n3340), .o (n3341) );
  buffer buf_n1187( .i (N263), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  assign n3807 = n1190 & n3688 ;
  assign n3808 = n3341 & ~n3807 ;
  buffer buf_n3809( .i (n3808), .o (n3809) );
  buffer buf_n3810( .i (n3809), .o (n3810) );
  buffer buf_n3811( .i (n3810), .o (n3811) );
  buffer buf_n3812( .i (n3811), .o (n3812) );
  buffer buf_n3813( .i (n3812), .o (n3813) );
  buffer buf_n3814( .i (n3813), .o (n3814) );
  buffer buf_n3815( .i (n3814), .o (n3815) );
  buffer buf_n3816( .i (n3815), .o (n3816) );
  buffer buf_n3817( .i (n3816), .o (n3817) );
  buffer buf_n3818( .i (n3817), .o (n3818) );
  buffer buf_n3819( .i (n3818), .o (n3819) );
  buffer buf_n3820( .i (n3819), .o (n3820) );
  buffer buf_n3821( .i (n3820), .o (n3821) );
  buffer buf_n3822( .i (n3821), .o (n3822) );
  buffer buf_n3823( .i (n3822), .o (n3823) );
  buffer buf_n3824( .i (n3823), .o (n3824) );
  buffer buf_n3825( .i (n3824), .o (n3825) );
  buffer buf_n3826( .i (n3825), .o (n3826) );
  buffer buf_n3827( .i (n3826), .o (n3827) );
  buffer buf_n3828( .i (n3827), .o (n3828) );
  buffer buf_n3829( .i (n3828), .o (n3829) );
  buffer buf_n3830( .i (n3829), .o (n3830) );
  buffer buf_n3831( .i (n3830), .o (n3831) );
  buffer buf_n3832( .i (n3831), .o (n3832) );
  buffer buf_n3833( .i (n3832), .o (n3833) );
  buffer buf_n3834( .i (n3833), .o (n3834) );
  buffer buf_n3835( .i (n3834), .o (n3835) );
  buffer buf_n3836( .i (n3835), .o (n3836) );
  buffer buf_n3837( .i (n3836), .o (n3837) );
  buffer buf_n3838( .i (n3837), .o (n3838) );
  buffer buf_n3839( .i (n3838), .o (n3839) );
  buffer buf_n3840( .i (n3839), .o (n3840) );
  buffer buf_n3841( .i (n3840), .o (n3841) );
  buffer buf_n3842( .i (n3841), .o (n3842) );
  buffer buf_n3843( .i (n3842), .o (n3843) );
  buffer buf_n3844( .i (n3843), .o (n3844) );
  buffer buf_n3845( .i (n3844), .o (n3845) );
  buffer buf_n3846( .i (n3845), .o (n3846) );
  buffer buf_n3847( .i (n3846), .o (n3847) );
  buffer buf_n3848( .i (n3847), .o (n3848) );
  buffer buf_n3849( .i (n3848), .o (n3849) );
  buffer buf_n3850( .i (n3849), .o (n3850) );
  buffer buf_n3851( .i (n3850), .o (n3851) );
  buffer buf_n3852( .i (n3851), .o (n3852) );
  buffer buf_n3853( .i (n3852), .o (n3853) );
  buffer buf_n3854( .i (n3853), .o (n3854) );
  buffer buf_n3855( .i (n3854), .o (n3855) );
  buffer buf_n3856( .i (n3855), .o (n3856) );
  buffer buf_n3857( .i (n3856), .o (n3857) );
  buffer buf_n3858( .i (n3857), .o (n3858) );
  buffer buf_n3859( .i (n3858), .o (n3859) );
  buffer buf_n3860( .i (n3859), .o (n3860) );
  buffer buf_n3861( .i (n3860), .o (n3861) );
  buffer buf_n3862( .i (n3861), .o (n3862) );
  buffer buf_n3863( .i (n3862), .o (n3863) );
  buffer buf_n3864( .i (n3863), .o (n3864) );
  buffer buf_n3342( .i (n3341), .o (n3342) );
  buffer buf_n3343( .i (n3342), .o (n3343) );
  buffer buf_n3344( .i (n3343), .o (n3344) );
  buffer buf_n3345( .i (n3344), .o (n3345) );
  buffer buf_n3346( .i (n3345), .o (n3346) );
  buffer buf_n3347( .i (n3346), .o (n3347) );
  buffer buf_n3348( .i (n3347), .o (n3348) );
  buffer buf_n3349( .i (n3348), .o (n3349) );
  buffer buf_n3350( .i (n3349), .o (n3350) );
  buffer buf_n3351( .i (n3350), .o (n3351) );
  buffer buf_n3352( .i (n3351), .o (n3352) );
  buffer buf_n3353( .i (n3352), .o (n3353) );
  buffer buf_n3354( .i (n3353), .o (n3354) );
  buffer buf_n3355( .i (n3354), .o (n3355) );
  buffer buf_n3356( .i (n3355), .o (n3356) );
  buffer buf_n3357( .i (n3356), .o (n3357) );
  buffer buf_n3358( .i (n3357), .o (n3358) );
  buffer buf_n3359( .i (n3358), .o (n3359) );
  buffer buf_n3360( .i (n3359), .o (n3360) );
  buffer buf_n3361( .i (n3360), .o (n3361) );
  buffer buf_n3362( .i (n3361), .o (n3362) );
  buffer buf_n3363( .i (n3362), .o (n3363) );
  buffer buf_n3364( .i (n3363), .o (n3364) );
  buffer buf_n3365( .i (n3364), .o (n3365) );
  buffer buf_n3366( .i (n3365), .o (n3366) );
  buffer buf_n3367( .i (n3366), .o (n3367) );
  buffer buf_n3368( .i (n3367), .o (n3368) );
  buffer buf_n3369( .i (n3368), .o (n3369) );
  buffer buf_n3370( .i (n3369), .o (n3370) );
  buffer buf_n3371( .i (n3370), .o (n3371) );
  buffer buf_n3372( .i (n3371), .o (n3372) );
  buffer buf_n3373( .i (n3372), .o (n3373) );
  buffer buf_n3374( .i (n3373), .o (n3374) );
  buffer buf_n3375( .i (n3374), .o (n3375) );
  buffer buf_n3376( .i (n3375), .o (n3376) );
  buffer buf_n3377( .i (n3376), .o (n3377) );
  buffer buf_n3378( .i (n3377), .o (n3378) );
  buffer buf_n3379( .i (n3378), .o (n3379) );
  buffer buf_n3380( .i (n3379), .o (n3380) );
  buffer buf_n3381( .i (n3380), .o (n3381) );
  buffer buf_n3382( .i (n3381), .o (n3382) );
  buffer buf_n3383( .i (n3382), .o (n3383) );
  buffer buf_n3384( .i (n3383), .o (n3384) );
  buffer buf_n3385( .i (n3384), .o (n3385) );
  buffer buf_n3386( .i (n3385), .o (n3386) );
  buffer buf_n3387( .i (n3386), .o (n3387) );
  buffer buf_n3388( .i (n3387), .o (n3388) );
  buffer buf_n3389( .i (n3388), .o (n3389) );
  buffer buf_n3390( .i (n3389), .o (n3390) );
  buffer buf_n3391( .i (n3390), .o (n3391) );
  buffer buf_n3392( .i (n3391), .o (n3392) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n3395( .i (n3394), .o (n3395) );
  buffer buf_n3396( .i (n3395), .o (n3396) );
  buffer buf_n3397( .i (n3396), .o (n3397) );
  buffer buf_n3398( .i (n3397), .o (n3398) );
  buffer buf_n3399( .i (n3398), .o (n3399) );
  buffer buf_n3400( .i (n3399), .o (n3400) );
  buffer buf_n3401( .i (n3400), .o (n3401) );
  buffer buf_n3402( .i (n3401), .o (n3402) );
  buffer buf_n3403( .i (n3402), .o (n3403) );
  buffer buf_n3404( .i (n3403), .o (n3404) );
  buffer buf_n3405( .i (n3404), .o (n3405) );
  buffer buf_n3406( .i (n3405), .o (n3406) );
  buffer buf_n3407( .i (n3406), .o (n3407) );
  buffer buf_n3408( .i (n3407), .o (n3408) );
  buffer buf_n3409( .i (n3408), .o (n3409) );
  buffer buf_n3410( .i (n3409), .o (n3410) );
  buffer buf_n3411( .i (n3410), .o (n3411) );
  buffer buf_n3412( .i (n3411), .o (n3412) );
  buffer buf_n3413( .i (n3412), .o (n3413) );
  buffer buf_n3414( .i (n3413), .o (n3414) );
  buffer buf_n3415( .i (n3414), .o (n3415) );
  buffer buf_n3416( .i (n3415), .o (n3416) );
  buffer buf_n3417( .i (n3416), .o (n3417) );
  buffer buf_n3418( .i (n3417), .o (n3418) );
  buffer buf_n3419( .i (n3418), .o (n3419) );
  buffer buf_n3420( .i (n3419), .o (n3420) );
  buffer buf_n3421( .i (n3420), .o (n3421) );
  buffer buf_n3422( .i (n3421), .o (n3422) );
  buffer buf_n3423( .i (n3422), .o (n3423) );
  buffer buf_n3424( .i (n3423), .o (n3424) );
  buffer buf_n3425( .i (n3424), .o (n3425) );
  buffer buf_n3426( .i (n3425), .o (n3426) );
  buffer buf_n3427( .i (n3426), .o (n3427) );
  buffer buf_n3428( .i (n3427), .o (n3428) );
  buffer buf_n3429( .i (n3428), .o (n3429) );
  buffer buf_n3430( .i (n3429), .o (n3430) );
  buffer buf_n3431( .i (n3430), .o (n3431) );
  buffer buf_n3432( .i (n3431), .o (n3432) );
  buffer buf_n3433( .i (n3432), .o (n3433) );
  buffer buf_n3434( .i (n3433), .o (n3434) );
  buffer buf_n3435( .i (n3434), .o (n3435) );
  buffer buf_n3436( .i (n3435), .o (n3436) );
  buffer buf_n3437( .i (n3436), .o (n3437) );
  buffer buf_n3438( .i (n3437), .o (n3438) );
  buffer buf_n3439( .i (n3438), .o (n3439) );
  buffer buf_n3440( .i (n3439), .o (n3440) );
  buffer buf_n3441( .i (n3440), .o (n3441) );
  buffer buf_n3442( .i (n3441), .o (n3442) );
  buffer buf_n3443( .i (n3442), .o (n3443) );
  buffer buf_n3444( .i (n3443), .o (n3444) );
  buffer buf_n3445( .i (n3444), .o (n3445) );
  buffer buf_n3446( .i (n3445), .o (n3446) );
  assign n3865 = n1240 & n3446 ;
  buffer buf_n3866( .i (n3865), .o (n3866) );
  assign n3867 = n3392 & n3866 ;
  buffer buf_n3868( .i (n3867), .o (n3868) );
  assign n3872 = n3392 | n3866 ;
  buffer buf_n3873( .i (n3872), .o (n3873) );
  assign n3876 = ~n3868 & n3873 ;
  buffer buf_n3877( .i (n3876), .o (n3877) );
  buffer buf_n1121( .i (N260), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  assign n3878 = N12 & N9 ;
  buffer buf_n3879( .i (n3878), .o (n3879) );
  buffer buf_n3880( .i (n3879), .o (n3880) );
  buffer buf_n3881( .i (n3880), .o (n3881) );
  buffer buf_n3882( .i (n3881), .o (n3882) );
  buffer buf_n3883( .i (n3882), .o (n3883) );
  buffer buf_n685( .i (N213), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  assign n3885 = n589 & ~n688 ;
  buffer buf_n3886( .i (n3885), .o (n3886) );
  assign n3889 = n3883 | n3886 ;
  buffer buf_n3890( .i (n3889), .o (n3890) );
  assign n3891 = n1128 | n3890 ;
  buffer buf_n3892( .i (n3891), .o (n3892) );
  buffer buf_n3893( .i (n3892), .o (n3893) );
  buffer buf_n1051( .i (N257), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n689( .i (N214), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n3894( .i (n588), .o (n3894) );
  assign n3895 = ~n692 & n3894 ;
  buffer buf_n3896( .i (n3895), .o (n3896) );
  assign n3899 = n3883 | n3896 ;
  buffer buf_n3900( .i (n3899), .o (n3900) );
  assign n3901 = n1058 | n3900 ;
  buffer buf_n3902( .i (n3901), .o (n3902) );
  assign n3912 = n1128 & n3890 ;
  buffer buf_n3913( .i (n3912), .o (n3913) );
  assign n3914 = n3902 | n3913 ;
  assign n3915 = n3893 & n3914 ;
  buffer buf_n3916( .i (n3915), .o (n3916) );
  buffer buf_n3917( .i (n3916), .o (n3917) );
  buffer buf_n3918( .i (n3917), .o (n3918) );
  buffer buf_n3919( .i (n3918), .o (n3919) );
  buffer buf_n3920( .i (n3919), .o (n3920) );
  buffer buf_n3921( .i (n3920), .o (n3921) );
  buffer buf_n3922( .i (n3921), .o (n3922) );
  buffer buf_n3923( .i (n3922), .o (n3923) );
  buffer buf_n3924( .i (n3923), .o (n3924) );
  buffer buf_n3925( .i (n3924), .o (n3925) );
  buffer buf_n3926( .i (n3925), .o (n3926) );
  buffer buf_n3927( .i (n3926), .o (n3927) );
  buffer buf_n3928( .i (n3927), .o (n3928) );
  buffer buf_n3929( .i (n3928), .o (n3929) );
  buffer buf_n3930( .i (n3929), .o (n3930) );
  buffer buf_n3931( .i (n3930), .o (n3931) );
  buffer buf_n3932( .i (n3931), .o (n3932) );
  buffer buf_n3933( .i (n3932), .o (n3933) );
  buffer buf_n3934( .i (n3933), .o (n3934) );
  buffer buf_n3935( .i (n3934), .o (n3935) );
  buffer buf_n3936( .i (n3935), .o (n3936) );
  buffer buf_n3937( .i (n3936), .o (n3937) );
  buffer buf_n3938( .i (n3937), .o (n3938) );
  buffer buf_n3939( .i (n3938), .o (n3939) );
  buffer buf_n3940( .i (n3939), .o (n3940) );
  buffer buf_n3941( .i (n3940), .o (n3941) );
  buffer buf_n3942( .i (n3941), .o (n3942) );
  buffer buf_n3943( .i (n3942), .o (n3943) );
  buffer buf_n3944( .i (n3943), .o (n3944) );
  buffer buf_n3945( .i (n3944), .o (n3945) );
  buffer buf_n3946( .i (n3945), .o (n3946) );
  buffer buf_n3947( .i (n3946), .o (n3947) );
  buffer buf_n3948( .i (n3947), .o (n3948) );
  buffer buf_n3949( .i (n3948), .o (n3949) );
  buffer buf_n3950( .i (n3949), .o (n3950) );
  buffer buf_n3951( .i (n3950), .o (n3951) );
  buffer buf_n3952( .i (n3951), .o (n3952) );
  buffer buf_n3953( .i (n3952), .o (n3953) );
  buffer buf_n282( .i (N106), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n693( .i (N215), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  assign n3954 = ~n696 & n3894 ;
  buffer buf_n3955( .i (n3954), .o (n3955) );
  assign n3958 = n3883 | n3955 ;
  buffer buf_n3959( .i (n3958), .o (n3959) );
  assign n3960 = n289 | n3959 ;
  buffer buf_n3961( .i (n3960), .o (n3961) );
  buffer buf_n3962( .i (n3961), .o (n3962) );
  buffer buf_n3963( .i (n3962), .o (n3963) );
  buffer buf_n3964( .i (n3963), .o (n3964) );
  buffer buf_n3965( .i (n3964), .o (n3965) );
  buffer buf_n3966( .i (n3965), .o (n3966) );
  assign n3967 = n289 & n3959 ;
  buffer buf_n3968( .i (n3967), .o (n3968) );
  buffer buf_n3969( .i (n3968), .o (n3969) );
  buffer buf_n3970( .i (n3969), .o (n3970) );
  buffer buf_n3971( .i (n3970), .o (n3971) );
  buffer buf_n3972( .i (n3971), .o (n3972) );
  buffer buf_n985( .i (N254), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n697( .i (N216), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  assign n3973 = ~n700 & n3894 ;
  buffer buf_n3974( .i (n3973), .o (n3974) );
  buffer buf_n3977( .i (n3882), .o (n3977) );
  assign n3978 = n3974 | n3977 ;
  buffer buf_n3979( .i (n3978), .o (n3979) );
  assign n3980 = n992 & n3979 ;
  buffer buf_n3981( .i (n3980), .o (n3981) );
  buffer buf_n3982( .i (n3981), .o (n3982) );
  buffer buf_n3983( .i (n3982), .o (n3983) );
  buffer buf_n919( .i (N251), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n679( .i (N209), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  assign n3984 = ~n682 & n3894 ;
  buffer buf_n3985( .i (n3984), .o (n3985) );
  assign n3986 = n3977 | n3985 ;
  buffer buf_n3987( .i (n3986), .o (n3987) );
  assign n3988 = n926 | n3987 ;
  buffer buf_n3989( .i (n3988), .o (n3989) );
  assign n4036 = n992 | n3979 ;
  buffer buf_n4037( .i (n4036), .o (n4037) );
  assign n4038 = n3989 & n4037 ;
  buffer buf_n4039( .i (n4038), .o (n4039) );
  assign n4040 = n3983 | n4039 ;
  buffer buf_n4041( .i (n4040), .o (n4041) );
  assign n4077 = n3972 | n4041 ;
  assign n4078 = n3966 & n4077 ;
  buffer buf_n4079( .i (n4078), .o (n4079) );
  buffer buf_n4080( .i (n4079), .o (n4080) );
  buffer buf_n4081( .i (n4080), .o (n4081) );
  buffer buf_n4082( .i (n4081), .o (n4082) );
  buffer buf_n4083( .i (n4082), .o (n4083) );
  buffer buf_n4084( .i (n4083), .o (n4084) );
  buffer buf_n4085( .i (n4084), .o (n4085) );
  buffer buf_n4086( .i (n4085), .o (n4086) );
  buffer buf_n4087( .i (n4086), .o (n4087) );
  buffer buf_n4088( .i (n4087), .o (n4088) );
  buffer buf_n4089( .i (n4088), .o (n4089) );
  buffer buf_n4090( .i (n4089), .o (n4090) );
  buffer buf_n4091( .i (n4090), .o (n4091) );
  buffer buf_n4092( .i (n4091), .o (n4092) );
  buffer buf_n4093( .i (n4092), .o (n4093) );
  buffer buf_n4094( .i (n4093), .o (n4094) );
  buffer buf_n4095( .i (n4094), .o (n4095) );
  buffer buf_n4096( .i (n4095), .o (n4096) );
  buffer buf_n4097( .i (n4096), .o (n4097) );
  buffer buf_n4098( .i (n4097), .o (n4098) );
  buffer buf_n4099( .i (n4098), .o (n4099) );
  buffer buf_n4100( .i (n4099), .o (n4100) );
  buffer buf_n4101( .i (n4100), .o (n4101) );
  buffer buf_n4102( .i (n4101), .o (n4102) );
  buffer buf_n4103( .i (n4102), .o (n4103) );
  buffer buf_n4104( .i (n4103), .o (n4104) );
  buffer buf_n4105( .i (n4104), .o (n4105) );
  buffer buf_n4106( .i (n4105), .o (n4106) );
  buffer buf_n4107( .i (n4106), .o (n4107) );
  buffer buf_n4108( .i (n4107), .o (n4108) );
  buffer buf_n4109( .i (n4108), .o (n4109) );
  buffer buf_n4110( .i (n4109), .o (n4110) );
  buffer buf_n4111( .i (n4110), .o (n4111) );
  assign n4113 = n1058 & n3900 ;
  buffer buf_n4114( .i (n4113), .o (n4114) );
  assign n4123 = n3902 & ~n4114 ;
  buffer buf_n4124( .i (n4123), .o (n4124) );
  buffer buf_n4125( .i (n4124), .o (n4125) );
  buffer buf_n4126( .i (n4125), .o (n4126) );
  buffer buf_n4127( .i (n4126), .o (n4127) );
  buffer buf_n4128( .i (n4127), .o (n4128) );
  buffer buf_n4129( .i (n4128), .o (n4129) );
  buffer buf_n4130( .i (n4129), .o (n4130) );
  buffer buf_n4131( .i (n4130), .o (n4131) );
  buffer buf_n4132( .i (n4131), .o (n4132) );
  buffer buf_n4133( .i (n4132), .o (n4133) );
  buffer buf_n4134( .i (n4133), .o (n4134) );
  buffer buf_n4135( .i (n4134), .o (n4135) );
  buffer buf_n4136( .i (n4135), .o (n4136) );
  buffer buf_n4137( .i (n4136), .o (n4137) );
  buffer buf_n4138( .i (n4137), .o (n4138) );
  buffer buf_n4139( .i (n4138), .o (n4139) );
  buffer buf_n4140( .i (n4139), .o (n4140) );
  buffer buf_n4141( .i (n4140), .o (n4141) );
  buffer buf_n4142( .i (n4141), .o (n4142) );
  buffer buf_n4143( .i (n4142), .o (n4143) );
  buffer buf_n4144( .i (n4143), .o (n4144) );
  buffer buf_n4145( .i (n4144), .o (n4145) );
  buffer buf_n4146( .i (n4145), .o (n4146) );
  buffer buf_n4147( .i (n4146), .o (n4147) );
  buffer buf_n4148( .i (n4147), .o (n4148) );
  buffer buf_n4149( .i (n4148), .o (n4149) );
  buffer buf_n4150( .i (n4149), .o (n4150) );
  buffer buf_n4151( .i (n4150), .o (n4151) );
  buffer buf_n4152( .i (n4151), .o (n4152) );
  buffer buf_n4153( .i (n4152), .o (n4153) );
  buffer buf_n4154( .i (n4153), .o (n4154) );
  buffer buf_n4155( .i (n4154), .o (n4155) );
  buffer buf_n4156( .i (n4155), .o (n4156) );
  buffer buf_n4157( .i (n4156), .o (n4157) );
  buffer buf_n4158( .i (n4157), .o (n4158) );
  buffer buf_n4159( .i (n4158), .o (n4159) );
  assign n4165 = n3892 & ~n3913 ;
  buffer buf_n4166( .i (n4165), .o (n4166) );
  buffer buf_n4167( .i (n4166), .o (n4167) );
  buffer buf_n4168( .i (n4167), .o (n4168) );
  buffer buf_n4169( .i (n4168), .o (n4169) );
  buffer buf_n4170( .i (n4169), .o (n4170) );
  buffer buf_n4171( .i (n4170), .o (n4171) );
  buffer buf_n4172( .i (n4171), .o (n4172) );
  buffer buf_n4173( .i (n4172), .o (n4173) );
  buffer buf_n4174( .i (n4173), .o (n4174) );
  buffer buf_n4175( .i (n4174), .o (n4175) );
  buffer buf_n4176( .i (n4175), .o (n4176) );
  buffer buf_n4177( .i (n4176), .o (n4177) );
  buffer buf_n4178( .i (n4177), .o (n4178) );
  buffer buf_n4179( .i (n4178), .o (n4179) );
  buffer buf_n4180( .i (n4179), .o (n4180) );
  buffer buf_n4181( .i (n4180), .o (n4181) );
  buffer buf_n4182( .i (n4181), .o (n4182) );
  buffer buf_n4183( .i (n4182), .o (n4183) );
  buffer buf_n4184( .i (n4183), .o (n4184) );
  buffer buf_n4185( .i (n4184), .o (n4185) );
  buffer buf_n4186( .i (n4185), .o (n4186) );
  buffer buf_n4187( .i (n4186), .o (n4187) );
  buffer buf_n4188( .i (n4187), .o (n4188) );
  buffer buf_n4189( .i (n4188), .o (n4189) );
  buffer buf_n4190( .i (n4189), .o (n4190) );
  buffer buf_n4191( .i (n4190), .o (n4191) );
  buffer buf_n4192( .i (n4191), .o (n4192) );
  buffer buf_n4193( .i (n4192), .o (n4193) );
  buffer buf_n4194( .i (n4193), .o (n4194) );
  buffer buf_n4195( .i (n4194), .o (n4195) );
  buffer buf_n4196( .i (n4195), .o (n4196) );
  buffer buf_n4197( .i (n4196), .o (n4197) );
  buffer buf_n4198( .i (n4197), .o (n4198) );
  buffer buf_n4199( .i (n4198), .o (n4199) );
  buffer buf_n4200( .i (n4199), .o (n4200) );
  buffer buf_n4201( .i (n4200), .o (n4201) );
  assign n4208 = n4159 & n4201 ;
  buffer buf_n4209( .i (n4208), .o (n4209) );
  assign n4211 = ~n4111 & n4209 ;
  assign n4212 = n3953 & ~n4211 ;
  buffer buf_n4210( .i (n4209), .o (n4210) );
  buffer buf_n1918( .i (N303), .o (n1918) );
  buffer buf_n1919( .i (n1918), .o (n1919) );
  buffer buf_n1920( .i (n1919), .o (n1920) );
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n3884( .i (n3883), .o (n3884) );
  buffer buf_n489( .i (N153), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n590( .i (n589), .o (n590) );
  assign n4213 = ~n493 & n590 ;
  buffer buf_n4214( .i (n4213), .o (n4214) );
  assign n4217 = n3884 | n4214 ;
  buffer buf_n4218( .i (n4217), .o (n4218) );
  assign n4219 = n1926 & n4218 ;
  buffer buf_n4220( .i (n4219), .o (n4220) );
  buffer buf_n4221( .i (n4220), .o (n4221) );
  buffer buf_n4222( .i (n4221), .o (n4222) );
  buffer buf_n4223( .i (n4222), .o (n4223) );
  buffer buf_n4224( .i (n4223), .o (n4224) );
  buffer buf_n4225( .i (n4224), .o (n4225) );
  buffer buf_n4226( .i (n4225), .o (n4226) );
  buffer buf_n4227( .i (n4226), .o (n4227) );
  buffer buf_n4228( .i (n4227), .o (n4228) );
  buffer buf_n4229( .i (n4228), .o (n4229) );
  buffer buf_n4230( .i (n4229), .o (n4230) );
  buffer buf_n4231( .i (n4230), .o (n4231) );
  buffer buf_n4232( .i (n4231), .o (n4232) );
  buffer buf_n4233( .i (n4232), .o (n4233) );
  buffer buf_n4234( .i (n4233), .o (n4234) );
  buffer buf_n4235( .i (n4234), .o (n4235) );
  buffer buf_n4236( .i (n4235), .o (n4236) );
  buffer buf_n4237( .i (n4236), .o (n4237) );
  buffer buf_n4238( .i (n4237), .o (n4238) );
  buffer buf_n4239( .i (n4238), .o (n4239) );
  buffer buf_n4240( .i (n4239), .o (n4240) );
  buffer buf_n4241( .i (n4240), .o (n4241) );
  buffer buf_n4242( .i (n4241), .o (n4242) );
  buffer buf_n4243( .i (n4242), .o (n4243) );
  buffer buf_n4244( .i (n4243), .o (n4244) );
  buffer buf_n4245( .i (n4244), .o (n4245) );
  buffer buf_n4246( .i (n4245), .o (n4246) );
  buffer buf_n4247( .i (n4246), .o (n4247) );
  buffer buf_n4248( .i (n4247), .o (n4248) );
  buffer buf_n4249( .i (n4248), .o (n4249) );
  buffer buf_n4250( .i (n4249), .o (n4250) );
  buffer buf_n4251( .i (n4250), .o (n4251) );
  buffer buf_n4252( .i (n4251), .o (n4252) );
  buffer buf_n4253( .i (n4252), .o (n4253) );
  buffer buf_n4254( .i (n4253), .o (n4254) );
  buffer buf_n4255( .i (n4254), .o (n4255) );
  assign n4256 = n1926 | n4218 ;
  buffer buf_n4257( .i (n4256), .o (n4257) );
  buffer buf_n4258( .i (n4257), .o (n4258) );
  buffer buf_n4259( .i (n4258), .o (n4259) );
  buffer buf_n4260( .i (n4259), .o (n4260) );
  buffer buf_n4261( .i (n4260), .o (n4261) );
  buffer buf_n4262( .i (n4261), .o (n4262) );
  buffer buf_n4263( .i (n4262), .o (n4263) );
  buffer buf_n4264( .i (n4263), .o (n4264) );
  buffer buf_n4265( .i (n4264), .o (n4265) );
  buffer buf_n4266( .i (n4265), .o (n4266) );
  buffer buf_n4267( .i (n4266), .o (n4267) );
  buffer buf_n4268( .i (n4267), .o (n4268) );
  buffer buf_n4269( .i (n4268), .o (n4269) );
  buffer buf_n4270( .i (n4269), .o (n4270) );
  buffer buf_n4271( .i (n4270), .o (n4271) );
  buffer buf_n4272( .i (n4271), .o (n4272) );
  buffer buf_n4273( .i (n4272), .o (n4273) );
  buffer buf_n4274( .i (n4273), .o (n4274) );
  buffer buf_n4275( .i (n4274), .o (n4275) );
  buffer buf_n4276( .i (n4275), .o (n4276) );
  buffer buf_n4277( .i (n4276), .o (n4277) );
  buffer buf_n4278( .i (n4277), .o (n4278) );
  buffer buf_n4279( .i (n4278), .o (n4279) );
  buffer buf_n4280( .i (n4279), .o (n4280) );
  buffer buf_n4281( .i (n4280), .o (n4281) );
  buffer buf_n4282( .i (n4281), .o (n4282) );
  buffer buf_n4283( .i (n4282), .o (n4283) );
  buffer buf_n4284( .i (n4283), .o (n4284) );
  buffer buf_n4285( .i (n4284), .o (n4285) );
  buffer buf_n4286( .i (n4285), .o (n4286) );
  buffer buf_n4287( .i (n4286), .o (n4287) );
  buffer buf_n4288( .i (n4287), .o (n4288) );
  buffer buf_n4289( .i (n4288), .o (n4289) );
  buffer buf_n4290( .i (n4289), .o (n4290) );
  buffer buf_n4291( .i (n4290), .o (n4291) );
  buffer buf_n1852( .i (N299), .o (n1852) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n494( .i (N154), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  assign n4292 = ~n498 & n590 ;
  buffer buf_n4293( .i (n4292), .o (n4293) );
  assign n4296 = n3884 | n4293 ;
  buffer buf_n4297( .i (n4296), .o (n4297) );
  assign n4298 = n1860 & n4297 ;
  buffer buf_n4299( .i (n4298), .o (n4299) );
  buffer buf_n4300( .i (n4299), .o (n4300) );
  buffer buf_n4301( .i (n4300), .o (n4301) );
  buffer buf_n4302( .i (n4301), .o (n4302) );
  buffer buf_n4303( .i (n4302), .o (n4303) );
  buffer buf_n4304( .i (n4303), .o (n4304) );
  assign n4305 = n1860 | n4297 ;
  buffer buf_n4306( .i (n4305), .o (n4306) );
  buffer buf_n4307( .i (n4306), .o (n4307) );
  buffer buf_n4308( .i (n4307), .o (n4308) );
  buffer buf_n4309( .i (n4308), .o (n4309) );
  buffer buf_n1786( .i (N296), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n499( .i (N155), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n4310( .i (n588), .o (n4310) );
  assign n4311 = ~n502 & n4310 ;
  buffer buf_n4312( .i (n4311), .o (n4312) );
  assign n4315 = n3977 | n4312 ;
  buffer buf_n4316( .i (n4315), .o (n4316) );
  assign n4317 = n1793 & n4316 ;
  buffer buf_n4318( .i (n4317), .o (n4318) );
  buffer buf_n4319( .i (n4318), .o (n4319) );
  buffer buf_n4320( .i (n4319), .o (n4320) );
  assign n4321 = n1793 | n4316 ;
  buffer buf_n4322( .i (n4321), .o (n4322) );
  buffer buf_n1720( .i (N293), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n503( .i (N156), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  assign n4326 = ~n506 & n4310 ;
  buffer buf_n4327( .i (n4326), .o (n4327) );
  assign n4330 = n3977 | n4327 ;
  buffer buf_n4331( .i (n4330), .o (n4331) );
  assign n4332 = n1727 | n4331 ;
  buffer buf_n4333( .i (n4332), .o (n4333) );
  assign n4367 = n4322 & n4333 ;
  buffer buf_n4368( .i (n4367), .o (n4368) );
  assign n4370 = n4320 | n4368 ;
  buffer buf_n4371( .i (n4370), .o (n4371) );
  assign n4401 = n4309 & n4371 ;
  buffer buf_n4402( .i (n4401), .o (n4402) );
  assign n4403 = n4304 | n4402 ;
  buffer buf_n4404( .i (n4403), .o (n4404) );
  buffer buf_n4369( .i (n4368), .o (n4369) );
  assign n4429 = n1727 & n4331 ;
  buffer buf_n4430( .i (n4429), .o (n4430) );
  buffer buf_n4431( .i (n4430), .o (n4431) );
  assign n4463 = n4319 | n4431 ;
  buffer buf_n4464( .i (n4463), .o (n4464) );
  assign n4465 = n4369 & ~n4464 ;
  buffer buf_n4466( .i (n4465), .o (n4466) );
  assign n4494 = ~n4299 & n4306 ;
  buffer buf_n4495( .i (n4494), .o (n4495) );
  buffer buf_n4496( .i (n4495), .o (n4496) );
  buffer buf_n4497( .i (n4496), .o (n4497) );
  assign n4528 = n4466 & n4497 ;
  buffer buf_n4529( .i (n4528), .o (n4529) );
  buffer buf_n4530( .i (n4529), .o (n4530) );
  assign n4531 = n4404 & ~n4530 ;
  buffer buf_n4532( .i (n4531), .o (n4532) );
  buffer buf_n4533( .i (n4532), .o (n4533) );
  buffer buf_n4534( .i (n4533), .o (n4534) );
  buffer buf_n4535( .i (n4534), .o (n4535) );
  buffer buf_n4536( .i (n4535), .o (n4536) );
  buffer buf_n4537( .i (n4536), .o (n4537) );
  buffer buf_n4538( .i (n4537), .o (n4538) );
  buffer buf_n4539( .i (n4538), .o (n4539) );
  buffer buf_n4540( .i (n4539), .o (n4540) );
  buffer buf_n4541( .i (n4540), .o (n4541) );
  buffer buf_n4542( .i (n4541), .o (n4542) );
  buffer buf_n4543( .i (n4542), .o (n4543) );
  buffer buf_n4544( .i (n4543), .o (n4544) );
  buffer buf_n4545( .i (n4544), .o (n4545) );
  buffer buf_n4546( .i (n4545), .o (n4546) );
  buffer buf_n4547( .i (n4546), .o (n4547) );
  buffer buf_n4548( .i (n4547), .o (n4548) );
  buffer buf_n4549( .i (n4548), .o (n4549) );
  buffer buf_n4550( .i (n4549), .o (n4550) );
  buffer buf_n4551( .i (n4550), .o (n4551) );
  buffer buf_n4552( .i (n4551), .o (n4552) );
  buffer buf_n4553( .i (n4552), .o (n4553) );
  buffer buf_n4554( .i (n4553), .o (n4554) );
  buffer buf_n4555( .i (n4554), .o (n4555) );
  buffer buf_n4405( .i (n4404), .o (n4405) );
  buffer buf_n4406( .i (n4405), .o (n4406) );
  buffer buf_n4407( .i (n4406), .o (n4407) );
  buffer buf_n4408( .i (n4407), .o (n4408) );
  buffer buf_n4409( .i (n4408), .o (n4409) );
  buffer buf_n4410( .i (n4409), .o (n4410) );
  buffer buf_n4411( .i (n4410), .o (n4411) );
  buffer buf_n4412( .i (n4411), .o (n4412) );
  buffer buf_n4413( .i (n4412), .o (n4413) );
  buffer buf_n4414( .i (n4413), .o (n4414) );
  buffer buf_n4415( .i (n4414), .o (n4415) );
  buffer buf_n4416( .i (n4415), .o (n4416) );
  buffer buf_n4417( .i (n4416), .o (n4417) );
  buffer buf_n4418( .i (n4417), .o (n4418) );
  buffer buf_n4419( .i (n4418), .o (n4419) );
  buffer buf_n4420( .i (n4419), .o (n4420) );
  buffer buf_n4421( .i (n4420), .o (n4421) );
  buffer buf_n4422( .i (n4421), .o (n4422) );
  buffer buf_n4423( .i (n4422), .o (n4423) );
  buffer buf_n4424( .i (n4423), .o (n4424) );
  buffer buf_n4425( .i (n4424), .o (n4425) );
  buffer buf_n4426( .i (n4425), .o (n4426) );
  buffer buf_n4427( .i (n4426), .o (n4427) );
  buffer buf_n4428( .i (n4427), .o (n4428) );
  buffer buf_n1650( .i (N289), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  buffer buf_n507( .i (N157), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  assign n4556 = ~n511 & n590 ;
  buffer buf_n4557( .i (n3882), .o (n4557) );
  assign n4558 = n4556 | n4557 ;
  buffer buf_n4559( .i (n4558), .o (n4559) );
  assign n4560 = n1657 & n4559 ;
  buffer buf_n4561( .i (n4560), .o (n4561) );
  buffer buf_n4562( .i (n4561), .o (n4562) );
  buffer buf_n4563( .i (n4562), .o (n4563) );
  buffer buf_n4564( .i (n4563), .o (n4564) );
  buffer buf_n4565( .i (n4564), .o (n4565) );
  buffer buf_n4566( .i (n4565), .o (n4566) );
  buffer buf_n4567( .i (n4566), .o (n4567) );
  buffer buf_n4568( .i (n4567), .o (n4568) );
  buffer buf_n4569( .i (n4568), .o (n4569) );
  buffer buf_n4570( .i (n4569), .o (n4570) );
  buffer buf_n4571( .i (n4570), .o (n4571) );
  buffer buf_n4572( .i (n4571), .o (n4572) );
  buffer buf_n4573( .i (n4572), .o (n4573) );
  buffer buf_n4574( .i (n4573), .o (n4574) );
  buffer buf_n4575( .i (n4574), .o (n4575) );
  assign n4576 = n1657 | n4559 ;
  buffer buf_n4577( .i (n4576), .o (n4577) );
  buffer buf_n4578( .i (n4577), .o (n4578) );
  buffer buf_n4579( .i (n4578), .o (n4579) );
  buffer buf_n4580( .i (n4579), .o (n4580) );
  buffer buf_n4581( .i (n4580), .o (n4581) );
  buffer buf_n4582( .i (n4581), .o (n4582) );
  buffer buf_n4583( .i (n4582), .o (n4583) );
  buffer buf_n4584( .i (n4583), .o (n4584) );
  buffer buf_n4585( .i (n4584), .o (n4585) );
  buffer buf_n4586( .i (n4585), .o (n4586) );
  buffer buf_n4587( .i (n4586), .o (n4587) );
  buffer buf_n4588( .i (n4587), .o (n4588) );
  buffer buf_n1584( .i (N286), .o (n1584) );
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n399( .i (N135), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  assign n4589 = n402 & ~n4310 ;
  buffer buf_n4590( .i (n4589), .o (n4590) );
  buffer buf_n512( .i (N158), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  assign n4591 = n515 & n4310 ;
  buffer buf_n4592( .i (n4591), .o (n4592) );
  assign n4593 = n4590 | n4592 ;
  buffer buf_n4594( .i (n4593), .o (n4594) );
  assign n4595 = n1591 & ~n4594 ;
  buffer buf_n4596( .i (n4595), .o (n4596) );
  buffer buf_n4597( .i (n4596), .o (n4597) );
  buffer buf_n4598( .i (n4597), .o (n4598) );
  buffer buf_n4599( .i (n4598), .o (n4599) );
  buffer buf_n4600( .i (n4599), .o (n4600) );
  buffer buf_n4601( .i (n4600), .o (n4601) );
  buffer buf_n4602( .i (n4601), .o (n4602) );
  buffer buf_n4603( .i (n4602), .o (n4603) );
  buffer buf_n4604( .i (n4603), .o (n4604) );
  buffer buf_n4605( .i (n4604), .o (n4605) );
  assign n4606 = ~n1591 & n4594 ;
  buffer buf_n4607( .i (n4606), .o (n4607) );
  buffer buf_n4608( .i (n4607), .o (n4608) );
  buffer buf_n4609( .i (n4608), .o (n4609) );
  buffer buf_n4610( .i (n4609), .o (n4610) );
  buffer buf_n4611( .i (n4610), .o (n4611) );
  buffer buf_n4612( .i (n4611), .o (n4612) );
  buffer buf_n4613( .i (n4612), .o (n4613) );
  buffer buf_n4614( .i (n4613), .o (n4614) );
  buffer buf_n4615( .i (n4614), .o (n4615) );
  buffer buf_n1518( .i (N283), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n1522( .i (n1521), .o (n1522) );
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n411( .i (N144), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n4616( .i (n588), .o (n4616) );
  assign n4617 = n414 & ~n4616 ;
  buffer buf_n4618( .i (n4617), .o (n4618) );
  buffer buf_n516( .i (N159), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  assign n4619 = n519 & n4616 ;
  buffer buf_n4620( .i (n4619), .o (n4620) );
  assign n4621 = n4618 | n4620 ;
  buffer buf_n4622( .i (n4621), .o (n4622) );
  assign n4623 = ~n1525 & n4622 ;
  buffer buf_n4624( .i (n4623), .o (n4624) );
  buffer buf_n4625( .i (n4624), .o (n4625) );
  buffer buf_n4626( .i (n4625), .o (n4626) );
  buffer buf_n4627( .i (n4626), .o (n4627) );
  buffer buf_n4628( .i (n4627), .o (n4628) );
  buffer buf_n4629( .i (n4628), .o (n4629) );
  assign n4630 = n1525 & ~n4622 ;
  buffer buf_n4631( .i (n4630), .o (n4631) );
  buffer buf_n4632( .i (n4631), .o (n4632) );
  buffer buf_n4633( .i (n4632), .o (n4633) );
  buffer buf_n4634( .i (n4633), .o (n4634) );
  buffer buf_n4635( .i (n4634), .o (n4635) );
  buffer buf_n1452( .i (N280), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  buffer buf_n1455( .i (n1454), .o (n1455) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n403( .i (N138), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  assign n4636 = n406 & ~n4616 ;
  buffer buf_n4637( .i (n4636), .o (n4637) );
  buffer buf_n520( .i (N160), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  assign n4638 = n523 & n4616 ;
  buffer buf_n4639( .i (n4638), .o (n4639) );
  assign n4640 = n4637 | n4639 ;
  buffer buf_n4641( .i (n4640), .o (n4641) );
  assign n4642 = ~n1459 & n4641 ;
  buffer buf_n4643( .i (n4642), .o (n4643) );
  buffer buf_n4644( .i (n4643), .o (n4644) );
  buffer buf_n4645( .i (n4644), .o (n4645) );
  buffer buf_n1386( .i (N277), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n415( .i (N147), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n4646( .i (n587), .o (n4646) );
  buffer buf_n4647( .i (n4646), .o (n4647) );
  assign n4648 = n418 & ~n4647 ;
  buffer buf_n4649( .i (n4648), .o (n4649) );
  buffer buf_n485( .i (N151), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  assign n4650 = n488 & n4647 ;
  buffer buf_n4651( .i (n4650), .o (n4651) );
  assign n4652 = n4649 | n4651 ;
  buffer buf_n4653( .i (n4652), .o (n4653) );
  assign n4654 = ~n1393 & n4653 ;
  buffer buf_n4655( .i (n4654), .o (n4655) );
  assign n4691 = n1459 & ~n4641 ;
  buffer buf_n4692( .i (n4691), .o (n4692) );
  assign n4693 = n4655 & ~n4692 ;
  buffer buf_n4694( .i (n4693), .o (n4694) );
  assign n4695 = n4645 | n4694 ;
  buffer buf_n4696( .i (n4695), .o (n4696) );
  assign n4723 = ~n4635 & n4696 ;
  assign n4724 = n4629 | n4723 ;
  buffer buf_n4725( .i (n4724), .o (n4725) );
  buffer buf_n4726( .i (n4725), .o (n4726) );
  assign n4750 = n4615 | n4726 ;
  assign n4751 = ~n4605 & n4750 ;
  buffer buf_n4752( .i (n4751), .o (n4752) );
  assign n4774 = n4588 & ~n4752 ;
  buffer buf_n4775( .i (n4774), .o (n4775) );
  assign n4792 = n1393 & ~n4653 ;
  buffer buf_n4793( .i (n4792), .o (n4793) );
  assign n4794 = n4655 | n4793 ;
  buffer buf_n4795( .i (n4794), .o (n4795) );
  assign n4827 = n4643 | n4692 ;
  buffer buf_n4828( .i (n4827), .o (n4828) );
  assign n4864 = n4795 | n4828 ;
  buffer buf_n4865( .i (n4864), .o (n4865) );
  buffer buf_n4866( .i (n4865), .o (n4866) );
  buffer buf_n4867( .i (n4866), .o (n4867) );
  buffer buf_n4868( .i (n4867), .o (n4868) );
  buffer buf_n4869( .i (n4868), .o (n4869) );
  buffer buf_n4870( .i (n4869), .o (n4870) );
  buffer buf_n4871( .i (n4870), .o (n4871) );
  buffer buf_n4872( .i (n4871), .o (n4872) );
  assign n4891 = n4596 | n4607 ;
  buffer buf_n4892( .i (n4891), .o (n4892) );
  buffer buf_n4893( .i (n4892), .o (n4893) );
  buffer buf_n4894( .i (n4893), .o (n4894) );
  buffer buf_n4895( .i (n4894), .o (n4895) );
  buffer buf_n4896( .i (n4895), .o (n4896) );
  buffer buf_n4897( .i (n4896), .o (n4897) );
  buffer buf_n4898( .i (n4897), .o (n4898) );
  buffer buf_n4899( .i (n4898), .o (n4899) );
  assign n4924 = n4624 | n4631 ;
  buffer buf_n4925( .i (n4924), .o (n4925) );
  buffer buf_n4926( .i (n4925), .o (n4926) );
  buffer buf_n4927( .i (n4926), .o (n4927) );
  buffer buf_n4928( .i (n4927), .o (n4928) );
  buffer buf_n4929( .i (n4928), .o (n4929) );
  buffer buf_n4930( .i (n4929), .o (n4930) );
  buffer buf_n4931( .i (n4930), .o (n4931) );
  buffer buf_n4932( .i (n4931), .o (n4932) );
  assign n4956 = n4899 | n4932 ;
  buffer buf_n4957( .i (n4956), .o (n4957) );
  assign n4958 = n4872 | n4957 ;
  buffer buf_n4959( .i (n4958), .o (n4959) );
  assign n4961 = n4775 & n4959 ;
  assign n4962 = n4575 | n4961 ;
  buffer buf_n4963( .i (n4962), .o (n4963) );
  buffer buf_n4964( .i (n4963), .o (n4964) );
  buffer buf_n4965( .i (n4964), .o (n4965) );
  buffer buf_n4966( .i (n4965), .o (n4966) );
  buffer buf_n4967( .i (n4966), .o (n4967) );
  buffer buf_n4968( .i (n4967), .o (n4968) );
  buffer buf_n4969( .i (n4968), .o (n4969) );
  buffer buf_n4970( .i (n4969), .o (n4970) );
  buffer buf_n4971( .i (n4970), .o (n4971) );
  buffer buf_n4972( .i (n4971), .o (n4972) );
  buffer buf_n4973( .i (n4972), .o (n4973) );
  buffer buf_n4974( .i (n4973), .o (n4974) );
  buffer buf_n4975( .i (n4974), .o (n4975) );
  buffer buf_n4976( .i (n4975), .o (n4976) );
  buffer buf_n4977( .i (n4976), .o (n4977) );
  buffer buf_n4776( .i (n4775), .o (n4776) );
  buffer buf_n4777( .i (n4776), .o (n4777) );
  buffer buf_n4778( .i (n4777), .o (n4778) );
  buffer buf_n4779( .i (n4778), .o (n4779) );
  buffer buf_n4780( .i (n4779), .o (n4780) );
  buffer buf_n4781( .i (n4780), .o (n4781) );
  buffer buf_n4782( .i (n4781), .o (n4782) );
  buffer buf_n4783( .i (n4782), .o (n4783) );
  buffer buf_n4784( .i (n4783), .o (n4784) );
  buffer buf_n4785( .i (n4784), .o (n4785) );
  buffer buf_n4786( .i (n4785), .o (n4786) );
  buffer buf_n4787( .i (n4786), .o (n4787) );
  buffer buf_n4788( .i (n4787), .o (n4788) );
  buffer buf_n4789( .i (n4788), .o (n4789) );
  buffer buf_n4790( .i (n4789), .o (n4790) );
  buffer buf_n4791( .i (n4790), .o (n4791) );
  buffer buf_n3246( .i (N364), .o (n3246) );
  buffer buf_n3247( .i (n3246), .o (n3247) );
  buffer buf_n3248( .i (n3247), .o (n3248) );
  buffer buf_n3249( .i (n3248), .o (n3249) );
  buffer buf_n3250( .i (n3249), .o (n3250) );
  buffer buf_n3251( .i (n3250), .o (n3251) );
  buffer buf_n3252( .i (n3251), .o (n3252) );
  buffer buf_n3253( .i (n3252), .o (n3253) );
  buffer buf_n705( .i (N219), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  assign n4978 = n708 & n4647 ;
  buffer buf_n4979( .i (n4978), .o (n4979) );
  buffer buf_n3514( .i (N66), .o (n3514) );
  buffer buf_n3515( .i (n3514), .o (n3515) );
  buffer buf_n3516( .i (n3515), .o (n3516) );
  buffer buf_n3517( .i (n3516), .o (n3517) );
  assign n4980 = n3517 & ~n4647 ;
  buffer buf_n4981( .i (n4980), .o (n4981) );
  assign n4982 = n4979 | n4981 ;
  buffer buf_n4983( .i (n4982), .o (n4983) );
  assign n4984 = ~n3253 & n4983 ;
  buffer buf_n4985( .i (n4984), .o (n4985) );
  buffer buf_n4986( .i (n4985), .o (n4986) );
  buffer buf_n4987( .i (n4986), .o (n4987) );
  buffer buf_n4988( .i (n4987), .o (n4988) );
  buffer buf_n4989( .i (n4988), .o (n4989) );
  buffer buf_n4990( .i (n4989), .o (n4990) );
  buffer buf_n4991( .i (n4990), .o (n4991) );
  buffer buf_n4992( .i (n4991), .o (n4992) );
  buffer buf_n4993( .i (n4992), .o (n4993) );
  buffer buf_n4994( .i (n4993), .o (n4994) );
  buffer buf_n4995( .i (n4994), .o (n4995) );
  buffer buf_n4996( .i (n4995), .o (n4996) );
  buffer buf_n4997( .i (n4996), .o (n4997) );
  buffer buf_n4998( .i (n4997), .o (n4998) );
  buffer buf_n4999( .i (n4998), .o (n4999) );
  buffer buf_n5000( .i (n4999), .o (n5000) );
  buffer buf_n5001( .i (n5000), .o (n5001) );
  buffer buf_n5002( .i (n5001), .o (n5002) );
  buffer buf_n5003( .i (n5002), .o (n5003) );
  buffer buf_n5004( .i (n5003), .o (n5004) );
  buffer buf_n5005( .i (n5004), .o (n5005) );
  buffer buf_n5006( .i (n5005), .o (n5006) );
  buffer buf_n5007( .i (n5006), .o (n5007) );
  buffer buf_n5008( .i (n5007), .o (n5008) );
  buffer buf_n5009( .i (n5008), .o (n5009) );
  buffer buf_n5010( .i (n5009), .o (n5010) );
  buffer buf_n5011( .i (n5010), .o (n5011) );
  buffer buf_n5012( .i (n5011), .o (n5012) );
  assign n5013 = n3253 & ~n4983 ;
  buffer buf_n5014( .i (n5013), .o (n5014) );
  buffer buf_n5015( .i (n5014), .o (n5015) );
  buffer buf_n5016( .i (n5015), .o (n5016) );
  buffer buf_n5017( .i (n5016), .o (n5017) );
  buffer buf_n5018( .i (n5017), .o (n5018) );
  buffer buf_n5019( .i (n5018), .o (n5019) );
  buffer buf_n5020( .i (n5019), .o (n5020) );
  buffer buf_n5021( .i (n5020), .o (n5021) );
  buffer buf_n5022( .i (n5021), .o (n5022) );
  buffer buf_n5023( .i (n5022), .o (n5023) );
  buffer buf_n5024( .i (n5023), .o (n5024) );
  buffer buf_n5025( .i (n5024), .o (n5025) );
  buffer buf_n5026( .i (n5025), .o (n5026) );
  buffer buf_n5027( .i (n5026), .o (n5027) );
  buffer buf_n5028( .i (n5027), .o (n5028) );
  buffer buf_n5029( .i (n5028), .o (n5029) );
  buffer buf_n5030( .i (n5029), .o (n5030) );
  buffer buf_n5031( .i (n5030), .o (n5031) );
  buffer buf_n5032( .i (n5031), .o (n5032) );
  buffer buf_n5033( .i (n5032), .o (n5033) );
  buffer buf_n5034( .i (n5033), .o (n5034) );
  buffer buf_n5035( .i (n5034), .o (n5035) );
  buffer buf_n5036( .i (n5035), .o (n5036) );
  buffer buf_n5037( .i (n5036), .o (n5037) );
  buffer buf_n5038( .i (n5037), .o (n5038) );
  buffer buf_n5039( .i (n5038), .o (n5039) );
  buffer buf_n5040( .i (n5039), .o (n5040) );
  buffer buf_n3180( .i (N361), .o (n3180) );
  buffer buf_n3181( .i (n3180), .o (n3181) );
  buffer buf_n3182( .i (n3181), .o (n3182) );
  buffer buf_n3183( .i (n3182), .o (n3183) );
  buffer buf_n3184( .i (n3183), .o (n3184) );
  buffer buf_n3185( .i (n3184), .o (n3185) );
  buffer buf_n3186( .i (n3185), .o (n3186) );
  buffer buf_n3187( .i (n3186), .o (n3187) );
  buffer buf_n709( .i (N220), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n5041( .i (n4646), .o (n5041) );
  assign n5042 = n712 & n5041 ;
  buffer buf_n5043( .i (n5042), .o (n5043) );
  buffer buf_n3460( .i (N50), .o (n3460) );
  buffer buf_n3461( .i (n3460), .o (n3461) );
  buffer buf_n3462( .i (n3461), .o (n3462) );
  buffer buf_n3463( .i (n3462), .o (n3463) );
  assign n5044 = n3463 & ~n5041 ;
  buffer buf_n5045( .i (n5044), .o (n5045) );
  assign n5046 = n5043 | n5045 ;
  buffer buf_n5047( .i (n5046), .o (n5047) );
  assign n5048 = n3187 & ~n5047 ;
  buffer buf_n5049( .i (n5048), .o (n5049) );
  buffer buf_n5050( .i (n5049), .o (n5050) );
  buffer buf_n5051( .i (n5050), .o (n5051) );
  buffer buf_n5052( .i (n5051), .o (n5052) );
  buffer buf_n5053( .i (n5052), .o (n5053) );
  buffer buf_n5054( .i (n5053), .o (n5054) );
  assign n5056 = ~n3187 & n5047 ;
  buffer buf_n5057( .i (n5056), .o (n5057) );
  buffer buf_n5058( .i (n5057), .o (n5058) );
  buffer buf_n5059( .i (n5058), .o (n5059) );
  buffer buf_n5060( .i (n5059), .o (n5060) );
  buffer buf_n5061( .i (n5060), .o (n5061) );
  buffer buf_n3114( .i (N358), .o (n3114) );
  buffer buf_n3115( .i (n3114), .o (n3115) );
  buffer buf_n3116( .i (n3115), .o (n3116) );
  buffer buf_n3117( .i (n3116), .o (n3117) );
  buffer buf_n3118( .i (n3117), .o (n3118) );
  buffer buf_n3119( .i (n3118), .o (n3119) );
  buffer buf_n3120( .i (n3119), .o (n3120) );
  buffer buf_n3121( .i (n3120), .o (n3121) );
  buffer buf_n713( .i (N221), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  assign n5063 = n716 & n5041 ;
  buffer buf_n5064( .i (n5063), .o (n5064) );
  buffer buf_n2314( .i (N32), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  assign n5065 = n2317 & ~n5041 ;
  buffer buf_n5066( .i (n5065), .o (n5066) );
  assign n5067 = n5064 | n5066 ;
  buffer buf_n5068( .i (n5067), .o (n5068) );
  assign n5069 = n3121 & ~n5068 ;
  buffer buf_n5070( .i (n5069), .o (n5070) );
  buffer buf_n5071( .i (n5070), .o (n5071) );
  buffer buf_n5072( .i (n5071), .o (n5072) );
  assign n5073 = ~n3121 & n5068 ;
  buffer buf_n5074( .i (n5073), .o (n5074) );
  buffer buf_n3048( .i (N355), .o (n3048) );
  buffer buf_n3049( .i (n3048), .o (n3049) );
  buffer buf_n3050( .i (n3049), .o (n3050) );
  buffer buf_n3051( .i (n3050), .o (n3051) );
  buffer buf_n3052( .i (n3051), .o (n3052) );
  buffer buf_n3053( .i (n3052), .o (n3053) );
  buffer buf_n3054( .i (n3053), .o (n3054) );
  buffer buf_n3055( .i (n3054), .o (n3055) );
  buffer buf_n717( .i (N222), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n5076( .i (n4646), .o (n5076) );
  assign n5077 = n720 & n5076 ;
  buffer buf_n5078( .i (n5077), .o (n5078) );
  buffer buf_n2978( .i (N35), .o (n2978) );
  buffer buf_n2979( .i (n2978), .o (n2979) );
  buffer buf_n2980( .i (n2979), .o (n2980) );
  buffer buf_n2981( .i (n2980), .o (n2981) );
  assign n5079 = n2981 & ~n5076 ;
  buffer buf_n5080( .i (n5079), .o (n5080) );
  assign n5081 = n5078 | n5080 ;
  buffer buf_n5082( .i (n5081), .o (n5082) );
  assign n5083 = ~n3055 & n5082 ;
  buffer buf_n5084( .i (n5083), .o (n5084) );
  assign n5108 = n5074 | n5084 ;
  buffer buf_n5109( .i (n5108), .o (n5109) );
  assign n5110 = ~n5072 & n5109 ;
  buffer buf_n5111( .i (n5110), .o (n5111) );
  assign n5132 = n5061 | n5111 ;
  assign n5133 = ~n5054 & n5132 ;
  buffer buf_n5134( .i (n5133), .o (n5134) );
  buffer buf_n5055( .i (n5054), .o (n5055) );
  assign n5151 = n5070 | n5074 ;
  buffer buf_n5152( .i (n5151), .o (n5152) );
  buffer buf_n5153( .i (n5152), .o (n5153) );
  buffer buf_n5154( .i (n5153), .o (n5154) );
  buffer buf_n5085( .i (n5084), .o (n5085) );
  buffer buf_n5086( .i (n5085), .o (n5086) );
  assign n5177 = n3055 & ~n5082 ;
  buffer buf_n5178( .i (n5177), .o (n5178) );
  buffer buf_n5179( .i (n5178), .o (n5179) );
  buffer buf_n5180( .i (n5179), .o (n5180) );
  assign n5203 = n5086 | n5180 ;
  buffer buf_n5204( .i (n5203), .o (n5204) );
  assign n5227 = n5154 | n5204 ;
  buffer buf_n5228( .i (n5227), .o (n5228) );
  assign n5246 = n5055 | n5228 ;
  assign n5247 = ~n5134 & n5246 ;
  buffer buf_n5248( .i (n5247), .o (n5248) );
  buffer buf_n5249( .i (n5248), .o (n5249) );
  buffer buf_n5250( .i (n5249), .o (n5250) );
  buffer buf_n5251( .i (n5250), .o (n5251) );
  buffer buf_n5252( .i (n5251), .o (n5252) );
  buffer buf_n5253( .i (n5252), .o (n5253) );
  buffer buf_n5254( .i (n5253), .o (n5254) );
  buffer buf_n5255( .i (n5254), .o (n5255) );
  buffer buf_n5256( .i (n5255), .o (n5256) );
  buffer buf_n5257( .i (n5256), .o (n5257) );
  buffer buf_n5258( .i (n5257), .o (n5258) );
  buffer buf_n5259( .i (n5258), .o (n5259) );
  buffer buf_n5260( .i (n5259), .o (n5260) );
  buffer buf_n5261( .i (n5260), .o (n5261) );
  buffer buf_n5262( .i (n5261), .o (n5262) );
  buffer buf_n5263( .i (n5262), .o (n5263) );
  buffer buf_n5135( .i (n5134), .o (n5135) );
  buffer buf_n5136( .i (n5135), .o (n5136) );
  buffer buf_n5137( .i (n5136), .o (n5137) );
  buffer buf_n5138( .i (n5137), .o (n5138) );
  buffer buf_n5139( .i (n5138), .o (n5139) );
  buffer buf_n5140( .i (n5139), .o (n5140) );
  buffer buf_n5141( .i (n5140), .o (n5141) );
  buffer buf_n5142( .i (n5141), .o (n5142) );
  buffer buf_n5143( .i (n5142), .o (n5143) );
  buffer buf_n5144( .i (n5143), .o (n5144) );
  buffer buf_n5145( .i (n5144), .o (n5145) );
  buffer buf_n5146( .i (n5145), .o (n5146) );
  buffer buf_n5147( .i (n5146), .o (n5147) );
  buffer buf_n5148( .i (n5147), .o (n5148) );
  buffer buf_n5149( .i (n5148), .o (n5149) );
  buffer buf_n5150( .i (n5149), .o (n5150) );
  buffer buf_n2714( .i (N340), .o (n2714) );
  buffer buf_n2715( .i (n2714), .o (n2715) );
  buffer buf_n2716( .i (n2715), .o (n2716) );
  buffer buf_n2717( .i (n2716), .o (n2717) );
  buffer buf_n2718( .i (n2717), .o (n2718) );
  buffer buf_n2719( .i (n2718), .o (n2719) );
  buffer buf_n2720( .i (n2719), .o (n2720) );
  buffer buf_n2721( .i (n2720), .o (n2721) );
  buffer buf_n701( .i (N217), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  assign n5264 = n704 & n5076 ;
  buffer buf_n5265( .i (n5264), .o (n5265) );
  buffer buf_n376( .i (N118), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  assign n5266 = n379 & ~n5076 ;
  buffer buf_n5267( .i (n5266), .o (n5267) );
  assign n5268 = n5265 | n5267 ;
  buffer buf_n5269( .i (n5268), .o (n5269) );
  assign n5270 = ~n2721 & n5269 ;
  buffer buf_n5271( .i (n5270), .o (n5271) );
  buffer buf_n5272( .i (n5271), .o (n5272) );
  buffer buf_n5273( .i (n5272), .o (n5273) );
  buffer buf_n2780( .i (N343), .o (n2780) );
  buffer buf_n2781( .i (n2780), .o (n2781) );
  buffer buf_n2782( .i (n2781), .o (n2782) );
  buffer buf_n2783( .i (n2782), .o (n2783) );
  buffer buf_n2784( .i (n2783), .o (n2784) );
  buffer buf_n2785( .i (n2784), .o (n2785) );
  buffer buf_n2786( .i (n2785), .o (n2786) );
  buffer buf_n2787( .i (n2786), .o (n2787) );
  buffer buf_n733( .i (N226), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n5295( .i (n4646), .o (n5295) );
  assign n5296 = n736 & n5295 ;
  buffer buf_n5297( .i (n5296), .o (n5297) );
  buffer buf_n3604( .i (N97), .o (n3604) );
  buffer buf_n3605( .i (n3604), .o (n3605) );
  buffer buf_n3606( .i (n3605), .o (n3606) );
  buffer buf_n3607( .i (n3606), .o (n3607) );
  assign n5298 = n3607 & ~n5295 ;
  buffer buf_n5299( .i (n5298), .o (n5299) );
  assign n5300 = n5297 | n5299 ;
  buffer buf_n5301( .i (n5300), .o (n5301) );
  assign n5302 = n2787 & ~n5301 ;
  buffer buf_n5303( .i (n5302), .o (n5303) );
  buffer buf_n5304( .i (n5303), .o (n5304) );
  buffer buf_n5305( .i (n5304), .o (n5305) );
  assign n5306 = n5273 | n5305 ;
  buffer buf_n5307( .i (n5306), .o (n5307) );
  assign n5308 = n2721 & ~n5269 ;
  buffer buf_n5309( .i (n5308), .o (n5309) );
  assign n5329 = ~n2787 & n5301 ;
  buffer buf_n5330( .i (n5329), .o (n5330) );
  assign n5332 = n5309 | n5330 ;
  buffer buf_n5333( .i (n5332), .o (n5333) );
  buffer buf_n5334( .i (n5333), .o (n5334) );
  buffer buf_n5335( .i (n5334), .o (n5335) );
  assign n5336 = n5307 | n5335 ;
  buffer buf_n5337( .i (n5336), .o (n5337) );
  buffer buf_n2912( .i (N349), .o (n2912) );
  buffer buf_n2913( .i (n2912), .o (n2913) );
  buffer buf_n2914( .i (n2913), .o (n2914) );
  buffer buf_n2915( .i (n2914), .o (n2915) );
  buffer buf_n2916( .i (n2915), .o (n2916) );
  buffer buf_n2917( .i (n2916), .o (n2917) );
  buffer buf_n2918( .i (n2917), .o (n2918) );
  buffer buf_n2919( .i (n2918), .o (n2919) );
  buffer buf_n725( .i (N224), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  assign n5338 = n728 & n5295 ;
  buffer buf_n5339( .i (n5338), .o (n5339) );
  buffer buf_n380( .i (N121), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  assign n5340 = n383 & ~n5295 ;
  buffer buf_n5341( .i (n5340), .o (n5341) );
  assign n5342 = n5339 | n5341 ;
  buffer buf_n5343( .i (n5342), .o (n5343) );
  assign n5344 = n2919 & ~n5343 ;
  buffer buf_n5345( .i (n5344), .o (n5345) );
  assign n5354 = ~n2919 & n5343 ;
  buffer buf_n5355( .i (n5354), .o (n5355) );
  assign n5365 = n5345 | n5355 ;
  buffer buf_n5366( .i (n5365), .o (n5366) );
  buffer buf_n5367( .i (n5366), .o (n5367) );
  buffer buf_n5368( .i (n5367), .o (n5368) );
  buffer buf_n2846( .i (N346), .o (n2846) );
  buffer buf_n2847( .i (n2846), .o (n2847) );
  buffer buf_n2848( .i (n2847), .o (n2848) );
  buffer buf_n2849( .i (n2848), .o (n2849) );
  buffer buf_n2850( .i (n2849), .o (n2850) );
  buffer buf_n2851( .i (n2850), .o (n2851) );
  buffer buf_n2852( .i (n2851), .o (n2852) );
  buffer buf_n2853( .i (n2852), .o (n2853) );
  buffer buf_n729( .i (N225), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n5387( .i (n587), .o (n5387) );
  buffer buf_n5388( .i (n5387), .o (n5388) );
  assign n5389 = n732 & n5388 ;
  buffer buf_n5390( .i (n5389), .o (n5390) );
  buffer buf_n3600( .i (N94), .o (n3600) );
  buffer buf_n3601( .i (n3600), .o (n3601) );
  buffer buf_n3602( .i (n3601), .o (n3602) );
  buffer buf_n3603( .i (n3602), .o (n3603) );
  assign n5391 = n3603 & ~n5388 ;
  buffer buf_n5392( .i (n5391), .o (n5392) );
  assign n5393 = n5390 | n5392 ;
  buffer buf_n5394( .i (n5393), .o (n5394) );
  assign n5395 = n2853 & ~n5394 ;
  buffer buf_n5396( .i (n5395), .o (n5396) );
  assign n5401 = ~n2853 & n5394 ;
  buffer buf_n5402( .i (n5401), .o (n5402) );
  assign n5409 = n5396 | n5402 ;
  buffer buf_n5410( .i (n5409), .o (n5410) );
  buffer buf_n5411( .i (n5410), .o (n5411) );
  buffer buf_n5412( .i (n5411), .o (n5412) );
  assign n5435 = n5368 | n5412 ;
  buffer buf_n5436( .i (n5435), .o (n5436) );
  assign n5437 = n5337 | n5436 ;
  buffer buf_n5438( .i (n5437), .o (n5438) );
  buffer buf_n2982( .i (N352), .o (n2982) );
  buffer buf_n2983( .i (n2982), .o (n2983) );
  buffer buf_n2984( .i (n2983), .o (n2984) );
  buffer buf_n2985( .i (n2984), .o (n2985) );
  buffer buf_n2986( .i (n2985), .o (n2986) );
  buffer buf_n2987( .i (n2986), .o (n2987) );
  buffer buf_n2988( .i (n2987), .o (n2988) );
  buffer buf_n2989( .i (n2988), .o (n2989) );
  buffer buf_n721( .i (N223), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  assign n5450 = n724 & n5388 ;
  buffer buf_n5451( .i (n5450), .o (n5451) );
  buffer buf_n3455( .i (N47), .o (n3455) );
  buffer buf_n3456( .i (n3455), .o (n3456) );
  buffer buf_n3457( .i (n3456), .o (n3457) );
  buffer buf_n3458( .i (n3457), .o (n3458) );
  assign n5452 = n3458 & ~n5388 ;
  buffer buf_n5453( .i (n5452), .o (n5453) );
  assign n5454 = n5451 | n5453 ;
  buffer buf_n5455( .i (n5454), .o (n5455) );
  assign n5456 = ~n2989 & n5455 ;
  buffer buf_n5457( .i (n5456), .o (n5457) );
  assign n5470 = n2989 & ~n5455 ;
  buffer buf_n5471( .i (n5470), .o (n5471) );
  assign n5483 = n5457 | n5471 ;
  buffer buf_n5484( .i (n5483), .o (n5484) );
  buffer buf_n5485( .i (n5484), .o (n5485) );
  buffer buf_n5486( .i (n5485), .o (n5486) );
  buffer buf_n5487( .i (n5486), .o (n5487) );
  buffer buf_n5488( .i (n5487), .o (n5488) );
  buffer buf_n5489( .i (n5488), .o (n5489) );
  buffer buf_n5490( .i (n5489), .o (n5490) );
  assign n5494 = n5438 | n5490 ;
  buffer buf_n5495( .i (n5494), .o (n5495) );
  buffer buf_n5496( .i (n5495), .o (n5496) );
  buffer buf_n5497( .i (n5496), .o (n5497) );
  buffer buf_n5498( .i (n5497), .o (n5498) );
  buffer buf_n5499( .i (n5498), .o (n5499) );
  buffer buf_n5500( .i (n5499), .o (n5500) );
  buffer buf_n5501( .i (n5500), .o (n5501) );
  buffer buf_n5502( .i (n5501), .o (n5502) );
  buffer buf_n5503( .i (n5502), .o (n5503) );
  buffer buf_n5504( .i (n5503), .o (n5504) );
  buffer buf_n2582( .i (N334), .o (n2582) );
  buffer buf_n2583( .i (n2582), .o (n2583) );
  buffer buf_n2584( .i (n2583), .o (n2584) );
  buffer buf_n2585( .i (n2584), .o (n2585) );
  buffer buf_n2586( .i (n2585), .o (n2586) );
  buffer buf_n2587( .i (n2586), .o (n2587) );
  buffer buf_n2588( .i (n2587), .o (n2588) );
  buffer buf_n2589( .i (n2588), .o (n2589) );
  buffer buf_n749( .i (N231), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n5505( .i (n5387), .o (n5505) );
  assign n5506 = n752 & n5505 ;
  buffer buf_n5507( .i (n5506), .o (n5507) );
  buffer buf_n274( .i (N100), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  assign n5508 = n277 & ~n5505 ;
  buffer buf_n5509( .i (n5508), .o (n5509) );
  assign n5510 = n5507 | n5509 ;
  buffer buf_n5511( .i (n5510), .o (n5511) );
  assign n5512 = n2589 & ~n5511 ;
  buffer buf_n5513( .i (n5512), .o (n5513) );
  buffer buf_n5514( .i (n5513), .o (n5514) );
  buffer buf_n5515( .i (n5514), .o (n5515) );
  buffer buf_n5516( .i (n5515), .o (n5516) );
  buffer buf_n5517( .i (n5516), .o (n5517) );
  buffer buf_n5518( .i (n5517), .o (n5518) );
  buffer buf_n5519( .i (n5518), .o (n5519) );
  buffer buf_n5520( .i (n5519), .o (n5520) );
  assign n5521 = ~n2589 & n5511 ;
  buffer buf_n5522( .i (n5521), .o (n5522) );
  buffer buf_n5523( .i (n5522), .o (n5523) );
  buffer buf_n5524( .i (n5523), .o (n5524) );
  buffer buf_n5525( .i (n5524), .o (n5525) );
  buffer buf_n5526( .i (n5525), .o (n5526) );
  buffer buf_n5527( .i (n5526), .o (n5527) );
  buffer buf_n5528( .i (n5527), .o (n5528) );
  buffer buf_n2516( .i (N331), .o (n2516) );
  buffer buf_n2517( .i (n2516), .o (n2517) );
  buffer buf_n2518( .i (n2517), .o (n2518) );
  buffer buf_n2519( .i (n2518), .o (n2519) );
  buffer buf_n2520( .i (n2519), .o (n2520) );
  buffer buf_n2521( .i (n2520), .o (n2521) );
  buffer buf_n2522( .i (n2521), .o (n2522) );
  buffer buf_n2523( .i (n2522), .o (n2523) );
  buffer buf_n753( .i (N232), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  assign n5529 = n756 & n5505 ;
  buffer buf_n5530( .i (n5529), .o (n5530) );
  buffer buf_n384( .i (N124), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  assign n5531 = n387 & ~n5505 ;
  buffer buf_n5532( .i (n5531), .o (n5532) );
  assign n5533 = n5530 | n5532 ;
  buffer buf_n5534( .i (n5533), .o (n5534) );
  assign n5535 = n2523 & ~n5534 ;
  buffer buf_n5536( .i (n5535), .o (n5536) );
  buffer buf_n5537( .i (n5536), .o (n5537) );
  buffer buf_n5538( .i (n5537), .o (n5538) );
  buffer buf_n5539( .i (n5538), .o (n5539) );
  buffer buf_n5540( .i (n5539), .o (n5540) );
  assign n5541 = ~n2523 & n5534 ;
  buffer buf_n5542( .i (n5541), .o (n5542) );
  buffer buf_n5543( .i (n5542), .o (n5543) );
  buffer buf_n5544( .i (n5543), .o (n5544) );
  buffer buf_n5545( .i (n5544), .o (n5545) );
  buffer buf_n2450( .i (N328), .o (n2450) );
  buffer buf_n2451( .i (n2450), .o (n2451) );
  buffer buf_n2452( .i (n2451), .o (n2452) );
  buffer buf_n2453( .i (n2452), .o (n2453) );
  buffer buf_n2454( .i (n2453), .o (n2454) );
  buffer buf_n2455( .i (n2454), .o (n2455) );
  buffer buf_n2456( .i (n2455), .o (n2456) );
  buffer buf_n2457( .i (n2456), .o (n2457) );
  buffer buf_n757( .i (N233), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n5546( .i (n5387), .o (n5546) );
  assign n5547 = n760 & n5546 ;
  buffer buf_n5548( .i (n5547), .o (n5548) );
  buffer buf_n388( .i (N127), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  assign n5549 = n391 & ~n5546 ;
  buffer buf_n5550( .i (n5549), .o (n5550) );
  assign n5551 = n5548 | n5550 ;
  buffer buf_n5552( .i (n5551), .o (n5552) );
  assign n5553 = n2457 & ~n5552 ;
  buffer buf_n5554( .i (n5553), .o (n5554) );
  buffer buf_n5555( .i (n5554), .o (n5555) );
  assign n5556 = ~n2457 & n5552 ;
  buffer buf_n5557( .i (n5556), .o (n5557) );
  buffer buf_n2384( .i (N325), .o (n2384) );
  buffer buf_n2385( .i (n2384), .o (n2385) );
  buffer buf_n2386( .i (n2385), .o (n2386) );
  buffer buf_n2387( .i (n2386), .o (n2387) );
  buffer buf_n2388( .i (n2387), .o (n2388) );
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2391( .i (n2390), .o (n2391) );
  buffer buf_n761( .i (N234), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  assign n5559 = n764 & n5546 ;
  buffer buf_n5560( .i (n5559), .o (n5560) );
  buffer buf_n392( .i (N130), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  assign n5561 = n395 & ~n5546 ;
  buffer buf_n5562( .i (n5561), .o (n5562) );
  assign n5563 = n5560 | n5562 ;
  buffer buf_n5564( .i (n5563), .o (n5564) );
  assign n5565 = ~n2391 & n5564 ;
  buffer buf_n5566( .i (n5565), .o (n5566) );
  assign n5585 = n5557 | n5566 ;
  assign n5586 = ~n5555 & n5585 ;
  buffer buf_n5587( .i (n5586), .o (n5587) );
  assign n5604 = n5545 | n5587 ;
  assign n5605 = ~n5540 & n5604 ;
  buffer buf_n5606( .i (n5605), .o (n5606) );
  assign n5618 = n5528 | n5606 ;
  assign n5619 = ~n5520 & n5618 ;
  buffer buf_n5620( .i (n5619), .o (n5620) );
  buffer buf_n5621( .i (n5620), .o (n5621) );
  buffer buf_n5622( .i (n5621), .o (n5622) );
  buffer buf_n5623( .i (n5622), .o (n5623) );
  buffer buf_n5624( .i (n5623), .o (n5624) );
  buffer buf_n5625( .i (n5624), .o (n5625) );
  buffer buf_n5626( .i (n5625), .o (n5626) );
  buffer buf_n5627( .i (n5626), .o (n5627) );
  buffer buf_n5628( .i (n5627), .o (n5628) );
  buffer buf_n3322( .i (n3321), .o (n3322) );
  buffer buf_n3323( .i (n3322), .o (n3323) );
  buffer buf_n3324( .i (n3323), .o (n3324) );
  buffer buf_n3325( .i (n3324), .o (n3325) );
  buffer buf_n3326( .i (n3325), .o (n3326) );
  buffer buf_n3327( .i (n3326), .o (n3327) );
  buffer buf_n3328( .i (n3327), .o (n3328) );
  buffer buf_n3329( .i (n3328), .o (n3329) );
  buffer buf_n3330( .i (n3329), .o (n3330) );
  buffer buf_n3331( .i (n3330), .o (n3331) );
  buffer buf_n3332( .i (n3331), .o (n3332) );
  buffer buf_n3333( .i (n3332), .o (n3333) );
  buffer buf_n2318( .i (N322), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n2321( .i (n2320), .o (n2321) );
  buffer buf_n2322( .i (n2321), .o (n2322) );
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2325( .i (n2324), .o (n2325) );
  buffer buf_n765( .i (N235), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n5629( .i (n5387), .o (n5629) );
  assign n5630 = n768 & n5629 ;
  buffer buf_n5631( .i (n5630), .o (n5631) );
  buffer buf_n278( .i (N103), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  assign n5632 = n281 & ~n5629 ;
  buffer buf_n5633( .i (n5632), .o (n5633) );
  assign n5634 = n5631 | n5633 ;
  buffer buf_n5635( .i (n5634), .o (n5635) );
  assign n5636 = ~n2325 & n5635 ;
  buffer buf_n5637( .i (n5636), .o (n5637) );
  buffer buf_n5638( .i (n5637), .o (n5638) );
  buffer buf_n5639( .i (n5638), .o (n5639) );
  buffer buf_n5640( .i (n5639), .o (n5640) );
  buffer buf_n5641( .i (n5640), .o (n5641) );
  buffer buf_n5642( .i (n5641), .o (n5642) );
  buffer buf_n5643( .i (n5642), .o (n5643) );
  buffer buf_n5644( .i (n5643), .o (n5644) );
  buffer buf_n5645( .i (n5644), .o (n5645) );
  buffer buf_n5646( .i (n5645), .o (n5646) );
  buffer buf_n5647( .i (n5646), .o (n5647) );
  assign n5650 = n2325 & ~n5635 ;
  buffer buf_n5651( .i (n5650), .o (n5651) );
  buffer buf_n5652( .i (n5651), .o (n5652) );
  buffer buf_n5653( .i (n5652), .o (n5653) );
  buffer buf_n5654( .i (n5653), .o (n5654) );
  buffer buf_n5655( .i (n5654), .o (n5655) );
  buffer buf_n5656( .i (n5655), .o (n5656) );
  buffer buf_n5657( .i (n5656), .o (n5657) );
  buffer buf_n5658( .i (n5657), .o (n5658) );
  buffer buf_n5659( .i (n5658), .o (n5659) );
  buffer buf_n5660( .i (n5659), .o (n5660) );
  buffer buf_n2248( .i (N319), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  buffer buf_n2250( .i (n2249), .o (n2250) );
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n769( .i (N236), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  assign n5663 = n772 & n5629 ;
  buffer buf_n5664( .i (n5663), .o (n5664) );
  buffer buf_n745( .i (N23), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  assign n5665 = n748 & ~n5629 ;
  buffer buf_n5666( .i (n5665), .o (n5666) );
  assign n5667 = n5664 | n5666 ;
  buffer buf_n5668( .i (n5667), .o (n5668) );
  assign n5669 = n2255 & ~n5668 ;
  buffer buf_n5670( .i (n5669), .o (n5670) );
  buffer buf_n5671( .i (n5670), .o (n5671) );
  buffer buf_n5672( .i (n5671), .o (n5672) );
  buffer buf_n5673( .i (n5672), .o (n5673) );
  buffer buf_n5674( .i (n5673), .o (n5674) );
  buffer buf_n5675( .i (n5674), .o (n5675) );
  buffer buf_n5676( .i (n5675), .o (n5676) );
  buffer buf_n5677( .i (n5676), .o (n5677) );
  assign n5680 = ~n2255 & n5668 ;
  buffer buf_n5681( .i (n5680), .o (n5681) );
  buffer buf_n5682( .i (n5681), .o (n5682) );
  buffer buf_n5683( .i (n5682), .o (n5683) );
  buffer buf_n5684( .i (n5683), .o (n5684) );
  buffer buf_n5685( .i (n5684), .o (n5685) );
  buffer buf_n5686( .i (n5685), .o (n5686) );
  buffer buf_n2182( .i (N316), .o (n2182) );
  buffer buf_n2183( .i (n2182), .o (n2183) );
  buffer buf_n2184( .i (n2183), .o (n2184) );
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  buffer buf_n2187( .i (n2186), .o (n2187) );
  buffer buf_n2188( .i (n2187), .o (n2188) );
  buffer buf_n2189( .i (n2188), .o (n2189) );
  buffer buf_n773( .i (N237), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n5687( .i (n587), .o (n5687) );
  buffer buf_n5688( .i (n5687), .o (n5688) );
  assign n5689 = n776 & n5688 ;
  buffer buf_n5690( .i (n5689), .o (n5690) );
  buffer buf_n1117( .i (N26), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  assign n5691 = n1120 & ~n5688 ;
  buffer buf_n5692( .i (n5691), .o (n5692) );
  assign n5693 = n5690 | n5692 ;
  buffer buf_n5694( .i (n5693), .o (n5694) );
  assign n5695 = n2189 & ~n5694 ;
  buffer buf_n5696( .i (n5695), .o (n5696) );
  buffer buf_n5697( .i (n5696), .o (n5697) );
  buffer buf_n5698( .i (n5697), .o (n5698) );
  buffer buf_n5699( .i (n5698), .o (n5699) );
  buffer buf_n3612( .i (n3611), .o (n3612) );
  buffer buf_n3613( .i (n3612), .o (n3613) );
  buffer buf_n2116( .i (N313), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  buffer buf_n2119( .i (n2118), .o (n2119) );
  buffer buf_n2120( .i (n2119), .o (n2120) );
  buffer buf_n2121( .i (n2120), .o (n2121) );
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n777( .i (N238), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  assign n5700 = n780 & n5688 ;
  buffer buf_n5701( .i (n5700), .o (n5701) );
  buffer buf_n1716( .i (N29), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n1719( .i (n1718), .o (n1719) );
  assign n5702 = n1719 & ~n5688 ;
  buffer buf_n5703( .i (n5702), .o (n5703) );
  assign n5704 = n5701 | n5703 ;
  buffer buf_n5705( .i (n5704), .o (n5705) );
  assign n5706 = n2123 & ~n5705 ;
  buffer buf_n5707( .i (n5706), .o (n5707) );
  assign n5711 = n3613 & ~n5707 ;
  buffer buf_n5712( .i (n5711), .o (n5712) );
  assign n5713 = ~n2189 & n5694 ;
  buffer buf_n5714( .i (n5713), .o (n5714) );
  assign n5715 = ~n2123 & n5705 ;
  buffer buf_n5716( .i (n5715), .o (n5716) );
  assign n5719 = n5714 | n5716 ;
  buffer buf_n5720( .i (n5719), .o (n5720) );
  assign n5721 = n5712 | n5720 ;
  assign n5722 = ~n5699 & n5721 ;
  buffer buf_n5723( .i (n5722), .o (n5723) );
  assign n5727 = n5686 | n5723 ;
  buffer buf_n5728( .i (n5727), .o (n5728) );
  assign n5730 = ~n5677 & n5728 ;
  buffer buf_n5731( .i (n5730), .o (n5731) );
  assign n5732 = ~n5660 & n5731 ;
  assign n5733 = n5647 | n5732 ;
  buffer buf_n5734( .i (n5733), .o (n5734) );
  assign n5735 = n3333 | n5734 ;
  buffer buf_n5736( .i (n5735), .o (n5736) );
  buffer buf_n5648( .i (n5647), .o (n5648) );
  buffer buf_n5649( .i (n5648), .o (n5649) );
  buffer buf_n5661( .i (n5660), .o (n5661) );
  buffer buf_n5662( .i (n5661), .o (n5662) );
  assign n5737 = n5696 | n5714 ;
  buffer buf_n5738( .i (n5737), .o (n5738) );
  buffer buf_n5739( .i (n5738), .o (n5739) );
  buffer buf_n5740( .i (n5739), .o (n5740) );
  buffer buf_n3627( .i (n3626), .o (n3627) );
  buffer buf_n3628( .i (n3627), .o (n3628) );
  assign n5742 = n5707 | n5716 ;
  buffer buf_n5743( .i (n5742), .o (n5743) );
  assign n5746 = n3628 | n5743 ;
  buffer buf_n5747( .i (n5746), .o (n5747) );
  assign n5748 = n5740 | n5747 ;
  buffer buf_n5749( .i (n5748), .o (n5749) );
  assign n5750 = n5670 | n5681 ;
  buffer buf_n5751( .i (n5750), .o (n5751) );
  buffer buf_n5752( .i (n5751), .o (n5752) );
  buffer buf_n5753( .i (n5752), .o (n5753) );
  buffer buf_n5754( .i (n5753), .o (n5754) );
  buffer buf_n5755( .i (n5754), .o (n5755) );
  assign n5760 = n5749 | n5755 ;
  buffer buf_n5761( .i (n5760), .o (n5761) );
  buffer buf_n5762( .i (n5761), .o (n5762) );
  assign n5763 = ~n5731 & n5762 ;
  buffer buf_n5764( .i (n5763), .o (n5764) );
  assign n5765 = n5662 | n5764 ;
  assign n5766 = ~n5649 & n5765 ;
  buffer buf_n5767( .i (n5766), .o (n5767) );
  assign n5768 = n5736 & ~n5767 ;
  buffer buf_n5769( .i (n5768), .o (n5769) );
  assign n5771 = n5554 | n5557 ;
  buffer buf_n5772( .i (n5771), .o (n5772) );
  buffer buf_n5773( .i (n5772), .o (n5773) );
  buffer buf_n5567( .i (n5566), .o (n5567) );
  assign n5791 = n2391 & ~n5564 ;
  buffer buf_n5792( .i (n5791), .o (n5792) );
  buffer buf_n5793( .i (n5792), .o (n5793) );
  assign n5809 = n5567 | n5793 ;
  buffer buf_n5810( .i (n5809), .o (n5810) );
  assign n5825 = n5773 | n5810 ;
  buffer buf_n5826( .i (n5825), .o (n5826) );
  assign n5827 = n5536 | n5542 ;
  buffer buf_n5828( .i (n5827), .o (n5828) );
  buffer buf_n5829( .i (n5828), .o (n5829) );
  assign n5848 = n5513 | n5522 ;
  buffer buf_n5849( .i (n5848), .o (n5849) );
  buffer buf_n5850( .i (n5849), .o (n5850) );
  assign n5867 = n5829 | n5850 ;
  buffer buf_n5868( .i (n5867), .o (n5868) );
  assign n5869 = n5826 | n5868 ;
  buffer buf_n5870( .i (n5869), .o (n5870) );
  buffer buf_n5871( .i (n5870), .o (n5871) );
  buffer buf_n5872( .i (n5871), .o (n5872) );
  buffer buf_n5873( .i (n5872), .o (n5873) );
  buffer buf_n5874( .i (n5873), .o (n5874) );
  buffer buf_n5875( .i (n5874), .o (n5875) );
  buffer buf_n5876( .i (n5875), .o (n5876) );
  buffer buf_n5877( .i (n5876), .o (n5877) );
  buffer buf_n5878( .i (n5877), .o (n5878) );
  buffer buf_n5879( .i (n5878), .o (n5879) );
  assign n5880 = n5769 & ~n5879 ;
  assign n5881 = n5628 | n5880 ;
  buffer buf_n5882( .i (n5881), .o (n5882) );
  assign n5885 = ~n5504 & n5882 ;
  buffer buf_n5886( .i (n5885), .o (n5886) );
  buffer buf_n5458( .i (n5457), .o (n5458) );
  buffer buf_n5459( .i (n5458), .o (n5459) );
  buffer buf_n5460( .i (n5459), .o (n5460) );
  buffer buf_n5461( .i (n5460), .o (n5461) );
  buffer buf_n5462( .i (n5461), .o (n5462) );
  buffer buf_n5463( .i (n5462), .o (n5463) );
  buffer buf_n5464( .i (n5463), .o (n5464) );
  buffer buf_n5465( .i (n5464), .o (n5465) );
  buffer buf_n5466( .i (n5465), .o (n5466) );
  buffer buf_n5467( .i (n5466), .o (n5467) );
  buffer buf_n5468( .i (n5467), .o (n5468) );
  buffer buf_n5469( .i (n5468), .o (n5469) );
  buffer buf_n5472( .i (n5471), .o (n5472) );
  buffer buf_n5473( .i (n5472), .o (n5473) );
  buffer buf_n5474( .i (n5473), .o (n5474) );
  buffer buf_n5475( .i (n5474), .o (n5475) );
  buffer buf_n5476( .i (n5475), .o (n5476) );
  buffer buf_n5477( .i (n5476), .o (n5477) );
  buffer buf_n5478( .i (n5477), .o (n5478) );
  buffer buf_n5479( .i (n5478), .o (n5479) );
  buffer buf_n5480( .i (n5479), .o (n5480) );
  buffer buf_n5481( .i (n5480), .o (n5481) );
  buffer buf_n5482( .i (n5481), .o (n5482) );
  buffer buf_n5356( .i (n5355), .o (n5356) );
  buffer buf_n5357( .i (n5356), .o (n5357) );
  buffer buf_n5358( .i (n5357), .o (n5358) );
  buffer buf_n5359( .i (n5358), .o (n5359) );
  buffer buf_n5360( .i (n5359), .o (n5360) );
  buffer buf_n5361( .i (n5360), .o (n5361) );
  buffer buf_n5362( .i (n5361), .o (n5362) );
  buffer buf_n5363( .i (n5362), .o (n5363) );
  buffer buf_n5364( .i (n5363), .o (n5364) );
  buffer buf_n5346( .i (n5345), .o (n5346) );
  buffer buf_n5347( .i (n5346), .o (n5347) );
  buffer buf_n5348( .i (n5347), .o (n5348) );
  buffer buf_n5349( .i (n5348), .o (n5349) );
  buffer buf_n5350( .i (n5349), .o (n5350) );
  buffer buf_n5351( .i (n5350), .o (n5351) );
  buffer buf_n5352( .i (n5351), .o (n5352) );
  buffer buf_n5353( .i (n5352), .o (n5353) );
  buffer buf_n5403( .i (n5402), .o (n5403) );
  buffer buf_n5404( .i (n5403), .o (n5404) );
  buffer buf_n5405( .i (n5404), .o (n5405) );
  buffer buf_n5406( .i (n5405), .o (n5406) );
  buffer buf_n5407( .i (n5406), .o (n5407) );
  buffer buf_n5408( .i (n5407), .o (n5408) );
  buffer buf_n5397( .i (n5396), .o (n5397) );
  buffer buf_n5398( .i (n5397), .o (n5398) );
  buffer buf_n5399( .i (n5398), .o (n5399) );
  buffer buf_n5400( .i (n5399), .o (n5400) );
  buffer buf_n5331( .i (n5330), .o (n5331) );
  assign n5887 = n5272 | n5331 ;
  assign n5888 = ~n5305 & n5887 ;
  buffer buf_n5889( .i (n5888), .o (n5889) );
  assign n5910 = ~n5400 & n5889 ;
  buffer buf_n5911( .i (n5910), .o (n5911) );
  assign n5912 = n5408 | n5911 ;
  buffer buf_n5913( .i (n5912), .o (n5913) );
  assign n5926 = ~n5353 & n5913 ;
  assign n5927 = n5364 | n5926 ;
  buffer buf_n5928( .i (n5927), .o (n5928) );
  assign n5929 = ~n5482 & n5928 ;
  assign n5930 = n5469 | n5929 ;
  buffer buf_n5931( .i (n5930), .o (n5931) );
  buffer buf_n5932( .i (n5931), .o (n5932) );
  buffer buf_n5933( .i (n5932), .o (n5933) );
  buffer buf_n5934( .i (n5933), .o (n5934) );
  buffer buf_n5935( .i (n5934), .o (n5935) );
  buffer buf_n5936( .i (n5935), .o (n5936) );
  buffer buf_n5937( .i (n5936), .o (n5937) );
  buffer buf_n5938( .i (n5937), .o (n5938) );
  assign n5939 = n5886 | n5938 ;
  buffer buf_n5940( .i (n5939), .o (n5940) );
  assign n5944 = n5150 | n5940 ;
  assign n5945 = ~n5263 & n5944 ;
  buffer buf_n5946( .i (n5945), .o (n5946) );
  assign n5947 = ~n5040 & n5946 ;
  assign n5948 = n5012 | n5947 ;
  buffer buf_n5949( .i (n5948), .o (n5949) );
  assign n5954 = n4791 & ~n5949 ;
  assign n5955 = n4977 | n5954 ;
  buffer buf_n5956( .i (n5955), .o (n5956) );
  assign n5962 = n4428 & n5956 ;
  assign n5963 = n4555 | n5962 ;
  buffer buf_n5964( .i (n5963), .o (n5964) );
  assign n5965 = n4291 & n5964 ;
  assign n5966 = n4255 | n5965 ;
  buffer buf_n5967( .i (n5966), .o (n5967) );
  assign n5974 = n3961 & ~n3968 ;
  buffer buf_n5975( .i (n5974), .o (n5975) );
  buffer buf_n5976( .i (n5975), .o (n5976) );
  buffer buf_n5977( .i (n5976), .o (n5977) );
  assign n6015 = n926 & n3987 ;
  buffer buf_n6016( .i (n6015), .o (n6016) );
  assign n6017 = n3989 & ~n6016 ;
  buffer buf_n6018( .i (n6017), .o (n6018) );
  assign n6061 = ~n3981 & n4037 ;
  buffer buf_n6062( .i (n6061), .o (n6062) );
  assign n6109 = n6018 & n6062 ;
  buffer buf_n6110( .i (n6109), .o (n6110) );
  assign n6145 = n5977 & n6110 ;
  buffer buf_n6146( .i (n6145), .o (n6146) );
  buffer buf_n6147( .i (n6146), .o (n6147) );
  buffer buf_n6148( .i (n6147), .o (n6148) );
  buffer buf_n6149( .i (n6148), .o (n6149) );
  buffer buf_n6150( .i (n6149), .o (n6150) );
  buffer buf_n6151( .i (n6150), .o (n6151) );
  buffer buf_n6152( .i (n6151), .o (n6152) );
  buffer buf_n6153( .i (n6152), .o (n6153) );
  buffer buf_n6154( .i (n6153), .o (n6154) );
  buffer buf_n6155( .i (n6154), .o (n6155) );
  buffer buf_n6156( .i (n6155), .o (n6156) );
  buffer buf_n6157( .i (n6156), .o (n6157) );
  buffer buf_n6158( .i (n6157), .o (n6158) );
  buffer buf_n6159( .i (n6158), .o (n6159) );
  buffer buf_n6160( .i (n6159), .o (n6160) );
  buffer buf_n6161( .i (n6160), .o (n6161) );
  buffer buf_n6162( .i (n6161), .o (n6162) );
  buffer buf_n6163( .i (n6162), .o (n6163) );
  buffer buf_n6164( .i (n6163), .o (n6164) );
  buffer buf_n6165( .i (n6164), .o (n6165) );
  buffer buf_n6166( .i (n6165), .o (n6166) );
  buffer buf_n6167( .i (n6166), .o (n6167) );
  buffer buf_n6168( .i (n6167), .o (n6168) );
  buffer buf_n6169( .i (n6168), .o (n6169) );
  buffer buf_n6170( .i (n6169), .o (n6170) );
  buffer buf_n6171( .i (n6170), .o (n6171) );
  buffer buf_n6172( .i (n6171), .o (n6172) );
  buffer buf_n6173( .i (n6172), .o (n6173) );
  buffer buf_n6174( .i (n6173), .o (n6174) );
  buffer buf_n6175( .i (n6174), .o (n6175) );
  buffer buf_n6176( .i (n6175), .o (n6176) );
  buffer buf_n6177( .i (n6176), .o (n6177) );
  buffer buf_n6178( .i (n6177), .o (n6178) );
  assign n6179 = ~n5967 & n6178 ;
  buffer buf_n6180( .i (n6179), .o (n6180) );
  assign n6181 = n4210 & n6180 ;
  assign n6182 = n4212 & ~n6181 ;
  buffer buf_n6183( .i (n6182), .o (n6183) );
  buffer buf_n6184( .i (n6183), .o (n6184) );
  buffer buf_n6185( .i (n6184), .o (n6185) );
  buffer buf_n6186( .i (n6185), .o (n6186) );
  buffer buf_n6187( .i (n6186), .o (n6187) );
  buffer buf_n6188( .i (n6187), .o (n6188) );
  buffer buf_n6189( .i (n6188), .o (n6189) );
  buffer buf_n6190( .i (n6189), .o (n6190) );
  assign n6191 = n3877 | n6190 ;
  buffer buf_n6192( .i (n6191), .o (n6192) );
  assign n6193 = ~n3864 & n6192 ;
  assign n6194 = n3806 | n6193 ;
  buffer buf_n6195( .i (n6194), .o (n6195) );
  buffer buf_n6196( .i (n6195), .o (n6196) );
  buffer buf_n852( .i (N245), .o (n852) );
  buffer buf_n1319( .i (N271), .o (n1319) );
  assign n6197 = n852 & n1319 ;
  buffer buf_n6198( .i (n6197), .o (n6198) );
  assign n6199 = ~n3338 & n3394 ;
  assign n6200 = ~n6198 & n6199 ;
  buffer buf_n6201( .i (n6200), .o (n6201) );
  buffer buf_n6202( .i (n6201), .o (n6202) );
  buffer buf_n6203( .i (n6202), .o (n6203) );
  buffer buf_n6204( .i (n6203), .o (n6204) );
  buffer buf_n6205( .i (n6204), .o (n6205) );
  buffer buf_n6206( .i (n6205), .o (n6206) );
  buffer buf_n6207( .i (n6206), .o (n6207) );
  buffer buf_n6208( .i (n6207), .o (n6208) );
  buffer buf_n6209( .i (n6208), .o (n6209) );
  buffer buf_n6210( .i (n6209), .o (n6210) );
  buffer buf_n6211( .i (n6210), .o (n6211) );
  buffer buf_n6212( .i (n6211), .o (n6212) );
  buffer buf_n6213( .i (n6212), .o (n6213) );
  buffer buf_n6214( .i (n6213), .o (n6214) );
  buffer buf_n6215( .i (n6214), .o (n6215) );
  buffer buf_n6216( .i (n6215), .o (n6216) );
  buffer buf_n6217( .i (n6216), .o (n6217) );
  buffer buf_n6218( .i (n6217), .o (n6218) );
  buffer buf_n6219( .i (n6218), .o (n6219) );
  buffer buf_n6220( .i (n6219), .o (n6220) );
  buffer buf_n6221( .i (n6220), .o (n6221) );
  buffer buf_n6222( .i (n6221), .o (n6222) );
  buffer buf_n6223( .i (n6222), .o (n6223) );
  buffer buf_n6224( .i (n6223), .o (n6224) );
  buffer buf_n6225( .i (n6224), .o (n6225) );
  buffer buf_n3464( .i (N53), .o (n3464) );
  buffer buf_n3465( .i (n3464), .o (n3465) );
  buffer buf_n3466( .i (n3465), .o (n3466) );
  buffer buf_n3467( .i (n3466), .o (n3467) );
  buffer buf_n6226( .i (n5687), .o (n6226) );
  assign n6227 = n3467 & ~n6226 ;
  assign n6228 = ~n2387 & n6226 ;
  assign n6229 = n6227 | n6228 ;
  buffer buf_n6230( .i (n6229), .o (n6230) );
  buffer buf_n6231( .i (n6230), .o (n6231) );
  buffer buf_n655( .i (N203), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  assign n6232 = n658 & n6226 ;
  buffer buf_n6233( .i (n6232), .o (n6233) );
  assign n6234 = n5562 | n6233 ;
  buffer buf_n6235( .i (n6234), .o (n6235) );
  assign n6236 = n6231 | n6235 ;
  buffer buf_n6237( .i (n6236), .o (n6237) );
  buffer buf_n6238( .i (n6237), .o (n6238) );
  buffer buf_n6239( .i (n6238), .o (n6239) );
  buffer buf_n6240( .i (n6239), .o (n6240) );
  buffer buf_n6241( .i (n6240), .o (n6241) );
  buffer buf_n3527( .i (N73), .o (n3527) );
  buffer buf_n3528( .i (n3527), .o (n3528) );
  buffer buf_n3529( .i (n3528), .o (n3529) );
  buffer buf_n3530( .i (n3529), .o (n3530) );
  assign n6242 = n3530 & ~n6226 ;
  buffer buf_n6243( .i (n5687), .o (n6243) );
  assign n6244 = ~n2321 & n6243 ;
  assign n6245 = n6242 | n6244 ;
  buffer buf_n6246( .i (n6245), .o (n6246) );
  buffer buf_n6247( .i (n6246), .o (n6247) );
  buffer buf_n659( .i (N204), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  assign n6248 = n662 & n6243 ;
  buffer buf_n6249( .i (n6248), .o (n6249) );
  assign n6250 = n5633 | n6249 ;
  buffer buf_n6251( .i (n6250), .o (n6251) );
  assign n6252 = n6247 & n6251 ;
  buffer buf_n6253( .i (n6252), .o (n6253) );
  buffer buf_n6254( .i (n6253), .o (n6254) );
  buffer buf_n6255( .i (n6254), .o (n6255) );
  buffer buf_n6256( .i (n6255), .o (n6256) );
  buffer buf_n3531( .i (N74), .o (n3531) );
  buffer buf_n3532( .i (n3531), .o (n3532) );
  buffer buf_n3533( .i (n3532), .o (n3533) );
  buffer buf_n3534( .i (n3533), .o (n3534) );
  buffer buf_n3535( .i (n3534), .o (n3535) );
  assign n6257 = ~n590 & n3535 ;
  buffer buf_n6258( .i (n6243), .o (n6258) );
  assign n6259 = ~n2120 & n6258 ;
  assign n6260 = n6257 | n6259 ;
  buffer buf_n6261( .i (n6260), .o (n6261) );
  buffer buf_n671( .i (N207), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  assign n6262 = n674 & n6243 ;
  buffer buf_n6263( .i (n6262), .o (n6263) );
  assign n6264 = n5703 | n6263 ;
  buffer buf_n6265( .i (n6264), .o (n6265) );
  assign n6266 = n6261 & n6265 ;
  buffer buf_n3522( .i (N70), .o (n3522) );
  buffer buf_n3523( .i (n3522), .o (n3523) );
  buffer buf_n3524( .i (n3523), .o (n3524) );
  buffer buf_n3525( .i (n3524), .o (n3525) );
  buffer buf_n3526( .i (n3525), .o (n3526) );
  buffer buf_n3594( .i (N89), .o (n3594) );
  buffer buf_n3595( .i (n3594), .o (n3595) );
  buffer buf_n3596( .i (n3595), .o (n3596) );
  buffer buf_n3597( .i (n3596), .o (n3597) );
  buffer buf_n3598( .i (n3597), .o (n3598) );
  assign n6267 = n3526 | n3598 ;
  assign n6268 = n3609 & n6267 ;
  buffer buf_n3599( .i (n3598), .o (n3599) );
  buffer buf_n6269( .i (n5687), .o (n6269) );
  assign n6270 = n3525 | n6269 ;
  buffer buf_n6271( .i (n6270), .o (n6271) );
  assign n6272 = n3599 & n6271 ;
  assign n6273 = n6268 | n6272 ;
  buffer buf_n6274( .i (n6273), .o (n6274) );
  assign n6275 = n6266 | n6274 ;
  buffer buf_n3540( .i (N76), .o (n3540) );
  buffer buf_n3541( .i (n3540), .o (n3541) );
  buffer buf_n3542( .i (n3541), .o (n3542) );
  buffer buf_n3543( .i (n3542), .o (n3543) );
  buffer buf_n3544( .i (n3543), .o (n3544) );
  assign n6276 = n3544 & ~n6258 ;
  assign n6277 = ~n2186 & n6258 ;
  assign n6278 = n6276 | n6277 ;
  buffer buf_n6279( .i (n6278), .o (n6279) );
  buffer buf_n667( .i (N206), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  assign n6280 = n670 & n6269 ;
  buffer buf_n6281( .i (n6280), .o (n6281) );
  assign n6282 = n5692 | n6281 ;
  buffer buf_n6283( .i (n6282), .o (n6283) );
  assign n6284 = n6279 | n6283 ;
  assign n6285 = n6261 | n6265 ;
  assign n6286 = n6284 & n6285 ;
  assign n6287 = n6275 & n6286 ;
  assign n6288 = n6279 & n6283 ;
  buffer buf_n3536( .i (N75), .o (n3536) );
  buffer buf_n3537( .i (n3536), .o (n3537) );
  buffer buf_n3538( .i (n3537), .o (n3538) );
  buffer buf_n3539( .i (n3538), .o (n3539) );
  assign n6289 = n3539 & ~n6269 ;
  assign n6290 = ~n2251 & n6269 ;
  assign n6291 = n6289 | n6290 ;
  buffer buf_n6292( .i (n6291), .o (n6292) );
  buffer buf_n6293( .i (n6292), .o (n6293) );
  buffer buf_n663( .i (N205), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n6296( .i (n586), .o (n6296) );
  buffer buf_n6297( .i (n6296), .o (n6297) );
  buffer buf_n6298( .i (n6297), .o (n6298) );
  assign n6299 = n666 & n6298 ;
  buffer buf_n6300( .i (n6299), .o (n6300) );
  assign n6301 = n5666 | n6300 ;
  buffer buf_n6302( .i (n6301), .o (n6302) );
  assign n6303 = n6293 & n6302 ;
  assign n6304 = n6288 | n6303 ;
  buffer buf_n6305( .i (n6304), .o (n6305) );
  assign n6306 = n6287 | n6305 ;
  assign n6307 = n6247 | n6251 ;
  assign n6308 = n6293 | n6302 ;
  assign n6309 = n6307 & n6308 ;
  buffer buf_n6310( .i (n6309), .o (n6310) );
  buffer buf_n6311( .i (n6310), .o (n6311) );
  assign n6312 = n6306 & n6311 ;
  assign n6313 = n6256 | n6312 ;
  assign n6314 = n6241 & n6313 ;
  buffer buf_n3468( .i (N54), .o (n3468) );
  buffer buf_n3469( .i (n3468), .o (n3469) );
  buffer buf_n3470( .i (n3469), .o (n3470) );
  buffer buf_n3471( .i (n3470), .o (n3471) );
  assign n6315 = n3471 & ~n6298 ;
  assign n6316 = ~n2453 & n6298 ;
  assign n6317 = n6315 | n6316 ;
  buffer buf_n6318( .i (n6317), .o (n6318) );
  buffer buf_n6319( .i (n6318), .o (n6319) );
  buffer buf_n651( .i (N202), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  assign n6322 = n654 & n6298 ;
  buffer buf_n6323( .i (n6322), .o (n6323) );
  assign n6324 = n5550 | n6323 ;
  buffer buf_n6325( .i (n6324), .o (n6325) );
  assign n6326 = n6319 & n6325 ;
  assign n6327 = n6231 & n6235 ;
  assign n6328 = n6326 | n6327 ;
  buffer buf_n6329( .i (n6328), .o (n6329) );
  buffer buf_n6330( .i (n6329), .o (n6330) );
  buffer buf_n6331( .i (n6330), .o (n6331) );
  buffer buf_n6332( .i (n6331), .o (n6332) );
  buffer buf_n6333( .i (n6332), .o (n6333) );
  assign n6334 = n6314 | n6333 ;
  buffer buf_n3476( .i (N56), .o (n3476) );
  buffer buf_n3477( .i (n3476), .o (n3477) );
  buffer buf_n3478( .i (n3477), .o (n3478) );
  buffer buf_n3479( .i (n3478), .o (n3479) );
  buffer buf_n6335( .i (n6297), .o (n6335) );
  assign n6336 = n3479 & ~n6335 ;
  assign n6337 = ~n2585 & n6335 ;
  assign n6338 = n6336 | n6337 ;
  buffer buf_n6339( .i (n6338), .o (n6339) );
  buffer buf_n6340( .i (n6339), .o (n6340) );
  buffer buf_n643( .i (N200), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  assign n6341 = n646 & n6335 ;
  buffer buf_n6342( .i (n6341), .o (n6342) );
  assign n6343 = n5509 | n6342 ;
  buffer buf_n6344( .i (n6343), .o (n6344) );
  assign n6345 = n6340 | n6344 ;
  buffer buf_n6346( .i (n6345), .o (n6346) );
  buffer buf_n3472( .i (N55), .o (n3472) );
  buffer buf_n3473( .i (n3472), .o (n3473) );
  buffer buf_n3474( .i (n3473), .o (n3474) );
  buffer buf_n3475( .i (n3474), .o (n3475) );
  assign n6347 = n3475 & ~n6335 ;
  buffer buf_n6348( .i (n6297), .o (n6348) );
  assign n6349 = ~n2519 & n6348 ;
  assign n6350 = n6347 | n6349 ;
  buffer buf_n6351( .i (n6350), .o (n6351) );
  buffer buf_n6352( .i (n6351), .o (n6352) );
  buffer buf_n647( .i (N201), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  assign n6353 = n650 & n6348 ;
  buffer buf_n6354( .i (n6353), .o (n6354) );
  assign n6355 = n5532 | n6354 ;
  buffer buf_n6356( .i (n6355), .o (n6356) );
  assign n6357 = n6352 & n6356 ;
  buffer buf_n6358( .i (n6357), .o (n6358) );
  assign n6359 = n6346 & ~n6358 ;
  assign n6360 = n6319 | n6325 ;
  assign n6361 = n6352 | n6356 ;
  assign n6362 = n6360 & n6361 ;
  buffer buf_n6363( .i (n6362), .o (n6363) );
  assign n6364 = n6359 & n6363 ;
  buffer buf_n6365( .i (n6364), .o (n6365) );
  buffer buf_n6366( .i (n6365), .o (n6366) );
  buffer buf_n6367( .i (n6366), .o (n6367) );
  buffer buf_n6368( .i (n6367), .o (n6368) );
  assign n6369 = n6334 & n6368 ;
  assign n6370 = n6346 & n6358 ;
  assign n6371 = n6340 & n6344 ;
  buffer buf_n3545( .i (N77), .o (n3545) );
  buffer buf_n3546( .i (n3545), .o (n3546) );
  buffer buf_n3547( .i (n3546), .o (n3547) );
  buffer buf_n3548( .i (n3547), .o (n3548) );
  assign n6372 = n3548 & ~n6348 ;
  assign n6373 = ~n2717 & n6348 ;
  assign n6374 = n6372 | n6373 ;
  buffer buf_n6375( .i (n6374), .o (n6375) );
  buffer buf_n6376( .i (n6375), .o (n6376) );
  buffer buf_n599( .i (N187), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n6377( .i (n6297), .o (n6377) );
  assign n6378 = n602 & n6377 ;
  buffer buf_n6379( .i (n6378), .o (n6379) );
  assign n6380 = n5267 | n6379 ;
  buffer buf_n6381( .i (n6380), .o (n6381) );
  assign n6382 = n6376 & n6381 ;
  assign n6383 = n6371 | n6382 ;
  buffer buf_n6384( .i (n6383), .o (n6384) );
  assign n6385 = n6370 | n6384 ;
  buffer buf_n6386( .i (n6385), .o (n6386) );
  buffer buf_n6387( .i (n6386), .o (n6387) );
  buffer buf_n6388( .i (n6387), .o (n6388) );
  buffer buf_n6389( .i (n6388), .o (n6389) );
  buffer buf_n6390( .i (n6389), .o (n6390) );
  assign n6391 = n6369 | n6390 ;
  buffer buf_n3562( .i (N81), .o (n3562) );
  buffer buf_n3563( .i (n3562), .o (n3563) );
  buffer buf_n3564( .i (n3563), .o (n3564) );
  buffer buf_n3565( .i (n3564), .o (n3565) );
  assign n6392 = n3565 & ~n6377 ;
  assign n6393 = ~n2915 & n6377 ;
  assign n6394 = n6392 | n6393 ;
  buffer buf_n6395( .i (n6394), .o (n6395) );
  buffer buf_n6396( .i (n6395), .o (n6396) );
  buffer buf_n623( .i (N194), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  assign n6397 = n626 & n6377 ;
  buffer buf_n6398( .i (n6397), .o (n6398) );
  assign n6399 = n5341 | n6398 ;
  buffer buf_n6400( .i (n6399), .o (n6400) );
  assign n6401 = n6396 & n6400 ;
  buffer buf_n3558( .i (N80), .o (n3558) );
  buffer buf_n3559( .i (n3558), .o (n3559) );
  buffer buf_n3560( .i (n3559), .o (n3560) );
  buffer buf_n3561( .i (n3560), .o (n3561) );
  buffer buf_n6402( .i (n6296), .o (n6402) );
  buffer buf_n6403( .i (n6402), .o (n6403) );
  assign n6404 = n3561 & ~n6403 ;
  assign n6405 = ~n2985 & n6403 ;
  assign n6406 = n6404 | n6405 ;
  buffer buf_n6407( .i (n6406), .o (n6407) );
  buffer buf_n6408( .i (n6407), .o (n6408) );
  buffer buf_n619( .i (N193), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  assign n6409 = n622 & n6403 ;
  buffer buf_n6410( .i (n6409), .o (n6410) );
  assign n6411 = n5453 | n6410 ;
  buffer buf_n6412( .i (n6411), .o (n6412) );
  assign n6413 = n6408 & n6412 ;
  assign n6414 = n6401 | n6413 ;
  buffer buf_n6415( .i (n6414), .o (n6415) );
  buffer buf_n6416( .i (n6415), .o (n6416) );
  buffer buf_n3485( .i (N59), .o (n3485) );
  buffer buf_n3486( .i (n3485), .o (n3486) );
  buffer buf_n3487( .i (n3486), .o (n3487) );
  buffer buf_n3488( .i (n3487), .o (n3488) );
  buffer buf_n3489( .i (n3488), .o (n3489) );
  assign n6417 = n3489 & ~n6258 ;
  buffer buf_n6418( .i (n6403), .o (n6418) );
  assign n6419 = ~n2850 & n6418 ;
  assign n6420 = n6417 | n6419 ;
  buffer buf_n6421( .i (n6420), .o (n6421) );
  buffer buf_n627( .i (N195), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n6422( .i (n6402), .o (n6422) );
  assign n6423 = n630 & n6422 ;
  buffer buf_n6424( .i (n6423), .o (n6424) );
  assign n6425 = n5392 | n6424 ;
  buffer buf_n6426( .i (n6425), .o (n6426) );
  assign n6427 = n6421 | n6426 ;
  buffer buf_n6428( .i (n6427), .o (n6428) );
  buffer buf_n6429( .i (n6428), .o (n6429) );
  assign n6430 = n6396 | n6400 ;
  buffer buf_n6431( .i (n6430), .o (n6431) );
  assign n6432 = n6408 | n6412 ;
  buffer buf_n6433( .i (n6432), .o (n6433) );
  assign n6435 = n6431 & n6433 ;
  assign n6436 = n6429 & n6435 ;
  assign n6437 = ~n6416 & n6436 ;
  buffer buf_n6438( .i (n6437), .o (n6438) );
  buffer buf_n3549( .i (N78), .o (n3549) );
  buffer buf_n3550( .i (n3549), .o (n3550) );
  buffer buf_n3551( .i (n3550), .o (n3551) );
  buffer buf_n3552( .i (n3551), .o (n3552) );
  buffer buf_n3553( .i (n3552), .o (n3553) );
  assign n6439 = n3553 & ~n6418 ;
  assign n6440 = ~n2784 & n6418 ;
  assign n6441 = n6439 | n6440 ;
  buffer buf_n6442( .i (n6441), .o (n6442) );
  buffer buf_n631( .i (N196), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  assign n6443 = n634 & n6422 ;
  buffer buf_n6444( .i (n6443), .o (n6444) );
  assign n6445 = n5299 | n6444 ;
  buffer buf_n6446( .i (n6445), .o (n6446) );
  assign n6447 = n6442 & n6446 ;
  assign n6448 = n6421 & n6426 ;
  assign n6449 = n6447 | n6448 ;
  buffer buf_n6450( .i (n6449), .o (n6450) );
  assign n6454 = n6376 | n6381 ;
  assign n6455 = n6442 | n6446 ;
  assign n6456 = n6454 & n6455 ;
  buffer buf_n6457( .i (n6456), .o (n6457) );
  assign n6458 = ~n6450 & n6457 ;
  buffer buf_n6459( .i (n6458), .o (n6459) );
  buffer buf_n6460( .i (n6459), .o (n6460) );
  assign n6461 = n6438 & n6460 ;
  buffer buf_n6462( .i (n6461), .o (n6462) );
  buffer buf_n6463( .i (n6462), .o (n6463) );
  buffer buf_n6464( .i (n6463), .o (n6464) );
  assign n6465 = n6391 & n6464 ;
  buffer buf_n6451( .i (n6450), .o (n6451) );
  buffer buf_n6452( .i (n6451), .o (n6452) );
  buffer buf_n6453( .i (n6452), .o (n6453) );
  assign n6466 = n6438 & n6453 ;
  buffer buf_n6434( .i (n6433), .o (n6434) );
  assign n6467 = n6415 & n6434 ;
  buffer buf_n6468( .i (n6467), .o (n6468) );
  buffer buf_n6469( .i (n6468), .o (n6469) );
  buffer buf_n6470( .i (n6469), .o (n6470) );
  assign n6471 = n6466 | n6470 ;
  buffer buf_n6472( .i (n6471), .o (n6472) );
  buffer buf_n6473( .i (n6472), .o (n6473) );
  buffer buf_n6474( .i (n6473), .o (n6474) );
  assign n6475 = n6465 | n6474 ;
  buffer buf_n3498( .i (N62), .o (n3498) );
  buffer buf_n3499( .i (n3498), .o (n3499) );
  buffer buf_n3500( .i (n3499), .o (n3500) );
  buffer buf_n3501( .i (n3500), .o (n3501) );
  assign n6476 = n3501 & ~n6422 ;
  assign n6477 = ~n3249 & n6422 ;
  assign n6478 = n6476 | n6477 ;
  buffer buf_n6479( .i (n6478), .o (n6479) );
  buffer buf_n6480( .i (n6479), .o (n6480) );
  buffer buf_n603( .i (N189), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n6481( .i (n6402), .o (n6481) );
  assign n6482 = n606 & n6481 ;
  buffer buf_n6483( .i (n6482), .o (n6483) );
  assign n6484 = n4981 | n6483 ;
  buffer buf_n6485( .i (n6484), .o (n6485) );
  assign n6486 = n6480 | n6485 ;
  buffer buf_n6487( .i (n6486), .o (n6487) );
  buffer buf_n3494( .i (N61), .o (n3494) );
  buffer buf_n3495( .i (n3494), .o (n3495) );
  buffer buf_n3496( .i (n3495), .o (n3496) );
  buffer buf_n3497( .i (n3496), .o (n3497) );
  assign n6488 = n3497 & ~n6481 ;
  assign n6489 = ~n3183 & n6481 ;
  assign n6490 = n6488 | n6489 ;
  buffer buf_n6491( .i (n6490), .o (n6491) );
  buffer buf_n6492( .i (n6491), .o (n6492) );
  buffer buf_n607( .i (N190), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  assign n6493 = n610 & n6481 ;
  buffer buf_n6494( .i (n6493), .o (n6494) );
  assign n6495 = n5045 | n6494 ;
  buffer buf_n6496( .i (n6495), .o (n6496) );
  assign n6497 = n6492 & n6496 ;
  buffer buf_n6498( .i (n6497), .o (n6498) );
  assign n6499 = n6487 & ~n6498 ;
  assign n6500 = n6480 & n6485 ;
  buffer buf_n6501( .i (n6500), .o (n6501) );
  assign n6503 = n6492 | n6496 ;
  buffer buf_n6504( .i (n6503), .o (n6504) );
  assign n6505 = ~n6501 & n6504 ;
  assign n6506 = n6499 & n6505 ;
  buffer buf_n6507( .i (n6506), .o (n6507) );
  buffer buf_n3490( .i (N60), .o (n3490) );
  buffer buf_n3491( .i (n3490), .o (n3491) );
  buffer buf_n3492( .i (n3491), .o (n3492) );
  buffer buf_n3493( .i (n3492), .o (n3493) );
  buffer buf_n6508( .i (n6402), .o (n6508) );
  assign n6509 = n3493 & ~n6508 ;
  assign n6510 = ~n3117 & n6508 ;
  assign n6511 = n6509 | n6510 ;
  buffer buf_n6512( .i (n6511), .o (n6512) );
  buffer buf_n6513( .i (n6512), .o (n6513) );
  buffer buf_n611( .i (N191), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  assign n6514 = n614 & n6508 ;
  buffer buf_n6515( .i (n6514), .o (n6515) );
  assign n6516 = n5066 | n6515 ;
  buffer buf_n6517( .i (n6516), .o (n6517) );
  assign n6518 = n6513 & n6517 ;
  buffer buf_n3554( .i (N79), .o (n3554) );
  buffer buf_n3555( .i (n3554), .o (n3555) );
  buffer buf_n3556( .i (n3555), .o (n3556) );
  buffer buf_n3557( .i (n3556), .o (n3557) );
  assign n6519 = n3557 & ~n6508 ;
  buffer buf_n6520( .i (n6296), .o (n6520) );
  buffer buf_n6521( .i (n6520), .o (n6521) );
  assign n6522 = ~n3051 & n6521 ;
  assign n6523 = n6519 | n6522 ;
  buffer buf_n6524( .i (n6523), .o (n6524) );
  buffer buf_n6525( .i (n6524), .o (n6525) );
  buffer buf_n615( .i (N192), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  assign n6526 = n618 & n6521 ;
  buffer buf_n6527( .i (n6526), .o (n6527) );
  assign n6528 = n5080 | n6527 ;
  buffer buf_n6529( .i (n6528), .o (n6529) );
  assign n6530 = n6525 & n6529 ;
  assign n6531 = n6518 | n6530 ;
  buffer buf_n6532( .i (n6531), .o (n6532) );
  assign n6533 = n6513 | n6517 ;
  buffer buf_n6534( .i (n6533), .o (n6534) );
  assign n6536 = n6525 | n6529 ;
  buffer buf_n6537( .i (n6536), .o (n6537) );
  assign n6538 = n6534 & n6537 ;
  assign n6539 = ~n6532 & n6538 ;
  buffer buf_n6540( .i (n6539), .o (n6540) );
  assign n6541 = n6507 & n6540 ;
  buffer buf_n6542( .i (n6541), .o (n6542) );
  buffer buf_n6543( .i (n6542), .o (n6543) );
  buffer buf_n6544( .i (n6543), .o (n6544) );
  buffer buf_n6545( .i (n6544), .o (n6545) );
  buffer buf_n6546( .i (n6545), .o (n6546) );
  buffer buf_n6547( .i (n6546), .o (n6547) );
  assign n6548 = n6475 & n6547 ;
  buffer buf_n6535( .i (n6534), .o (n6535) );
  assign n6549 = n6532 & n6535 ;
  buffer buf_n6550( .i (n6549), .o (n6550) );
  assign n6551 = n6507 & n6550 ;
  buffer buf_n6502( .i (n6501), .o (n6502) );
  assign n6552 = n6487 & n6498 ;
  assign n6553 = n6502 | n6552 ;
  buffer buf_n6554( .i (n6553), .o (n6554) );
  buffer buf_n6555( .i (n6554), .o (n6555) );
  assign n6556 = n6551 | n6555 ;
  buffer buf_n6557( .i (n6556), .o (n6557) );
  buffer buf_n6558( .i (n6557), .o (n6558) );
  buffer buf_n6559( .i (n6558), .o (n6559) );
  buffer buf_n6560( .i (n6559), .o (n6560) );
  buffer buf_n6561( .i (n6560), .o (n6561) );
  buffer buf_n6562( .i (n6561), .o (n6562) );
  assign n6563 = n6548 | n6562 ;
  buffer buf_n6564( .i (n6563), .o (n6564) );
  buffer buf_n3506( .i (N64), .o (n3506) );
  buffer buf_n3507( .i (n3506), .o (n3507) );
  buffer buf_n3508( .i (n3507), .o (n3508) );
  buffer buf_n3509( .i (n3508), .o (n3509) );
  assign n6608 = n3509 & ~n6521 ;
  assign n6609 = ~n1653 & n6521 ;
  assign n6610 = n6608 | n6609 ;
  buffer buf_n6611( .i (n6610), .o (n6611) );
  buffer buf_n574( .i (N177), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n6612( .i (n6520), .o (n6612) );
  assign n6613 = ~n577 & n6612 ;
  assign n6614 = n3882 | n6613 ;
  buffer buf_n6615( .i (n6614), .o (n6615) );
  assign n6617 = n6611 & ~n6615 ;
  buffer buf_n6618( .i (n6617), .o (n6618) );
  buffer buf_n3578( .i (N85), .o (n3578) );
  buffer buf_n3579( .i (n3578), .o (n3579) );
  buffer buf_n3580( .i (n3579), .o (n3580) );
  buffer buf_n3581( .i (n3580), .o (n3581) );
  assign n6619 = n3581 & ~n6612 ;
  assign n6620 = ~n1587 & n6612 ;
  assign n6621 = n6619 | n6620 ;
  buffer buf_n6622( .i (n6621), .o (n6622) );
  buffer buf_n6623( .i (n6622), .o (n6623) );
  buffer buf_n578( .i (N178), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  assign n6624 = n581 & n6612 ;
  buffer buf_n6625( .i (n6624), .o (n6625) );
  assign n6626 = n4590 | n6625 ;
  buffer buf_n6627( .i (n6626), .o (n6627) );
  assign n6628 = n6623 & n6627 ;
  assign n6629 = n6618 | n6628 ;
  buffer buf_n6630( .i (n6629), .o (n6630) );
  assign n6631 = ~n6611 & n6615 ;
  buffer buf_n6632( .i (n6631), .o (n6632) );
  assign n6635 = n6623 | n6627 ;
  assign n6636 = ~n6632 & n6635 ;
  buffer buf_n6637( .i (n6636), .o (n6637) );
  assign n6638 = ~n6630 & n6637 ;
  buffer buf_n6639( .i (n6638), .o (n6639) );
  buffer buf_n3574( .i (N84), .o (n3574) );
  buffer buf_n3575( .i (n3574), .o (n3575) );
  buffer buf_n3576( .i (n3575), .o (n3576) );
  buffer buf_n3577( .i (n3576), .o (n3577) );
  buffer buf_n6640( .i (n6520), .o (n6640) );
  assign n6641 = n3577 & ~n6640 ;
  assign n6642 = ~n1521 & n6640 ;
  assign n6643 = n6641 | n6642 ;
  buffer buf_n6644( .i (n6643), .o (n6644) );
  buffer buf_n6645( .i (n6644), .o (n6645) );
  buffer buf_n582( .i (N179), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  assign n6648 = n585 & n6640 ;
  buffer buf_n6649( .i (n6648), .o (n6649) );
  assign n6650 = n4618 | n6649 ;
  buffer buf_n6651( .i (n6650), .o (n6651) );
  assign n6652 = n6645 & n6651 ;
  buffer buf_n3570( .i (N83), .o (n3570) );
  buffer buf_n3571( .i (n3570), .o (n3571) );
  buffer buf_n3572( .i (n3571), .o (n3572) );
  buffer buf_n3573( .i (n3572), .o (n3573) );
  assign n6653 = n3573 & ~n6640 ;
  buffer buf_n6654( .i (n6520), .o (n6654) );
  assign n6655 = ~n1455 & n6654 ;
  assign n6656 = n6653 | n6655 ;
  buffer buf_n6657( .i (n6656), .o (n6657) );
  buffer buf_n6658( .i (n6657), .o (n6658) );
  buffer buf_n591( .i (N180), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  assign n6661 = n594 & n6654 ;
  buffer buf_n6662( .i (n6661), .o (n6662) );
  assign n6663 = n4637 | n6662 ;
  buffer buf_n6664( .i (n6663), .o (n6664) );
  assign n6665 = n6658 & n6664 ;
  assign n6666 = n6652 | n6665 ;
  buffer buf_n6667( .i (n6666), .o (n6667) );
  assign n6668 = n6645 | n6651 ;
  buffer buf_n6669( .i (n6668), .o (n6669) );
  assign n6671 = n6658 | n6664 ;
  buffer buf_n6672( .i (n6671), .o (n6672) );
  assign n6673 = n6669 & n6672 ;
  assign n6674 = ~n6667 & n6673 ;
  buffer buf_n6675( .i (n6674), .o (n6675) );
  assign n6676 = n6639 & n6675 ;
  buffer buf_n6677( .i (n6676), .o (n6677) );
  buffer buf_n3510( .i (N65), .o (n3510) );
  buffer buf_n3511( .i (n3510), .o (n3511) );
  buffer buf_n3512( .i (n3511), .o (n3512) );
  buffer buf_n3513( .i (n3512), .o (n3513) );
  assign n6678 = n3513 & ~n6654 ;
  assign n6679 = ~n1389 & n6654 ;
  assign n6680 = n6678 | n6679 ;
  buffer buf_n6681( .i (n6680), .o (n6681) );
  buffer buf_n6682( .i (n6681), .o (n6682) );
  buffer buf_n554( .i (N171), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n6683( .i (n6296), .o (n6683) );
  buffer buf_n6684( .i (n6683), .o (n6684) );
  assign n6685 = n557 & n6684 ;
  buffer buf_n6686( .i (n6685), .o (n6686) );
  assign n6687 = n4649 | n6686 ;
  buffer buf_n6688( .i (n6687), .o (n6688) );
  assign n6689 = n6682 & n6688 ;
  buffer buf_n6690( .i (n6689), .o (n6690) );
  assign n6696 = n6682 | n6688 ;
  buffer buf_n6697( .i (n6696), .o (n6697) );
  assign n6698 = ~n6690 & n6697 ;
  buffer buf_n6699( .i (n6698), .o (n6699) );
  buffer buf_n6700( .i (n6699), .o (n6700) );
  buffer buf_n6701( .i (n6700), .o (n6701) );
  buffer buf_n6702( .i (n6701), .o (n6702) );
  assign n6703 = n6677 & n6702 ;
  buffer buf_n6704( .i (n6703), .o (n6704) );
  buffer buf_n6705( .i (n6704), .o (n6705) );
  buffer buf_n6706( .i (n6705), .o (n6706) );
  buffer buf_n6707( .i (n6706), .o (n6707) );
  buffer buf_n6708( .i (n6707), .o (n6708) );
  buffer buf_n6709( .i (n6708), .o (n6709) );
  buffer buf_n6710( .i (n6709), .o (n6710) );
  assign n6711 = n6564 & n6710 ;
  buffer buf_n6691( .i (n6690), .o (n6691) );
  buffer buf_n6692( .i (n6691), .o (n6692) );
  buffer buf_n6693( .i (n6692), .o (n6693) );
  buffer buf_n6694( .i (n6693), .o (n6694) );
  buffer buf_n6695( .i (n6694), .o (n6695) );
  assign n6712 = n6677 & n6695 ;
  buffer buf_n6670( .i (n6669), .o (n6670) );
  assign n6713 = n6667 & n6670 ;
  buffer buf_n6714( .i (n6713), .o (n6714) );
  assign n6715 = n6639 & n6714 ;
  buffer buf_n6633( .i (n6632), .o (n6633) );
  buffer buf_n6634( .i (n6633), .o (n6634) );
  assign n6716 = n6630 & ~n6634 ;
  buffer buf_n6717( .i (n6716), .o (n6717) );
  buffer buf_n6718( .i (n6717), .o (n6718) );
  assign n6719 = n6715 | n6718 ;
  buffer buf_n6720( .i (n6719), .o (n6720) );
  assign n6721 = n6712 | n6720 ;
  buffer buf_n6722( .i (n6721), .o (n6722) );
  buffer buf_n6723( .i (n6722), .o (n6723) );
  buffer buf_n6724( .i (n6723), .o (n6724) );
  buffer buf_n6725( .i (n6724), .o (n6725) );
  buffer buf_n6726( .i (n6725), .o (n6726) );
  buffer buf_n6727( .i (n6726), .o (n6727) );
  buffer buf_n6728( .i (n6727), .o (n6728) );
  assign n6729 = n6711 | n6728 ;
  buffer buf_n348( .i (N109), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  assign n6730 = n351 & ~n6684 ;
  assign n6731 = ~n1855 & n6684 ;
  assign n6732 = n6730 | n6731 ;
  buffer buf_n6733( .i (n6732), .o (n6733) );
  buffer buf_n6734( .i (n6733), .o (n6734) );
  buffer buf_n562( .i (N174), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  assign n6735 = ~n565 & n6684 ;
  buffer buf_n6736( .i (n6735), .o (n6736) );
  assign n6739 = n4557 | n6736 ;
  buffer buf_n6740( .i (n6739), .o (n6740) );
  assign n6741 = n6734 & ~n6740 ;
  buffer buf_n352( .i (N110), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n6742( .i (n6683), .o (n6742) );
  assign n6743 = n355 & ~n6742 ;
  assign n6744 = ~n1921 & n6742 ;
  assign n6745 = n6743 | n6744 ;
  buffer buf_n6746( .i (n6745), .o (n6746) );
  buffer buf_n6747( .i (n6746), .o (n6747) );
  buffer buf_n558( .i (N173), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  assign n6748 = ~n561 & n6742 ;
  buffer buf_n6749( .i (n6748), .o (n6749) );
  assign n6752 = n4557 | n6749 ;
  buffer buf_n6753( .i (n6752), .o (n6753) );
  assign n6754 = n6747 & ~n6753 ;
  assign n6755 = n6741 | n6754 ;
  buffer buf_n6756( .i (n6755), .o (n6756) );
  assign n6757 = ~n6734 & n6740 ;
  buffer buf_n6758( .i (n6757), .o (n6758) );
  assign n6759 = ~n6747 & n6753 ;
  buffer buf_n6760( .i (n6759), .o (n6760) );
  assign n6762 = n6758 | n6760 ;
  assign n6763 = n6756 | n6762 ;
  buffer buf_n6764( .i (n6763), .o (n6764) );
  buffer buf_n3582( .i (N86), .o (n3582) );
  buffer buf_n3583( .i (n3582), .o (n3583) );
  buffer buf_n3584( .i (n3583), .o (n3584) );
  buffer buf_n3585( .i (n3584), .o (n3585) );
  assign n6765 = n3585 & ~n6742 ;
  buffer buf_n6766( .i (n6683), .o (n6766) );
  assign n6767 = ~n1789 & n6766 ;
  assign n6768 = n6765 | n6767 ;
  buffer buf_n6769( .i (n6768), .o (n6769) );
  buffer buf_n6770( .i (n6769), .o (n6770) );
  buffer buf_n566( .i (N175), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  assign n6771 = ~n569 & n6766 ;
  buffer buf_n6772( .i (n6771), .o (n6772) );
  assign n6775 = n4557 | n6772 ;
  buffer buf_n6776( .i (n6775), .o (n6776) );
  assign n6777 = n6770 & ~n6776 ;
  buffer buf_n3502( .i (N63), .o (n3502) );
  buffer buf_n3503( .i (n3502), .o (n3503) );
  buffer buf_n3504( .i (n3503), .o (n3504) );
  buffer buf_n3505( .i (n3504), .o (n3505) );
  assign n6778 = n3505 & ~n6766 ;
  assign n6779 = ~n1723 & n6766 ;
  assign n6780 = n6778 | n6779 ;
  buffer buf_n6781( .i (n6780), .o (n6781) );
  buffer buf_n6782( .i (n6781), .o (n6782) );
  buffer buf_n570( .i (N176), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n6783( .i (n6683), .o (n6783) );
  assign n6784 = ~n573 & n6783 ;
  buffer buf_n6785( .i (n6784), .o (n6785) );
  buffer buf_n6788( .i (n3881), .o (n6788) );
  buffer buf_n6789( .i (n6788), .o (n6789) );
  assign n6790 = n6785 | n6789 ;
  buffer buf_n6791( .i (n6790), .o (n6791) );
  assign n6792 = n6782 & ~n6791 ;
  assign n6793 = n6777 | n6792 ;
  buffer buf_n6794( .i (n6793), .o (n6794) );
  assign n6795 = ~n6770 & n6776 ;
  buffer buf_n6796( .i (n6795), .o (n6796) );
  assign n6798 = ~n6782 & n6791 ;
  buffer buf_n6799( .i (n6798), .o (n6799) );
  assign n6800 = n6796 | n6799 ;
  assign n6801 = n6794 | n6800 ;
  buffer buf_n6802( .i (n6801), .o (n6802) );
  assign n6803 = n6764 | n6802 ;
  buffer buf_n6804( .i (n6803), .o (n6804) );
  buffer buf_n6805( .i (n6804), .o (n6805) );
  buffer buf_n6806( .i (n6805), .o (n6806) );
  buffer buf_n6807( .i (n6806), .o (n6807) );
  buffer buf_n6808( .i (n6807), .o (n6808) );
  buffer buf_n6809( .i (n6808), .o (n6809) );
  buffer buf_n6810( .i (n6809), .o (n6810) );
  buffer buf_n6811( .i (n6810), .o (n6811) );
  buffer buf_n6812( .i (n6811), .o (n6812) );
  buffer buf_n6813( .i (n6812), .o (n6813) );
  buffer buf_n6814( .i (n6813), .o (n6814) );
  assign n6815 = n6729 & ~n6814 ;
  buffer buf_n6797( .i (n6796), .o (n6797) );
  assign n6816 = n6794 & ~n6797 ;
  buffer buf_n6817( .i (n6816), .o (n6817) );
  assign n6818 = ~n6764 & n6817 ;
  buffer buf_n6761( .i (n6760), .o (n6761) );
  assign n6819 = n6756 & ~n6761 ;
  buffer buf_n6820( .i (n6819), .o (n6820) );
  buffer buf_n6821( .i (n6820), .o (n6821) );
  assign n6822 = n6818 | n6821 ;
  buffer buf_n6823( .i (n6822), .o (n6823) );
  buffer buf_n6824( .i (n6823), .o (n6824) );
  buffer buf_n6825( .i (n6824), .o (n6825) );
  buffer buf_n6826( .i (n6825), .o (n6826) );
  buffer buf_n6827( .i (n6826), .o (n6827) );
  buffer buf_n6828( .i (n6827), .o (n6828) );
  buffer buf_n6829( .i (n6828), .o (n6829) );
  buffer buf_n6830( .i (n6829), .o (n6830) );
  buffer buf_n6831( .i (n6830), .o (n6831) );
  buffer buf_n6832( .i (n6831), .o (n6832) );
  buffer buf_n6833( .i (n6832), .o (n6833) );
  assign n6834 = n6815 | n6833 ;
  buffer buf_n3586( .i (N87), .o (n3586) );
  buffer buf_n3587( .i (n3586), .o (n3587) );
  buffer buf_n3588( .i (n3587), .o (n3588) );
  buffer buf_n3589( .i (n3588), .o (n3589) );
  assign n6835 = n3589 & ~n6783 ;
  assign n6836 = ~n285 & n6783 ;
  assign n6837 = n6835 | n6836 ;
  buffer buf_n6838( .i (n6837), .o (n6838) );
  buffer buf_n6839( .i (n6838), .o (n6839) );
  buffer buf_n540( .i (N168), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  assign n6840 = ~n543 & n6783 ;
  buffer buf_n6841( .i (n6840), .o (n6841) );
  assign n6844 = n6789 | n6841 ;
  buffer buf_n6845( .i (n6844), .o (n6845) );
  assign n6846 = ~n6839 & n6845 ;
  buffer buf_n6847( .i (n6846), .o (n6847) );
  buffer buf_n6848( .i (n6847), .o (n6848) );
  buffer buf_n6849( .i (n6848), .o (n6849) );
  buffer buf_n3590( .i (N88), .o (n3590) );
  buffer buf_n3591( .i (n3590), .o (n3591) );
  buffer buf_n3592( .i (n3591), .o (n3592) );
  buffer buf_n3593( .i (n3592), .o (n3593) );
  buffer buf_n6850( .i (n586), .o (n6850) );
  buffer buf_n6851( .i (n6850), .o (n6851) );
  buffer buf_n6852( .i (n6851), .o (n6852) );
  assign n6853 = n3593 & ~n6852 ;
  assign n6854 = ~n1124 & n6852 ;
  assign n6855 = n6853 | n6854 ;
  buffer buf_n6856( .i (n6855), .o (n6856) );
  buffer buf_n6857( .i (n6856), .o (n6857) );
  buffer buf_n532( .i (N166), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  assign n6858 = ~n535 & n6852 ;
  buffer buf_n6859( .i (n6858), .o (n6859) );
  assign n6862 = n6789 | n6859 ;
  buffer buf_n6863( .i (n6862), .o (n6863) );
  assign n6864 = ~n6857 & n6863 ;
  buffer buf_n6865( .i (n6864), .o (n6865) );
  assign n6867 = n6857 & ~n6863 ;
  buffer buf_n6868( .i (n6867), .o (n6868) );
  assign n6869 = n6865 | n6868 ;
  buffer buf_n360( .i (N112), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  assign n6870 = n363 & ~n6852 ;
  buffer buf_n6871( .i (n6851), .o (n6871) );
  assign n6872 = ~n1054 & n6871 ;
  assign n6873 = n6870 | n6872 ;
  buffer buf_n6874( .i (n6873), .o (n6874) );
  buffer buf_n6875( .i (n6874), .o (n6875) );
  buffer buf_n536( .i (N167), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  assign n6876 = ~n539 & n6871 ;
  buffer buf_n6877( .i (n6876), .o (n6877) );
  assign n6880 = n6789 | n6877 ;
  buffer buf_n6881( .i (n6880), .o (n6881) );
  assign n6882 = n6875 & ~n6881 ;
  buffer buf_n6883( .i (n6882), .o (n6883) );
  assign n6884 = ~n6875 & n6881 ;
  buffer buf_n6885( .i (n6884), .o (n6885) );
  assign n6886 = n6883 | n6885 ;
  assign n6887 = n6869 | n6886 ;
  assign n6888 = n6849 | n6887 ;
  buffer buf_n6889( .i (n6888), .o (n6889) );
  buffer buf_n364( .i (N113), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  assign n6890 = n367 & ~n6871 ;
  assign n6891 = ~n922 & n6871 ;
  assign n6892 = n6890 | n6891 ;
  buffer buf_n6893( .i (n6892), .o (n6893) );
  assign n6894 = ~n3884 & n6893 ;
  buffer buf_n6895( .i (n6894), .o (n6895) );
  buffer buf_n356( .i (N111), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n6896( .i (n6851), .o (n6896) );
  assign n6897 = n359 & ~n6896 ;
  assign n6898 = ~n988 & n6896 ;
  assign n6899 = n6897 | n6898 ;
  buffer buf_n6900( .i (n6899), .o (n6900) );
  buffer buf_n6901( .i (n6900), .o (n6901) );
  buffer buf_n544( .i (N169), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  assign n6902 = ~n547 & n6896 ;
  buffer buf_n6903( .i (n6902), .o (n6903) );
  buffer buf_n6906( .i (n6788), .o (n6906) );
  assign n6907 = n6903 | n6906 ;
  buffer buf_n6908( .i (n6907), .o (n6908) );
  assign n6909 = n6901 & ~n6908 ;
  assign n6910 = n6895 | n6909 ;
  buffer buf_n6911( .i (n6910), .o (n6911) );
  buffer buf_n6912( .i (n6911), .o (n6912) );
  assign n6913 = n3884 & ~n6893 ;
  buffer buf_n6914( .i (n6913), .o (n6914) );
  buffer buf_n6915( .i (n6914), .o (n6915) );
  buffer buf_n6916( .i (n6915), .o (n6916) );
  assign n6917 = n6839 & ~n6845 ;
  buffer buf_n6918( .i (n6917), .o (n6918) );
  assign n6921 = ~n6901 & n6908 ;
  buffer buf_n6922( .i (n6921), .o (n6922) );
  assign n6924 = n6918 | n6922 ;
  assign n6925 = n6916 | n6924 ;
  assign n6926 = n6912 | n6925 ;
  buffer buf_n6927( .i (n6926), .o (n6927) );
  assign n6928 = n6889 | n6927 ;
  buffer buf_n6929( .i (n6928), .o (n6929) );
  buffer buf_n6930( .i (n6929), .o (n6930) );
  buffer buf_n6931( .i (n6930), .o (n6931) );
  buffer buf_n6932( .i (n6931), .o (n6932) );
  buffer buf_n6933( .i (n6932), .o (n6933) );
  buffer buf_n6934( .i (n6933), .o (n6934) );
  buffer buf_n6935( .i (n6934), .o (n6935) );
  buffer buf_n6936( .i (n6935), .o (n6936) );
  buffer buf_n6937( .i (n6936), .o (n6937) );
  buffer buf_n6938( .i (n6937), .o (n6938) );
  buffer buf_n6939( .i (n6938), .o (n6939) );
  buffer buf_n6940( .i (n6939), .o (n6940) );
  assign n6941 = n6834 & ~n6940 ;
  buffer buf_n6919( .i (n6918), .o (n6919) );
  buffer buf_n6920( .i (n6919), .o (n6920) );
  buffer buf_n6923( .i (n6922), .o (n6923) );
  assign n6942 = n6911 & ~n6923 ;
  assign n6943 = n6920 | n6942 ;
  buffer buf_n6944( .i (n6943), .o (n6944) );
  assign n6945 = ~n6889 & n6944 ;
  assign n6946 = n852 | n1319 ;
  buffer buf_n6947( .i (n6946), .o (n6947) );
  assign n6949 = n3395 & ~n6947 ;
  assign n6950 = n3340 & ~n6949 ;
  buffer buf_n6951( .i (n6950), .o (n6951) );
  buffer buf_n6952( .i (n6951), .o (n6952) );
  buffer buf_n6953( .i (n6952), .o (n6953) );
  buffer buf_n6954( .i (n6953), .o (n6954) );
  buffer buf_n6955( .i (n6954), .o (n6955) );
  buffer buf_n6956( .i (n6955), .o (n6956) );
  buffer buf_n6957( .i (n6956), .o (n6957) );
  buffer buf_n6866( .i (n6865), .o (n6866) );
  assign n6958 = n6868 | n6883 ;
  assign n6959 = ~n6866 & n6958 ;
  assign n6960 = n6957 | n6959 ;
  buffer buf_n6961( .i (n6960), .o (n6961) );
  buffer buf_n6962( .i (n6961), .o (n6962) );
  assign n6963 = n6945 | n6962 ;
  buffer buf_n6964( .i (n6963), .o (n6964) );
  buffer buf_n6965( .i (n6964), .o (n6965) );
  buffer buf_n6966( .i (n6965), .o (n6966) );
  buffer buf_n6967( .i (n6966), .o (n6967) );
  buffer buf_n6968( .i (n6967), .o (n6968) );
  buffer buf_n6969( .i (n6968), .o (n6969) );
  buffer buf_n6970( .i (n6969), .o (n6970) );
  buffer buf_n6971( .i (n6970), .o (n6971) );
  buffer buf_n6972( .i (n6971), .o (n6972) );
  buffer buf_n6973( .i (n6972), .o (n6973) );
  buffer buf_n6974( .i (n6973), .o (n6974) );
  buffer buf_n6975( .i (n6974), .o (n6975) );
  assign n6976 = n6941 | n6975 ;
  assign n6977 = ~n6225 & n6976 ;
  buffer buf_n6978( .i (n6977), .o (n6978) );
  buffer buf_n6979( .i (n6978), .o (n6979) );
  buffer buf_n6980( .i (n6979), .o (n6980) );
  buffer buf_n6981( .i (n6980), .o (n6981) );
  buffer buf_n6982( .i (n6981), .o (n6982) );
  buffer buf_n6983( .i (n6982), .o (n6983) );
  buffer buf_n6984( .i (n6983), .o (n6984) );
  buffer buf_n6985( .i (n6984), .o (n6985) );
  buffer buf_n6986( .i (n6985), .o (n6986) );
  buffer buf_n6987( .i (n6986), .o (n6987) );
  buffer buf_n6988( .i (n6987), .o (n6988) );
  buffer buf_n6989( .i (n6988), .o (n6989) );
  buffer buf_n6990( .i (n6989), .o (n6990) );
  buffer buf_n6991( .i (n6990), .o (n6991) );
  buffer buf_n6992( .i (n6991), .o (n6992) );
  buffer buf_n6993( .i (n6992), .o (n6993) );
  buffer buf_n6994( .i (n6993), .o (n6994) );
  buffer buf_n6995( .i (n6994), .o (n6995) );
  buffer buf_n6996( .i (n6995), .o (n6996) );
  buffer buf_n6997( .i (n6996), .o (n6997) );
  buffer buf_n6998( .i (n6997), .o (n6998) );
  buffer buf_n6999( .i (n6998), .o (n6999) );
  buffer buf_n7000( .i (n6999), .o (n7000) );
  buffer buf_n7001( .i (n7000), .o (n7001) );
  buffer buf_n7002( .i (n7001), .o (n7002) );
  buffer buf_n7003( .i (n7002), .o (n7003) );
  buffer buf_n7004( .i (n7003), .o (n7004) );
  buffer buf_n7005( .i (n7004), .o (n7005) );
  buffer buf_n7006( .i (n7005), .o (n7006) );
  buffer buf_n7007( .i (n7006), .o (n7007) );
  buffer buf_n7008( .i (n7007), .o (n7008) );
  buffer buf_n7009( .i (n7008), .o (n7009) );
  buffer buf_n7010( .i (n7009), .o (n7010) );
  buffer buf_n7011( .i (n7010), .o (n7011) );
  buffer buf_n7012( .i (n7011), .o (n7012) );
  buffer buf_n7013( .i (n7012), .o (n7013) );
  assign n7014 = n5637 | n5651 ;
  buffer buf_n7015( .i (n7014), .o (n7015) );
  buffer buf_n7016( .i (n7015), .o (n7016) );
  buffer buf_n7017( .i (n7016), .o (n7017) );
  buffer buf_n7018( .i (n7017), .o (n7018) );
  buffer buf_n7019( .i (n7018), .o (n7019) );
  buffer buf_n7020( .i (n7019), .o (n7020) );
  buffer buf_n7021( .i (n7020), .o (n7021) );
  buffer buf_n7022( .i (n7021), .o (n7022) );
  buffer buf_n7023( .i (n7022), .o (n7023) );
  buffer buf_n7024( .i (n7023), .o (n7024) );
  buffer buf_n5678( .i (n5677), .o (n5678) );
  buffer buf_n5679( .i (n5678), .o (n5679) );
  buffer buf_n5729( .i (n5728), .o (n5729) );
  assign n7025 = n3327 & ~n5749 ;
  buffer buf_n7026( .i (n7025), .o (n7026) );
  assign n7027 = n5729 | n7026 ;
  assign n7028 = ~n5679 & n7027 ;
  buffer buf_n7029( .i (n7028), .o (n7029) );
  assign n7030 = ~n7024 & n7029 ;
  assign n7031 = n7024 & ~n7029 ;
  assign n7032 = n7030 | n7031 ;
  buffer buf_n7033( .i (n7032), .o (n7033) );
  buffer buf_n7034( .i (n7033), .o (n7034) );
  buffer buf_n7035( .i (n7034), .o (n7035) );
  buffer buf_n7036( .i (n7035), .o (n7036) );
  buffer buf_n7037( .i (n7036), .o (n7037) );
  buffer buf_n7038( .i (n7037), .o (n7038) );
  buffer buf_n7039( .i (n7038), .o (n7039) );
  buffer buf_n7040( .i (n7039), .o (n7040) );
  buffer buf_n7041( .i (n7040), .o (n7041) );
  buffer buf_n7042( .i (n7041), .o (n7042) );
  buffer buf_n7043( .i (n7042), .o (n7043) );
  buffer buf_n7044( .i (n7043), .o (n7044) );
  buffer buf_n7045( .i (n7044), .o (n7045) );
  buffer buf_n7046( .i (n7045), .o (n7046) );
  buffer buf_n7047( .i (n7046), .o (n7047) );
  buffer buf_n7048( .i (n7047), .o (n7048) );
  buffer buf_n7049( .i (n7048), .o (n7049) );
  buffer buf_n7050( .i (n7049), .o (n7050) );
  buffer buf_n7051( .i (n7050), .o (n7051) );
  buffer buf_n7052( .i (n7051), .o (n7052) );
  buffer buf_n7053( .i (n7052), .o (n7053) );
  buffer buf_n7054( .i (n7053), .o (n7054) );
  buffer buf_n7055( .i (n7054), .o (n7055) );
  buffer buf_n7056( .i (n7055), .o (n7056) );
  buffer buf_n7057( .i (n7056), .o (n7057) );
  buffer buf_n7058( .i (n7057), .o (n7058) );
  buffer buf_n7059( .i (n7058), .o (n7059) );
  buffer buf_n7060( .i (n7059), .o (n7060) );
  buffer buf_n7061( .i (n7060), .o (n7061) );
  buffer buf_n7062( .i (n7061), .o (n7062) );
  buffer buf_n7063( .i (n7062), .o (n7063) );
  buffer buf_n7064( .i (n7063), .o (n7064) );
  buffer buf_n7065( .i (n7064), .o (n7065) );
  buffer buf_n7066( .i (n7065), .o (n7066) );
  buffer buf_n7067( .i (n7066), .o (n7067) );
  buffer buf_n7068( .i (n7067), .o (n7068) );
  buffer buf_n7069( .i (n7068), .o (n7069) );
  buffer buf_n7070( .i (n7069), .o (n7070) );
  buffer buf_n7071( .i (n7070), .o (n7071) );
  buffer buf_n7072( .i (n7071), .o (n7072) );
  buffer buf_n7073( .i (n7072), .o (n7073) );
  buffer buf_n7074( .i (n7073), .o (n7074) );
  buffer buf_n7075( .i (n7074), .o (n7075) );
  buffer buf_n5756( .i (n5755), .o (n5756) );
  buffer buf_n5757( .i (n5756), .o (n5757) );
  buffer buf_n5758( .i (n5757), .o (n5758) );
  buffer buf_n5759( .i (n5758), .o (n5759) );
  buffer buf_n5724( .i (n5723), .o (n5724) );
  buffer buf_n5725( .i (n5724), .o (n5725) );
  buffer buf_n5726( .i (n5725), .o (n5726) );
  assign n7076 = n5726 | n7026 ;
  buffer buf_n7077( .i (n7076), .o (n7077) );
  assign n7078 = n5759 & n7077 ;
  assign n7079 = n5759 | n7077 ;
  assign n7080 = ~n7078 & n7079 ;
  buffer buf_n7081( .i (n7080), .o (n7081) );
  buffer buf_n7082( .i (n7081), .o (n7082) );
  buffer buf_n7083( .i (n7082), .o (n7083) );
  buffer buf_n7084( .i (n7083), .o (n7084) );
  buffer buf_n7085( .i (n7084), .o (n7085) );
  buffer buf_n7086( .i (n7085), .o (n7086) );
  buffer buf_n7087( .i (n7086), .o (n7087) );
  buffer buf_n7088( .i (n7087), .o (n7088) );
  buffer buf_n7089( .i (n7088), .o (n7089) );
  buffer buf_n7090( .i (n7089), .o (n7090) );
  buffer buf_n7091( .i (n7090), .o (n7091) );
  buffer buf_n7092( .i (n7091), .o (n7092) );
  buffer buf_n7093( .i (n7092), .o (n7093) );
  buffer buf_n7094( .i (n7093), .o (n7094) );
  buffer buf_n7095( .i (n7094), .o (n7095) );
  buffer buf_n7096( .i (n7095), .o (n7096) );
  buffer buf_n7097( .i (n7096), .o (n7097) );
  buffer buf_n7098( .i (n7097), .o (n7098) );
  buffer buf_n7099( .i (n7098), .o (n7099) );
  buffer buf_n7100( .i (n7099), .o (n7100) );
  buffer buf_n7101( .i (n7100), .o (n7101) );
  buffer buf_n7102( .i (n7101), .o (n7102) );
  buffer buf_n7103( .i (n7102), .o (n7103) );
  buffer buf_n7104( .i (n7103), .o (n7104) );
  buffer buf_n7105( .i (n7104), .o (n7105) );
  buffer buf_n7106( .i (n7105), .o (n7106) );
  buffer buf_n7107( .i (n7106), .o (n7107) );
  buffer buf_n7108( .i (n7107), .o (n7108) );
  buffer buf_n7109( .i (n7108), .o (n7109) );
  buffer buf_n7110( .i (n7109), .o (n7110) );
  buffer buf_n7111( .i (n7110), .o (n7111) );
  buffer buf_n7112( .i (n7111), .o (n7112) );
  buffer buf_n7113( .i (n7112), .o (n7113) );
  buffer buf_n7114( .i (n7113), .o (n7114) );
  buffer buf_n7115( .i (n7114), .o (n7115) );
  buffer buf_n7116( .i (n7115), .o (n7116) );
  buffer buf_n7117( .i (n7116), .o (n7117) );
  buffer buf_n7118( .i (n7117), .o (n7118) );
  buffer buf_n7119( .i (n7118), .o (n7119) );
  buffer buf_n7120( .i (n7119), .o (n7120) );
  buffer buf_n7121( .i (n7120), .o (n7121) );
  buffer buf_n7122( .i (n7121), .o (n7122) );
  buffer buf_n7123( .i (n7122), .o (n7123) );
  buffer buf_n7124( .i (n7123), .o (n7124) );
  buffer buf_n5741( .i (n5740), .o (n5741) );
  buffer buf_n5708( .i (n5707), .o (n5708) );
  buffer buf_n5709( .i (n5708), .o (n5709) );
  buffer buf_n5710( .i (n5709), .o (n5710) );
  assign n7125 = n3613 | n5716 ;
  buffer buf_n7126( .i (n7125), .o (n7126) );
  assign n7127 = n3630 | n7126 ;
  assign n7128 = ~n5710 & n7127 ;
  buffer buf_n7129( .i (n7128), .o (n7129) );
  assign n7130 = n5741 & n7129 ;
  assign n7131 = n5741 | n7129 ;
  assign n7132 = ~n7130 & n7131 ;
  buffer buf_n7133( .i (n7132), .o (n7133) );
  buffer buf_n7134( .i (n7133), .o (n7134) );
  buffer buf_n7135( .i (n7134), .o (n7135) );
  buffer buf_n7136( .i (n7135), .o (n7136) );
  buffer buf_n7137( .i (n7136), .o (n7137) );
  buffer buf_n7138( .i (n7137), .o (n7138) );
  buffer buf_n7139( .i (n7138), .o (n7139) );
  buffer buf_n7140( .i (n7139), .o (n7140) );
  buffer buf_n7141( .i (n7140), .o (n7141) );
  buffer buf_n7142( .i (n7141), .o (n7142) );
  buffer buf_n7143( .i (n7142), .o (n7143) );
  buffer buf_n7144( .i (n7143), .o (n7144) );
  buffer buf_n7145( .i (n7144), .o (n7145) );
  buffer buf_n7146( .i (n7145), .o (n7146) );
  buffer buf_n7147( .i (n7146), .o (n7147) );
  buffer buf_n7148( .i (n7147), .o (n7148) );
  buffer buf_n7149( .i (n7148), .o (n7149) );
  buffer buf_n7150( .i (n7149), .o (n7150) );
  buffer buf_n7151( .i (n7150), .o (n7151) );
  buffer buf_n7152( .i (n7151), .o (n7152) );
  buffer buf_n7153( .i (n7152), .o (n7153) );
  buffer buf_n7154( .i (n7153), .o (n7154) );
  buffer buf_n7155( .i (n7154), .o (n7155) );
  buffer buf_n7156( .i (n7155), .o (n7156) );
  buffer buf_n7157( .i (n7156), .o (n7157) );
  buffer buf_n7158( .i (n7157), .o (n7158) );
  buffer buf_n7159( .i (n7158), .o (n7159) );
  buffer buf_n7160( .i (n7159), .o (n7160) );
  buffer buf_n7161( .i (n7160), .o (n7161) );
  buffer buf_n7162( .i (n7161), .o (n7162) );
  buffer buf_n7163( .i (n7162), .o (n7163) );
  buffer buf_n7164( .i (n7163), .o (n7164) );
  buffer buf_n7165( .i (n7164), .o (n7165) );
  buffer buf_n7166( .i (n7165), .o (n7166) );
  buffer buf_n7167( .i (n7166), .o (n7167) );
  buffer buf_n7168( .i (n7167), .o (n7168) );
  buffer buf_n7169( .i (n7168), .o (n7169) );
  buffer buf_n7170( .i (n7169), .o (n7170) );
  buffer buf_n7171( .i (n7170), .o (n7171) );
  buffer buf_n7172( .i (n7171), .o (n7172) );
  buffer buf_n7173( .i (n7172), .o (n7173) );
  buffer buf_n7174( .i (n7173), .o (n7174) );
  buffer buf_n7175( .i (n7174), .o (n7175) );
  buffer buf_n7176( .i (n7175), .o (n7176) );
  buffer buf_n7177( .i (n7176), .o (n7177) );
  buffer buf_n7178( .i (n7177), .o (n7178) );
  buffer buf_n7179( .i (n7178), .o (n7179) );
  buffer buf_n7180( .i (n7179), .o (n7180) );
  buffer buf_n7181( .i (n7180), .o (n7181) );
  buffer buf_n5744( .i (n5743), .o (n5744) );
  buffer buf_n5745( .i (n5744), .o (n5745) );
  buffer buf_n3614( .i (n3613), .o (n3614) );
  buffer buf_n3615( .i (n3614), .o (n3615) );
  assign n7182 = n3615 | n3630 ;
  buffer buf_n7183( .i (n7182), .o (n7183) );
  assign n7184 = n5745 | n7183 ;
  assign n7185 = n5745 & n7183 ;
  assign n7186 = n7184 & ~n7185 ;
  buffer buf_n7187( .i (n7186), .o (n7187) );
  buffer buf_n7188( .i (n7187), .o (n7188) );
  buffer buf_n7189( .i (n7188), .o (n7189) );
  buffer buf_n7190( .i (n7189), .o (n7190) );
  buffer buf_n7191( .i (n7190), .o (n7191) );
  buffer buf_n7192( .i (n7191), .o (n7192) );
  buffer buf_n7193( .i (n7192), .o (n7193) );
  buffer buf_n7194( .i (n7193), .o (n7194) );
  buffer buf_n7195( .i (n7194), .o (n7195) );
  buffer buf_n7196( .i (n7195), .o (n7196) );
  buffer buf_n7197( .i (n7196), .o (n7197) );
  buffer buf_n7198( .i (n7197), .o (n7198) );
  buffer buf_n7199( .i (n7198), .o (n7199) );
  buffer buf_n7200( .i (n7199), .o (n7200) );
  buffer buf_n7201( .i (n7200), .o (n7201) );
  buffer buf_n7202( .i (n7201), .o (n7202) );
  buffer buf_n7203( .i (n7202), .o (n7203) );
  buffer buf_n7204( .i (n7203), .o (n7204) );
  buffer buf_n7205( .i (n7204), .o (n7205) );
  buffer buf_n7206( .i (n7205), .o (n7206) );
  buffer buf_n7207( .i (n7206), .o (n7207) );
  buffer buf_n7208( .i (n7207), .o (n7208) );
  buffer buf_n7209( .i (n7208), .o (n7209) );
  buffer buf_n7210( .i (n7209), .o (n7210) );
  buffer buf_n7211( .i (n7210), .o (n7211) );
  buffer buf_n7212( .i (n7211), .o (n7212) );
  buffer buf_n7213( .i (n7212), .o (n7213) );
  buffer buf_n7214( .i (n7213), .o (n7214) );
  buffer buf_n7215( .i (n7214), .o (n7215) );
  buffer buf_n7216( .i (n7215), .o (n7216) );
  buffer buf_n7217( .i (n7216), .o (n7217) );
  buffer buf_n7218( .i (n7217), .o (n7218) );
  buffer buf_n7219( .i (n7218), .o (n7219) );
  buffer buf_n7220( .i (n7219), .o (n7220) );
  buffer buf_n7221( .i (n7220), .o (n7221) );
  buffer buf_n7222( .i (n7221), .o (n7222) );
  buffer buf_n7223( .i (n7222), .o (n7223) );
  buffer buf_n7224( .i (n7223), .o (n7224) );
  buffer buf_n7225( .i (n7224), .o (n7225) );
  buffer buf_n7226( .i (n7225), .o (n7226) );
  buffer buf_n7227( .i (n7226), .o (n7227) );
  buffer buf_n7228( .i (n7227), .o (n7228) );
  buffer buf_n7229( .i (n7228), .o (n7229) );
  buffer buf_n7230( .i (n7229), .o (n7230) );
  buffer buf_n7231( .i (n7230), .o (n7231) );
  buffer buf_n7232( .i (n7231), .o (n7232) );
  buffer buf_n7233( .i (n7232), .o (n7233) );
  buffer buf_n7234( .i (n7233), .o (n7234) );
  buffer buf_n7235( .i (n7234), .o (n7235) );
  buffer buf_n7236( .i (n7235), .o (n7236) );
  buffer buf_n5851( .i (n5850), .o (n5851) );
  buffer buf_n5852( .i (n5851), .o (n5852) );
  buffer buf_n5853( .i (n5852), .o (n5853) );
  buffer buf_n5854( .i (n5853), .o (n5854) );
  buffer buf_n5855( .i (n5854), .o (n5855) );
  buffer buf_n5856( .i (n5855), .o (n5856) );
  buffer buf_n5857( .i (n5856), .o (n5857) );
  buffer buf_n5858( .i (n5857), .o (n5858) );
  buffer buf_n5859( .i (n5858), .o (n5859) );
  buffer buf_n5860( .i (n5859), .o (n5860) );
  buffer buf_n5861( .i (n5860), .o (n5861) );
  buffer buf_n5862( .i (n5861), .o (n5862) );
  buffer buf_n5863( .i (n5862), .o (n5863) );
  buffer buf_n5864( .i (n5863), .o (n5864) );
  buffer buf_n5865( .i (n5864), .o (n5865) );
  buffer buf_n5866( .i (n5865), .o (n5866) );
  buffer buf_n5607( .i (n5606), .o (n5607) );
  buffer buf_n5608( .i (n5607), .o (n5608) );
  buffer buf_n5609( .i (n5608), .o (n5609) );
  buffer buf_n5610( .i (n5609), .o (n5610) );
  buffer buf_n5611( .i (n5610), .o (n5611) );
  buffer buf_n5612( .i (n5611), .o (n5612) );
  buffer buf_n5613( .i (n5612), .o (n5613) );
  buffer buf_n5614( .i (n5613), .o (n5614) );
  buffer buf_n5615( .i (n5614), .o (n5615) );
  buffer buf_n5616( .i (n5615), .o (n5616) );
  buffer buf_n5617( .i (n5616), .o (n5617) );
  buffer buf_n5830( .i (n5829), .o (n5830) );
  buffer buf_n5831( .i (n5830), .o (n5831) );
  assign n7237 = n5826 | n5831 ;
  buffer buf_n7238( .i (n7237), .o (n7238) );
  buffer buf_n7239( .i (n7238), .o (n7239) );
  buffer buf_n7240( .i (n7239), .o (n7240) );
  buffer buf_n7241( .i (n7240), .o (n7241) );
  buffer buf_n7242( .i (n7241), .o (n7242) );
  buffer buf_n7243( .i (n7242), .o (n7243) );
  buffer buf_n7244( .i (n7243), .o (n7244) );
  buffer buf_n7245( .i (n7244), .o (n7245) );
  buffer buf_n7246( .i (n7245), .o (n7246) );
  buffer buf_n7247( .i (n7246), .o (n7247) );
  assign n7248 = n5769 & ~n7247 ;
  assign n7249 = n5617 | n7248 ;
  buffer buf_n7250( .i (n7249), .o (n7250) );
  assign n7251 = n5866 | n7250 ;
  assign n7252 = n5866 & n7250 ;
  assign n7253 = n7251 & ~n7252 ;
  buffer buf_n7254( .i (n7253), .o (n7254) );
  buffer buf_n7255( .i (n7254), .o (n7255) );
  buffer buf_n7256( .i (n7255), .o (n7256) );
  buffer buf_n7257( .i (n7256), .o (n7257) );
  buffer buf_n7258( .i (n7257), .o (n7258) );
  buffer buf_n7259( .i (n7258), .o (n7259) );
  buffer buf_n7260( .i (n7259), .o (n7260) );
  buffer buf_n7261( .i (n7260), .o (n7261) );
  buffer buf_n7262( .i (n7261), .o (n7262) );
  buffer buf_n7263( .i (n7262), .o (n7263) );
  buffer buf_n7264( .i (n7263), .o (n7264) );
  buffer buf_n7265( .i (n7264), .o (n7265) );
  buffer buf_n7266( .i (n7265), .o (n7266) );
  buffer buf_n7267( .i (n7266), .o (n7267) );
  buffer buf_n7268( .i (n7267), .o (n7268) );
  buffer buf_n7269( .i (n7268), .o (n7269) );
  buffer buf_n7270( .i (n7269), .o (n7270) );
  buffer buf_n7271( .i (n7270), .o (n7271) );
  buffer buf_n7272( .i (n7271), .o (n7272) );
  buffer buf_n7273( .i (n7272), .o (n7273) );
  buffer buf_n7274( .i (n7273), .o (n7274) );
  buffer buf_n7275( .i (n7274), .o (n7275) );
  buffer buf_n7276( .i (n7275), .o (n7276) );
  buffer buf_n7277( .i (n7276), .o (n7277) );
  buffer buf_n7278( .i (n7277), .o (n7278) );
  buffer buf_n7279( .i (n7278), .o (n7279) );
  buffer buf_n7280( .i (n7279), .o (n7280) );
  buffer buf_n7281( .i (n7280), .o (n7281) );
  buffer buf_n7282( .i (n7281), .o (n7282) );
  buffer buf_n7283( .i (n7282), .o (n7283) );
  buffer buf_n7284( .i (n7283), .o (n7284) );
  buffer buf_n7285( .i (n7284), .o (n7285) );
  buffer buf_n7286( .i (n7285), .o (n7286) );
  buffer buf_n7287( .i (n7286), .o (n7287) );
  buffer buf_n7288( .i (n7287), .o (n7288) );
  buffer buf_n5832( .i (n5831), .o (n5832) );
  buffer buf_n5833( .i (n5832), .o (n5833) );
  buffer buf_n5834( .i (n5833), .o (n5834) );
  buffer buf_n5835( .i (n5834), .o (n5835) );
  buffer buf_n5836( .i (n5835), .o (n5836) );
  buffer buf_n5837( .i (n5836), .o (n5837) );
  buffer buf_n5838( .i (n5837), .o (n5838) );
  buffer buf_n5839( .i (n5838), .o (n5839) );
  buffer buf_n5840( .i (n5839), .o (n5840) );
  buffer buf_n5841( .i (n5840), .o (n5841) );
  buffer buf_n5842( .i (n5841), .o (n5842) );
  buffer buf_n5843( .i (n5842), .o (n5843) );
  buffer buf_n5844( .i (n5843), .o (n5844) );
  buffer buf_n5845( .i (n5844), .o (n5845) );
  buffer buf_n5846( .i (n5845), .o (n5846) );
  buffer buf_n5847( .i (n5846), .o (n5847) );
  buffer buf_n5588( .i (n5587), .o (n5588) );
  buffer buf_n5589( .i (n5588), .o (n5589) );
  buffer buf_n5590( .i (n5589), .o (n5590) );
  buffer buf_n5591( .i (n5590), .o (n5591) );
  buffer buf_n5592( .i (n5591), .o (n5592) );
  buffer buf_n5593( .i (n5592), .o (n5593) );
  buffer buf_n5594( .i (n5593), .o (n5594) );
  buffer buf_n5595( .i (n5594), .o (n5595) );
  buffer buf_n5596( .i (n5595), .o (n5596) );
  buffer buf_n5597( .i (n5596), .o (n5597) );
  buffer buf_n5598( .i (n5597), .o (n5598) );
  buffer buf_n5599( .i (n5598), .o (n5599) );
  buffer buf_n5600( .i (n5599), .o (n5600) );
  buffer buf_n5601( .i (n5600), .o (n5601) );
  buffer buf_n5602( .i (n5601), .o (n5602) );
  buffer buf_n5603( .i (n5602), .o (n5603) );
  buffer buf_n5774( .i (n5773), .o (n5774) );
  buffer buf_n5775( .i (n5774), .o (n5775) );
  buffer buf_n5776( .i (n5775), .o (n5776) );
  buffer buf_n5777( .i (n5776), .o (n5777) );
  buffer buf_n5778( .i (n5777), .o (n5778) );
  buffer buf_n5779( .i (n5778), .o (n5779) );
  buffer buf_n5780( .i (n5779), .o (n5780) );
  buffer buf_n5781( .i (n5780), .o (n5781) );
  buffer buf_n5782( .i (n5781), .o (n5782) );
  buffer buf_n5783( .i (n5782), .o (n5783) );
  buffer buf_n5784( .i (n5783), .o (n5784) );
  buffer buf_n5785( .i (n5784), .o (n5785) );
  buffer buf_n5786( .i (n5785), .o (n5786) );
  buffer buf_n5787( .i (n5786), .o (n5787) );
  buffer buf_n5788( .i (n5787), .o (n5788) );
  buffer buf_n5794( .i (n5793), .o (n5794) );
  buffer buf_n5795( .i (n5794), .o (n5795) );
  buffer buf_n5796( .i (n5795), .o (n5796) );
  buffer buf_n5797( .i (n5796), .o (n5797) );
  buffer buf_n5798( .i (n5797), .o (n5798) );
  buffer buf_n5799( .i (n5798), .o (n5799) );
  buffer buf_n5800( .i (n5799), .o (n5800) );
  buffer buf_n5801( .i (n5800), .o (n5801) );
  buffer buf_n5802( .i (n5801), .o (n5802) );
  buffer buf_n5803( .i (n5802), .o (n5803) );
  buffer buf_n5804( .i (n5803), .o (n5804) );
  buffer buf_n5805( .i (n5804), .o (n5805) );
  buffer buf_n5806( .i (n5805), .o (n5806) );
  buffer buf_n5807( .i (n5806), .o (n5807) );
  buffer buf_n5808( .i (n5807), .o (n5808) );
  assign n7289 = n5769 & ~n5808 ;
  buffer buf_n7290( .i (n7289), .o (n7290) );
  assign n7291 = ~n5788 & n7290 ;
  assign n7292 = n5603 | n7291 ;
  buffer buf_n7293( .i (n7292), .o (n7293) );
  assign n7294 = n5847 | n7293 ;
  assign n7295 = n5847 & n7293 ;
  assign n7296 = n7294 & ~n7295 ;
  buffer buf_n7297( .i (n7296), .o (n7297) );
  buffer buf_n7298( .i (n7297), .o (n7298) );
  buffer buf_n7299( .i (n7298), .o (n7299) );
  buffer buf_n7300( .i (n7299), .o (n7300) );
  buffer buf_n7301( .i (n7300), .o (n7301) );
  buffer buf_n7302( .i (n7301), .o (n7302) );
  buffer buf_n7303( .i (n7302), .o (n7303) );
  buffer buf_n7304( .i (n7303), .o (n7304) );
  buffer buf_n7305( .i (n7304), .o (n7305) );
  buffer buf_n7306( .i (n7305), .o (n7306) );
  buffer buf_n7307( .i (n7306), .o (n7307) );
  buffer buf_n7308( .i (n7307), .o (n7308) );
  buffer buf_n7309( .i (n7308), .o (n7309) );
  buffer buf_n7310( .i (n7309), .o (n7310) );
  buffer buf_n7311( .i (n7310), .o (n7311) );
  buffer buf_n7312( .i (n7311), .o (n7312) );
  buffer buf_n7313( .i (n7312), .o (n7313) );
  buffer buf_n7314( .i (n7313), .o (n7314) );
  buffer buf_n7315( .i (n7314), .o (n7315) );
  buffer buf_n7316( .i (n7315), .o (n7316) );
  buffer buf_n7317( .i (n7316), .o (n7317) );
  buffer buf_n7318( .i (n7317), .o (n7318) );
  buffer buf_n7319( .i (n7318), .o (n7319) );
  buffer buf_n7320( .i (n7319), .o (n7320) );
  buffer buf_n7321( .i (n7320), .o (n7321) );
  buffer buf_n7322( .i (n7321), .o (n7322) );
  buffer buf_n7323( .i (n7322), .o (n7323) );
  buffer buf_n7324( .i (n7323), .o (n7324) );
  buffer buf_n7325( .i (n7324), .o (n7325) );
  buffer buf_n7326( .i (n7325), .o (n7326) );
  buffer buf_n7327( .i (n7326), .o (n7327) );
  buffer buf_n7328( .i (n7327), .o (n7328) );
  buffer buf_n7329( .i (n7328), .o (n7329) );
  buffer buf_n5789( .i (n5788), .o (n5789) );
  buffer buf_n5790( .i (n5789), .o (n5790) );
  buffer buf_n5568( .i (n5567), .o (n5568) );
  buffer buf_n5569( .i (n5568), .o (n5569) );
  buffer buf_n5570( .i (n5569), .o (n5570) );
  buffer buf_n5571( .i (n5570), .o (n5571) );
  buffer buf_n5572( .i (n5571), .o (n5572) );
  buffer buf_n5573( .i (n5572), .o (n5573) );
  buffer buf_n5574( .i (n5573), .o (n5574) );
  buffer buf_n5575( .i (n5574), .o (n5575) );
  buffer buf_n5576( .i (n5575), .o (n5576) );
  buffer buf_n5577( .i (n5576), .o (n5577) );
  buffer buf_n5578( .i (n5577), .o (n5578) );
  buffer buf_n5579( .i (n5578), .o (n5579) );
  buffer buf_n5580( .i (n5579), .o (n5580) );
  buffer buf_n5581( .i (n5580), .o (n5581) );
  buffer buf_n5582( .i (n5581), .o (n5582) );
  buffer buf_n5583( .i (n5582), .o (n5583) );
  buffer buf_n5584( .i (n5583), .o (n5584) );
  assign n7330 = n5584 | n7290 ;
  buffer buf_n7331( .i (n7330), .o (n7331) );
  assign n7332 = n5790 | n7331 ;
  assign n7333 = n5790 & n7331 ;
  assign n7334 = n7332 & ~n7333 ;
  buffer buf_n7335( .i (n7334), .o (n7335) );
  buffer buf_n7336( .i (n7335), .o (n7336) );
  buffer buf_n7337( .i (n7336), .o (n7337) );
  buffer buf_n7338( .i (n7337), .o (n7338) );
  buffer buf_n7339( .i (n7338), .o (n7339) );
  buffer buf_n7340( .i (n7339), .o (n7340) );
  buffer buf_n7341( .i (n7340), .o (n7341) );
  buffer buf_n7342( .i (n7341), .o (n7342) );
  buffer buf_n7343( .i (n7342), .o (n7343) );
  buffer buf_n7344( .i (n7343), .o (n7344) );
  buffer buf_n7345( .i (n7344), .o (n7345) );
  buffer buf_n7346( .i (n7345), .o (n7346) );
  buffer buf_n7347( .i (n7346), .o (n7347) );
  buffer buf_n7348( .i (n7347), .o (n7348) );
  buffer buf_n7349( .i (n7348), .o (n7349) );
  buffer buf_n7350( .i (n7349), .o (n7350) );
  buffer buf_n7351( .i (n7350), .o (n7351) );
  buffer buf_n7352( .i (n7351), .o (n7352) );
  buffer buf_n7353( .i (n7352), .o (n7353) );
  buffer buf_n7354( .i (n7353), .o (n7354) );
  buffer buf_n7355( .i (n7354), .o (n7355) );
  buffer buf_n7356( .i (n7355), .o (n7356) );
  buffer buf_n7357( .i (n7356), .o (n7357) );
  buffer buf_n7358( .i (n7357), .o (n7358) );
  buffer buf_n7359( .i (n7358), .o (n7359) );
  buffer buf_n7360( .i (n7359), .o (n7360) );
  buffer buf_n7361( .i (n7360), .o (n7361) );
  buffer buf_n7362( .i (n7361), .o (n7362) );
  buffer buf_n7363( .i (n7362), .o (n7363) );
  buffer buf_n7364( .i (n7363), .o (n7364) );
  buffer buf_n7365( .i (n7364), .o (n7365) );
  buffer buf_n7366( .i (n7365), .o (n7366) );
  buffer buf_n7367( .i (n7366), .o (n7367) );
  buffer buf_n7368( .i (n7367), .o (n7368) );
  buffer buf_n5770( .i (n5769), .o (n5770) );
  buffer buf_n5811( .i (n5810), .o (n5811) );
  buffer buf_n5812( .i (n5811), .o (n5812) );
  buffer buf_n5813( .i (n5812), .o (n5813) );
  buffer buf_n5814( .i (n5813), .o (n5814) );
  buffer buf_n5815( .i (n5814), .o (n5815) );
  buffer buf_n5816( .i (n5815), .o (n5816) );
  buffer buf_n5817( .i (n5816), .o (n5817) );
  buffer buf_n5818( .i (n5817), .o (n5818) );
  buffer buf_n5819( .i (n5818), .o (n5819) );
  buffer buf_n5820( .i (n5819), .o (n5820) );
  buffer buf_n5821( .i (n5820), .o (n5821) );
  buffer buf_n5822( .i (n5821), .o (n5822) );
  buffer buf_n5823( .i (n5822), .o (n5823) );
  buffer buf_n5824( .i (n5823), .o (n5824) );
  assign n7369 = n5770 & n5824 ;
  assign n7370 = n5770 | n5824 ;
  assign n7371 = ~n7369 & n7370 ;
  buffer buf_n7372( .i (n7371), .o (n7372) );
  buffer buf_n7373( .i (n7372), .o (n7373) );
  buffer buf_n7374( .i (n7373), .o (n7374) );
  buffer buf_n7375( .i (n7374), .o (n7375) );
  buffer buf_n7376( .i (n7375), .o (n7376) );
  buffer buf_n7377( .i (n7376), .o (n7377) );
  buffer buf_n7378( .i (n7377), .o (n7378) );
  buffer buf_n7379( .i (n7378), .o (n7379) );
  buffer buf_n7380( .i (n7379), .o (n7380) );
  buffer buf_n7381( .i (n7380), .o (n7381) );
  buffer buf_n7382( .i (n7381), .o (n7382) );
  buffer buf_n7383( .i (n7382), .o (n7383) );
  buffer buf_n7384( .i (n7383), .o (n7384) );
  buffer buf_n7385( .i (n7384), .o (n7385) );
  buffer buf_n7386( .i (n7385), .o (n7386) );
  buffer buf_n7387( .i (n7386), .o (n7387) );
  buffer buf_n7388( .i (n7387), .o (n7388) );
  buffer buf_n7389( .i (n7388), .o (n7389) );
  buffer buf_n7390( .i (n7389), .o (n7390) );
  buffer buf_n7391( .i (n7390), .o (n7391) );
  buffer buf_n7392( .i (n7391), .o (n7392) );
  buffer buf_n7393( .i (n7392), .o (n7393) );
  buffer buf_n7394( .i (n7393), .o (n7394) );
  buffer buf_n7395( .i (n7394), .o (n7395) );
  buffer buf_n7396( .i (n7395), .o (n7396) );
  buffer buf_n7397( .i (n7396), .o (n7397) );
  buffer buf_n7398( .i (n7397), .o (n7398) );
  buffer buf_n7399( .i (n7398), .o (n7399) );
  buffer buf_n7400( .i (n7399), .o (n7400) );
  buffer buf_n7401( .i (n7400), .o (n7401) );
  buffer buf_n7402( .i (n7401), .o (n7402) );
  buffer buf_n7403( .i (n7402), .o (n7403) );
  buffer buf_n7404( .i (n7403), .o (n7404) );
  buffer buf_n7405( .i (n7404), .o (n7405) );
  buffer buf_n7406( .i (n7405), .o (n7406) );
  buffer buf_n7407( .i (n7406), .o (n7407) );
  buffer buf_n7408( .i (n7407), .o (n7408) );
  buffer buf_n4215( .i (n4214), .o (n4215) );
  buffer buf_n4216( .i (n4215), .o (n4216) );
  assign n7409 = n4216 & ~n4297 ;
  buffer buf_n4294( .i (n4293), .o (n4294) );
  buffer buf_n4295( .i (n4294), .o (n4295) );
  assign n7410 = ~n4218 & n4295 ;
  assign n7411 = n7409 | n7410 ;
  buffer buf_n7412( .i (n7411), .o (n7412) );
  buffer buf_n7413( .i (n7412), .o (n7413) );
  buffer buf_n7414( .i (n7413), .o (n7414) );
  buffer buf_n4313( .i (n4312), .o (n4313) );
  buffer buf_n4314( .i (n4313), .o (n4314) );
  assign n7415 = n4314 & ~n4331 ;
  buffer buf_n4328( .i (n4327), .o (n4328) );
  buffer buf_n4329( .i (n4328), .o (n4329) );
  assign n7416 = ~n4316 & n4329 ;
  assign n7417 = n7415 | n7416 ;
  buffer buf_n7418( .i (n7417), .o (n7418) );
  buffer buf_n407( .i (N141), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  assign n7419 = n410 & ~n6896 ;
  buffer buf_n7420( .i (n7419), .o (n7420) );
  buffer buf_n524( .i (N161), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n7421( .i (n6851), .o (n7421) );
  assign n7422 = n527 & n7421 ;
  buffer buf_n7423( .i (n7422), .o (n7423) );
  assign n7424 = n7420 | n7423 ;
  buffer buf_n7425( .i (n7424), .o (n7425) );
  assign n7426 = n4653 | n7425 ;
  assign n7427 = n4653 & n7425 ;
  assign n7428 = n7426 & ~n7427 ;
  buffer buf_n7429( .i (n7428), .o (n7429) );
  assign n7430 = n7418 | n7429 ;
  assign n7431 = n7418 & n7429 ;
  assign n7432 = n7430 & ~n7431 ;
  buffer buf_n7433( .i (n7432), .o (n7433) );
  assign n7434 = n7414 & ~n7433 ;
  assign n7435 = ~n7414 & n7433 ;
  assign n7436 = n7434 | n7435 ;
  buffer buf_n7437( .i (n7436), .o (n7437) );
  assign n7438 = n4559 & ~n4594 ;
  assign n7439 = ~n4559 & n4594 ;
  assign n7440 = n7438 | n7439 ;
  buffer buf_n7441( .i (n7440), .o (n7441) );
  assign n7442 = n4622 & n4641 ;
  assign n7443 = n4622 | n4641 ;
  assign n7444 = ~n7442 & n7443 ;
  buffer buf_n7445( .i (n7444), .o (n7445) );
  assign n7446 = n7441 & n7445 ;
  assign n7447 = n7441 | n7445 ;
  assign n7448 = ~n7446 & n7447 ;
  buffer buf_n7449( .i (n7448), .o (n7449) );
  buffer buf_n7450( .i (n7449), .o (n7450) );
  buffer buf_n7451( .i (n7450), .o (n7451) );
  buffer buf_n7452( .i (n7451), .o (n7452) );
  assign n7453 = ~n7437 & n7452 ;
  buffer buf_n7454( .i (n7453), .o (n7454) );
  assign n7455 = n3985 & ~n6906 ;
  buffer buf_n7456( .i (n7455), .o (n7456) );
  buffer buf_n7457( .i (n7456), .o (n7457) );
  buffer buf_n7458( .i (n7457), .o (n7458) );
  buffer buf_n7459( .i (n7458), .o (n7459) );
  buffer buf_n3887( .i (n3886), .o (n3887) );
  buffer buf_n3888( .i (n3887), .o (n3888) );
  assign n7460 = n3888 & ~n3900 ;
  buffer buf_n3897( .i (n3896), .o (n3897) );
  buffer buf_n3898( .i (n3897), .o (n3898) );
  assign n7461 = ~n3890 & n3898 ;
  assign n7462 = n7460 | n7461 ;
  buffer buf_n7463( .i (n7462), .o (n7463) );
  assign n7464 = n7459 | n7463 ;
  assign n7465 = n7459 & n7463 ;
  assign n7466 = n7464 & ~n7465 ;
  buffer buf_n7467( .i (n7466), .o (n7467) );
  buffer buf_n3956( .i (n3955), .o (n3956) );
  buffer buf_n3957( .i (n3956), .o (n3957) );
  assign n7468 = n3957 & ~n3979 ;
  buffer buf_n3975( .i (n3974), .o (n3975) );
  buffer buf_n3976( .i (n3975), .o (n3976) );
  assign n7469 = ~n3959 & n3976 ;
  assign n7470 = n7468 | n7469 ;
  buffer buf_n7471( .i (n7470), .o (n7471) );
  assign n7472 = ~n3881 & n7421 ;
  buffer buf_n7473( .i (n7472), .o (n7473) );
  buffer buf_n683( .i (N211), .o (n683) );
  buffer buf_n684( .i (N212), .o (n684) );
  assign n7474 = n683 | n684 ;
  assign n7475 = n683 & n684 ;
  assign n7476 = n7474 & ~n7475 ;
  buffer buf_n7477( .i (n7476), .o (n7477) );
  buffer buf_n7478( .i (n7477), .o (n7478) );
  buffer buf_n7479( .i (n7478), .o (n7479) );
  assign n7480 = n7473 & n7479 ;
  buffer buf_n7481( .i (n7480), .o (n7481) );
  buffer buf_n7482( .i (n7481), .o (n7482) );
  buffer buf_n7483( .i (n7482), .o (n7483) );
  buffer buf_n7484( .i (n7483), .o (n7484) );
  assign n7485 = ~n7471 & n7484 ;
  assign n7486 = n7471 & ~n7484 ;
  assign n7487 = n7485 | n7486 ;
  buffer buf_n7488( .i (n7487), .o (n7488) );
  assign n7489 = n7467 | n7488 ;
  assign n7490 = n7467 & n7488 ;
  assign n7491 = n7489 & ~n7490 ;
  buffer buf_n7492( .i (n7491), .o (n7492) );
  buffer buf_n7493( .i (n7492), .o (n7493) );
  assign n7494 = n7437 & ~n7452 ;
  assign n7495 = n7493 | n7494 ;
  assign n7496 = n7454 | n7495 ;
  buffer buf_n741( .i (N229), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  assign n7497 = n744 & n7421 ;
  buffer buf_n7498( .i (n7497), .o (n7498) );
  assign n7499 = n3609 | n7498 ;
  buffer buf_n7500( .i (n7499), .o (n7500) );
  assign n7501 = ~n5534 & n7500 ;
  assign n7502 = n5534 & ~n7500 ;
  assign n7503 = n7501 | n7502 ;
  buffer buf_n7504( .i (n7503), .o (n7504) );
  assign n7505 = n5511 & ~n5668 ;
  assign n7506 = ~n5511 & n5668 ;
  assign n7507 = n7505 | n7506 ;
  buffer buf_n7508( .i (n7507), .o (n7508) );
  assign n7509 = ~n7504 & n7508 ;
  assign n7510 = n7504 & ~n7508 ;
  assign n7511 = n7509 | n7510 ;
  buffer buf_n7512( .i (n7511), .o (n7512) );
  buffer buf_n7513( .i (n7512), .o (n7513) );
  buffer buf_n7514( .i (n7513), .o (n7514) );
  buffer buf_n7515( .i (n7514), .o (n7515) );
  assign n7516 = ~n5635 & n5694 ;
  assign n7517 = n5635 & ~n5694 ;
  assign n7518 = n7516 | n7517 ;
  buffer buf_n7519( .i (n7518), .o (n7519) );
  buffer buf_n7520( .i (n7519), .o (n7520) );
  buffer buf_n7521( .i (n7520), .o (n7521) );
  buffer buf_n7522( .i (n7521), .o (n7522) );
  assign n7523 = n5552 & ~n5564 ;
  assign n7524 = ~n5552 & n5564 ;
  assign n7525 = n7523 | n7524 ;
  buffer buf_n7526( .i (n7525), .o (n7526) );
  buffer buf_n781( .i (N239), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  assign n7527 = n784 & n7421 ;
  buffer buf_n7528( .i (n7527), .o (n7528) );
  buffer buf_n3451( .i (N44), .o (n3451) );
  buffer buf_n3452( .i (n3451), .o (n3452) );
  buffer buf_n3453( .i (n3452), .o (n3453) );
  buffer buf_n3454( .i (n3453), .o (n3454) );
  buffer buf_n7529( .i (n6850), .o (n7529) );
  buffer buf_n7530( .i (n7529), .o (n7530) );
  assign n7531 = n3454 & ~n7530 ;
  buffer buf_n7532( .i (n7531), .o (n7532) );
  assign n7533 = n7528 | n7532 ;
  buffer buf_n7534( .i (n7533), .o (n7534) );
  assign n7535 = n5705 | n7534 ;
  assign n7536 = n5705 & n7534 ;
  assign n7537 = n7535 & ~n7536 ;
  buffer buf_n7538( .i (n7537), .o (n7538) );
  assign n7539 = n7526 & ~n7538 ;
  assign n7540 = ~n7526 & n7538 ;
  assign n7541 = n7539 | n7540 ;
  buffer buf_n7542( .i (n7541), .o (n7542) );
  assign n7543 = n7522 | n7542 ;
  assign n7544 = n7522 & n7542 ;
  assign n7545 = n7543 & ~n7544 ;
  buffer buf_n7546( .i (n7545), .o (n7546) );
  assign n7547 = ~n7515 & n7546 ;
  assign n7548 = n7515 & ~n7546 ;
  assign n7549 = n7547 | n7548 ;
  assign n7550 = ~n5343 & n5455 ;
  assign n7551 = n5343 & ~n5455 ;
  assign n7552 = n7550 | n7551 ;
  buffer buf_n7553( .i (n7552), .o (n7553) );
  assign n7554 = n5301 & n5394 ;
  assign n7555 = n5301 | n5394 ;
  assign n7556 = ~n7554 & n7555 ;
  buffer buf_n7557( .i (n7556), .o (n7557) );
  assign n7558 = n7553 & ~n7557 ;
  assign n7559 = ~n7553 & n7557 ;
  assign n7560 = n7558 | n7559 ;
  buffer buf_n7561( .i (n7560), .o (n7561) );
  buffer buf_n7562( .i (n7561), .o (n7562) );
  buffer buf_n7563( .i (n7562), .o (n7563) );
  buffer buf_n7564( .i (n7563), .o (n7564) );
  buffer buf_n737( .i (N227), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  assign n7565 = n740 & n7530 ;
  buffer buf_n7566( .i (n7565), .o (n7566) );
  buffer buf_n372( .i (N115), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  assign n7567 = n375 & ~n7530 ;
  buffer buf_n7568( .i (n7567), .o (n7568) );
  assign n7569 = n7566 | n7568 ;
  buffer buf_n7570( .i (n7569), .o (n7570) );
  assign n7571 = n5269 | n7570 ;
  assign n7572 = n5269 & n7570 ;
  assign n7573 = n7571 & ~n7572 ;
  buffer buf_n7574( .i (n7573), .o (n7574) );
  buffer buf_n7575( .i (n7574), .o (n7575) );
  buffer buf_n7576( .i (n7575), .o (n7576) );
  buffer buf_n7577( .i (n7576), .o (n7577) );
  assign n7578 = n4983 & ~n5047 ;
  assign n7579 = ~n4983 & n5047 ;
  assign n7580 = n7578 | n7579 ;
  buffer buf_n7581( .i (n7580), .o (n7581) );
  assign n7582 = n5068 & n5082 ;
  assign n7583 = n5068 | n5082 ;
  assign n7584 = ~n7582 & n7583 ;
  buffer buf_n7585( .i (n7584), .o (n7585) );
  assign n7586 = n7581 | n7585 ;
  assign n7587 = n7581 & n7585 ;
  assign n7588 = n7586 & ~n7587 ;
  buffer buf_n7589( .i (n7588), .o (n7589) );
  assign n7590 = ~n7577 & n7589 ;
  assign n7591 = n7577 & ~n7589 ;
  assign n7592 = n7590 | n7591 ;
  buffer buf_n7593( .i (n7592), .o (n7593) );
  assign n7594 = n7564 & ~n7593 ;
  assign n7595 = ~n7564 & n7593 ;
  assign n7596 = n7594 | n7595 ;
  assign n7597 = n7549 & n7596 ;
  assign n7598 = ~n7496 & n7597 ;
  buffer buf_n7599( .i (n7598), .o (n7599) );
  buffer buf_n7600( .i (n7599), .o (n7600) );
  buffer buf_n7601( .i (n7600), .o (n7601) );
  buffer buf_n7602( .i (n7601), .o (n7602) );
  buffer buf_n7603( .i (n7602), .o (n7603) );
  buffer buf_n7604( .i (n7603), .o (n7604) );
  buffer buf_n7605( .i (n7604), .o (n7605) );
  buffer buf_n7606( .i (n7605), .o (n7606) );
  buffer buf_n7607( .i (n7606), .o (n7607) );
  buffer buf_n7608( .i (n7607), .o (n7608) );
  buffer buf_n7609( .i (n7608), .o (n7609) );
  buffer buf_n7610( .i (n7609), .o (n7610) );
  buffer buf_n7611( .i (n7610), .o (n7611) );
  buffer buf_n7612( .i (n7611), .o (n7612) );
  buffer buf_n7613( .i (n7612), .o (n7613) );
  buffer buf_n7614( .i (n7613), .o (n7614) );
  buffer buf_n7615( .i (n7614), .o (n7615) );
  buffer buf_n7616( .i (n7615), .o (n7616) );
  buffer buf_n7617( .i (n7616), .o (n7617) );
  buffer buf_n7618( .i (n7617), .o (n7618) );
  buffer buf_n7619( .i (n7618), .o (n7619) );
  buffer buf_n7620( .i (n7619), .o (n7620) );
  buffer buf_n7621( .i (n7620), .o (n7621) );
  buffer buf_n7622( .i (n7621), .o (n7622) );
  buffer buf_n7623( .i (n7622), .o (n7623) );
  buffer buf_n7624( .i (n7623), .o (n7624) );
  buffer buf_n7625( .i (n7624), .o (n7625) );
  buffer buf_n7626( .i (n7625), .o (n7626) );
  buffer buf_n7627( .i (n7626), .o (n7627) );
  buffer buf_n7628( .i (n7627), .o (n7628) );
  buffer buf_n7629( .i (n7628), .o (n7629) );
  buffer buf_n7630( .i (n7629), .o (n7630) );
  buffer buf_n7631( .i (n7630), .o (n7631) );
  buffer buf_n7632( .i (n7631), .o (n7632) );
  buffer buf_n7633( .i (n7632), .o (n7633) );
  buffer buf_n7634( .i (n7633), .o (n7634) );
  buffer buf_n7635( .i (n7634), .o (n7635) );
  buffer buf_n7636( .i (n7635), .o (n7636) );
  buffer buf_n7637( .i (n7636), .o (n7637) );
  buffer buf_n7638( .i (n7637), .o (n7638) );
  buffer buf_n7639( .i (n7638), .o (n7639) );
  buffer buf_n7640( .i (n7639), .o (n7640) );
  buffer buf_n7641( .i (n7640), .o (n7641) );
  buffer buf_n7642( .i (n7641), .o (n7642) );
  buffer buf_n7643( .i (n7642), .o (n7643) );
  buffer buf_n368( .i (N114), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  assign n7644 = n371 & ~n7530 ;
  buffer buf_n853( .i (N248), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n7645( .i (n7529), .o (n7645) );
  assign n7646 = ~n856 & n7645 ;
  assign n7647 = n7644 | n7646 ;
  buffer buf_n7648( .i (n7647), .o (n7648) );
  assign n7649 = n6893 & n7648 ;
  assign n7650 = n6893 | n7648 ;
  assign n7651 = ~n7649 & n7650 ;
  buffer buf_n7652( .i (n7651), .o (n7652) );
  assign n7653 = n6856 & ~n6874 ;
  assign n7654 = ~n6856 & n6874 ;
  assign n7655 = n7653 | n7654 ;
  buffer buf_n7656( .i (n7655), .o (n7656) );
  assign n7657 = ~n7652 & n7656 ;
  assign n7658 = n7652 & ~n7656 ;
  assign n7659 = n7657 | n7658 ;
  buffer buf_n7660( .i (n7659), .o (n7660) );
  assign n7661 = n6838 & n6900 ;
  assign n7662 = n6838 | n6900 ;
  assign n7663 = ~n7661 & n7662 ;
  buffer buf_n7664( .i (n7663), .o (n7664) );
  assign n7665 = n1188 & ~n1254 ;
  assign n7666 = ~n1188 & n1254 ;
  assign n7667 = n7665 | n7666 ;
  assign n7668 = n7645 & n7667 ;
  buffer buf_n6948( .i (n6947), .o (n6948) );
  assign n7669 = n6198 | n7529 ;
  assign n7670 = n6948 & ~n7669 ;
  assign n7671 = n7668 | n7670 ;
  buffer buf_n7672( .i (n7671), .o (n7672) );
  buffer buf_n7673( .i (n7672), .o (n7673) );
  buffer buf_n7674( .i (n7673), .o (n7674) );
  buffer buf_n7675( .i (n7674), .o (n7675) );
  assign n7676 = ~n7664 & n7675 ;
  assign n7677 = n7664 & ~n7675 ;
  assign n7678 = n7676 | n7677 ;
  buffer buf_n7679( .i (n7678), .o (n7679) );
  assign n7680 = ~n7660 & n7679 ;
  assign n7681 = n7660 & ~n7679 ;
  assign n7682 = n7680 | n7681 ;
  buffer buf_n7683( .i (n7682), .o (n7683) );
  buffer buf_n7684( .i (n7683), .o (n7684) );
  buffer buf_n7685( .i (n7684), .o (n7685) );
  assign n7686 = n2054 & n6418 ;
  assign n7687 = n6271 & ~n7686 ;
  buffer buf_n7688( .i (n7687), .o (n7688) );
  buffer buf_n3518( .i (N69), .o (n3518) );
  buffer buf_n3519( .i (n3518), .o (n3519) );
  buffer buf_n3520( .i (n3519), .o (n3520) );
  buffer buf_n3521( .i (n3520), .o (n3521) );
  assign n7689 = n3521 & ~n7645 ;
  buffer buf_n1984( .i (N307), .o (n1984) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n1986( .i (n1985), .o (n1986) );
  buffer buf_n1987( .i (n1986), .o (n1987) );
  assign n7690 = ~n1987 & n7645 ;
  assign n7691 = n7689 | n7690 ;
  buffer buf_n7692( .i (n7691), .o (n7692) );
  buffer buf_n7693( .i (n7692), .o (n7693) );
  assign n7694 = n7688 & n7693 ;
  assign n7695 = n7688 | n7693 ;
  assign n7696 = ~n7694 & n7695 ;
  buffer buf_n7697( .i (n7696), .o (n7697) );
  assign n7698 = n6261 & n6279 ;
  assign n7699 = n6261 | n6279 ;
  assign n7700 = ~n7698 & n7699 ;
  buffer buf_n7701( .i (n7700), .o (n7701) );
  assign n7702 = n7697 & ~n7701 ;
  assign n7703 = ~n7697 & n7701 ;
  assign n7704 = n7702 | n7703 ;
  buffer buf_n7705( .i (n7704), .o (n7705) );
  buffer buf_n7706( .i (n7705), .o (n7706) );
  buffer buf_n7707( .i (n7706), .o (n7707) );
  buffer buf_n6320( .i (n6319), .o (n6320) );
  buffer buf_n6321( .i (n6320), .o (n6321) );
  assign n7708 = n6339 & ~n6351 ;
  assign n7709 = ~n6339 & n6351 ;
  assign n7710 = n7708 | n7709 ;
  buffer buf_n7711( .i (n7710), .o (n7711) );
  assign n7712 = n6321 & ~n7711 ;
  assign n7713 = ~n6321 & n7711 ;
  assign n7714 = n7712 | n7713 ;
  buffer buf_n7715( .i (n7714), .o (n7715) );
  buffer buf_n6294( .i (n6293), .o (n6294) );
  buffer buf_n6295( .i (n6294), .o (n6295) );
  assign n7716 = n6230 & n6246 ;
  assign n7717 = n6230 | n6246 ;
  assign n7718 = ~n7716 & n7717 ;
  buffer buf_n7719( .i (n7718), .o (n7719) );
  assign n7720 = n6295 & n7719 ;
  assign n7721 = n6295 | n7719 ;
  assign n7722 = ~n7720 & n7721 ;
  buffer buf_n7723( .i (n7722), .o (n7723) );
  assign n7724 = ~n7715 & n7723 ;
  assign n7725 = n7715 & ~n7723 ;
  assign n7726 = n7724 | n7725 ;
  buffer buf_n7727( .i (n7726), .o (n7727) );
  assign n7728 = ~n7707 & n7727 ;
  assign n7729 = n7707 & ~n7727 ;
  assign n7730 = n7728 | n7729 ;
  assign n7731 = n7685 & n7730 ;
  assign n7732 = n6395 & n6407 ;
  assign n7733 = n6395 | n6407 ;
  assign n7734 = ~n7732 & n7733 ;
  buffer buf_n7735( .i (n7734), .o (n7735) );
  assign n7736 = n6479 & ~n6491 ;
  assign n7737 = ~n6479 & n6491 ;
  assign n7738 = n7736 | n7737 ;
  buffer buf_n7739( .i (n7738), .o (n7739) );
  assign n7740 = n7735 | n7739 ;
  assign n7741 = n7735 & n7739 ;
  assign n7742 = n7740 & ~n7741 ;
  buffer buf_n7743( .i (n7742), .o (n7743) );
  assign n7744 = n6421 & n6442 ;
  assign n7745 = n6421 | n6442 ;
  assign n7746 = ~n7744 & n7745 ;
  buffer buf_n7747( .i (n7746), .o (n7747) );
  buffer buf_n7748( .i (n7747), .o (n7748) );
  buffer buf_n7749( .i (n7748), .o (n7749) );
  assign n7750 = ~n7743 & n7749 ;
  assign n7751 = n7743 & ~n7749 ;
  assign n7752 = n7750 | n7751 ;
  buffer buf_n7753( .i (n7752), .o (n7753) );
  assign n7754 = n6512 & n6524 ;
  assign n7755 = n6512 | n6524 ;
  assign n7756 = ~n7754 & n7755 ;
  buffer buf_n7757( .i (n7756), .o (n7757) );
  buffer buf_n3481( .i (N58), .o (n3481) );
  buffer buf_n3482( .i (n3481), .o (n3482) );
  buffer buf_n3483( .i (n3482), .o (n3483) );
  buffer buf_n3484( .i (n3483), .o (n3484) );
  buffer buf_n7758( .i (n7529), .o (n7758) );
  assign n7759 = n3484 & ~n7758 ;
  buffer buf_n2648( .i (N337), .o (n2648) );
  buffer buf_n2649( .i (n2648), .o (n2649) );
  buffer buf_n2650( .i (n2649), .o (n2650) );
  buffer buf_n2651( .i (n2650), .o (n2651) );
  assign n7760 = ~n2651 & n7758 ;
  assign n7761 = n7759 | n7760 ;
  buffer buf_n7762( .i (n7761), .o (n7762) );
  assign n7763 = n6375 & n7762 ;
  assign n7764 = n6375 | n7762 ;
  assign n7765 = ~n7763 & n7764 ;
  buffer buf_n7766( .i (n7765), .o (n7766) );
  assign n7767 = n7757 | n7766 ;
  assign n7768 = n7757 & n7766 ;
  assign n7769 = n7767 & ~n7768 ;
  buffer buf_n7770( .i (n7769), .o (n7770) );
  buffer buf_n7771( .i (n7770), .o (n7771) );
  buffer buf_n7772( .i (n7771), .o (n7772) );
  buffer buf_n7773( .i (n7772), .o (n7773) );
  assign n7774 = n7753 & ~n7773 ;
  assign n7775 = ~n7753 & n7773 ;
  assign n7776 = n7774 | n7775 ;
  assign n7777 = n6611 & n6622 ;
  assign n7778 = n6611 | n6622 ;
  assign n7779 = ~n7777 & n7778 ;
  buffer buf_n7780( .i (n7779), .o (n7780) );
  assign n7781 = ~n6733 & n6746 ;
  assign n7782 = n6733 & ~n6746 ;
  assign n7783 = n7781 | n7782 ;
  buffer buf_n7784( .i (n7783), .o (n7784) );
  assign n7785 = ~n7780 & n7784 ;
  assign n7786 = n7780 & ~n7784 ;
  assign n7787 = n7785 | n7786 ;
  buffer buf_n7788( .i (n7787), .o (n7788) );
  buffer buf_n7789( .i (n7788), .o (n7789) );
  buffer buf_n7790( .i (n7789), .o (n7790) );
  buffer buf_n7791( .i (n7790), .o (n7791) );
  buffer buf_n6646( .i (n6645), .o (n6646) );
  buffer buf_n6647( .i (n6646), .o (n6647) );
  buffer buf_n3566( .i (N82), .o (n3566) );
  buffer buf_n3567( .i (n3566), .o (n3567) );
  buffer buf_n3568( .i (n3567), .o (n3568) );
  buffer buf_n3569( .i (n3568), .o (n3569) );
  assign n7792 = n3569 & ~n7758 ;
  buffer buf_n1320( .i (N274), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  assign n7793 = ~n1323 & n7758 ;
  assign n7794 = n7792 | n7793 ;
  buffer buf_n7795( .i (n7794), .o (n7795) );
  assign n7796 = n6681 & ~n7795 ;
  assign n7797 = ~n6681 & n7795 ;
  assign n7798 = n7796 | n7797 ;
  buffer buf_n7799( .i (n7798), .o (n7799) );
  assign n7800 = n6647 | n7799 ;
  assign n7801 = n6647 & n7799 ;
  assign n7802 = n7800 & ~n7801 ;
  buffer buf_n7803( .i (n7802), .o (n7803) );
  buffer buf_n6659( .i (n6658), .o (n6659) );
  buffer buf_n6660( .i (n6659), .o (n6660) );
  assign n7804 = n6769 & ~n6781 ;
  assign n7805 = ~n6769 & n6781 ;
  assign n7806 = n7804 | n7805 ;
  buffer buf_n7807( .i (n7806), .o (n7807) );
  assign n7808 = n6660 & n7807 ;
  assign n7809 = n6660 | n7807 ;
  assign n7810 = ~n7808 & n7809 ;
  buffer buf_n7811( .i (n7810), .o (n7811) );
  assign n7812 = n7803 & n7811 ;
  assign n7813 = n7803 | n7811 ;
  assign n7814 = ~n7812 & n7813 ;
  buffer buf_n7815( .i (n7814), .o (n7815) );
  assign n7816 = n7791 & n7815 ;
  assign n7817 = n7791 | n7815 ;
  assign n7818 = ~n7816 & n7817 ;
  assign n7819 = n7776 & n7818 ;
  assign n7820 = n7731 & n7819 ;
  buffer buf_n7821( .i (n7820), .o (n7821) );
  buffer buf_n7822( .i (n7821), .o (n7822) );
  buffer buf_n7823( .i (n7822), .o (n7823) );
  buffer buf_n7824( .i (n7823), .o (n7824) );
  buffer buf_n7825( .i (n7824), .o (n7825) );
  buffer buf_n7826( .i (n7825), .o (n7826) );
  buffer buf_n7827( .i (n7826), .o (n7827) );
  buffer buf_n7828( .i (n7827), .o (n7828) );
  buffer buf_n7829( .i (n7828), .o (n7829) );
  buffer buf_n7830( .i (n7829), .o (n7830) );
  buffer buf_n7831( .i (n7830), .o (n7831) );
  buffer buf_n7832( .i (n7831), .o (n7832) );
  buffer buf_n7833( .i (n7832), .o (n7833) );
  buffer buf_n7834( .i (n7833), .o (n7834) );
  buffer buf_n7835( .i (n7834), .o (n7835) );
  buffer buf_n7836( .i (n7835), .o (n7836) );
  buffer buf_n7837( .i (n7836), .o (n7837) );
  buffer buf_n7838( .i (n7837), .o (n7838) );
  buffer buf_n7839( .i (n7838), .o (n7839) );
  buffer buf_n7840( .i (n7839), .o (n7840) );
  buffer buf_n7841( .i (n7840), .o (n7841) );
  buffer buf_n7842( .i (n7841), .o (n7842) );
  buffer buf_n7843( .i (n7842), .o (n7843) );
  buffer buf_n7844( .i (n7843), .o (n7844) );
  buffer buf_n7845( .i (n7844), .o (n7845) );
  buffer buf_n7846( .i (n7845), .o (n7846) );
  buffer buf_n7847( .i (n7846), .o (n7847) );
  buffer buf_n7848( .i (n7847), .o (n7848) );
  buffer buf_n7849( .i (n7848), .o (n7849) );
  buffer buf_n7850( .i (n7849), .o (n7850) );
  buffer buf_n7851( .i (n7850), .o (n7851) );
  buffer buf_n7852( .i (n7851), .o (n7852) );
  buffer buf_n7853( .i (n7852), .o (n7853) );
  buffer buf_n7854( .i (n7853), .o (n7854) );
  buffer buf_n7855( .i (n7854), .o (n7855) );
  buffer buf_n7856( .i (n7855), .o (n7856) );
  buffer buf_n7857( .i (n7856), .o (n7857) );
  buffer buf_n7858( .i (n7857), .o (n7858) );
  buffer buf_n7859( .i (n7858), .o (n7859) );
  buffer buf_n7860( .i (n7859), .o (n7860) );
  buffer buf_n7861( .i (n7860), .o (n7861) );
  buffer buf_n7862( .i (n7861), .o (n7862) );
  buffer buf_n7863( .i (n7862), .o (n7863) );
  buffer buf_n7864( .i (n7863), .o (n7864) );
  buffer buf_n7865( .i (n7864), .o (n7865) );
  buffer buf_n7866( .i (n7865), .o (n7866) );
  buffer buf_n548( .i (N170), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  assign n7867 = ~n553 & n7473 ;
  buffer buf_n7868( .i (n7867), .o (n7868) );
  buffer buf_n7869( .i (n7868), .o (n7869) );
  buffer buf_n7870( .i (n7869), .o (n7870) );
  buffer buf_n7871( .i (n7870), .o (n7871) );
  buffer buf_n6860( .i (n6859), .o (n6860) );
  buffer buf_n6861( .i (n6860), .o (n6861) );
  assign n7872 = n6861 & ~n6881 ;
  buffer buf_n6878( .i (n6877), .o (n6878) );
  buffer buf_n6879( .i (n6878), .o (n6879) );
  assign n7873 = ~n6863 & n6879 ;
  assign n7874 = n7872 | n7873 ;
  buffer buf_n7875( .i (n7874), .o (n7875) );
  assign n7876 = ~n7871 & n7875 ;
  assign n7877 = n7871 & ~n7875 ;
  assign n7878 = n7876 | n7877 ;
  buffer buf_n7879( .i (n7878), .o (n7879) );
  buffer buf_n6842( .i (n6841), .o (n6842) );
  buffer buf_n6843( .i (n6842), .o (n6843) );
  assign n7880 = n6843 & ~n6908 ;
  buffer buf_n6904( .i (n6903), .o (n6904) );
  buffer buf_n6905( .i (n6904), .o (n6905) );
  assign n7881 = ~n6845 & n6905 ;
  assign n7882 = n7880 | n7881 ;
  buffer buf_n7883( .i (n7882), .o (n7883) );
  buffer buf_n530( .i (N164), .o (n530) );
  buffer buf_n531( .i (N165), .o (n531) );
  assign n7884 = ~n530 & n531 ;
  assign n7885 = n530 & ~n531 ;
  assign n7886 = n7884 | n7885 ;
  buffer buf_n7887( .i (n7886), .o (n7887) );
  buffer buf_n7888( .i (n7887), .o (n7888) );
  buffer buf_n7889( .i (n7888), .o (n7889) );
  assign n7890 = n7473 & n7889 ;
  buffer buf_n7891( .i (n7890), .o (n7891) );
  buffer buf_n7892( .i (n7891), .o (n7892) );
  buffer buf_n7893( .i (n7892), .o (n7893) );
  buffer buf_n7894( .i (n7893), .o (n7894) );
  assign n7895 = n7883 | n7894 ;
  assign n7896 = n7883 & n7894 ;
  assign n7897 = n7895 & ~n7896 ;
  buffer buf_n7898( .i (n7897), .o (n7898) );
  assign n7899 = n7879 | n7898 ;
  assign n7900 = n7879 & n7898 ;
  assign n7901 = n7899 & ~n7900 ;
  buffer buf_n7902( .i (n7901), .o (n7902) );
  buffer buf_n7903( .i (n7902), .o (n7903) );
  buffer buf_n7904( .i (n7903), .o (n7904) );
  assign n7905 = n6426 & n6446 ;
  assign n7906 = n6426 | n6446 ;
  assign n7907 = ~n7905 & n7906 ;
  buffer buf_n7908( .i (n7907), .o (n7908) );
  buffer buf_n7909( .i (n7908), .o (n7909) );
  buffer buf_n7910( .i (n7909), .o (n7910) );
  buffer buf_n7911( .i (n7910), .o (n7911) );
  assign n7912 = n6485 & ~n6496 ;
  assign n7913 = ~n6485 & n6496 ;
  assign n7914 = n7912 | n7913 ;
  buffer buf_n7915( .i (n7914), .o (n7915) );
  assign n7916 = n6517 & n6529 ;
  assign n7917 = n6517 | n6529 ;
  assign n7918 = ~n7916 & n7917 ;
  buffer buf_n7919( .i (n7918), .o (n7919) );
  assign n7920 = ~n7915 & n7919 ;
  assign n7921 = n7915 & ~n7919 ;
  assign n7922 = n7920 | n7921 ;
  buffer buf_n7923( .i (n7922), .o (n7923) );
  assign n7924 = n7911 & n7923 ;
  assign n7925 = n7911 | n7923 ;
  assign n7926 = ~n7924 & n7925 ;
  buffer buf_n7927( .i (n7926), .o (n7927) );
  assign n7928 = n6400 & n6412 ;
  assign n7929 = n6400 | n6412 ;
  assign n7930 = ~n7928 & n7929 ;
  buffer buf_n7931( .i (n7930), .o (n7931) );
  buffer buf_n635( .i (N197), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n7932( .i (n6850), .o (n7932) );
  buffer buf_n7933( .i (n7932), .o (n7933) );
  assign n7934 = n638 & n7933 ;
  buffer buf_n7935( .i (n7934), .o (n7935) );
  assign n7936 = n7568 | n7935 ;
  buffer buf_n7937( .i (n7936), .o (n7937) );
  assign n7938 = n6381 | n7937 ;
  assign n7939 = n6381 & n7937 ;
  assign n7940 = n7938 & ~n7939 ;
  buffer buf_n7941( .i (n7940), .o (n7941) );
  assign n7942 = ~n7931 & n7941 ;
  assign n7943 = n7931 & ~n7941 ;
  assign n7944 = n7942 | n7943 ;
  buffer buf_n7945( .i (n7944), .o (n7945) );
  buffer buf_n7946( .i (n7945), .o (n7946) );
  buffer buf_n7947( .i (n7946), .o (n7947) );
  buffer buf_n7948( .i (n7947), .o (n7948) );
  assign n7949 = n7927 | n7948 ;
  assign n7950 = n7927 & n7948 ;
  assign n7951 = n7949 & ~n7950 ;
  assign n7952 = ~n7904 & n7951 ;
  buffer buf_n595( .i (N181), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  assign n7953 = n598 & n7933 ;
  buffer buf_n7954( .i (n7953), .o (n7954) );
  assign n7955 = n7420 | n7954 ;
  buffer buf_n7956( .i (n7955), .o (n7956) );
  assign n7957 = n6688 & ~n7956 ;
  assign n7958 = ~n6688 & n7956 ;
  assign n7959 = n7957 | n7958 ;
  buffer buf_n7960( .i (n7959), .o (n7960) );
  buffer buf_n7961( .i (n7960), .o (n7961) );
  buffer buf_n7962( .i (n7961), .o (n7962) );
  buffer buf_n7963( .i (n7962), .o (n7963) );
  buffer buf_n6750( .i (n6749), .o (n6750) );
  buffer buf_n6751( .i (n6750), .o (n6751) );
  assign n7964 = ~n6740 & n6751 ;
  buffer buf_n6737( .i (n6736), .o (n6737) );
  buffer buf_n6738( .i (n6737), .o (n6738) );
  assign n7965 = n6738 & ~n6753 ;
  assign n7966 = n7964 | n7965 ;
  buffer buf_n7967( .i (n7966), .o (n7967) );
  buffer buf_n6773( .i (n6772), .o (n6773) );
  buffer buf_n6774( .i (n6773), .o (n6774) );
  assign n7968 = n6774 & ~n6791 ;
  buffer buf_n6786( .i (n6785), .o (n6786) );
  buffer buf_n6787( .i (n6786), .o (n6787) );
  assign n7969 = ~n6776 & n6787 ;
  assign n7970 = n7968 | n7969 ;
  buffer buf_n7971( .i (n7970), .o (n7971) );
  assign n7972 = n7967 | n7971 ;
  assign n7973 = n7967 & n7971 ;
  assign n7974 = n7972 & ~n7973 ;
  buffer buf_n7975( .i (n7974), .o (n7975) );
  assign n7976 = ~n7963 & n7975 ;
  assign n7977 = n7963 & ~n7975 ;
  assign n7978 = n7976 | n7977 ;
  buffer buf_n7979( .i (n7978), .o (n7979) );
  buffer buf_n6616( .i (n6615), .o (n6616) );
  assign n7980 = n6616 & n6627 ;
  assign n7981 = n6616 | n6627 ;
  assign n7982 = ~n7980 & n7981 ;
  buffer buf_n7983( .i (n7982), .o (n7983) );
  assign n7984 = n6651 & n6664 ;
  assign n7985 = n6651 | n6664 ;
  assign n7986 = ~n7984 & n7985 ;
  buffer buf_n7987( .i (n7986), .o (n7987) );
  assign n7988 = ~n7983 & n7987 ;
  assign n7989 = n7983 & ~n7987 ;
  assign n7990 = n7988 | n7989 ;
  buffer buf_n7991( .i (n7990), .o (n7991) );
  buffer buf_n7992( .i (n7991), .o (n7992) );
  buffer buf_n7993( .i (n7992), .o (n7993) );
  buffer buf_n7994( .i (n7993), .o (n7994) );
  assign n7995 = ~n7979 & n7994 ;
  assign n7996 = n7979 & ~n7994 ;
  assign n7997 = n7995 | n7996 ;
  buffer buf_n675( .i (N208), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  assign n7998 = n678 & n7933 ;
  buffer buf_n7999( .i (n7998), .o (n7999) );
  assign n8000 = n7532 | n7999 ;
  buffer buf_n8001( .i (n8000), .o (n8001) );
  buffer buf_n639( .i (N198), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  assign n8002 = n642 & n7933 ;
  buffer buf_n8003( .i (n8002), .o (n8003) );
  assign n8004 = n3609 | n8003 ;
  buffer buf_n8005( .i (n8004), .o (n8005) );
  assign n8006 = n8001 | n8005 ;
  assign n8007 = n8001 & n8005 ;
  assign n8008 = n8006 & ~n8007 ;
  buffer buf_n8009( .i (n8008), .o (n8009) );
  buffer buf_n8010( .i (n8009), .o (n8010) );
  buffer buf_n8011( .i (n8010), .o (n8011) );
  buffer buf_n8012( .i (n8011), .o (n8012) );
  assign n8013 = n6265 & n6283 ;
  assign n8014 = n6265 | n6283 ;
  assign n8015 = ~n8013 & n8014 ;
  buffer buf_n8016( .i (n8015), .o (n8016) );
  assign n8017 = n6251 & ~n6302 ;
  assign n8018 = ~n6251 & n6302 ;
  assign n8019 = n8017 | n8018 ;
  buffer buf_n8020( .i (n8019), .o (n8020) );
  assign n8021 = n8016 | n8020 ;
  assign n8022 = n8016 & n8020 ;
  assign n8023 = n8021 & ~n8022 ;
  buffer buf_n8024( .i (n8023), .o (n8024) );
  assign n8025 = n8012 | n8024 ;
  assign n8026 = n8012 & n8024 ;
  assign n8027 = n8025 & ~n8026 ;
  buffer buf_n8028( .i (n8027), .o (n8028) );
  assign n8029 = n6344 & ~n6356 ;
  assign n8030 = ~n6344 & n6356 ;
  assign n8031 = n8029 | n8030 ;
  buffer buf_n8032( .i (n8031), .o (n8032) );
  assign n8033 = n6235 & n6325 ;
  assign n8034 = n6235 | n6325 ;
  assign n8035 = ~n8033 & n8034 ;
  buffer buf_n8036( .i (n8035), .o (n8036) );
  assign n8037 = n8032 | n8036 ;
  assign n8038 = n8032 & n8036 ;
  assign n8039 = n8037 & ~n8038 ;
  buffer buf_n8040( .i (n8039), .o (n8040) );
  buffer buf_n8041( .i (n8040), .o (n8041) );
  buffer buf_n8042( .i (n8041), .o (n8042) );
  buffer buf_n8043( .i (n8042), .o (n8043) );
  assign n8044 = n8028 & n8043 ;
  assign n8045 = n8028 | n8043 ;
  assign n8046 = ~n8044 & n8045 ;
  assign n8047 = ~n7997 & n8046 ;
  assign n8048 = n7952 & n8047 ;
  buffer buf_n8049( .i (n8048), .o (n8049) );
  buffer buf_n8050( .i (n8049), .o (n8050) );
  buffer buf_n8051( .i (n8050), .o (n8051) );
  buffer buf_n8052( .i (n8051), .o (n8052) );
  buffer buf_n8053( .i (n8052), .o (n8053) );
  buffer buf_n8054( .i (n8053), .o (n8054) );
  buffer buf_n8055( .i (n8054), .o (n8055) );
  buffer buf_n8056( .i (n8055), .o (n8056) );
  buffer buf_n8057( .i (n8056), .o (n8057) );
  buffer buf_n8058( .i (n8057), .o (n8058) );
  buffer buf_n8059( .i (n8058), .o (n8059) );
  buffer buf_n8060( .i (n8059), .o (n8060) );
  buffer buf_n8061( .i (n8060), .o (n8061) );
  buffer buf_n8062( .i (n8061), .o (n8062) );
  buffer buf_n8063( .i (n8062), .o (n8063) );
  buffer buf_n8064( .i (n8063), .o (n8064) );
  buffer buf_n8065( .i (n8064), .o (n8065) );
  buffer buf_n8066( .i (n8065), .o (n8066) );
  buffer buf_n8067( .i (n8066), .o (n8067) );
  buffer buf_n8068( .i (n8067), .o (n8068) );
  buffer buf_n8069( .i (n8068), .o (n8069) );
  buffer buf_n8070( .i (n8069), .o (n8070) );
  buffer buf_n8071( .i (n8070), .o (n8071) );
  buffer buf_n8072( .i (n8071), .o (n8072) );
  buffer buf_n8073( .i (n8072), .o (n8073) );
  buffer buf_n8074( .i (n8073), .o (n8074) );
  buffer buf_n8075( .i (n8074), .o (n8075) );
  buffer buf_n8076( .i (n8075), .o (n8076) );
  buffer buf_n8077( .i (n8076), .o (n8077) );
  buffer buf_n8078( .i (n8077), .o (n8078) );
  buffer buf_n8079( .i (n8078), .o (n8079) );
  buffer buf_n8080( .i (n8079), .o (n8080) );
  buffer buf_n8081( .i (n8080), .o (n8081) );
  buffer buf_n8082( .i (n8081), .o (n8082) );
  buffer buf_n8083( .i (n8082), .o (n8083) );
  buffer buf_n8084( .i (n8083), .o (n8084) );
  buffer buf_n8085( .i (n8084), .o (n8085) );
  buffer buf_n8086( .i (n8085), .o (n8086) );
  buffer buf_n8087( .i (n8086), .o (n8087) );
  buffer buf_n8088( .i (n8087), .o (n8088) );
  buffer buf_n8089( .i (n8088), .o (n8089) );
  buffer buf_n8090( .i (n8089), .o (n8090) );
  buffer buf_n8091( .i (n8090), .o (n8091) );
  buffer buf_n8092( .i (n8091), .o (n8092) );
  buffer buf_n8093( .i (n8092), .o (n8093) );
  buffer buf_n4796( .i (n4795), .o (n4796) );
  buffer buf_n4797( .i (n4796), .o (n4797) );
  buffer buf_n4798( .i (n4797), .o (n4798) );
  buffer buf_n4799( .i (n4798), .o (n4799) );
  buffer buf_n4800( .i (n4799), .o (n4800) );
  buffer buf_n4801( .i (n4800), .o (n4801) );
  buffer buf_n4802( .i (n4801), .o (n4802) );
  buffer buf_n4803( .i (n4802), .o (n4803) );
  buffer buf_n4804( .i (n4803), .o (n4804) );
  buffer buf_n4805( .i (n4804), .o (n4805) );
  buffer buf_n4806( .i (n4805), .o (n4806) );
  buffer buf_n4807( .i (n4806), .o (n4807) );
  buffer buf_n4808( .i (n4807), .o (n4808) );
  buffer buf_n4809( .i (n4808), .o (n4809) );
  buffer buf_n4810( .i (n4809), .o (n4810) );
  buffer buf_n4811( .i (n4810), .o (n4811) );
  buffer buf_n4812( .i (n4811), .o (n4812) );
  buffer buf_n4813( .i (n4812), .o (n4813) );
  buffer buf_n4814( .i (n4813), .o (n4814) );
  buffer buf_n4815( .i (n4814), .o (n4815) );
  buffer buf_n4816( .i (n4815), .o (n4816) );
  buffer buf_n4817( .i (n4816), .o (n4817) );
  buffer buf_n4818( .i (n4817), .o (n4818) );
  buffer buf_n4819( .i (n4818), .o (n4819) );
  buffer buf_n4820( .i (n4819), .o (n4820) );
  buffer buf_n4821( .i (n4820), .o (n4821) );
  buffer buf_n4822( .i (n4821), .o (n4822) );
  buffer buf_n4823( .i (n4822), .o (n4823) );
  buffer buf_n4824( .i (n4823), .o (n4824) );
  buffer buf_n4825( .i (n4824), .o (n4825) );
  buffer buf_n4826( .i (n4825), .o (n4826) );
  buffer buf_n5950( .i (n5949), .o (n5950) );
  buffer buf_n5951( .i (n5950), .o (n5951) );
  buffer buf_n5952( .i (n5951), .o (n5952) );
  buffer buf_n5953( .i (n5952), .o (n5953) );
  assign n8094 = ~n4826 & n5953 ;
  buffer buf_n8095( .i (n8094), .o (n8095) );
  assign n8096 = n4826 & ~n5953 ;
  buffer buf_n8097( .i (n8096), .o (n8097) );
  assign n8098 = n8095 | n8097 ;
  buffer buf_n8099( .i (n8098), .o (n8099) );
  buffer buf_n8100( .i (n8099), .o (n8100) );
  buffer buf_n8101( .i (n8100), .o (n8101) );
  buffer buf_n8102( .i (n8101), .o (n8102) );
  buffer buf_n8103( .i (n8102), .o (n8103) );
  buffer buf_n8104( .i (n8103), .o (n8104) );
  buffer buf_n8105( .i (n8104), .o (n8105) );
  buffer buf_n8106( .i (n8105), .o (n8106) );
  buffer buf_n8107( .i (n8106), .o (n8107) );
  buffer buf_n8108( .i (n8107), .o (n8108) );
  buffer buf_n8109( .i (n8108), .o (n8109) );
  buffer buf_n8110( .i (n8109), .o (n8110) );
  buffer buf_n8111( .i (n8110), .o (n8111) );
  buffer buf_n8112( .i (n8111), .o (n8112) );
  buffer buf_n8113( .i (n8112), .o (n8113) );
  buffer buf_n8114( .i (n8113), .o (n8114) );
  buffer buf_n8115( .i (n8114), .o (n8115) );
  buffer buf_n8116( .i (n8115), .o (n8116) );
  buffer buf_n8117( .i (n8116), .o (n8117) );
  buffer buf_n8118( .i (n8117), .o (n8118) );
  buffer buf_n5968( .i (n5967), .o (n5968) );
  buffer buf_n5969( .i (n5968), .o (n5969) );
  buffer buf_n5970( .i (n5969), .o (n5970) );
  buffer buf_n5971( .i (n5970), .o (n5971) );
  buffer buf_n5972( .i (n5971), .o (n5972) );
  buffer buf_n5973( .i (n5972), .o (n5973) );
  buffer buf_n6019( .i (n6018), .o (n6019) );
  buffer buf_n6020( .i (n6019), .o (n6020) );
  buffer buf_n6021( .i (n6020), .o (n6021) );
  buffer buf_n6022( .i (n6021), .o (n6022) );
  buffer buf_n6023( .i (n6022), .o (n6023) );
  buffer buf_n6024( .i (n6023), .o (n6024) );
  buffer buf_n6025( .i (n6024), .o (n6025) );
  buffer buf_n6026( .i (n6025), .o (n6026) );
  buffer buf_n6027( .i (n6026), .o (n6027) );
  buffer buf_n6028( .i (n6027), .o (n6028) );
  buffer buf_n6029( .i (n6028), .o (n6029) );
  buffer buf_n6030( .i (n6029), .o (n6030) );
  buffer buf_n6031( .i (n6030), .o (n6031) );
  buffer buf_n6032( .i (n6031), .o (n6032) );
  buffer buf_n6033( .i (n6032), .o (n6033) );
  buffer buf_n6034( .i (n6033), .o (n6034) );
  buffer buf_n6035( .i (n6034), .o (n6035) );
  buffer buf_n6036( .i (n6035), .o (n6036) );
  buffer buf_n6037( .i (n6036), .o (n6037) );
  buffer buf_n6038( .i (n6037), .o (n6038) );
  buffer buf_n6039( .i (n6038), .o (n6039) );
  buffer buf_n6040( .i (n6039), .o (n6040) );
  buffer buf_n6041( .i (n6040), .o (n6041) );
  buffer buf_n6042( .i (n6041), .o (n6042) );
  buffer buf_n6043( .i (n6042), .o (n6043) );
  buffer buf_n6044( .i (n6043), .o (n6044) );
  buffer buf_n6045( .i (n6044), .o (n6045) );
  buffer buf_n6046( .i (n6045), .o (n6046) );
  buffer buf_n6047( .i (n6046), .o (n6047) );
  buffer buf_n6048( .i (n6047), .o (n6048) );
  buffer buf_n6049( .i (n6048), .o (n6049) );
  buffer buf_n6050( .i (n6049), .o (n6050) );
  buffer buf_n6051( .i (n6050), .o (n6051) );
  buffer buf_n6052( .i (n6051), .o (n6052) );
  buffer buf_n6053( .i (n6052), .o (n6053) );
  buffer buf_n6054( .i (n6053), .o (n6054) );
  buffer buf_n6055( .i (n6054), .o (n6055) );
  buffer buf_n6056( .i (n6055), .o (n6056) );
  buffer buf_n6057( .i (n6056), .o (n6057) );
  buffer buf_n6058( .i (n6057), .o (n6058) );
  buffer buf_n6059( .i (n6058), .o (n6059) );
  buffer buf_n6060( .i (n6059), .o (n6060) );
  assign n8119 = ~n5973 & n6060 ;
  buffer buf_n8120( .i (n8119), .o (n8120) );
  assign n8121 = n5973 & ~n6060 ;
  buffer buf_n8122( .i (n8121), .o (n8122) );
  assign n8123 = n8120 | n8122 ;
  buffer buf_n8124( .i (n8123), .o (n8124) );
  buffer buf_n8125( .i (n8124), .o (n8125) );
  buffer buf_n8126( .i (n8125), .o (n8126) );
  buffer buf_n8127( .i (n8126), .o (n8127) );
  buffer buf_n8128( .i (n8127), .o (n8128) );
  buffer buf_n8129( .i (n8128), .o (n8129) );
  buffer buf_n8130( .i (n8129), .o (n8130) );
  buffer buf_n8131( .i (n8130), .o (n8131) );
  buffer buf_n8132( .i (n8131), .o (n8132) );
  buffer buf_n6565( .i (n6564), .o (n6565) );
  buffer buf_n6566( .i (n6565), .o (n6566) );
  buffer buf_n6567( .i (n6566), .o (n6567) );
  buffer buf_n6568( .i (n6567), .o (n6568) );
  buffer buf_n6569( .i (n6568), .o (n6569) );
  buffer buf_n6570( .i (n6569), .o (n6570) );
  buffer buf_n6571( .i (n6570), .o (n6571) );
  buffer buf_n6572( .i (n6571), .o (n6572) );
  buffer buf_n6573( .i (n6572), .o (n6573) );
  buffer buf_n6574( .i (n6573), .o (n6574) );
  buffer buf_n6575( .i (n6574), .o (n6575) );
  buffer buf_n6576( .i (n6575), .o (n6576) );
  buffer buf_n6577( .i (n6576), .o (n6577) );
  buffer buf_n6578( .i (n6577), .o (n6578) );
  buffer buf_n6579( .i (n6578), .o (n6579) );
  buffer buf_n6580( .i (n6579), .o (n6580) );
  buffer buf_n6581( .i (n6580), .o (n6581) );
  buffer buf_n6582( .i (n6581), .o (n6582) );
  buffer buf_n6583( .i (n6582), .o (n6583) );
  buffer buf_n6584( .i (n6583), .o (n6584) );
  buffer buf_n6585( .i (n6584), .o (n6585) );
  buffer buf_n6586( .i (n6585), .o (n6586) );
  buffer buf_n6587( .i (n6586), .o (n6587) );
  buffer buf_n6588( .i (n6587), .o (n6588) );
  buffer buf_n6589( .i (n6588), .o (n6589) );
  buffer buf_n6590( .i (n6589), .o (n6590) );
  buffer buf_n6591( .i (n6590), .o (n6591) );
  buffer buf_n6592( .i (n6591), .o (n6592) );
  buffer buf_n6593( .i (n6592), .o (n6593) );
  buffer buf_n6594( .i (n6593), .o (n6594) );
  buffer buf_n6595( .i (n6594), .o (n6595) );
  buffer buf_n6596( .i (n6595), .o (n6596) );
  buffer buf_n6597( .i (n6596), .o (n6597) );
  buffer buf_n6598( .i (n6597), .o (n6598) );
  buffer buf_n6599( .i (n6598), .o (n6599) );
  buffer buf_n6600( .i (n6599), .o (n6600) );
  buffer buf_n6601( .i (n6600), .o (n6601) );
  buffer buf_n6602( .i (n6601), .o (n6602) );
  buffer buf_n6603( .i (n6602), .o (n6603) );
  buffer buf_n6604( .i (n6603), .o (n6604) );
  buffer buf_n6605( .i (n6604), .o (n6605) );
  buffer buf_n6606( .i (n6605), .o (n6606) );
  buffer buf_n6607( .i (n6606), .o (n6607) );
  assign n8133 = ~n4561 & n4577 ;
  buffer buf_n8134( .i (n8133), .o (n8134) );
  buffer buf_n8135( .i (n8134), .o (n8135) );
  buffer buf_n8136( .i (n8135), .o (n8136) );
  buffer buf_n8137( .i (n8136), .o (n8137) );
  buffer buf_n8138( .i (n8137), .o (n8138) );
  buffer buf_n8139( .i (n8138), .o (n8139) );
  buffer buf_n8140( .i (n8139), .o (n8140) );
  buffer buf_n8141( .i (n8140), .o (n8141) );
  buffer buf_n8142( .i (n8141), .o (n8142) );
  buffer buf_n8143( .i (n8142), .o (n8143) );
  buffer buf_n8144( .i (n8143), .o (n8144) );
  buffer buf_n8145( .i (n8144), .o (n8145) );
  buffer buf_n8146( .i (n8145), .o (n8146) );
  buffer buf_n8147( .i (n8146), .o (n8147) );
  buffer buf_n8148( .i (n8147), .o (n8148) );
  buffer buf_n8149( .i (n8148), .o (n8149) );
  buffer buf_n8150( .i (n8149), .o (n8150) );
  buffer buf_n8151( .i (n8150), .o (n8151) );
  buffer buf_n8152( .i (n8151), .o (n8152) );
  buffer buf_n8153( .i (n8152), .o (n8153) );
  buffer buf_n8154( .i (n8153), .o (n8154) );
  buffer buf_n8155( .i (n8154), .o (n8155) );
  buffer buf_n8156( .i (n8155), .o (n8156) );
  buffer buf_n8157( .i (n8156), .o (n8157) );
  buffer buf_n8158( .i (n8157), .o (n8158) );
  buffer buf_n8159( .i (n8158), .o (n8159) );
  buffer buf_n8160( .i (n8159), .o (n8160) );
  buffer buf_n8161( .i (n8160), .o (n8161) );
  buffer buf_n8162( .i (n8161), .o (n8162) );
  buffer buf_n8163( .i (n8162), .o (n8163) );
  buffer buf_n8164( .i (n8163), .o (n8164) );
  buffer buf_n8165( .i (n8164), .o (n8165) );
  buffer buf_n8166( .i (n8165), .o (n8166) );
  buffer buf_n4753( .i (n4752), .o (n4753) );
  buffer buf_n4754( .i (n4753), .o (n4754) );
  buffer buf_n4755( .i (n4754), .o (n4755) );
  buffer buf_n4756( .i (n4755), .o (n4756) );
  buffer buf_n4757( .i (n4756), .o (n4757) );
  buffer buf_n4758( .i (n4757), .o (n4758) );
  buffer buf_n4759( .i (n4758), .o (n4759) );
  buffer buf_n4760( .i (n4759), .o (n4760) );
  buffer buf_n4761( .i (n4760), .o (n4761) );
  buffer buf_n4762( .i (n4761), .o (n4762) );
  buffer buf_n4763( .i (n4762), .o (n4763) );
  buffer buf_n4764( .i (n4763), .o (n4764) );
  buffer buf_n4765( .i (n4764), .o (n4765) );
  buffer buf_n4766( .i (n4765), .o (n4766) );
  buffer buf_n4767( .i (n4766), .o (n4767) );
  buffer buf_n4768( .i (n4767), .o (n4768) );
  buffer buf_n4769( .i (n4768), .o (n4769) );
  buffer buf_n4770( .i (n4769), .o (n4770) );
  buffer buf_n4771( .i (n4770), .o (n4771) );
  buffer buf_n4772( .i (n4771), .o (n4772) );
  buffer buf_n4773( .i (n4772), .o (n4773) );
  buffer buf_n4900( .i (n4899), .o (n4900) );
  buffer buf_n4901( .i (n4900), .o (n4901) );
  buffer buf_n4902( .i (n4901), .o (n4902) );
  buffer buf_n4903( .i (n4902), .o (n4903) );
  buffer buf_n4904( .i (n4903), .o (n4904) );
  buffer buf_n4905( .i (n4904), .o (n4905) );
  buffer buf_n4906( .i (n4905), .o (n4906) );
  buffer buf_n4907( .i (n4906), .o (n4907) );
  buffer buf_n4908( .i (n4907), .o (n4908) );
  buffer buf_n4909( .i (n4908), .o (n4909) );
  buffer buf_n4910( .i (n4909), .o (n4910) );
  buffer buf_n4911( .i (n4910), .o (n4911) );
  buffer buf_n4912( .i (n4911), .o (n4912) );
  buffer buf_n4913( .i (n4912), .o (n4913) );
  buffer buf_n4914( .i (n4913), .o (n4914) );
  buffer buf_n4915( .i (n4914), .o (n4915) );
  buffer buf_n4916( .i (n4915), .o (n4916) );
  buffer buf_n4917( .i (n4916), .o (n4917) );
  buffer buf_n4918( .i (n4917), .o (n4918) );
  buffer buf_n4919( .i (n4918), .o (n4919) );
  buffer buf_n4920( .i (n4919), .o (n4920) );
  buffer buf_n4921( .i (n4920), .o (n4921) );
  assign n8167 = n4865 | n4927 ;
  buffer buf_n8168( .i (n8167), .o (n8168) );
  buffer buf_n8169( .i (n8168), .o (n8169) );
  buffer buf_n8170( .i (n8169), .o (n8170) );
  buffer buf_n8171( .i (n8170), .o (n8171) );
  buffer buf_n8172( .i (n8171), .o (n8172) );
  buffer buf_n8173( .i (n8172), .o (n8173) );
  buffer buf_n8174( .i (n8173), .o (n8174) );
  buffer buf_n8175( .i (n8174), .o (n8175) );
  buffer buf_n8176( .i (n8175), .o (n8176) );
  buffer buf_n8177( .i (n8176), .o (n8177) );
  buffer buf_n8178( .i (n8177), .o (n8178) );
  buffer buf_n8179( .i (n8178), .o (n8179) );
  buffer buf_n8180( .i (n8179), .o (n8180) );
  buffer buf_n8181( .i (n8180), .o (n8181) );
  buffer buf_n8182( .i (n8181), .o (n8182) );
  buffer buf_n8183( .i (n8182), .o (n8183) );
  buffer buf_n8184( .i (n8183), .o (n8184) );
  buffer buf_n8185( .i (n8184), .o (n8185) );
  buffer buf_n8186( .i (n8185), .o (n8186) );
  buffer buf_n8187( .i (n8186), .o (n8187) );
  buffer buf_n8188( .i (n8187), .o (n8188) );
  buffer buf_n8189( .i (n8188), .o (n8189) );
  buffer buf_n8190( .i (n8189), .o (n8190) );
  buffer buf_n8191( .i (n8190), .o (n8191) );
  assign n8192 = n5949 & ~n8191 ;
  buffer buf_n8193( .i (n8192), .o (n8193) );
  assign n8194 = ~n4921 & n8193 ;
  assign n8195 = n4773 | n8194 ;
  buffer buf_n8196( .i (n8195), .o (n8196) );
  assign n8197 = n8166 & ~n8196 ;
  assign n8198 = ~n8166 & n8196 ;
  assign n8199 = n8197 | n8198 ;
  buffer buf_n8200( .i (n8199), .o (n8200) );
  buffer buf_n8201( .i (n8200), .o (n8201) );
  buffer buf_n8202( .i (n8201), .o (n8202) );
  buffer buf_n8203( .i (n8202), .o (n8203) );
  buffer buf_n8204( .i (n8203), .o (n8204) );
  buffer buf_n8205( .i (n8204), .o (n8205) );
  buffer buf_n8206( .i (n8205), .o (n8206) );
  buffer buf_n8207( .i (n8206), .o (n8207) );
  buffer buf_n8208( .i (n8207), .o (n8208) );
  buffer buf_n8209( .i (n8208), .o (n8209) );
  buffer buf_n8210( .i (n8209), .o (n8210) );
  buffer buf_n8211( .i (n8210), .o (n8211) );
  buffer buf_n8212( .i (n8211), .o (n8212) );
  buffer buf_n8213( .i (n8212), .o (n8213) );
  buffer buf_n8214( .i (n8213), .o (n8214) );
  buffer buf_n8215( .i (n8214), .o (n8215) );
  buffer buf_n8216( .i (n8215), .o (n8216) );
  buffer buf_n8217( .i (n8216), .o (n8217) );
  buffer buf_n8218( .i (n8217), .o (n8218) );
  buffer buf_n8219( .i (n8218), .o (n8219) );
  buffer buf_n4922( .i (n4921), .o (n4922) );
  buffer buf_n4923( .i (n4922), .o (n4923) );
  buffer buf_n4727( .i (n4726), .o (n4727) );
  buffer buf_n4728( .i (n4727), .o (n4728) );
  buffer buf_n4729( .i (n4728), .o (n4729) );
  buffer buf_n4730( .i (n4729), .o (n4730) );
  buffer buf_n4731( .i (n4730), .o (n4731) );
  buffer buf_n4732( .i (n4731), .o (n4732) );
  buffer buf_n4733( .i (n4732), .o (n4733) );
  buffer buf_n4734( .i (n4733), .o (n4734) );
  buffer buf_n4735( .i (n4734), .o (n4735) );
  buffer buf_n4736( .i (n4735), .o (n4736) );
  buffer buf_n4737( .i (n4736), .o (n4737) );
  buffer buf_n4738( .i (n4737), .o (n4738) );
  buffer buf_n4739( .i (n4738), .o (n4739) );
  buffer buf_n4740( .i (n4739), .o (n4740) );
  buffer buf_n4741( .i (n4740), .o (n4741) );
  buffer buf_n4742( .i (n4741), .o (n4742) );
  buffer buf_n4743( .i (n4742), .o (n4743) );
  buffer buf_n4744( .i (n4743), .o (n4744) );
  buffer buf_n4745( .i (n4744), .o (n4745) );
  buffer buf_n4746( .i (n4745), .o (n4746) );
  buffer buf_n4747( .i (n4746), .o (n4747) );
  buffer buf_n4748( .i (n4747), .o (n4748) );
  buffer buf_n4749( .i (n4748), .o (n4749) );
  assign n8220 = n4749 | n8193 ;
  buffer buf_n8221( .i (n8220), .o (n8221) );
  assign n8222 = n4923 | n8221 ;
  assign n8223 = n4923 & n8221 ;
  assign n8224 = n8222 & ~n8223 ;
  buffer buf_n8225( .i (n8224), .o (n8225) );
  buffer buf_n8226( .i (n8225), .o (n8226) );
  buffer buf_n8227( .i (n8226), .o (n8227) );
  buffer buf_n8228( .i (n8227), .o (n8228) );
  buffer buf_n8229( .i (n8228), .o (n8229) );
  buffer buf_n8230( .i (n8229), .o (n8230) );
  buffer buf_n8231( .i (n8230), .o (n8231) );
  buffer buf_n8232( .i (n8231), .o (n8232) );
  buffer buf_n8233( .i (n8232), .o (n8233) );
  buffer buf_n8234( .i (n8233), .o (n8234) );
  buffer buf_n8235( .i (n8234), .o (n8235) );
  buffer buf_n8236( .i (n8235), .o (n8236) );
  buffer buf_n8237( .i (n8236), .o (n8237) );
  buffer buf_n8238( .i (n8237), .o (n8238) );
  buffer buf_n8239( .i (n8238), .o (n8239) );
  buffer buf_n8240( .i (n8239), .o (n8240) );
  buffer buf_n8241( .i (n8240), .o (n8241) );
  buffer buf_n8242( .i (n8241), .o (n8242) );
  buffer buf_n8243( .i (n8242), .o (n8243) );
  buffer buf_n8244( .i (n8243), .o (n8244) );
  buffer buf_n8245( .i (n8244), .o (n8245) );
  buffer buf_n4933( .i (n4932), .o (n4933) );
  buffer buf_n4934( .i (n4933), .o (n4934) );
  buffer buf_n4935( .i (n4934), .o (n4935) );
  buffer buf_n4936( .i (n4935), .o (n4936) );
  buffer buf_n4937( .i (n4936), .o (n4937) );
  buffer buf_n4938( .i (n4937), .o (n4938) );
  buffer buf_n4939( .i (n4938), .o (n4939) );
  buffer buf_n4940( .i (n4939), .o (n4940) );
  buffer buf_n4941( .i (n4940), .o (n4941) );
  buffer buf_n4942( .i (n4941), .o (n4942) );
  buffer buf_n4943( .i (n4942), .o (n4943) );
  buffer buf_n4944( .i (n4943), .o (n4944) );
  buffer buf_n4945( .i (n4944), .o (n4945) );
  buffer buf_n4946( .i (n4945), .o (n4946) );
  buffer buf_n4947( .i (n4946), .o (n4947) );
  buffer buf_n4948( .i (n4947), .o (n4948) );
  buffer buf_n4949( .i (n4948), .o (n4949) );
  buffer buf_n4950( .i (n4949), .o (n4950) );
  buffer buf_n4951( .i (n4950), .o (n4951) );
  buffer buf_n4952( .i (n4951), .o (n4952) );
  buffer buf_n4953( .i (n4952), .o (n4953) );
  buffer buf_n4954( .i (n4953), .o (n4954) );
  buffer buf_n4955( .i (n4954), .o (n4955) );
  buffer buf_n4697( .i (n4696), .o (n4697) );
  buffer buf_n4698( .i (n4697), .o (n4698) );
  buffer buf_n4699( .i (n4698), .o (n4699) );
  buffer buf_n4700( .i (n4699), .o (n4700) );
  buffer buf_n4701( .i (n4700), .o (n4701) );
  buffer buf_n4702( .i (n4701), .o (n4702) );
  buffer buf_n4703( .i (n4702), .o (n4703) );
  buffer buf_n4704( .i (n4703), .o (n4704) );
  buffer buf_n4705( .i (n4704), .o (n4705) );
  buffer buf_n4706( .i (n4705), .o (n4706) );
  buffer buf_n4707( .i (n4706), .o (n4707) );
  buffer buf_n4708( .i (n4707), .o (n4708) );
  buffer buf_n4709( .i (n4708), .o (n4709) );
  buffer buf_n4710( .i (n4709), .o (n4710) );
  buffer buf_n4711( .i (n4710), .o (n4711) );
  buffer buf_n4712( .i (n4711), .o (n4712) );
  buffer buf_n4713( .i (n4712), .o (n4713) );
  buffer buf_n4714( .i (n4713), .o (n4714) );
  buffer buf_n4715( .i (n4714), .o (n4715) );
  buffer buf_n4716( .i (n4715), .o (n4716) );
  buffer buf_n4717( .i (n4716), .o (n4717) );
  buffer buf_n4718( .i (n4717), .o (n4718) );
  buffer buf_n4719( .i (n4718), .o (n4719) );
  buffer buf_n4720( .i (n4719), .o (n4720) );
  buffer buf_n4721( .i (n4720), .o (n4721) );
  buffer buf_n4722( .i (n4721), .o (n4722) );
  buffer buf_n4873( .i (n4872), .o (n4873) );
  buffer buf_n4874( .i (n4873), .o (n4874) );
  buffer buf_n4875( .i (n4874), .o (n4875) );
  buffer buf_n4876( .i (n4875), .o (n4876) );
  buffer buf_n4877( .i (n4876), .o (n4877) );
  buffer buf_n4878( .i (n4877), .o (n4878) );
  buffer buf_n4879( .i (n4878), .o (n4879) );
  buffer buf_n4880( .i (n4879), .o (n4880) );
  buffer buf_n4881( .i (n4880), .o (n4881) );
  buffer buf_n4882( .i (n4881), .o (n4882) );
  buffer buf_n4883( .i (n4882), .o (n4883) );
  buffer buf_n4884( .i (n4883), .o (n4884) );
  buffer buf_n4885( .i (n4884), .o (n4885) );
  buffer buf_n4886( .i (n4885), .o (n4886) );
  buffer buf_n4887( .i (n4886), .o (n4887) );
  buffer buf_n4888( .i (n4887), .o (n4888) );
  buffer buf_n4889( .i (n4888), .o (n4889) );
  buffer buf_n4890( .i (n4889), .o (n4890) );
  assign n8246 = ~n4890 & n5949 ;
  assign n8247 = n4722 | n8246 ;
  buffer buf_n8248( .i (n8247), .o (n8248) );
  assign n8249 = n4955 & n8248 ;
  assign n8250 = n4955 | n8248 ;
  assign n8251 = ~n8249 & n8250 ;
  buffer buf_n8252( .i (n8251), .o (n8252) );
  buffer buf_n8253( .i (n8252), .o (n8253) );
  buffer buf_n8254( .i (n8253), .o (n8254) );
  buffer buf_n8255( .i (n8254), .o (n8255) );
  buffer buf_n8256( .i (n8255), .o (n8256) );
  buffer buf_n8257( .i (n8256), .o (n8257) );
  buffer buf_n8258( .i (n8257), .o (n8258) );
  buffer buf_n8259( .i (n8258), .o (n8259) );
  buffer buf_n8260( .i (n8259), .o (n8260) );
  buffer buf_n8261( .i (n8260), .o (n8261) );
  buffer buf_n8262( .i (n8261), .o (n8262) );
  buffer buf_n8263( .i (n8262), .o (n8263) );
  buffer buf_n8264( .i (n8263), .o (n8264) );
  buffer buf_n8265( .i (n8264), .o (n8265) );
  buffer buf_n8266( .i (n8265), .o (n8266) );
  buffer buf_n8267( .i (n8266), .o (n8267) );
  buffer buf_n8268( .i (n8267), .o (n8268) );
  buffer buf_n8269( .i (n8268), .o (n8269) );
  buffer buf_n8270( .i (n8269), .o (n8270) );
  buffer buf_n8271( .i (n8270), .o (n8271) );
  buffer buf_n8272( .i (n8271), .o (n8272) );
  buffer buf_n8273( .i (n8272), .o (n8273) );
  buffer buf_n4829( .i (n4828), .o (n4829) );
  buffer buf_n4830( .i (n4829), .o (n4830) );
  buffer buf_n4831( .i (n4830), .o (n4831) );
  buffer buf_n4832( .i (n4831), .o (n4832) );
  buffer buf_n4833( .i (n4832), .o (n4833) );
  buffer buf_n4834( .i (n4833), .o (n4834) );
  buffer buf_n4835( .i (n4834), .o (n4835) );
  buffer buf_n4836( .i (n4835), .o (n4836) );
  buffer buf_n4837( .i (n4836), .o (n4837) );
  buffer buf_n4838( .i (n4837), .o (n4838) );
  buffer buf_n4839( .i (n4838), .o (n4839) );
  buffer buf_n4840( .i (n4839), .o (n4840) );
  buffer buf_n4841( .i (n4840), .o (n4841) );
  buffer buf_n4842( .i (n4841), .o (n4842) );
  buffer buf_n4843( .i (n4842), .o (n4843) );
  buffer buf_n4844( .i (n4843), .o (n4844) );
  buffer buf_n4845( .i (n4844), .o (n4845) );
  buffer buf_n4846( .i (n4845), .o (n4846) );
  buffer buf_n4847( .i (n4846), .o (n4847) );
  buffer buf_n4848( .i (n4847), .o (n4848) );
  buffer buf_n4849( .i (n4848), .o (n4849) );
  buffer buf_n4850( .i (n4849), .o (n4850) );
  buffer buf_n4851( .i (n4850), .o (n4851) );
  buffer buf_n4852( .i (n4851), .o (n4852) );
  buffer buf_n4853( .i (n4852), .o (n4853) );
  buffer buf_n4854( .i (n4853), .o (n4854) );
  buffer buf_n4855( .i (n4854), .o (n4855) );
  buffer buf_n4856( .i (n4855), .o (n4856) );
  buffer buf_n4857( .i (n4856), .o (n4857) );
  buffer buf_n4858( .i (n4857), .o (n4858) );
  buffer buf_n4859( .i (n4858), .o (n4859) );
  buffer buf_n4860( .i (n4859), .o (n4860) );
  buffer buf_n4861( .i (n4860), .o (n4861) );
  buffer buf_n4862( .i (n4861), .o (n4862) );
  buffer buf_n4863( .i (n4862), .o (n4863) );
  buffer buf_n4656( .i (n4655), .o (n4656) );
  buffer buf_n4657( .i (n4656), .o (n4657) );
  buffer buf_n4658( .i (n4657), .o (n4658) );
  buffer buf_n4659( .i (n4658), .o (n4659) );
  buffer buf_n4660( .i (n4659), .o (n4660) );
  buffer buf_n4661( .i (n4660), .o (n4661) );
  buffer buf_n4662( .i (n4661), .o (n4662) );
  buffer buf_n4663( .i (n4662), .o (n4663) );
  buffer buf_n4664( .i (n4663), .o (n4664) );
  buffer buf_n4665( .i (n4664), .o (n4665) );
  buffer buf_n4666( .i (n4665), .o (n4666) );
  buffer buf_n4667( .i (n4666), .o (n4667) );
  buffer buf_n4668( .i (n4667), .o (n4668) );
  buffer buf_n4669( .i (n4668), .o (n4669) );
  buffer buf_n4670( .i (n4669), .o (n4670) );
  buffer buf_n4671( .i (n4670), .o (n4671) );
  buffer buf_n4672( .i (n4671), .o (n4672) );
  buffer buf_n4673( .i (n4672), .o (n4673) );
  buffer buf_n4674( .i (n4673), .o (n4674) );
  buffer buf_n4675( .i (n4674), .o (n4675) );
  buffer buf_n4676( .i (n4675), .o (n4676) );
  buffer buf_n4677( .i (n4676), .o (n4677) );
  buffer buf_n4678( .i (n4677), .o (n4678) );
  buffer buf_n4679( .i (n4678), .o (n4679) );
  buffer buf_n4680( .i (n4679), .o (n4680) );
  buffer buf_n4681( .i (n4680), .o (n4681) );
  buffer buf_n4682( .i (n4681), .o (n4682) );
  buffer buf_n4683( .i (n4682), .o (n4683) );
  buffer buf_n4684( .i (n4683), .o (n4684) );
  buffer buf_n4685( .i (n4684), .o (n4685) );
  buffer buf_n4686( .i (n4685), .o (n4686) );
  buffer buf_n4687( .i (n4686), .o (n4687) );
  buffer buf_n4688( .i (n4687), .o (n4688) );
  buffer buf_n4689( .i (n4688), .o (n4689) );
  buffer buf_n4690( .i (n4689), .o (n4690) );
  assign n8274 = n4690 | n8095 ;
  buffer buf_n8275( .i (n8274), .o (n8275) );
  assign n8276 = n4863 | n8275 ;
  assign n8277 = n4863 & n8275 ;
  assign n8278 = n8276 & ~n8277 ;
  buffer buf_n8279( .i (n8278), .o (n8279) );
  buffer buf_n8280( .i (n8279), .o (n8280) );
  buffer buf_n8281( .i (n8280), .o (n8281) );
  buffer buf_n8282( .i (n8281), .o (n8282) );
  buffer buf_n8283( .i (n8282), .o (n8283) );
  buffer buf_n8284( .i (n8283), .o (n8284) );
  buffer buf_n8285( .i (n8284), .o (n8285) );
  buffer buf_n8286( .i (n8285), .o (n8286) );
  buffer buf_n8287( .i (n8286), .o (n8287) );
  buffer buf_n8288( .i (n8287), .o (n8288) );
  buffer buf_n8289( .i (n8288), .o (n8289) );
  buffer buf_n8290( .i (n8289), .o (n8290) );
  buffer buf_n8291( .i (n8290), .o (n8291) );
  buffer buf_n8292( .i (n8291), .o (n8292) );
  buffer buf_n8293( .i (n8292), .o (n8293) );
  buffer buf_n8294( .i (n8293), .o (n8294) );
  buffer buf_n8295( .i (n8294), .o (n8295) );
  buffer buf_n4202( .i (n4201), .o (n4202) );
  buffer buf_n4203( .i (n4202), .o (n4203) );
  buffer buf_n4204( .i (n4203), .o (n4204) );
  buffer buf_n4205( .i (n4204), .o (n4205) );
  buffer buf_n4206( .i (n4205), .o (n4206) );
  buffer buf_n4207( .i (n4206), .o (n4207) );
  buffer buf_n3903( .i (n3902), .o (n3903) );
  buffer buf_n3904( .i (n3903), .o (n3904) );
  buffer buf_n3905( .i (n3904), .o (n3905) );
  buffer buf_n3906( .i (n3905), .o (n3906) );
  buffer buf_n3907( .i (n3906), .o (n3907) );
  buffer buf_n3908( .i (n3907), .o (n3908) );
  buffer buf_n3909( .i (n3908), .o (n3909) );
  buffer buf_n3910( .i (n3909), .o (n3910) );
  buffer buf_n3911( .i (n3910), .o (n3911) );
  buffer buf_n4115( .i (n4114), .o (n4115) );
  buffer buf_n4116( .i (n4115), .o (n4116) );
  buffer buf_n4117( .i (n4116), .o (n4117) );
  buffer buf_n4118( .i (n4117), .o (n4118) );
  buffer buf_n4119( .i (n4118), .o (n4119) );
  buffer buf_n4120( .i (n4119), .o (n4120) );
  buffer buf_n4121( .i (n4120), .o (n4121) );
  buffer buf_n4122( .i (n4121), .o (n4122) );
  assign n8296 = n4080 | n4122 ;
  assign n8297 = n3911 & n8296 ;
  buffer buf_n8298( .i (n8297), .o (n8298) );
  buffer buf_n8299( .i (n8298), .o (n8299) );
  buffer buf_n8300( .i (n8299), .o (n8300) );
  buffer buf_n8301( .i (n8300), .o (n8301) );
  buffer buf_n8302( .i (n8301), .o (n8302) );
  buffer buf_n8303( .i (n8302), .o (n8303) );
  buffer buf_n8304( .i (n8303), .o (n8304) );
  buffer buf_n8305( .i (n8304), .o (n8305) );
  buffer buf_n8306( .i (n8305), .o (n8306) );
  buffer buf_n8307( .i (n8306), .o (n8307) );
  buffer buf_n8308( .i (n8307), .o (n8308) );
  buffer buf_n8309( .i (n8308), .o (n8309) );
  buffer buf_n8310( .i (n8309), .o (n8310) );
  buffer buf_n8311( .i (n8310), .o (n8311) );
  buffer buf_n8312( .i (n8311), .o (n8312) );
  buffer buf_n8313( .i (n8312), .o (n8313) );
  buffer buf_n8314( .i (n8313), .o (n8314) );
  buffer buf_n8315( .i (n8314), .o (n8315) );
  buffer buf_n8316( .i (n8315), .o (n8316) );
  buffer buf_n8317( .i (n8316), .o (n8317) );
  buffer buf_n8318( .i (n8317), .o (n8318) );
  buffer buf_n8319( .i (n8318), .o (n8319) );
  buffer buf_n8320( .i (n8319), .o (n8320) );
  buffer buf_n8321( .i (n8320), .o (n8321) );
  buffer buf_n8322( .i (n8321), .o (n8322) );
  buffer buf_n8323( .i (n8322), .o (n8323) );
  buffer buf_n8324( .i (n8323), .o (n8324) );
  buffer buf_n8325( .i (n8324), .o (n8325) );
  buffer buf_n8326( .i (n8325), .o (n8326) );
  buffer buf_n8327( .i (n8326), .o (n8327) );
  buffer buf_n8328( .i (n8327), .o (n8328) );
  buffer buf_n4160( .i (n4159), .o (n4160) );
  buffer buf_n4161( .i (n4160), .o (n4161) );
  buffer buf_n4162( .i (n4161), .o (n4162) );
  assign n8329 = n4162 & n6180 ;
  assign n8330 = n8328 & ~n8329 ;
  buffer buf_n8331( .i (n8330), .o (n8331) );
  assign n8332 = n4207 & n8331 ;
  assign n8333 = n4207 | n8331 ;
  assign n8334 = ~n8332 & n8333 ;
  buffer buf_n8335( .i (n8334), .o (n8335) );
  buffer buf_n8336( .i (n8335), .o (n8336) );
  buffer buf_n8337( .i (n8336), .o (n8337) );
  buffer buf_n8338( .i (n8337), .o (n8338) );
  buffer buf_n8339( .i (n8338), .o (n8339) );
  buffer buf_n8340( .i (n8339), .o (n8340) );
  buffer buf_n8341( .i (n8340), .o (n8341) );
  buffer buf_n8342( .i (n8341), .o (n8342) );
  buffer buf_n8343( .i (n8342), .o (n8343) );
  buffer buf_n8344( .i (n8343), .o (n8344) );
  buffer buf_n8345( .i (n8344), .o (n8345) );
  buffer buf_n4163( .i (n4162), .o (n4163) );
  buffer buf_n4164( .i (n4163), .o (n4164) );
  buffer buf_n4112( .i (n4111), .o (n4112) );
  assign n8346 = n4112 & ~n6180 ;
  buffer buf_n8347( .i (n8346), .o (n8347) );
  assign n8348 = n4164 | n8347 ;
  assign n8349 = n4164 & n8347 ;
  assign n8350 = n8348 & ~n8349 ;
  buffer buf_n8351( .i (n8350), .o (n8351) );
  buffer buf_n8352( .i (n8351), .o (n8352) );
  buffer buf_n8353( .i (n8352), .o (n8353) );
  buffer buf_n8354( .i (n8353), .o (n8354) );
  buffer buf_n8355( .i (n8354), .o (n8355) );
  buffer buf_n8356( .i (n8355), .o (n8356) );
  buffer buf_n8357( .i (n8356), .o (n8357) );
  buffer buf_n8358( .i (n8357), .o (n8358) );
  buffer buf_n8359( .i (n8358), .o (n8359) );
  buffer buf_n8360( .i (n8359), .o (n8360) );
  buffer buf_n8361( .i (n8360), .o (n8361) );
  buffer buf_n8362( .i (n8361), .o (n8362) );
  buffer buf_n5978( .i (n5977), .o (n5978) );
  buffer buf_n5979( .i (n5978), .o (n5979) );
  buffer buf_n5980( .i (n5979), .o (n5980) );
  buffer buf_n5981( .i (n5980), .o (n5981) );
  buffer buf_n5982( .i (n5981), .o (n5982) );
  buffer buf_n5983( .i (n5982), .o (n5983) );
  buffer buf_n5984( .i (n5983), .o (n5984) );
  buffer buf_n5985( .i (n5984), .o (n5985) );
  buffer buf_n5986( .i (n5985), .o (n5986) );
  buffer buf_n5987( .i (n5986), .o (n5987) );
  buffer buf_n5988( .i (n5987), .o (n5988) );
  buffer buf_n5989( .i (n5988), .o (n5989) );
  buffer buf_n5990( .i (n5989), .o (n5990) );
  buffer buf_n5991( .i (n5990), .o (n5991) );
  buffer buf_n5992( .i (n5991), .o (n5992) );
  buffer buf_n5993( .i (n5992), .o (n5993) );
  buffer buf_n5994( .i (n5993), .o (n5994) );
  buffer buf_n5995( .i (n5994), .o (n5995) );
  buffer buf_n5996( .i (n5995), .o (n5996) );
  buffer buf_n5997( .i (n5996), .o (n5997) );
  buffer buf_n5998( .i (n5997), .o (n5998) );
  buffer buf_n5999( .i (n5998), .o (n5999) );
  buffer buf_n6000( .i (n5999), .o (n6000) );
  buffer buf_n6001( .i (n6000), .o (n6001) );
  buffer buf_n6002( .i (n6001), .o (n6002) );
  buffer buf_n6003( .i (n6002), .o (n6003) );
  buffer buf_n6004( .i (n6003), .o (n6004) );
  buffer buf_n6005( .i (n6004), .o (n6005) );
  buffer buf_n6006( .i (n6005), .o (n6006) );
  buffer buf_n6007( .i (n6006), .o (n6007) );
  buffer buf_n6008( .i (n6007), .o (n6008) );
  buffer buf_n6009( .i (n6008), .o (n6009) );
  buffer buf_n6010( .i (n6009), .o (n6010) );
  buffer buf_n6011( .i (n6010), .o (n6011) );
  buffer buf_n6012( .i (n6011), .o (n6012) );
  buffer buf_n6013( .i (n6012), .o (n6013) );
  buffer buf_n6014( .i (n6013), .o (n6014) );
  buffer buf_n4042( .i (n4041), .o (n4042) );
  buffer buf_n4043( .i (n4042), .o (n4043) );
  buffer buf_n4044( .i (n4043), .o (n4044) );
  buffer buf_n4045( .i (n4044), .o (n4045) );
  buffer buf_n4046( .i (n4045), .o (n4046) );
  buffer buf_n4047( .i (n4046), .o (n4047) );
  buffer buf_n4048( .i (n4047), .o (n4048) );
  buffer buf_n4049( .i (n4048), .o (n4049) );
  buffer buf_n4050( .i (n4049), .o (n4050) );
  buffer buf_n4051( .i (n4050), .o (n4051) );
  buffer buf_n4052( .i (n4051), .o (n4052) );
  buffer buf_n4053( .i (n4052), .o (n4053) );
  buffer buf_n4054( .i (n4053), .o (n4054) );
  buffer buf_n4055( .i (n4054), .o (n4055) );
  buffer buf_n4056( .i (n4055), .o (n4056) );
  buffer buf_n4057( .i (n4056), .o (n4057) );
  buffer buf_n4058( .i (n4057), .o (n4058) );
  buffer buf_n4059( .i (n4058), .o (n4059) );
  buffer buf_n4060( .i (n4059), .o (n4060) );
  buffer buf_n4061( .i (n4060), .o (n4061) );
  buffer buf_n4062( .i (n4061), .o (n4062) );
  buffer buf_n4063( .i (n4062), .o (n4063) );
  buffer buf_n4064( .i (n4063), .o (n4064) );
  buffer buf_n4065( .i (n4064), .o (n4065) );
  buffer buf_n4066( .i (n4065), .o (n4066) );
  buffer buf_n4067( .i (n4066), .o (n4067) );
  buffer buf_n4068( .i (n4067), .o (n4068) );
  buffer buf_n4069( .i (n4068), .o (n4069) );
  buffer buf_n4070( .i (n4069), .o (n4070) );
  buffer buf_n4071( .i (n4070), .o (n4071) );
  buffer buf_n4072( .i (n4071), .o (n4072) );
  buffer buf_n4073( .i (n4072), .o (n4073) );
  buffer buf_n4074( .i (n4073), .o (n4074) );
  buffer buf_n4075( .i (n4074), .o (n4075) );
  buffer buf_n4076( .i (n4075), .o (n4076) );
  buffer buf_n6111( .i (n6110), .o (n6111) );
  buffer buf_n6112( .i (n6111), .o (n6112) );
  buffer buf_n6113( .i (n6112), .o (n6113) );
  buffer buf_n6114( .i (n6113), .o (n6114) );
  buffer buf_n6115( .i (n6114), .o (n6115) );
  buffer buf_n6116( .i (n6115), .o (n6116) );
  buffer buf_n6117( .i (n6116), .o (n6117) );
  buffer buf_n6118( .i (n6117), .o (n6118) );
  buffer buf_n6119( .i (n6118), .o (n6119) );
  buffer buf_n6120( .i (n6119), .o (n6120) );
  buffer buf_n6121( .i (n6120), .o (n6121) );
  buffer buf_n6122( .i (n6121), .o (n6122) );
  buffer buf_n6123( .i (n6122), .o (n6123) );
  buffer buf_n6124( .i (n6123), .o (n6124) );
  buffer buf_n6125( .i (n6124), .o (n6125) );
  buffer buf_n6126( .i (n6125), .o (n6126) );
  buffer buf_n6127( .i (n6126), .o (n6127) );
  buffer buf_n6128( .i (n6127), .o (n6128) );
  buffer buf_n6129( .i (n6128), .o (n6129) );
  buffer buf_n6130( .i (n6129), .o (n6130) );
  buffer buf_n6131( .i (n6130), .o (n6131) );
  buffer buf_n6132( .i (n6131), .o (n6132) );
  buffer buf_n6133( .i (n6132), .o (n6133) );
  buffer buf_n6134( .i (n6133), .o (n6134) );
  buffer buf_n6135( .i (n6134), .o (n6135) );
  buffer buf_n6136( .i (n6135), .o (n6136) );
  buffer buf_n6137( .i (n6136), .o (n6137) );
  buffer buf_n6138( .i (n6137), .o (n6138) );
  buffer buf_n6139( .i (n6138), .o (n6139) );
  buffer buf_n6140( .i (n6139), .o (n6140) );
  buffer buf_n6141( .i (n6140), .o (n6141) );
  buffer buf_n6142( .i (n6141), .o (n6142) );
  buffer buf_n6143( .i (n6142), .o (n6143) );
  buffer buf_n6144( .i (n6143), .o (n6144) );
  assign n8363 = ~n5967 & n6144 ;
  assign n8364 = n4076 & ~n8363 ;
  buffer buf_n8365( .i (n8364), .o (n8365) );
  assign n8366 = n6014 | n8365 ;
  assign n8367 = n6014 & n8365 ;
  assign n8368 = n8366 & ~n8367 ;
  buffer buf_n8369( .i (n8368), .o (n8369) );
  buffer buf_n8370( .i (n8369), .o (n8370) );
  buffer buf_n8371( .i (n8370), .o (n8371) );
  buffer buf_n8372( .i (n8371), .o (n8372) );
  buffer buf_n8373( .i (n8372), .o (n8373) );
  buffer buf_n8374( .i (n8373), .o (n8374) );
  buffer buf_n8375( .i (n8374), .o (n8375) );
  buffer buf_n8376( .i (n8375), .o (n8376) );
  buffer buf_n8377( .i (n8376), .o (n8377) );
  buffer buf_n8378( .i (n8377), .o (n8378) );
  buffer buf_n8379( .i (n8378), .o (n8379) );
  buffer buf_n8380( .i (n8379), .o (n8380) );
  buffer buf_n8381( .i (n8380), .o (n8381) );
  buffer buf_n6063( .i (n6062), .o (n6063) );
  buffer buf_n6064( .i (n6063), .o (n6064) );
  buffer buf_n6065( .i (n6064), .o (n6065) );
  buffer buf_n6066( .i (n6065), .o (n6066) );
  buffer buf_n6067( .i (n6066), .o (n6067) );
  buffer buf_n6068( .i (n6067), .o (n6068) );
  buffer buf_n6069( .i (n6068), .o (n6069) );
  buffer buf_n6070( .i (n6069), .o (n6070) );
  buffer buf_n6071( .i (n6070), .o (n6071) );
  buffer buf_n6072( .i (n6071), .o (n6072) );
  buffer buf_n6073( .i (n6072), .o (n6073) );
  buffer buf_n6074( .i (n6073), .o (n6074) );
  buffer buf_n6075( .i (n6074), .o (n6075) );
  buffer buf_n6076( .i (n6075), .o (n6076) );
  buffer buf_n6077( .i (n6076), .o (n6077) );
  buffer buf_n6078( .i (n6077), .o (n6078) );
  buffer buf_n6079( .i (n6078), .o (n6079) );
  buffer buf_n6080( .i (n6079), .o (n6080) );
  buffer buf_n6081( .i (n6080), .o (n6081) );
  buffer buf_n6082( .i (n6081), .o (n6082) );
  buffer buf_n6083( .i (n6082), .o (n6083) );
  buffer buf_n6084( .i (n6083), .o (n6084) );
  buffer buf_n6085( .i (n6084), .o (n6085) );
  buffer buf_n6086( .i (n6085), .o (n6086) );
  buffer buf_n6087( .i (n6086), .o (n6087) );
  buffer buf_n6088( .i (n6087), .o (n6088) );
  buffer buf_n6089( .i (n6088), .o (n6089) );
  buffer buf_n6090( .i (n6089), .o (n6090) );
  buffer buf_n6091( .i (n6090), .o (n6091) );
  buffer buf_n6092( .i (n6091), .o (n6092) );
  buffer buf_n6093( .i (n6092), .o (n6093) );
  buffer buf_n6094( .i (n6093), .o (n6094) );
  buffer buf_n6095( .i (n6094), .o (n6095) );
  buffer buf_n6096( .i (n6095), .o (n6096) );
  buffer buf_n6097( .i (n6096), .o (n6097) );
  buffer buf_n6098( .i (n6097), .o (n6098) );
  buffer buf_n6099( .i (n6098), .o (n6099) );
  buffer buf_n6100( .i (n6099), .o (n6100) );
  buffer buf_n6101( .i (n6100), .o (n6101) );
  buffer buf_n6102( .i (n6101), .o (n6102) );
  buffer buf_n6103( .i (n6102), .o (n6103) );
  buffer buf_n6104( .i (n6103), .o (n6104) );
  buffer buf_n6105( .i (n6104), .o (n6105) );
  buffer buf_n6106( .i (n6105), .o (n6106) );
  buffer buf_n6107( .i (n6106), .o (n6107) );
  buffer buf_n6108( .i (n6107), .o (n6108) );
  buffer buf_n3990( .i (n3989), .o (n3990) );
  buffer buf_n3991( .i (n3990), .o (n3991) );
  buffer buf_n3992( .i (n3991), .o (n3992) );
  buffer buf_n3993( .i (n3992), .o (n3993) );
  buffer buf_n3994( .i (n3993), .o (n3994) );
  buffer buf_n3995( .i (n3994), .o (n3995) );
  buffer buf_n3996( .i (n3995), .o (n3996) );
  buffer buf_n3997( .i (n3996), .o (n3997) );
  buffer buf_n3998( .i (n3997), .o (n3998) );
  buffer buf_n3999( .i (n3998), .o (n3999) );
  buffer buf_n4000( .i (n3999), .o (n4000) );
  buffer buf_n4001( .i (n4000), .o (n4001) );
  buffer buf_n4002( .i (n4001), .o (n4002) );
  buffer buf_n4003( .i (n4002), .o (n4003) );
  buffer buf_n4004( .i (n4003), .o (n4004) );
  buffer buf_n4005( .i (n4004), .o (n4005) );
  buffer buf_n4006( .i (n4005), .o (n4006) );
  buffer buf_n4007( .i (n4006), .o (n4007) );
  buffer buf_n4008( .i (n4007), .o (n4008) );
  buffer buf_n4009( .i (n4008), .o (n4009) );
  buffer buf_n4010( .i (n4009), .o (n4010) );
  buffer buf_n4011( .i (n4010), .o (n4011) );
  buffer buf_n4012( .i (n4011), .o (n4012) );
  buffer buf_n4013( .i (n4012), .o (n4013) );
  buffer buf_n4014( .i (n4013), .o (n4014) );
  buffer buf_n4015( .i (n4014), .o (n4015) );
  buffer buf_n4016( .i (n4015), .o (n4016) );
  buffer buf_n4017( .i (n4016), .o (n4017) );
  buffer buf_n4018( .i (n4017), .o (n4018) );
  buffer buf_n4019( .i (n4018), .o (n4019) );
  buffer buf_n4020( .i (n4019), .o (n4020) );
  buffer buf_n4021( .i (n4020), .o (n4021) );
  buffer buf_n4022( .i (n4021), .o (n4022) );
  buffer buf_n4023( .i (n4022), .o (n4023) );
  buffer buf_n4024( .i (n4023), .o (n4024) );
  buffer buf_n4025( .i (n4024), .o (n4025) );
  buffer buf_n4026( .i (n4025), .o (n4026) );
  buffer buf_n4027( .i (n4026), .o (n4027) );
  buffer buf_n4028( .i (n4027), .o (n4028) );
  buffer buf_n4029( .i (n4028), .o (n4029) );
  buffer buf_n4030( .i (n4029), .o (n4030) );
  buffer buf_n4031( .i (n4030), .o (n4031) );
  buffer buf_n4032( .i (n4031), .o (n4032) );
  buffer buf_n4033( .i (n4032), .o (n4033) );
  buffer buf_n4034( .i (n4033), .o (n4034) );
  buffer buf_n4035( .i (n4034), .o (n4035) );
  assign n8382 = n4035 & ~n8120 ;
  buffer buf_n8383( .i (n8382), .o (n8383) );
  assign n8384 = ~n6108 & n8383 ;
  assign n8385 = n6108 & ~n8383 ;
  assign n8386 = n8384 | n8385 ;
  buffer buf_n8387( .i (n8386), .o (n8387) );
  buffer buf_n8388( .i (n8387), .o (n8388) );
  buffer buf_n8389( .i (n8388), .o (n8389) );
  buffer buf_n8390( .i (n8389), .o (n8390) );
  buffer buf_n8391( .i (n8390), .o (n8391) );
  buffer buf_n8392( .i (n8391), .o (n8392) );
  assign n8393 = N150 & N184 ;
  assign n8394 = N228 & N240 ;
  assign n8395 = n8393 & n8394 ;
  buffer buf_n8396( .i (n8395), .o (n8396) );
  assign n8460 = N152 & N210 ;
  assign n8461 = N218 & N230 ;
  assign n8462 = n8460 & n8461 ;
  buffer buf_n8463( .i (n8462), .o (n8463) );
  assign n8527 = n8396 & n8463 ;
  assign n8528 = N182 & N183 ;
  assign n8529 = N185 & N186 ;
  assign n8530 = n8528 & n8529 ;
  buffer buf_n8531( .i (n8530), .o (n8531) );
  assign n8595 = N162 & N172 ;
  assign n8596 = N188 & N199 ;
  assign n8597 = n8595 & n8596 ;
  buffer buf_n8598( .i (n8597), .o (n8598) );
  assign n8662 = n8531 & n8598 ;
  assign n8663 = n8527 & n8662 ;
  buffer buf_n8664( .i (n8663), .o (n8664) );
  buffer buf_n8665( .i (n8664), .o (n8665) );
  buffer buf_n8666( .i (n8665), .o (n8666) );
  buffer buf_n8667( .i (n8666), .o (n8667) );
  buffer buf_n8668( .i (n8667), .o (n8668) );
  buffer buf_n8669( .i (n8668), .o (n8669) );
  buffer buf_n8670( .i (n8669), .o (n8670) );
  buffer buf_n8671( .i (n8670), .o (n8671) );
  buffer buf_n8672( .i (n8671), .o (n8672) );
  buffer buf_n8673( .i (n8672), .o (n8673) );
  buffer buf_n8674( .i (n8673), .o (n8674) );
  buffer buf_n8675( .i (n8674), .o (n8675) );
  buffer buf_n8676( .i (n8675), .o (n8676) );
  buffer buf_n8677( .i (n8676), .o (n8677) );
  buffer buf_n8678( .i (n8677), .o (n8678) );
  buffer buf_n8679( .i (n8678), .o (n8679) );
  buffer buf_n8680( .i (n8679), .o (n8680) );
  assign n8681 = n7599 & n8680 ;
  assign n8682 = n7822 & n8049 ;
  assign n8683 = n8681 & n8682 ;
  buffer buf_n8684( .i (n8683), .o (n8684) );
  buffer buf_n8685( .i (n8684), .o (n8685) );
  buffer buf_n8686( .i (n8685), .o (n8686) );
  buffer buf_n8687( .i (n8686), .o (n8687) );
  buffer buf_n8688( .i (n8687), .o (n8688) );
  buffer buf_n8689( .i (n8688), .o (n8689) );
  buffer buf_n8690( .i (n8689), .o (n8690) );
  buffer buf_n8691( .i (n8690), .o (n8691) );
  buffer buf_n8692( .i (n8691), .o (n8692) );
  buffer buf_n8693( .i (n8692), .o (n8693) );
  buffer buf_n8694( .i (n8693), .o (n8694) );
  buffer buf_n8695( .i (n8694), .o (n8695) );
  buffer buf_n8696( .i (n8695), .o (n8696) );
  buffer buf_n8697( .i (n8696), .o (n8697) );
  buffer buf_n8698( .i (n8697), .o (n8698) );
  buffer buf_n8699( .i (n8698), .o (n8699) );
  buffer buf_n8700( .i (n8699), .o (n8700) );
  buffer buf_n8701( .i (n8700), .o (n8701) );
  buffer buf_n8702( .i (n8701), .o (n8702) );
  buffer buf_n8703( .i (n8702), .o (n8703) );
  buffer buf_n8704( .i (n8703), .o (n8704) );
  buffer buf_n8705( .i (n8704), .o (n8705) );
  buffer buf_n8706( .i (n8705), .o (n8706) );
  buffer buf_n8707( .i (n8706), .o (n8707) );
  buffer buf_n8708( .i (n8707), .o (n8708) );
  buffer buf_n8709( .i (n8708), .o (n8709) );
  buffer buf_n8710( .i (n8709), .o (n8710) );
  buffer buf_n8711( .i (n8710), .o (n8711) );
  buffer buf_n8712( .i (n8711), .o (n8712) );
  buffer buf_n8713( .i (n8712), .o (n8713) );
  buffer buf_n8714( .i (n8713), .o (n8714) );
  buffer buf_n8715( .i (n8714), .o (n8715) );
  buffer buf_n8716( .i (n8715), .o (n8716) );
  buffer buf_n8717( .i (n8716), .o (n8717) );
  buffer buf_n8718( .i (n8717), .o (n8718) );
  buffer buf_n8719( .i (n8718), .o (n8719) );
  buffer buf_n8720( .i (n8719), .o (n8720) );
  buffer buf_n8721( .i (n8720), .o (n8721) );
  buffer buf_n8722( .i (n8721), .o (n8722) );
  buffer buf_n8723( .i (n8722), .o (n8723) );
  buffer buf_n8724( .i (n8723), .o (n8724) );
  buffer buf_n8725( .i (n8724), .o (n8725) );
  assign n8726 = ~n4220 & n4257 ;
  buffer buf_n8727( .i (n8726), .o (n8727) );
  buffer buf_n8728( .i (n8727), .o (n8728) );
  buffer buf_n8729( .i (n8728), .o (n8729) );
  buffer buf_n8730( .i (n8729), .o (n8730) );
  buffer buf_n8731( .i (n8730), .o (n8731) );
  buffer buf_n8732( .i (n8731), .o (n8732) );
  buffer buf_n8733( .i (n8732), .o (n8733) );
  buffer buf_n8734( .i (n8733), .o (n8734) );
  buffer buf_n8735( .i (n8734), .o (n8735) );
  buffer buf_n8736( .i (n8735), .o (n8736) );
  buffer buf_n8737( .i (n8736), .o (n8737) );
  buffer buf_n8738( .i (n8737), .o (n8738) );
  buffer buf_n8739( .i (n8738), .o (n8739) );
  buffer buf_n8740( .i (n8739), .o (n8740) );
  buffer buf_n8741( .i (n8740), .o (n8741) );
  buffer buf_n8742( .i (n8741), .o (n8742) );
  buffer buf_n8743( .i (n8742), .o (n8743) );
  buffer buf_n8744( .i (n8743), .o (n8744) );
  buffer buf_n8745( .i (n8744), .o (n8745) );
  buffer buf_n8746( .i (n8745), .o (n8746) );
  buffer buf_n8747( .i (n8746), .o (n8747) );
  buffer buf_n8748( .i (n8747), .o (n8748) );
  buffer buf_n8749( .i (n8748), .o (n8749) );
  buffer buf_n8750( .i (n8749), .o (n8750) );
  buffer buf_n8751( .i (n8750), .o (n8751) );
  buffer buf_n8752( .i (n8751), .o (n8752) );
  buffer buf_n8753( .i (n8752), .o (n8753) );
  buffer buf_n8754( .i (n8753), .o (n8754) );
  buffer buf_n8755( .i (n8754), .o (n8755) );
  buffer buf_n8756( .i (n8755), .o (n8756) );
  buffer buf_n8757( .i (n8756), .o (n8757) );
  buffer buf_n8758( .i (n8757), .o (n8758) );
  buffer buf_n8759( .i (n8758), .o (n8759) );
  assign n8760 = n5964 | n8759 ;
  assign n8761 = n5964 & n8759 ;
  assign n8762 = n8760 & ~n8761 ;
  buffer buf_n8763( .i (n8762), .o (n8763) );
  buffer buf_n8764( .i (n8763), .o (n8764) );
  buffer buf_n8765( .i (n8764), .o (n8765) );
  buffer buf_n8766( .i (n8765), .o (n8766) );
  buffer buf_n8767( .i (n8766), .o (n8767) );
  buffer buf_n8768( .i (n8767), .o (n8768) );
  buffer buf_n8769( .i (n8768), .o (n8769) );
  buffer buf_n8770( .i (n8769), .o (n8770) );
  buffer buf_n8771( .i (n8770), .o (n8771) );
  buffer buf_n8772( .i (n8771), .o (n8772) );
  buffer buf_n8773( .i (n8772), .o (n8773) );
  buffer buf_n8774( .i (n8773), .o (n8774) );
  buffer buf_n8775( .i (n8774), .o (n8775) );
  buffer buf_n8776( .i (n8775), .o (n8776) );
  buffer buf_n8777( .i (n8776), .o (n8777) );
  buffer buf_n8778( .i (n8777), .o (n8778) );
  buffer buf_n8779( .i (n8778), .o (n8779) );
  buffer buf_n8780( .i (n8779), .o (n8780) );
  buffer buf_n8781( .i (n8780), .o (n8781) );
  buffer buf_n4498( .i (n4497), .o (n4498) );
  buffer buf_n4499( .i (n4498), .o (n4499) );
  buffer buf_n4500( .i (n4499), .o (n4500) );
  buffer buf_n4501( .i (n4500), .o (n4501) );
  buffer buf_n4502( .i (n4501), .o (n4502) );
  buffer buf_n4503( .i (n4502), .o (n4503) );
  buffer buf_n4504( .i (n4503), .o (n4504) );
  buffer buf_n4505( .i (n4504), .o (n4505) );
  buffer buf_n4506( .i (n4505), .o (n4506) );
  buffer buf_n4507( .i (n4506), .o (n4507) );
  buffer buf_n4508( .i (n4507), .o (n4508) );
  buffer buf_n4509( .i (n4508), .o (n4509) );
  buffer buf_n4510( .i (n4509), .o (n4510) );
  buffer buf_n4511( .i (n4510), .o (n4511) );
  buffer buf_n4512( .i (n4511), .o (n4512) );
  buffer buf_n4513( .i (n4512), .o (n4513) );
  buffer buf_n4514( .i (n4513), .o (n4514) );
  buffer buf_n4515( .i (n4514), .o (n4515) );
  buffer buf_n4516( .i (n4515), .o (n4516) );
  buffer buf_n4517( .i (n4516), .o (n4517) );
  buffer buf_n4518( .i (n4517), .o (n4518) );
  buffer buf_n4519( .i (n4518), .o (n4519) );
  buffer buf_n4520( .i (n4519), .o (n4520) );
  buffer buf_n4521( .i (n4520), .o (n4521) );
  buffer buf_n4522( .i (n4521), .o (n4522) );
  buffer buf_n4523( .i (n4522), .o (n4523) );
  buffer buf_n4524( .i (n4523), .o (n4524) );
  buffer buf_n4525( .i (n4524), .o (n4525) );
  buffer buf_n4526( .i (n4525), .o (n4526) );
  buffer buf_n4527( .i (n4526), .o (n4527) );
  buffer buf_n4372( .i (n4371), .o (n4372) );
  buffer buf_n4373( .i (n4372), .o (n4373) );
  buffer buf_n4374( .i (n4373), .o (n4374) );
  buffer buf_n4375( .i (n4374), .o (n4375) );
  buffer buf_n4376( .i (n4375), .o (n4376) );
  buffer buf_n4377( .i (n4376), .o (n4377) );
  buffer buf_n4378( .i (n4377), .o (n4378) );
  buffer buf_n4379( .i (n4378), .o (n4379) );
  buffer buf_n4380( .i (n4379), .o (n4380) );
  buffer buf_n4381( .i (n4380), .o (n4381) );
  buffer buf_n4382( .i (n4381), .o (n4382) );
  buffer buf_n4383( .i (n4382), .o (n4383) );
  buffer buf_n4384( .i (n4383), .o (n4384) );
  buffer buf_n4385( .i (n4384), .o (n4385) );
  buffer buf_n4386( .i (n4385), .o (n4386) );
  buffer buf_n4387( .i (n4386), .o (n4387) );
  buffer buf_n4388( .i (n4387), .o (n4388) );
  buffer buf_n4389( .i (n4388), .o (n4389) );
  buffer buf_n4390( .i (n4389), .o (n4390) );
  buffer buf_n4391( .i (n4390), .o (n4391) );
  buffer buf_n4392( .i (n4391), .o (n4392) );
  buffer buf_n4393( .i (n4392), .o (n4393) );
  buffer buf_n4394( .i (n4393), .o (n4394) );
  buffer buf_n4395( .i (n4394), .o (n4395) );
  buffer buf_n4396( .i (n4395), .o (n4396) );
  buffer buf_n4397( .i (n4396), .o (n4397) );
  buffer buf_n4398( .i (n4397), .o (n4398) );
  buffer buf_n4399( .i (n4398), .o (n4399) );
  buffer buf_n4400( .i (n4399), .o (n4400) );
  buffer buf_n4467( .i (n4466), .o (n4467) );
  buffer buf_n4468( .i (n4467), .o (n4468) );
  buffer buf_n4469( .i (n4468), .o (n4469) );
  buffer buf_n4470( .i (n4469), .o (n4470) );
  buffer buf_n4471( .i (n4470), .o (n4471) );
  buffer buf_n4472( .i (n4471), .o (n4472) );
  buffer buf_n4473( .i (n4472), .o (n4473) );
  buffer buf_n4474( .i (n4473), .o (n4474) );
  buffer buf_n4475( .i (n4474), .o (n4475) );
  buffer buf_n4476( .i (n4475), .o (n4476) );
  buffer buf_n4477( .i (n4476), .o (n4477) );
  buffer buf_n4478( .i (n4477), .o (n4478) );
  buffer buf_n4479( .i (n4478), .o (n4479) );
  buffer buf_n4480( .i (n4479), .o (n4480) );
  buffer buf_n4481( .i (n4480), .o (n4481) );
  buffer buf_n4482( .i (n4481), .o (n4482) );
  buffer buf_n4483( .i (n4482), .o (n4483) );
  buffer buf_n4484( .i (n4483), .o (n4484) );
  buffer buf_n4485( .i (n4484), .o (n4485) );
  buffer buf_n4486( .i (n4485), .o (n4486) );
  buffer buf_n4487( .i (n4486), .o (n4487) );
  buffer buf_n4488( .i (n4487), .o (n4488) );
  buffer buf_n4489( .i (n4488), .o (n4489) );
  buffer buf_n4490( .i (n4489), .o (n4490) );
  buffer buf_n4491( .i (n4490), .o (n4491) );
  buffer buf_n4492( .i (n4491), .o (n4492) );
  buffer buf_n4493( .i (n4492), .o (n4493) );
  assign n8782 = n4493 & ~n5956 ;
  assign n8783 = n4400 & ~n8782 ;
  buffer buf_n8784( .i (n8783), .o (n8784) );
  assign n8785 = n4527 & n8784 ;
  assign n8786 = n4527 | n8784 ;
  assign n8787 = ~n8785 & n8786 ;
  buffer buf_n8788( .i (n8787), .o (n8788) );
  buffer buf_n8789( .i (n8788), .o (n8789) );
  buffer buf_n8790( .i (n8789), .o (n8790) );
  buffer buf_n8791( .i (n8790), .o (n8791) );
  buffer buf_n8792( .i (n8791), .o (n8792) );
  buffer buf_n8793( .i (n8792), .o (n8793) );
  buffer buf_n8794( .i (n8793), .o (n8794) );
  buffer buf_n8795( .i (n8794), .o (n8795) );
  buffer buf_n8796( .i (n8795), .o (n8796) );
  buffer buf_n8797( .i (n8796), .o (n8797) );
  buffer buf_n8798( .i (n8797), .o (n8798) );
  buffer buf_n8799( .i (n8798), .o (n8799) );
  buffer buf_n8800( .i (n8799), .o (n8800) );
  buffer buf_n8801( .i (n8800), .o (n8801) );
  buffer buf_n8802( .i (n8801), .o (n8802) );
  buffer buf_n8803( .i (n8802), .o (n8803) );
  buffer buf_n8804( .i (n8803), .o (n8804) );
  buffer buf_n8805( .i (n8804), .o (n8805) );
  buffer buf_n8806( .i (n8805), .o (n8806) );
  assign n8807 = ~n4318 & n4322 ;
  buffer buf_n8808( .i (n8807), .o (n8808) );
  buffer buf_n8809( .i (n8808), .o (n8809) );
  buffer buf_n8810( .i (n8809), .o (n8810) );
  buffer buf_n8811( .i (n8810), .o (n8811) );
  buffer buf_n8812( .i (n8811), .o (n8812) );
  buffer buf_n8813( .i (n8812), .o (n8813) );
  buffer buf_n8814( .i (n8813), .o (n8814) );
  buffer buf_n8815( .i (n8814), .o (n8815) );
  buffer buf_n8816( .i (n8815), .o (n8816) );
  buffer buf_n8817( .i (n8816), .o (n8817) );
  buffer buf_n8818( .i (n8817), .o (n8818) );
  buffer buf_n8819( .i (n8818), .o (n8819) );
  buffer buf_n8820( .i (n8819), .o (n8820) );
  buffer buf_n8821( .i (n8820), .o (n8821) );
  buffer buf_n8822( .i (n8821), .o (n8822) );
  buffer buf_n8823( .i (n8822), .o (n8823) );
  buffer buf_n8824( .i (n8823), .o (n8824) );
  buffer buf_n8825( .i (n8824), .o (n8825) );
  buffer buf_n8826( .i (n8825), .o (n8826) );
  buffer buf_n8827( .i (n8826), .o (n8827) );
  buffer buf_n8828( .i (n8827), .o (n8828) );
  buffer buf_n8829( .i (n8828), .o (n8829) );
  buffer buf_n8830( .i (n8829), .o (n8830) );
  buffer buf_n8831( .i (n8830), .o (n8831) );
  buffer buf_n8832( .i (n8831), .o (n8832) );
  buffer buf_n8833( .i (n8832), .o (n8833) );
  buffer buf_n8834( .i (n8833), .o (n8834) );
  buffer buf_n8835( .i (n8834), .o (n8835) );
  buffer buf_n8836( .i (n8835), .o (n8836) );
  buffer buf_n8837( .i (n8836), .o (n8837) );
  buffer buf_n8838( .i (n8837), .o (n8838) );
  buffer buf_n8839( .i (n8838), .o (n8839) );
  buffer buf_n8840( .i (n8839), .o (n8840) );
  buffer buf_n8841( .i (n8840), .o (n8841) );
  buffer buf_n4334( .i (n4333), .o (n4334) );
  buffer buf_n4335( .i (n4334), .o (n4335) );
  buffer buf_n4336( .i (n4335), .o (n4336) );
  buffer buf_n4337( .i (n4336), .o (n4337) );
  buffer buf_n4338( .i (n4337), .o (n4338) );
  buffer buf_n4339( .i (n4338), .o (n4339) );
  buffer buf_n4340( .i (n4339), .o (n4340) );
  buffer buf_n4341( .i (n4340), .o (n4341) );
  buffer buf_n4342( .i (n4341), .o (n4342) );
  buffer buf_n4343( .i (n4342), .o (n4343) );
  buffer buf_n4344( .i (n4343), .o (n4344) );
  buffer buf_n4345( .i (n4344), .o (n4345) );
  buffer buf_n4346( .i (n4345), .o (n4346) );
  buffer buf_n4347( .i (n4346), .o (n4347) );
  buffer buf_n4348( .i (n4347), .o (n4348) );
  buffer buf_n4349( .i (n4348), .o (n4349) );
  buffer buf_n4350( .i (n4349), .o (n4350) );
  buffer buf_n4351( .i (n4350), .o (n4351) );
  buffer buf_n4352( .i (n4351), .o (n4352) );
  buffer buf_n4353( .i (n4352), .o (n4353) );
  buffer buf_n4354( .i (n4353), .o (n4354) );
  buffer buf_n4355( .i (n4354), .o (n4355) );
  buffer buf_n4356( .i (n4355), .o (n4356) );
  buffer buf_n4357( .i (n4356), .o (n4357) );
  buffer buf_n4358( .i (n4357), .o (n4358) );
  buffer buf_n4359( .i (n4358), .o (n4359) );
  buffer buf_n4360( .i (n4359), .o (n4360) );
  buffer buf_n4361( .i (n4360), .o (n4361) );
  buffer buf_n4362( .i (n4361), .o (n4362) );
  buffer buf_n4363( .i (n4362), .o (n4363) );
  buffer buf_n4364( .i (n4363), .o (n4364) );
  buffer buf_n4365( .i (n4364), .o (n4365) );
  buffer buf_n4366( .i (n4365), .o (n4366) );
  buffer buf_n4432( .i (n4431), .o (n4432) );
  buffer buf_n4433( .i (n4432), .o (n4433) );
  buffer buf_n4434( .i (n4433), .o (n4434) );
  buffer buf_n4435( .i (n4434), .o (n4435) );
  buffer buf_n4436( .i (n4435), .o (n4436) );
  buffer buf_n4437( .i (n4436), .o (n4437) );
  buffer buf_n4438( .i (n4437), .o (n4438) );
  buffer buf_n4439( .i (n4438), .o (n4439) );
  buffer buf_n4440( .i (n4439), .o (n4440) );
  buffer buf_n4441( .i (n4440), .o (n4441) );
  buffer buf_n4442( .i (n4441), .o (n4442) );
  buffer buf_n4443( .i (n4442), .o (n4443) );
  buffer buf_n4444( .i (n4443), .o (n4444) );
  buffer buf_n4445( .i (n4444), .o (n4445) );
  buffer buf_n4446( .i (n4445), .o (n4446) );
  buffer buf_n4447( .i (n4446), .o (n4447) );
  buffer buf_n4448( .i (n4447), .o (n4448) );
  buffer buf_n4449( .i (n4448), .o (n4449) );
  buffer buf_n4450( .i (n4449), .o (n4450) );
  buffer buf_n4451( .i (n4450), .o (n4451) );
  buffer buf_n4452( .i (n4451), .o (n4452) );
  buffer buf_n4453( .i (n4452), .o (n4453) );
  buffer buf_n4454( .i (n4453), .o (n4454) );
  buffer buf_n4455( .i (n4454), .o (n4455) );
  buffer buf_n4456( .i (n4455), .o (n4456) );
  buffer buf_n4457( .i (n4456), .o (n4457) );
  buffer buf_n4458( .i (n4457), .o (n4458) );
  buffer buf_n4459( .i (n4458), .o (n4459) );
  buffer buf_n4460( .i (n4459), .o (n4460) );
  buffer buf_n4461( .i (n4460), .o (n4461) );
  buffer buf_n4462( .i (n4461), .o (n4462) );
  assign n8842 = n4462 | n5956 ;
  assign n8843 = n4366 & n8842 ;
  buffer buf_n8844( .i (n8843), .o (n8844) );
  assign n8845 = n8841 & ~n8844 ;
  assign n8846 = ~n8841 & n8844 ;
  assign n8847 = n8845 | n8846 ;
  buffer buf_n8848( .i (n8847), .o (n8848) );
  buffer buf_n8849( .i (n8848), .o (n8849) );
  buffer buf_n8850( .i (n8849), .o (n8850) );
  buffer buf_n8851( .i (n8850), .o (n8851) );
  buffer buf_n8852( .i (n8851), .o (n8852) );
  buffer buf_n8853( .i (n8852), .o (n8853) );
  buffer buf_n8854( .i (n8853), .o (n8854) );
  buffer buf_n8855( .i (n8854), .o (n8855) );
  buffer buf_n8856( .i (n8855), .o (n8856) );
  buffer buf_n8857( .i (n8856), .o (n8857) );
  buffer buf_n8858( .i (n8857), .o (n8858) );
  buffer buf_n8859( .i (n8858), .o (n8859) );
  buffer buf_n8860( .i (n8859), .o (n8860) );
  buffer buf_n8861( .i (n8860), .o (n8861) );
  buffer buf_n8862( .i (n8861), .o (n8862) );
  buffer buf_n8863( .i (n8862), .o (n8863) );
  buffer buf_n8864( .i (n8863), .o (n8864) );
  buffer buf_n8865( .i (n8864), .o (n8865) );
  buffer buf_n8866( .i (n8865), .o (n8866) );
  buffer buf_n5957( .i (n5956), .o (n5957) );
  buffer buf_n5958( .i (n5957), .o (n5958) );
  buffer buf_n5959( .i (n5958), .o (n5959) );
  buffer buf_n5960( .i (n5959), .o (n5960) );
  buffer buf_n5961( .i (n5960), .o (n5961) );
  assign n8867 = n4335 & ~n4432 ;
  buffer buf_n8868( .i (n8867), .o (n8868) );
  buffer buf_n8869( .i (n8868), .o (n8869) );
  buffer buf_n8870( .i (n8869), .o (n8870) );
  buffer buf_n8871( .i (n8870), .o (n8871) );
  buffer buf_n8872( .i (n8871), .o (n8872) );
  buffer buf_n8873( .i (n8872), .o (n8873) );
  buffer buf_n8874( .i (n8873), .o (n8874) );
  buffer buf_n8875( .i (n8874), .o (n8875) );
  buffer buf_n8876( .i (n8875), .o (n8876) );
  buffer buf_n8877( .i (n8876), .o (n8877) );
  buffer buf_n8878( .i (n8877), .o (n8878) );
  buffer buf_n8879( .i (n8878), .o (n8879) );
  buffer buf_n8880( .i (n8879), .o (n8880) );
  buffer buf_n8881( .i (n8880), .o (n8881) );
  buffer buf_n8882( .i (n8881), .o (n8882) );
  buffer buf_n8883( .i (n8882), .o (n8883) );
  buffer buf_n8884( .i (n8883), .o (n8884) );
  buffer buf_n8885( .i (n8884), .o (n8885) );
  buffer buf_n8886( .i (n8885), .o (n8886) );
  buffer buf_n8887( .i (n8886), .o (n8887) );
  buffer buf_n8888( .i (n8887), .o (n8888) );
  buffer buf_n8889( .i (n8888), .o (n8889) );
  buffer buf_n8890( .i (n8889), .o (n8890) );
  buffer buf_n8891( .i (n8890), .o (n8891) );
  buffer buf_n8892( .i (n8891), .o (n8892) );
  buffer buf_n8893( .i (n8892), .o (n8893) );
  buffer buf_n8894( .i (n8893), .o (n8894) );
  buffer buf_n8895( .i (n8894), .o (n8895) );
  buffer buf_n8896( .i (n8895), .o (n8896) );
  buffer buf_n8897( .i (n8896), .o (n8897) );
  buffer buf_n8898( .i (n8897), .o (n8898) );
  buffer buf_n8899( .i (n8898), .o (n8899) );
  buffer buf_n8900( .i (n8899), .o (n8900) );
  buffer buf_n8901( .i (n8900), .o (n8901) );
  assign n8902 = ~n5961 & n8901 ;
  assign n8903 = n5961 & ~n8901 ;
  assign n8904 = n8902 | n8903 ;
  buffer buf_n8905( .i (n8904), .o (n8905) );
  buffer buf_n8906( .i (n8905), .o (n8906) );
  buffer buf_n8907( .i (n8906), .o (n8907) );
  buffer buf_n8908( .i (n8907), .o (n8908) );
  buffer buf_n8909( .i (n8908), .o (n8909) );
  buffer buf_n8910( .i (n8909), .o (n8910) );
  buffer buf_n8911( .i (n8910), .o (n8911) );
  buffer buf_n8912( .i (n8911), .o (n8912) );
  buffer buf_n8913( .i (n8912), .o (n8913) );
  buffer buf_n8914( .i (n8913), .o (n8914) );
  buffer buf_n8915( .i (n8914), .o (n8915) );
  buffer buf_n8916( .i (n8915), .o (n8916) );
  buffer buf_n8917( .i (n8916), .o (n8917) );
  buffer buf_n8918( .i (n8917), .o (n8918) );
  buffer buf_n8919( .i (n8918), .o (n8919) );
  buffer buf_n8920( .i (n8919), .o (n8920) );
  buffer buf_n8921( .i (n8920), .o (n8921) );
  buffer buf_n5883( .i (n5882), .o (n5883) );
  buffer buf_n5884( .i (n5883), .o (n5884) );
  buffer buf_n5274( .i (n5273), .o (n5274) );
  buffer buf_n5275( .i (n5274), .o (n5275) );
  buffer buf_n5276( .i (n5275), .o (n5276) );
  buffer buf_n5277( .i (n5276), .o (n5277) );
  buffer buf_n5278( .i (n5277), .o (n5278) );
  buffer buf_n5279( .i (n5278), .o (n5279) );
  buffer buf_n5280( .i (n5279), .o (n5280) );
  buffer buf_n5281( .i (n5280), .o (n5281) );
  buffer buf_n5282( .i (n5281), .o (n5282) );
  buffer buf_n5283( .i (n5282), .o (n5283) );
  buffer buf_n5284( .i (n5283), .o (n5284) );
  buffer buf_n5285( .i (n5284), .o (n5285) );
  buffer buf_n5286( .i (n5285), .o (n5286) );
  buffer buf_n5287( .i (n5286), .o (n5287) );
  buffer buf_n5288( .i (n5287), .o (n5288) );
  buffer buf_n5289( .i (n5288), .o (n5289) );
  buffer buf_n5290( .i (n5289), .o (n5290) );
  buffer buf_n5310( .i (n5309), .o (n5310) );
  buffer buf_n5311( .i (n5310), .o (n5311) );
  buffer buf_n5312( .i (n5311), .o (n5312) );
  buffer buf_n5313( .i (n5312), .o (n5313) );
  buffer buf_n5314( .i (n5313), .o (n5314) );
  buffer buf_n5315( .i (n5314), .o (n5315) );
  buffer buf_n5316( .i (n5315), .o (n5316) );
  buffer buf_n5317( .i (n5316), .o (n5317) );
  buffer buf_n5318( .i (n5317), .o (n5318) );
  buffer buf_n5319( .i (n5318), .o (n5319) );
  buffer buf_n5320( .i (n5319), .o (n5320) );
  buffer buf_n5321( .i (n5320), .o (n5321) );
  buffer buf_n5322( .i (n5321), .o (n5322) );
  buffer buf_n5323( .i (n5322), .o (n5323) );
  buffer buf_n5324( .i (n5323), .o (n5324) );
  buffer buf_n5325( .i (n5324), .o (n5325) );
  buffer buf_n5326( .i (n5325), .o (n5326) );
  buffer buf_n5327( .i (n5326), .o (n5327) );
  buffer buf_n5328( .i (n5327), .o (n5328) );
  assign n8922 = n5290 | n5328 ;
  buffer buf_n8923( .i (n8922), .o (n8923) );
  assign n8924 = n5884 & ~n8923 ;
  buffer buf_n8925( .i (n8924), .o (n8925) );
  assign n8926 = ~n5884 & n8923 ;
  buffer buf_n8927( .i (n8926), .o (n8927) );
  assign n8928 = n8925 | n8927 ;
  buffer buf_n8929( .i (n8928), .o (n8929) );
  buffer buf_n8930( .i (n8929), .o (n8930) );
  buffer buf_n8931( .i (n8930), .o (n8931) );
  buffer buf_n8932( .i (n8931), .o (n8932) );
  buffer buf_n8933( .i (n8932), .o (n8933) );
  buffer buf_n8934( .i (n8933), .o (n8934) );
  buffer buf_n8935( .i (n8934), .o (n8935) );
  buffer buf_n8936( .i (n8935), .o (n8936) );
  buffer buf_n8937( .i (n8936), .o (n8937) );
  buffer buf_n8938( .i (n8937), .o (n8938) );
  buffer buf_n8939( .i (n8938), .o (n8939) );
  buffer buf_n8940( .i (n8939), .o (n8940) );
  buffer buf_n8941( .i (n8940), .o (n8941) );
  buffer buf_n8942( .i (n8941), .o (n8942) );
  buffer buf_n8943( .i (n8942), .o (n8943) );
  buffer buf_n8944( .i (n8943), .o (n8944) );
  buffer buf_n8945( .i (n8944), .o (n8945) );
  buffer buf_n8946( .i (n8945), .o (n8946) );
  buffer buf_n8947( .i (n8946), .o (n8947) );
  buffer buf_n8948( .i (n8947), .o (n8948) );
  buffer buf_n8949( .i (n8948), .o (n8949) );
  buffer buf_n8950( .i (n8949), .o (n8950) );
  buffer buf_n8951( .i (n8950), .o (n8951) );
  buffer buf_n8952( .i (n8951), .o (n8952) );
  buffer buf_n8953( .i (n8952), .o (n8953) );
  buffer buf_n8954( .i (n8953), .o (n8954) );
  buffer buf_n8955( .i (n8954), .o (n8955) );
  buffer buf_n8956( .i (n8955), .o (n8956) );
  buffer buf_n8957( .i (n8956), .o (n8957) );
  buffer buf_n8958( .i (n8957), .o (n8958) );
  buffer buf_n8959( .i (n8958), .o (n8959) );
  buffer buf_n8960( .i (n8959), .o (n8960) );
  buffer buf_n3689( .i (n3688), .o (n3689) );
  buffer buf_n3690( .i (n3689), .o (n3690) );
  buffer buf_n3691( .i (n3690), .o (n3691) );
  buffer buf_n3692( .i (n3691), .o (n3692) );
  buffer buf_n3693( .i (n3692), .o (n3693) );
  buffer buf_n3694( .i (n3693), .o (n3694) );
  buffer buf_n3695( .i (n3694), .o (n3695) );
  buffer buf_n3696( .i (n3695), .o (n3696) );
  buffer buf_n3697( .i (n3696), .o (n3697) );
  buffer buf_n3698( .i (n3697), .o (n3698) );
  buffer buf_n3699( .i (n3698), .o (n3699) );
  buffer buf_n3700( .i (n3699), .o (n3700) );
  buffer buf_n3701( .i (n3700), .o (n3701) );
  buffer buf_n3702( .i (n3701), .o (n3702) );
  buffer buf_n3703( .i (n3702), .o (n3703) );
  buffer buf_n3704( .i (n3703), .o (n3704) );
  buffer buf_n3705( .i (n3704), .o (n3705) );
  buffer buf_n3706( .i (n3705), .o (n3706) );
  buffer buf_n3707( .i (n3706), .o (n3707) );
  buffer buf_n3708( .i (n3707), .o (n3708) );
  buffer buf_n3709( .i (n3708), .o (n3709) );
  buffer buf_n3710( .i (n3709), .o (n3710) );
  buffer buf_n3711( .i (n3710), .o (n3711) );
  buffer buf_n3712( .i (n3711), .o (n3712) );
  buffer buf_n3713( .i (n3712), .o (n3713) );
  buffer buf_n3714( .i (n3713), .o (n3714) );
  buffer buf_n3715( .i (n3714), .o (n3715) );
  buffer buf_n3716( .i (n3715), .o (n3716) );
  buffer buf_n3717( .i (n3716), .o (n3717) );
  buffer buf_n3718( .i (n3717), .o (n3718) );
  buffer buf_n3719( .i (n3718), .o (n3719) );
  buffer buf_n3720( .i (n3719), .o (n3720) );
  buffer buf_n3721( .i (n3720), .o (n3721) );
  buffer buf_n3722( .i (n3721), .o (n3722) );
  buffer buf_n3723( .i (n3722), .o (n3723) );
  buffer buf_n3724( .i (n3723), .o (n3724) );
  buffer buf_n3725( .i (n3724), .o (n3725) );
  buffer buf_n3726( .i (n3725), .o (n3726) );
  buffer buf_n3727( .i (n3726), .o (n3727) );
  buffer buf_n3728( .i (n3727), .o (n3728) );
  buffer buf_n3729( .i (n3728), .o (n3729) );
  buffer buf_n3730( .i (n3729), .o (n3730) );
  buffer buf_n3731( .i (n3730), .o (n3731) );
  buffer buf_n3732( .i (n3731), .o (n3732) );
  buffer buf_n3733( .i (n3732), .o (n3733) );
  buffer buf_n3734( .i (n3733), .o (n3734) );
  buffer buf_n3735( .i (n3734), .o (n3735) );
  buffer buf_n3736( .i (n3735), .o (n3736) );
  buffer buf_n3737( .i (n3736), .o (n3737) );
  buffer buf_n3738( .i (n3737), .o (n3738) );
  buffer buf_n3739( .i (n3738), .o (n3739) );
  buffer buf_n3740( .i (n3739), .o (n3740) );
  buffer buf_n3741( .i (n3740), .o (n3741) );
  buffer buf_n3742( .i (n3741), .o (n3742) );
  buffer buf_n3743( .i (n3742), .o (n3743) );
  buffer buf_n3744( .i (n3743), .o (n3744) );
  buffer buf_n3745( .i (n3744), .o (n3745) );
  buffer buf_n3746( .i (n3745), .o (n3746) );
  buffer buf_n3747( .i (n3746), .o (n3747) );
  buffer buf_n3869( .i (n3868), .o (n3869) );
  buffer buf_n3870( .i (n3869), .o (n3870) );
  assign n8961 = n3870 & n6190 ;
  buffer buf_n3874( .i (n3873), .o (n3874) );
  buffer buf_n3875( .i (n3874), .o (n3875) );
  assign n8962 = n3875 | n6190 ;
  assign n8963 = ~n8961 & n8962 ;
  buffer buf_n8964( .i (n8963), .o (n8964) );
  assign n8965 = n3747 & n8964 ;
  assign n8966 = n3747 | n8964 ;
  assign n8967 = ~n8965 & n8966 ;
  buffer buf_n8968( .i (n8967), .o (n8968) );
  assign n8969 = n3877 & n6190 ;
  buffer buf_n8970( .i (n8969), .o (n8970) );
  assign n8971 = n6192 & ~n8970 ;
  buffer buf_n8972( .i (n8971), .o (n8972) );
  buffer buf_n8973( .i (n8972), .o (n8973) );
  buffer buf_n8974( .i (n8973), .o (n8974) );
  buffer buf_n5439( .i (n5438), .o (n5439) );
  buffer buf_n5440( .i (n5439), .o (n5440) );
  buffer buf_n5441( .i (n5440), .o (n5441) );
  buffer buf_n5442( .i (n5441), .o (n5442) );
  buffer buf_n5443( .i (n5442), .o (n5443) );
  buffer buf_n5444( .i (n5443), .o (n5444) );
  buffer buf_n5445( .i (n5444), .o (n5445) );
  buffer buf_n5446( .i (n5445), .o (n5446) );
  buffer buf_n5447( .i (n5446), .o (n5447) );
  buffer buf_n5448( .i (n5447), .o (n5448) );
  buffer buf_n5449( .i (n5448), .o (n5449) );
  assign n8975 = ~n5449 & n5882 ;
  buffer buf_n5491( .i (n5490), .o (n5491) );
  buffer buf_n5492( .i (n5491), .o (n5492) );
  buffer buf_n5493( .i (n5492), .o (n5493) );
  assign n8976 = ~n5493 & n5928 ;
  assign n8977 = n5493 & ~n5928 ;
  assign n8978 = n8976 | n8977 ;
  buffer buf_n8979( .i (n8978), .o (n8979) );
  buffer buf_n8980( .i (n8979), .o (n8980) );
  buffer buf_n8981( .i (n8980), .o (n8981) );
  buffer buf_n8982( .i (n8981), .o (n8982) );
  buffer buf_n8983( .i (n8982), .o (n8983) );
  buffer buf_n8984( .i (n8983), .o (n8984) );
  buffer buf_n8985( .i (n8984), .o (n8985) );
  assign n8986 = ~n8975 & n8985 ;
  assign n8987 = n5886 | n8986 ;
  buffer buf_n8988( .i (n8987), .o (n8988) );
  buffer buf_n8989( .i (n8988), .o (n8989) );
  buffer buf_n8990( .i (n8989), .o (n8990) );
  buffer buf_n8991( .i (n8990), .o (n8991) );
  buffer buf_n8992( .i (n8991), .o (n8992) );
  buffer buf_n8993( .i (n8992), .o (n8993) );
  buffer buf_n8994( .i (n8993), .o (n8994) );
  buffer buf_n8995( .i (n8994), .o (n8995) );
  buffer buf_n8996( .i (n8995), .o (n8996) );
  buffer buf_n8997( .i (n8996), .o (n8997) );
  buffer buf_n8998( .i (n8997), .o (n8998) );
  buffer buf_n8999( .i (n8998), .o (n8999) );
  buffer buf_n9000( .i (n8999), .o (n9000) );
  buffer buf_n9001( .i (n9000), .o (n9001) );
  buffer buf_n9002( .i (n9001), .o (n9002) );
  buffer buf_n9003( .i (n9002), .o (n9003) );
  buffer buf_n9004( .i (n9003), .o (n9004) );
  buffer buf_n9005( .i (n9004), .o (n9005) );
  buffer buf_n9006( .i (n9005), .o (n9006) );
  buffer buf_n9007( .i (n9006), .o (n9007) );
  buffer buf_n9008( .i (n9007), .o (n9008) );
  buffer buf_n9009( .i (n9008), .o (n9009) );
  buffer buf_n9010( .i (n9009), .o (n9010) );
  buffer buf_n9011( .i (n9010), .o (n9011) );
  buffer buf_n9012( .i (n9011), .o (n9012) );
  buffer buf_n9013( .i (n9012), .o (n9013) );
  buffer buf_n9014( .i (n9013), .o (n9014) );
  buffer buf_n9015( .i (n9014), .o (n9015) );
  buffer buf_n9016( .i (n9015), .o (n9016) );
  buffer buf_n9017( .i (n9016), .o (n9017) );
  buffer buf_n9018( .i (n9017), .o (n9018) );
  buffer buf_n9019( .i (n9018), .o (n9019) );
  buffer buf_n9020( .i (n9019), .o (n9020) );
  buffer buf_n9021( .i (n9020), .o (n9021) );
  buffer buf_n5369( .i (n5368), .o (n5369) );
  buffer buf_n5370( .i (n5369), .o (n5370) );
  buffer buf_n5371( .i (n5370), .o (n5371) );
  buffer buf_n5372( .i (n5371), .o (n5372) );
  buffer buf_n5373( .i (n5372), .o (n5373) );
  buffer buf_n5374( .i (n5373), .o (n5374) );
  buffer buf_n5375( .i (n5374), .o (n5375) );
  buffer buf_n5376( .i (n5375), .o (n5376) );
  buffer buf_n5377( .i (n5376), .o (n5377) );
  buffer buf_n5378( .i (n5377), .o (n5378) );
  buffer buf_n5379( .i (n5378), .o (n5379) );
  buffer buf_n5380( .i (n5379), .o (n5380) );
  buffer buf_n5381( .i (n5380), .o (n5381) );
  buffer buf_n5382( .i (n5381), .o (n5382) );
  buffer buf_n5383( .i (n5382), .o (n5383) );
  buffer buf_n5384( .i (n5383), .o (n5384) );
  buffer buf_n5385( .i (n5384), .o (n5385) );
  buffer buf_n5386( .i (n5385), .o (n5386) );
  buffer buf_n5914( .i (n5913), .o (n5914) );
  buffer buf_n5915( .i (n5914), .o (n5915) );
  buffer buf_n5916( .i (n5915), .o (n5916) );
  buffer buf_n5917( .i (n5916), .o (n5917) );
  buffer buf_n5918( .i (n5917), .o (n5918) );
  buffer buf_n5919( .i (n5918), .o (n5919) );
  buffer buf_n5920( .i (n5919), .o (n5920) );
  buffer buf_n5921( .i (n5920), .o (n5921) );
  buffer buf_n5922( .i (n5921), .o (n5922) );
  buffer buf_n5923( .i (n5922), .o (n5923) );
  buffer buf_n5924( .i (n5923), .o (n5924) );
  buffer buf_n5925( .i (n5924), .o (n5925) );
  buffer buf_n5413( .i (n5412), .o (n5413) );
  buffer buf_n5414( .i (n5413), .o (n5414) );
  assign n9022 = n5337 | n5414 ;
  buffer buf_n9023( .i (n9022), .o (n9023) );
  buffer buf_n9024( .i (n9023), .o (n9024) );
  buffer buf_n9025( .i (n9024), .o (n9025) );
  buffer buf_n9026( .i (n9025), .o (n9026) );
  buffer buf_n9027( .i (n9026), .o (n9027) );
  buffer buf_n9028( .i (n9027), .o (n9028) );
  buffer buf_n9029( .i (n9028), .o (n9029) );
  buffer buf_n9030( .i (n9029), .o (n9030) );
  buffer buf_n9031( .i (n9030), .o (n9031) );
  buffer buf_n9032( .i (n9031), .o (n9032) );
  buffer buf_n9033( .i (n9032), .o (n9033) );
  buffer buf_n9034( .i (n9033), .o (n9034) );
  assign n9035 = n5882 & ~n9034 ;
  assign n9036 = n5925 | n9035 ;
  buffer buf_n9037( .i (n9036), .o (n9037) );
  assign n9038 = n5386 | n9037 ;
  assign n9039 = n5386 & n9037 ;
  assign n9040 = n9038 & ~n9039 ;
  buffer buf_n9041( .i (n9040), .o (n9041) );
  buffer buf_n9042( .i (n9041), .o (n9042) );
  buffer buf_n9043( .i (n9042), .o (n9043) );
  buffer buf_n9044( .i (n9043), .o (n9044) );
  buffer buf_n9045( .i (n9044), .o (n9045) );
  buffer buf_n9046( .i (n9045), .o (n9046) );
  buffer buf_n9047( .i (n9046), .o (n9047) );
  buffer buf_n9048( .i (n9047), .o (n9048) );
  buffer buf_n9049( .i (n9048), .o (n9049) );
  buffer buf_n9050( .i (n9049), .o (n9050) );
  buffer buf_n9051( .i (n9050), .o (n9051) );
  buffer buf_n9052( .i (n9051), .o (n9052) );
  buffer buf_n9053( .i (n9052), .o (n9053) );
  buffer buf_n9054( .i (n9053), .o (n9054) );
  buffer buf_n9055( .i (n9054), .o (n9055) );
  buffer buf_n9056( .i (n9055), .o (n9056) );
  buffer buf_n9057( .i (n9056), .o (n9057) );
  buffer buf_n9058( .i (n9057), .o (n9058) );
  buffer buf_n9059( .i (n9058), .o (n9059) );
  buffer buf_n9060( .i (n9059), .o (n9060) );
  buffer buf_n9061( .i (n9060), .o (n9061) );
  buffer buf_n9062( .i (n9061), .o (n9062) );
  buffer buf_n9063( .i (n9062), .o (n9063) );
  buffer buf_n9064( .i (n9063), .o (n9064) );
  buffer buf_n9065( .i (n9064), .o (n9065) );
  buffer buf_n9066( .i (n9065), .o (n9066) );
  buffer buf_n9067( .i (n9066), .o (n9067) );
  buffer buf_n9068( .i (n9067), .o (n9068) );
  buffer buf_n9069( .i (n9068), .o (n9069) );
  buffer buf_n9070( .i (n9069), .o (n9070) );
  buffer buf_n9071( .i (n9070), .o (n9071) );
  buffer buf_n9072( .i (n9071), .o (n9072) );
  buffer buf_n5415( .i (n5414), .o (n5415) );
  buffer buf_n5416( .i (n5415), .o (n5416) );
  buffer buf_n5417( .i (n5416), .o (n5417) );
  buffer buf_n5418( .i (n5417), .o (n5418) );
  buffer buf_n5419( .i (n5418), .o (n5419) );
  buffer buf_n5420( .i (n5419), .o (n5420) );
  buffer buf_n5421( .i (n5420), .o (n5421) );
  buffer buf_n5422( .i (n5421), .o (n5422) );
  buffer buf_n5423( .i (n5422), .o (n5423) );
  buffer buf_n5424( .i (n5423), .o (n5424) );
  buffer buf_n5425( .i (n5424), .o (n5425) );
  buffer buf_n5426( .i (n5425), .o (n5426) );
  buffer buf_n5427( .i (n5426), .o (n5427) );
  buffer buf_n5428( .i (n5427), .o (n5428) );
  buffer buf_n5429( .i (n5428), .o (n5429) );
  buffer buf_n5430( .i (n5429), .o (n5430) );
  buffer buf_n5431( .i (n5430), .o (n5431) );
  buffer buf_n5432( .i (n5431), .o (n5432) );
  buffer buf_n5433( .i (n5432), .o (n5433) );
  buffer buf_n5434( .i (n5433), .o (n5434) );
  buffer buf_n5890( .i (n5889), .o (n5890) );
  buffer buf_n5891( .i (n5890), .o (n5891) );
  buffer buf_n5892( .i (n5891), .o (n5892) );
  buffer buf_n5893( .i (n5892), .o (n5893) );
  buffer buf_n5894( .i (n5893), .o (n5894) );
  buffer buf_n5895( .i (n5894), .o (n5895) );
  buffer buf_n5896( .i (n5895), .o (n5896) );
  buffer buf_n5897( .i (n5896), .o (n5897) );
  buffer buf_n5898( .i (n5897), .o (n5898) );
  buffer buf_n5899( .i (n5898), .o (n5899) );
  buffer buf_n5900( .i (n5899), .o (n5900) );
  buffer buf_n5901( .i (n5900), .o (n5901) );
  buffer buf_n5902( .i (n5901), .o (n5902) );
  buffer buf_n5903( .i (n5902), .o (n5903) );
  buffer buf_n5904( .i (n5903), .o (n5904) );
  buffer buf_n5905( .i (n5904), .o (n5905) );
  buffer buf_n5906( .i (n5905), .o (n5906) );
  buffer buf_n5907( .i (n5906), .o (n5907) );
  buffer buf_n5908( .i (n5907), .o (n5908) );
  buffer buf_n5909( .i (n5908), .o (n5909) );
  assign n9073 = n5303 | n5330 ;
  buffer buf_n9074( .i (n9073), .o (n9074) );
  buffer buf_n9075( .i (n9074), .o (n9075) );
  buffer buf_n9076( .i (n9075), .o (n9076) );
  buffer buf_n9077( .i (n9076), .o (n9077) );
  buffer buf_n9078( .i (n9077), .o (n9078) );
  buffer buf_n9079( .i (n9078), .o (n9079) );
  buffer buf_n9080( .i (n9079), .o (n9080) );
  buffer buf_n9081( .i (n9080), .o (n9081) );
  buffer buf_n9082( .i (n9081), .o (n9082) );
  buffer buf_n9083( .i (n9082), .o (n9083) );
  buffer buf_n9084( .i (n9083), .o (n9084) );
  buffer buf_n9085( .i (n9084), .o (n9085) );
  buffer buf_n9086( .i (n9085), .o (n9086) );
  buffer buf_n9087( .i (n9086), .o (n9087) );
  buffer buf_n9088( .i (n9087), .o (n9088) );
  buffer buf_n9089( .i (n9088), .o (n9089) );
  buffer buf_n9090( .i (n9089), .o (n9090) );
  buffer buf_n9091( .i (n9090), .o (n9091) );
  buffer buf_n9092( .i (n9091), .o (n9092) );
  buffer buf_n9093( .i (n9092), .o (n9093) );
  buffer buf_n9094( .i (n9093), .o (n9094) );
  buffer buf_n9095( .i (n9094), .o (n9095) );
  assign n9098 = n8925 & ~n9095 ;
  assign n9099 = n5909 | n9098 ;
  buffer buf_n9100( .i (n9099), .o (n9100) );
  assign n9101 = n5434 & n9100 ;
  assign n9102 = n5434 | n9100 ;
  assign n9103 = ~n9101 & n9102 ;
  buffer buf_n9104( .i (n9103), .o (n9104) );
  buffer buf_n9105( .i (n9104), .o (n9105) );
  buffer buf_n9106( .i (n9105), .o (n9106) );
  buffer buf_n9107( .i (n9106), .o (n9107) );
  buffer buf_n9108( .i (n9107), .o (n9108) );
  buffer buf_n9109( .i (n9108), .o (n9109) );
  buffer buf_n9110( .i (n9109), .o (n9110) );
  buffer buf_n9111( .i (n9110), .o (n9111) );
  buffer buf_n9112( .i (n9111), .o (n9112) );
  buffer buf_n9113( .i (n9112), .o (n9113) );
  buffer buf_n9114( .i (n9113), .o (n9114) );
  buffer buf_n9115( .i (n9114), .o (n9115) );
  buffer buf_n9116( .i (n9115), .o (n9116) );
  buffer buf_n9117( .i (n9116), .o (n9117) );
  buffer buf_n9118( .i (n9117), .o (n9118) );
  buffer buf_n9119( .i (n9118), .o (n9119) );
  buffer buf_n9120( .i (n9119), .o (n9120) );
  buffer buf_n9121( .i (n9120), .o (n9121) );
  buffer buf_n9122( .i (n9121), .o (n9122) );
  buffer buf_n9123( .i (n9122), .o (n9123) );
  buffer buf_n9124( .i (n9123), .o (n9124) );
  buffer buf_n9125( .i (n9124), .o (n9125) );
  buffer buf_n9126( .i (n9125), .o (n9126) );
  buffer buf_n9127( .i (n9126), .o (n9127) );
  buffer buf_n9128( .i (n9127), .o (n9128) );
  buffer buf_n9129( .i (n9128), .o (n9129) );
  buffer buf_n9130( .i (n9129), .o (n9130) );
  buffer buf_n9131( .i (n9130), .o (n9131) );
  buffer buf_n9096( .i (n9095), .o (n9096) );
  buffer buf_n9097( .i (n9096), .o (n9097) );
  buffer buf_n5291( .i (n5290), .o (n5291) );
  buffer buf_n5292( .i (n5291), .o (n5292) );
  buffer buf_n5293( .i (n5292), .o (n5293) );
  buffer buf_n5294( .i (n5293), .o (n5294) );
  assign n9132 = n5294 | n8925 ;
  buffer buf_n9133( .i (n9132), .o (n9133) );
  assign n9134 = n9097 | n9133 ;
  assign n9135 = n9097 & n9133 ;
  assign n9136 = n9134 & ~n9135 ;
  buffer buf_n9137( .i (n9136), .o (n9137) );
  buffer buf_n9138( .i (n9137), .o (n9138) );
  buffer buf_n9139( .i (n9138), .o (n9139) );
  buffer buf_n9140( .i (n9139), .o (n9140) );
  buffer buf_n9141( .i (n9140), .o (n9141) );
  buffer buf_n9142( .i (n9141), .o (n9142) );
  buffer buf_n9143( .i (n9142), .o (n9143) );
  buffer buf_n9144( .i (n9143), .o (n9144) );
  buffer buf_n9145( .i (n9144), .o (n9145) );
  buffer buf_n9146( .i (n9145), .o (n9146) );
  buffer buf_n9147( .i (n9146), .o (n9147) );
  buffer buf_n9148( .i (n9147), .o (n9148) );
  buffer buf_n9149( .i (n9148), .o (n9149) );
  buffer buf_n9150( .i (n9149), .o (n9150) );
  buffer buf_n9151( .i (n9150), .o (n9151) );
  buffer buf_n9152( .i (n9151), .o (n9152) );
  buffer buf_n9153( .i (n9152), .o (n9153) );
  buffer buf_n9154( .i (n9153), .o (n9154) );
  buffer buf_n9155( .i (n9154), .o (n9155) );
  buffer buf_n9156( .i (n9155), .o (n9156) );
  buffer buf_n9157( .i (n9156), .o (n9157) );
  buffer buf_n9158( .i (n9157), .o (n9158) );
  buffer buf_n9159( .i (n9158), .o (n9159) );
  buffer buf_n9160( .i (n9159), .o (n9160) );
  buffer buf_n9161( .i (n9160), .o (n9161) );
  buffer buf_n9162( .i (n9161), .o (n9162) );
  buffer buf_n9163( .i (n9162), .o (n9163) );
  buffer buf_n9164( .i (n9163), .o (n9164) );
  buffer buf_n9165( .i (n9164), .o (n9165) );
  assign n9166 = n4985 | n5014 ;
  buffer buf_n9167( .i (n9166), .o (n9167) );
  buffer buf_n9168( .i (n9167), .o (n9168) );
  buffer buf_n9169( .i (n9168), .o (n9169) );
  buffer buf_n9170( .i (n9169), .o (n9170) );
  buffer buf_n9171( .i (n9170), .o (n9171) );
  buffer buf_n9172( .i (n9171), .o (n9172) );
  buffer buf_n9173( .i (n9172), .o (n9173) );
  buffer buf_n9174( .i (n9173), .o (n9174) );
  buffer buf_n9175( .i (n9174), .o (n9175) );
  buffer buf_n9176( .i (n9175), .o (n9176) );
  buffer buf_n9177( .i (n9176), .o (n9177) );
  buffer buf_n9178( .i (n9177), .o (n9178) );
  buffer buf_n9179( .i (n9178), .o (n9179) );
  buffer buf_n9180( .i (n9179), .o (n9180) );
  buffer buf_n9181( .i (n9180), .o (n9181) );
  buffer buf_n9182( .i (n9181), .o (n9182) );
  buffer buf_n9183( .i (n9182), .o (n9183) );
  buffer buf_n9184( .i (n9183), .o (n9184) );
  buffer buf_n9185( .i (n9184), .o (n9185) );
  buffer buf_n9186( .i (n9185), .o (n9186) );
  buffer buf_n9187( .i (n9186), .o (n9187) );
  buffer buf_n9188( .i (n9187), .o (n9188) );
  buffer buf_n9189( .i (n9188), .o (n9189) );
  buffer buf_n9190( .i (n9189), .o (n9190) );
  buffer buf_n9191( .i (n9190), .o (n9191) );
  assign n9192 = ~n5946 & n9191 ;
  assign n9193 = n5946 & ~n9191 ;
  assign n9194 = n9192 | n9193 ;
  buffer buf_n9195( .i (n9194), .o (n9195) );
  buffer buf_n9196( .i (n9195), .o (n9196) );
  buffer buf_n9197( .i (n9196), .o (n9197) );
  buffer buf_n9198( .i (n9197), .o (n9198) );
  buffer buf_n9199( .i (n9198), .o (n9199) );
  buffer buf_n9200( .i (n9199), .o (n9200) );
  buffer buf_n9201( .i (n9200), .o (n9201) );
  buffer buf_n9202( .i (n9201), .o (n9202) );
  buffer buf_n9203( .i (n9202), .o (n9203) );
  buffer buf_n9204( .i (n9203), .o (n9204) );
  buffer buf_n9205( .i (n9204), .o (n9205) );
  buffer buf_n9206( .i (n9205), .o (n9206) );
  buffer buf_n9207( .i (n9206), .o (n9207) );
  buffer buf_n9208( .i (n9207), .o (n9208) );
  buffer buf_n9209( .i (n9208), .o (n9209) );
  buffer buf_n9210( .i (n9209), .o (n9210) );
  buffer buf_n9211( .i (n9210), .o (n9211) );
  buffer buf_n9212( .i (n9211), .o (n9212) );
  buffer buf_n9213( .i (n9212), .o (n9213) );
  buffer buf_n9214( .i (n9213), .o (n9214) );
  buffer buf_n9215( .i (n9214), .o (n9215) );
  buffer buf_n9216( .i (n9215), .o (n9216) );
  buffer buf_n9217( .i (n9216), .o (n9217) );
  buffer buf_n9218( .i (n9217), .o (n9218) );
  buffer buf_n9219( .i (n9218), .o (n9219) );
  buffer buf_n9220( .i (n9219), .o (n9220) );
  buffer buf_n9221( .i (n9220), .o (n9221) );
  buffer buf_n9222( .i (n9221), .o (n9222) );
  assign n9223 = n5049 | n5057 ;
  buffer buf_n9224( .i (n9223), .o (n9224) );
  buffer buf_n9225( .i (n9224), .o (n9225) );
  buffer buf_n9226( .i (n9225), .o (n9226) );
  buffer buf_n9227( .i (n9226), .o (n9227) );
  buffer buf_n9228( .i (n9227), .o (n9228) );
  buffer buf_n9229( .i (n9228), .o (n9229) );
  buffer buf_n9230( .i (n9229), .o (n9230) );
  buffer buf_n9231( .i (n9230), .o (n9231) );
  buffer buf_n9232( .i (n9231), .o (n9232) );
  buffer buf_n9233( .i (n9232), .o (n9233) );
  buffer buf_n9234( .i (n9233), .o (n9234) );
  buffer buf_n9235( .i (n9234), .o (n9235) );
  buffer buf_n9236( .i (n9235), .o (n9236) );
  buffer buf_n9237( .i (n9236), .o (n9237) );
  buffer buf_n9238( .i (n9237), .o (n9238) );
  buffer buf_n9239( .i (n9238), .o (n9239) );
  buffer buf_n9240( .i (n9239), .o (n9240) );
  buffer buf_n9241( .i (n9240), .o (n9241) );
  buffer buf_n9242( .i (n9241), .o (n9242) );
  buffer buf_n9243( .i (n9242), .o (n9243) );
  buffer buf_n9244( .i (n9243), .o (n9244) );
  buffer buf_n9245( .i (n9244), .o (n9245) );
  buffer buf_n9246( .i (n9245), .o (n9246) );
  buffer buf_n9247( .i (n9246), .o (n9247) );
  buffer buf_n9248( .i (n9247), .o (n9248) );
  buffer buf_n5112( .i (n5111), .o (n5112) );
  buffer buf_n5113( .i (n5112), .o (n5113) );
  buffer buf_n5114( .i (n5113), .o (n5114) );
  buffer buf_n5115( .i (n5114), .o (n5115) );
  buffer buf_n5116( .i (n5115), .o (n5116) );
  buffer buf_n5117( .i (n5116), .o (n5117) );
  buffer buf_n5118( .i (n5117), .o (n5118) );
  buffer buf_n5119( .i (n5118), .o (n5119) );
  buffer buf_n5120( .i (n5119), .o (n5120) );
  buffer buf_n5121( .i (n5120), .o (n5121) );
  buffer buf_n5122( .i (n5121), .o (n5122) );
  buffer buf_n5123( .i (n5122), .o (n5123) );
  buffer buf_n5124( .i (n5123), .o (n5124) );
  buffer buf_n5125( .i (n5124), .o (n5125) );
  buffer buf_n5126( .i (n5125), .o (n5126) );
  buffer buf_n5127( .i (n5126), .o (n5127) );
  buffer buf_n5128( .i (n5127), .o (n5128) );
  buffer buf_n5129( .i (n5128), .o (n5129) );
  buffer buf_n5130( .i (n5129), .o (n5130) );
  buffer buf_n5131( .i (n5130), .o (n5131) );
  buffer buf_n5229( .i (n5228), .o (n5229) );
  buffer buf_n5230( .i (n5229), .o (n5230) );
  buffer buf_n5231( .i (n5230), .o (n5231) );
  buffer buf_n5232( .i (n5231), .o (n5232) );
  buffer buf_n5233( .i (n5232), .o (n5233) );
  buffer buf_n5234( .i (n5233), .o (n5234) );
  buffer buf_n5235( .i (n5234), .o (n5235) );
  buffer buf_n5236( .i (n5235), .o (n5236) );
  buffer buf_n5237( .i (n5236), .o (n5237) );
  buffer buf_n5238( .i (n5237), .o (n5238) );
  buffer buf_n5239( .i (n5238), .o (n5239) );
  buffer buf_n5240( .i (n5239), .o (n5240) );
  buffer buf_n5241( .i (n5240), .o (n5241) );
  buffer buf_n5242( .i (n5241), .o (n5242) );
  buffer buf_n5243( .i (n5242), .o (n5243) );
  buffer buf_n5244( .i (n5243), .o (n5244) );
  buffer buf_n5245( .i (n5244), .o (n5245) );
  assign n9249 = ~n5245 & n5940 ;
  assign n9250 = n5131 | n9249 ;
  buffer buf_n9251( .i (n9250), .o (n9251) );
  assign n9252 = n9248 | n9251 ;
  assign n9253 = n9248 & n9251 ;
  assign n9254 = n9252 & ~n9253 ;
  buffer buf_n9255( .i (n9254), .o (n9255) );
  buffer buf_n9256( .i (n9255), .o (n9256) );
  buffer buf_n9257( .i (n9256), .o (n9257) );
  buffer buf_n9258( .i (n9257), .o (n9258) );
  buffer buf_n9259( .i (n9258), .o (n9259) );
  buffer buf_n9260( .i (n9259), .o (n9260) );
  buffer buf_n9261( .i (n9260), .o (n9261) );
  buffer buf_n9262( .i (n9261), .o (n9262) );
  buffer buf_n9263( .i (n9262), .o (n9263) );
  buffer buf_n9264( .i (n9263), .o (n9264) );
  buffer buf_n9265( .i (n9264), .o (n9265) );
  buffer buf_n9266( .i (n9265), .o (n9266) );
  buffer buf_n9267( .i (n9266), .o (n9267) );
  buffer buf_n9268( .i (n9267), .o (n9268) );
  buffer buf_n9269( .i (n9268), .o (n9269) );
  buffer buf_n9270( .i (n9269), .o (n9270) );
  buffer buf_n9271( .i (n9270), .o (n9271) );
  buffer buf_n9272( .i (n9271), .o (n9272) );
  buffer buf_n9273( .i (n9272), .o (n9273) );
  buffer buf_n9274( .i (n9273), .o (n9274) );
  buffer buf_n9275( .i (n9274), .o (n9275) );
  buffer buf_n9276( .i (n9275), .o (n9276) );
  buffer buf_n9277( .i (n9276), .o (n9277) );
  buffer buf_n9278( .i (n9277), .o (n9278) );
  buffer buf_n9279( .i (n9278), .o (n9279) );
  buffer buf_n9280( .i (n9279), .o (n9280) );
  buffer buf_n9281( .i (n9280), .o (n9281) );
  buffer buf_n9282( .i (n9281), .o (n9282) );
  buffer buf_n5155( .i (n5154), .o (n5155) );
  buffer buf_n5156( .i (n5155), .o (n5156) );
  buffer buf_n5157( .i (n5156), .o (n5157) );
  buffer buf_n5158( .i (n5157), .o (n5158) );
  buffer buf_n5159( .i (n5158), .o (n5159) );
  buffer buf_n5160( .i (n5159), .o (n5160) );
  buffer buf_n5161( .i (n5160), .o (n5161) );
  buffer buf_n5162( .i (n5161), .o (n5162) );
  buffer buf_n5163( .i (n5162), .o (n5163) );
  buffer buf_n5164( .i (n5163), .o (n5164) );
  buffer buf_n5165( .i (n5164), .o (n5165) );
  buffer buf_n5166( .i (n5165), .o (n5166) );
  buffer buf_n5167( .i (n5166), .o (n5167) );
  buffer buf_n5168( .i (n5167), .o (n5168) );
  buffer buf_n5169( .i (n5168), .o (n5169) );
  buffer buf_n5170( .i (n5169), .o (n5170) );
  buffer buf_n5171( .i (n5170), .o (n5171) );
  buffer buf_n5172( .i (n5171), .o (n5172) );
  buffer buf_n5173( .i (n5172), .o (n5173) );
  buffer buf_n5174( .i (n5173), .o (n5174) );
  buffer buf_n5175( .i (n5174), .o (n5175) );
  buffer buf_n5176( .i (n5175), .o (n5176) );
  buffer buf_n5181( .i (n5180), .o (n5181) );
  buffer buf_n5182( .i (n5181), .o (n5182) );
  buffer buf_n5183( .i (n5182), .o (n5183) );
  buffer buf_n5184( .i (n5183), .o (n5184) );
  buffer buf_n5185( .i (n5184), .o (n5185) );
  buffer buf_n5186( .i (n5185), .o (n5186) );
  buffer buf_n5187( .i (n5186), .o (n5187) );
  buffer buf_n5188( .i (n5187), .o (n5188) );
  buffer buf_n5189( .i (n5188), .o (n5189) );
  buffer buf_n5190( .i (n5189), .o (n5190) );
  buffer buf_n5191( .i (n5190), .o (n5191) );
  buffer buf_n5192( .i (n5191), .o (n5192) );
  buffer buf_n5193( .i (n5192), .o (n5193) );
  buffer buf_n5194( .i (n5193), .o (n5194) );
  buffer buf_n5195( .i (n5194), .o (n5195) );
  buffer buf_n5196( .i (n5195), .o (n5196) );
  buffer buf_n5197( .i (n5196), .o (n5197) );
  buffer buf_n5198( .i (n5197), .o (n5198) );
  buffer buf_n5199( .i (n5198), .o (n5199) );
  buffer buf_n5200( .i (n5199), .o (n5200) );
  buffer buf_n5201( .i (n5200), .o (n5201) );
  buffer buf_n5202( .i (n5201), .o (n5202) );
  buffer buf_n5087( .i (n5086), .o (n5087) );
  buffer buf_n5088( .i (n5087), .o (n5088) );
  buffer buf_n5089( .i (n5088), .o (n5089) );
  buffer buf_n5090( .i (n5089), .o (n5090) );
  buffer buf_n5091( .i (n5090), .o (n5091) );
  buffer buf_n5092( .i (n5091), .o (n5092) );
  buffer buf_n5093( .i (n5092), .o (n5093) );
  buffer buf_n5094( .i (n5093), .o (n5094) );
  buffer buf_n5095( .i (n5094), .o (n5095) );
  buffer buf_n5096( .i (n5095), .o (n5096) );
  buffer buf_n5097( .i (n5096), .o (n5097) );
  buffer buf_n5098( .i (n5097), .o (n5098) );
  buffer buf_n5099( .i (n5098), .o (n5099) );
  buffer buf_n5100( .i (n5099), .o (n5100) );
  buffer buf_n5101( .i (n5100), .o (n5101) );
  buffer buf_n5102( .i (n5101), .o (n5102) );
  buffer buf_n5103( .i (n5102), .o (n5103) );
  buffer buf_n5104( .i (n5103), .o (n5104) );
  buffer buf_n5105( .i (n5104), .o (n5105) );
  buffer buf_n5106( .i (n5105), .o (n5106) );
  buffer buf_n5107( .i (n5106), .o (n5107) );
  assign n9283 = n5107 | n5940 ;
  assign n9284 = ~n5202 & n9283 ;
  buffer buf_n9285( .i (n9284), .o (n9285) );
  assign n9286 = n5176 & ~n9285 ;
  assign n9287 = ~n5176 & n9285 ;
  assign n9288 = n9286 | n9287 ;
  buffer buf_n9289( .i (n9288), .o (n9289) );
  buffer buf_n9290( .i (n9289), .o (n9290) );
  buffer buf_n9291( .i (n9290), .o (n9291) );
  buffer buf_n9292( .i (n9291), .o (n9292) );
  buffer buf_n9293( .i (n9292), .o (n9293) );
  buffer buf_n9294( .i (n9293), .o (n9294) );
  buffer buf_n9295( .i (n9294), .o (n9295) );
  buffer buf_n9296( .i (n9295), .o (n9296) );
  buffer buf_n9297( .i (n9296), .o (n9297) );
  buffer buf_n9298( .i (n9297), .o (n9298) );
  buffer buf_n9299( .i (n9298), .o (n9299) );
  buffer buf_n9300( .i (n9299), .o (n9300) );
  buffer buf_n9301( .i (n9300), .o (n9301) );
  buffer buf_n9302( .i (n9301), .o (n9302) );
  buffer buf_n9303( .i (n9302), .o (n9303) );
  buffer buf_n9304( .i (n9303), .o (n9304) );
  buffer buf_n9305( .i (n9304), .o (n9305) );
  buffer buf_n9306( .i (n9305), .o (n9306) );
  buffer buf_n9307( .i (n9306), .o (n9307) );
  buffer buf_n9308( .i (n9307), .o (n9308) );
  buffer buf_n9309( .i (n9308), .o (n9309) );
  buffer buf_n9310( .i (n9309), .o (n9310) );
  buffer buf_n9311( .i (n9310), .o (n9311) );
  buffer buf_n9312( .i (n9311), .o (n9312) );
  buffer buf_n9313( .i (n9312), .o (n9313) );
  buffer buf_n9314( .i (n9313), .o (n9314) );
  buffer buf_n9315( .i (n9314), .o (n9315) );
  buffer buf_n9316( .i (n9315), .o (n9316) );
  buffer buf_n5205( .i (n5204), .o (n5205) );
  buffer buf_n5206( .i (n5205), .o (n5206) );
  buffer buf_n5207( .i (n5206), .o (n5207) );
  buffer buf_n5208( .i (n5207), .o (n5208) );
  buffer buf_n5209( .i (n5208), .o (n5209) );
  buffer buf_n5210( .i (n5209), .o (n5210) );
  buffer buf_n5211( .i (n5210), .o (n5211) );
  buffer buf_n5212( .i (n5211), .o (n5212) );
  buffer buf_n5213( .i (n5212), .o (n5213) );
  buffer buf_n5214( .i (n5213), .o (n5214) );
  buffer buf_n5215( .i (n5214), .o (n5215) );
  buffer buf_n5216( .i (n5215), .o (n5216) );
  buffer buf_n5217( .i (n5216), .o (n5217) );
  buffer buf_n5218( .i (n5217), .o (n5218) );
  buffer buf_n5219( .i (n5218), .o (n5219) );
  buffer buf_n5220( .i (n5219), .o (n5220) );
  buffer buf_n5221( .i (n5220), .o (n5221) );
  buffer buf_n5222( .i (n5221), .o (n5222) );
  buffer buf_n5223( .i (n5222), .o (n5223) );
  buffer buf_n5224( .i (n5223), .o (n5224) );
  buffer buf_n5225( .i (n5224), .o (n5225) );
  buffer buf_n5226( .i (n5225), .o (n5226) );
  buffer buf_n5941( .i (n5940), .o (n5941) );
  buffer buf_n5942( .i (n5941), .o (n5942) );
  buffer buf_n5943( .i (n5942), .o (n5943) );
  assign n9317 = ~n5226 & n5943 ;
  assign n9318 = n5226 & ~n5943 ;
  assign n9319 = n9317 | n9318 ;
  buffer buf_n9320( .i (n9319), .o (n9320) );
  buffer buf_n9321( .i (n9320), .o (n9321) );
  buffer buf_n9322( .i (n9321), .o (n9322) );
  buffer buf_n9323( .i (n9322), .o (n9323) );
  buffer buf_n9324( .i (n9323), .o (n9324) );
  buffer buf_n9325( .i (n9324), .o (n9325) );
  buffer buf_n9326( .i (n9325), .o (n9326) );
  buffer buf_n9327( .i (n9326), .o (n9327) );
  buffer buf_n9328( .i (n9327), .o (n9328) );
  buffer buf_n9329( .i (n9328), .o (n9329) );
  buffer buf_n9330( .i (n9329), .o (n9330) );
  buffer buf_n9331( .i (n9330), .o (n9331) );
  buffer buf_n9332( .i (n9331), .o (n9332) );
  buffer buf_n9333( .i (n9332), .o (n9333) );
  buffer buf_n9334( .i (n9333), .o (n9334) );
  buffer buf_n9335( .i (n9334), .o (n9335) );
  buffer buf_n9336( .i (n9335), .o (n9336) );
  buffer buf_n9337( .i (n9336), .o (n9337) );
  buffer buf_n9338( .i (n9337), .o (n9338) );
  buffer buf_n9339( .i (n9338), .o (n9339) );
  buffer buf_n9340( .i (n9339), .o (n9340) );
  buffer buf_n9341( .i (n9340), .o (n9341) );
  buffer buf_n9342( .i (n9341), .o (n9342) );
  buffer buf_n9343( .i (n9342), .o (n9343) );
  buffer buf_n9344( .i (n9343), .o (n9344) );
  buffer buf_n9345( .i (n9344), .o (n9345) );
  buffer buf_n9346( .i (n9345), .o (n9346) );
  buffer buf_n9347( .i (n9346), .o (n9347) );
  buffer buf_n851( .i (N242), .o (n851) );
  buffer buf_n3459( .i (N5), .o (n3459) );
  assign n9348 = n851 & ~n3459 ;
  buffer buf_n9349( .i (n9348), .o (n9349) );
  buffer buf_n9350( .i (n9349), .o (n9350) );
  buffer buf_n9351( .i (n9350), .o (n9351) );
  buffer buf_n9352( .i (n9351), .o (n9352) );
  buffer buf_n9353( .i (n9352), .o (n9353) );
  buffer buf_n9354( .i (n9353), .o (n9354) );
  buffer buf_n9355( .i (n9354), .o (n9355) );
  buffer buf_n9356( .i (n9355), .o (n9356) );
  buffer buf_n9357( .i (n9356), .o (n9357) );
  buffer buf_n9358( .i (n9357), .o (n9358) );
  buffer buf_n9359( .i (n9358), .o (n9359) );
  buffer buf_n9360( .i (n9359), .o (n9360) );
  buffer buf_n9361( .i (n9360), .o (n9361) );
  buffer buf_n9362( .i (n9361), .o (n9362) );
  buffer buf_n9363( .i (n9362), .o (n9363) );
  buffer buf_n9364( .i (n9363), .o (n9364) );
  buffer buf_n9365( .i (n9364), .o (n9365) );
  buffer buf_n9366( .i (n9365), .o (n9366) );
  buffer buf_n9367( .i (n9366), .o (n9367) );
  buffer buf_n9368( .i (n9367), .o (n9368) );
  buffer buf_n9369( .i (n9368), .o (n9369) );
  buffer buf_n9370( .i (n9369), .o (n9370) );
  buffer buf_n9371( .i (n9370), .o (n9371) );
  buffer buf_n9372( .i (n9371), .o (n9372) );
  buffer buf_n9373( .i (n9372), .o (n9373) );
  buffer buf_n9374( .i (n9373), .o (n9374) );
  buffer buf_n9375( .i (n9374), .o (n9375) );
  buffer buf_n9376( .i (n9375), .o (n9376) );
  buffer buf_n9377( .i (n9376), .o (n9377) );
  buffer buf_n9378( .i (n9377), .o (n9378) );
  buffer buf_n9379( .i (n9378), .o (n9379) );
  buffer buf_n9380( .i (n9379), .o (n9380) );
  buffer buf_n9381( .i (n9380), .o (n9381) );
  buffer buf_n9382( .i (n9381), .o (n9382) );
  buffer buf_n9383( .i (n9382), .o (n9383) );
  buffer buf_n9384( .i (n9383), .o (n9384) );
  buffer buf_n9385( .i (n9384), .o (n9385) );
  buffer buf_n9386( .i (n9385), .o (n9386) );
  buffer buf_n9387( .i (n9386), .o (n9387) );
  buffer buf_n9388( .i (n9387), .o (n9388) );
  buffer buf_n9389( .i (n9388), .o (n9389) );
  buffer buf_n9390( .i (n9389), .o (n9390) );
  buffer buf_n9391( .i (n9390), .o (n9391) );
  buffer buf_n9392( .i (n9391), .o (n9392) );
  buffer buf_n9393( .i (n9392), .o (n9393) );
  buffer buf_n9394( .i (n9393), .o (n9394) );
  buffer buf_n9395( .i (n9394), .o (n9395) );
  buffer buf_n9396( .i (n9395), .o (n9396) );
  buffer buf_n9397( .i (n9396), .o (n9397) );
  buffer buf_n9398( .i (n9397), .o (n9398) );
  buffer buf_n9399( .i (n9398), .o (n9399) );
  buffer buf_n9400( .i (n9399), .o (n9400) );
  buffer buf_n9401( .i (n9400), .o (n9401) );
  buffer buf_n9402( .i (n9401), .o (n9402) );
  buffer buf_n9403( .i (n9402), .o (n9403) );
  buffer buf_n9404( .i (n9403), .o (n9404) );
  buffer buf_n9405( .i (n9404), .o (n9405) );
  buffer buf_n9406( .i (n9405), .o (n9406) );
  buffer buf_n9407( .i (n9406), .o (n9407) );
  buffer buf_n9408( .i (n9407), .o (n9408) );
  buffer buf_n9409( .i (n9408), .o (n9409) );
  buffer buf_n9410( .i (n9409), .o (n9410) );
  buffer buf_n9411( .i (n9410), .o (n9411) );
  buffer buf_n9412( .i (n9411), .o (n9412) );
  buffer buf_n419( .i (N15), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n396( .i (N133), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (N134), .o (n398) );
  assign n9413 = n398 & ~n3459 ;
  assign n9414 = n397 & n9413 ;
  buffer buf_n9415( .i (n9414), .o (n9415) );
  buffer buf_n9416( .i (n9415), .o (n9416) );
  buffer buf_n9417( .i (n9416), .o (n9417) );
  buffer buf_n9418( .i (n9417), .o (n9418) );
  buffer buf_n9419( .i (n9418), .o (n9419) );
  buffer buf_n9420( .i (n9419), .o (n9420) );
  buffer buf_n9421( .i (n9420), .o (n9421) );
  buffer buf_n9422( .i (n9421), .o (n9422) );
  buffer buf_n9423( .i (n9422), .o (n9423) );
  buffer buf_n9424( .i (n9423), .o (n9424) );
  buffer buf_n9425( .i (n9424), .o (n9425) );
  buffer buf_n9426( .i (n9425), .o (n9426) );
  buffer buf_n9427( .i (n9426), .o (n9427) );
  buffer buf_n9428( .i (n9427), .o (n9428) );
  buffer buf_n9429( .i (n9428), .o (n9429) );
  buffer buf_n9430( .i (n9429), .o (n9430) );
  buffer buf_n9431( .i (n9430), .o (n9431) );
  buffer buf_n9432( .i (n9431), .o (n9432) );
  buffer buf_n9433( .i (n9432), .o (n9433) );
  buffer buf_n9434( .i (n9433), .o (n9434) );
  buffer buf_n9435( .i (n9434), .o (n9435) );
  buffer buf_n9436( .i (n9435), .o (n9436) );
  buffer buf_n9437( .i (n9436), .o (n9437) );
  buffer buf_n9438( .i (n9437), .o (n9438) );
  buffer buf_n9439( .i (n9438), .o (n9439) );
  buffer buf_n9440( .i (n9439), .o (n9440) );
  buffer buf_n9441( .i (n9440), .o (n9441) );
  buffer buf_n9442( .i (n9441), .o (n9442) );
  buffer buf_n9443( .i (n9442), .o (n9443) );
  buffer buf_n9444( .i (n9443), .o (n9444) );
  buffer buf_n9445( .i (n9444), .o (n9445) );
  buffer buf_n9446( .i (n9445), .o (n9446) );
  buffer buf_n9447( .i (n9446), .o (n9447) );
  buffer buf_n9448( .i (n9447), .o (n9448) );
  buffer buf_n9449( .i (n9448), .o (n9449) );
  buffer buf_n9450( .i (n9449), .o (n9450) );
  buffer buf_n9451( .i (n9450), .o (n9451) );
  buffer buf_n9452( .i (n9451), .o (n9452) );
  buffer buf_n9453( .i (n9452), .o (n9453) );
  buffer buf_n9454( .i (n9453), .o (n9454) );
  buffer buf_n9455( .i (n9454), .o (n9455) );
  buffer buf_n9456( .i (n9455), .o (n9456) );
  buffer buf_n9457( .i (n9456), .o (n9457) );
  buffer buf_n9458( .i (n9457), .o (n9458) );
  buffer buf_n9459( .i (n9458), .o (n9459) );
  buffer buf_n9460( .i (n9459), .o (n9460) );
  buffer buf_n9461( .i (n9460), .o (n9461) );
  buffer buf_n9462( .i (n9461), .o (n9462) );
  buffer buf_n9463( .i (n9462), .o (n9463) );
  buffer buf_n9464( .i (n9463), .o (n9464) );
  buffer buf_n9465( .i (n9464), .o (n9465) );
  buffer buf_n9466( .i (n9465), .o (n9466) );
  buffer buf_n9467( .i (n9466), .o (n9467) );
  buffer buf_n9468( .i (n9467), .o (n9468) );
  buffer buf_n9469( .i (n9468), .o (n9469) );
  buffer buf_n9470( .i (n9469), .o (n9470) );
  buffer buf_n9471( .i (n9470), .o (n9471) );
  buffer buf_n9472( .i (n9471), .o (n9472) );
  buffer buf_n9473( .i (n9472), .o (n9473) );
  buffer buf_n9474( .i (n9473), .o (n9474) );
  buffer buf_n9475( .i (n9474), .o (n9475) );
  buffer buf_n9476( .i (n9475), .o (n9476) );
  buffer buf_n9477( .i (n9476), .o (n9477) );
  buffer buf_n4960( .i (n4959), .o (n4960) );
  assign n9478 = n4795 & n4828 ;
  buffer buf_n9479( .i (n9478), .o (n9479) );
  assign n9480 = n4865 & ~n9479 ;
  buffer buf_n9481( .i (n9480), .o (n9481) );
  buffer buf_n9482( .i (n9481), .o (n9482) );
  buffer buf_n9483( .i (n9482), .o (n9483) );
  buffer buf_n9484( .i (n9483), .o (n9484) );
  buffer buf_n9485( .i (n9484), .o (n9485) );
  buffer buf_n9486( .i (n9485), .o (n9486) );
  assign n9487 = n4752 & n9486 ;
  assign n9488 = n4752 | n9486 ;
  assign n9489 = ~n9487 & n9488 ;
  buffer buf_n9490( .i (n9489), .o (n9490) );
  assign n9491 = n4960 & ~n9490 ;
  buffer buf_n9492( .i (n9491), .o (n9492) );
  assign n9493 = ~n4726 & n8170 ;
  buffer buf_n9494( .i (n9493), .o (n9494) );
  assign n9495 = ~n4643 & n4793 ;
  assign n9496 = n4692 | n4793 ;
  assign n9497 = ~n9495 & n9496 ;
  buffer buf_n9498( .i (n9497), .o (n9498) );
  assign n9499 = n8135 & ~n9498 ;
  assign n9500 = ~n8135 & n9498 ;
  assign n9501 = n9499 | n9500 ;
  buffer buf_n9502( .i (n9501), .o (n9502) );
  buffer buf_n9503( .i (n9502), .o (n9503) );
  buffer buf_n9504( .i (n9503), .o (n9504) );
  buffer buf_n9505( .i (n9504), .o (n9505) );
  buffer buf_n9506( .i (n9505), .o (n9506) );
  assign n9507 = n9494 & ~n9506 ;
  assign n9508 = ~n9494 & n9506 ;
  assign n9509 = n9507 | n9508 ;
  buffer buf_n9510( .i (n9509), .o (n9510) );
  buffer buf_n9511( .i (n9510), .o (n9511) );
  buffer buf_n9512( .i (n9511), .o (n9512) );
  buffer buf_n9513( .i (n9512), .o (n9513) );
  assign n9514 = n9492 | n9513 ;
  assign n9515 = n9492 & n9513 ;
  assign n9516 = n9514 & ~n9515 ;
  buffer buf_n9517( .i (n9516), .o (n9517) );
  buffer buf_n9518( .i (n9517), .o (n9518) );
  buffer buf_n9519( .i (n9518), .o (n9519) );
  buffer buf_n9520( .i (n9519), .o (n9520) );
  buffer buf_n9521( .i (n9520), .o (n9521) );
  buffer buf_n9522( .i (n9521), .o (n9522) );
  buffer buf_n9523( .i (n9522), .o (n9523) );
  buffer buf_n9524( .i (n9523), .o (n9524) );
  buffer buf_n9525( .i (n9524), .o (n9525) );
  buffer buf_n9526( .i (n9525), .o (n9526) );
  buffer buf_n9527( .i (n9526), .o (n9527) );
  buffer buf_n9528( .i (n9527), .o (n9528) );
  buffer buf_n9529( .i (n9528), .o (n9529) );
  buffer buf_n9530( .i (n9529), .o (n9530) );
  buffer buf_n9531( .i (n9530), .o (n9531) );
  assign n9532 = n5953 & ~n9531 ;
  assign n9533 = n4643 | n4655 ;
  buffer buf_n9534( .i (n9533), .o (n9534) );
  assign n9535 = ~n4694 & n9534 ;
  buffer buf_n9536( .i (n9535), .o (n9536) );
  assign n9537 = n8136 & n9536 ;
  assign n9538 = n8136 | n9536 ;
  assign n9539 = ~n9537 & n9538 ;
  buffer buf_n9540( .i (n9539), .o (n9540) );
  buffer buf_n9541( .i (n9540), .o (n9541) );
  assign n9542 = n4726 | n9541 ;
  buffer buf_n9543( .i (n4725), .o (n9543) );
  assign n9544 = n9541 & n9543 ;
  assign n9545 = n9542 & ~n9544 ;
  buffer buf_n9546( .i (n9545), .o (n9546) );
  buffer buf_n9547( .i (n9546), .o (n9547) );
  buffer buf_n9548( .i (n9547), .o (n9548) );
  buffer buf_n9549( .i (n9548), .o (n9549) );
  assign n9550 = n9490 & n9549 ;
  assign n9551 = n9490 | n9549 ;
  assign n9552 = ~n9550 & n9551 ;
  buffer buf_n9553( .i (n9552), .o (n9553) );
  buffer buf_n9554( .i (n9553), .o (n9554) );
  buffer buf_n9555( .i (n9554), .o (n9555) );
  buffer buf_n9556( .i (n9555), .o (n9556) );
  buffer buf_n9557( .i (n9556), .o (n9557) );
  buffer buf_n9558( .i (n9557), .o (n9558) );
  buffer buf_n9559( .i (n9558), .o (n9559) );
  buffer buf_n9560( .i (n9559), .o (n9560) );
  buffer buf_n9561( .i (n9560), .o (n9561) );
  buffer buf_n9562( .i (n9561), .o (n9562) );
  buffer buf_n9563( .i (n9562), .o (n9563) );
  buffer buf_n9564( .i (n9563), .o (n9564) );
  buffer buf_n9565( .i (n9564), .o (n9565) );
  buffer buf_n9566( .i (n9565), .o (n9566) );
  buffer buf_n9567( .i (n9566), .o (n9567) );
  buffer buf_n9568( .i (n9567), .o (n9568) );
  buffer buf_n9569( .i (n9568), .o (n9569) );
  assign n9570 = ~n5953 & n9569 ;
  assign n9571 = n9532 | n9570 ;
  buffer buf_n9572( .i (n9571), .o (n9572) );
  assign n9573 = n4900 & n4933 ;
  assign n9574 = n4957 & ~n9573 ;
  buffer buf_n9575( .i (n9574), .o (n9575) );
  buffer buf_n9576( .i (n9575), .o (n9576) );
  buffer buf_n9577( .i (n9576), .o (n9577) );
  buffer buf_n9578( .i (n9577), .o (n9578) );
  buffer buf_n9579( .i (n9578), .o (n9579) );
  buffer buf_n9580( .i (n9579), .o (n9580) );
  buffer buf_n9581( .i (n9580), .o (n9581) );
  buffer buf_n9582( .i (n9581), .o (n9582) );
  buffer buf_n9583( .i (n9582), .o (n9583) );
  buffer buf_n9584( .i (n9583), .o (n9584) );
  buffer buf_n9585( .i (n9584), .o (n9585) );
  buffer buf_n9586( .i (n9585), .o (n9586) );
  buffer buf_n9587( .i (n9586), .o (n9587) );
  buffer buf_n9588( .i (n9587), .o (n9588) );
  buffer buf_n9589( .i (n9588), .o (n9589) );
  buffer buf_n9590( .i (n9589), .o (n9590) );
  buffer buf_n9591( .i (n9590), .o (n9591) );
  buffer buf_n9592( .i (n9591), .o (n9592) );
  buffer buf_n9593( .i (n9592), .o (n9593) );
  buffer buf_n9594( .i (n9593), .o (n9594) );
  buffer buf_n9595( .i (n9594), .o (n9595) );
  buffer buf_n9596( .i (n9595), .o (n9596) );
  buffer buf_n9597( .i (n9596), .o (n9597) );
  buffer buf_n9598( .i (n9597), .o (n9598) );
  assign n9599 = n9572 & ~n9598 ;
  assign n9600 = ~n9572 & n9598 ;
  assign n9601 = n9599 | n9600 ;
  buffer buf_n9602( .i (n9601), .o (n9602) );
  buffer buf_n9603( .i (n9602), .o (n9603) );
  assign n9604 = n4302 | n4371 ;
  buffer buf_n9605( .i (n9604), .o (n9605) );
  assign n9606 = ~n4402 & n9605 ;
  buffer buf_n9607( .i (n9606), .o (n9607) );
  buffer buf_n9608( .i (n9607), .o (n9608) );
  buffer buf_n4323( .i (n4322), .o (n4323) );
  buffer buf_n4324( .i (n4323), .o (n4324) );
  buffer buf_n4325( .i (n4324), .o (n4325) );
  assign n9609 = n4325 & ~n4464 ;
  assign n9610 = n4432 & ~n8808 ;
  buffer buf_n9611( .i (n9610), .o (n9611) );
  assign n9612 = n9609 | n9611 ;
  buffer buf_n9613( .i (n9612), .o (n9613) );
  assign n9614 = ~n4495 & n8727 ;
  assign n9615 = n4495 & ~n8727 ;
  assign n9616 = n9614 | n9615 ;
  buffer buf_n9617( .i (n9616), .o (n9617) );
  assign n9618 = n9613 | n9617 ;
  assign n9619 = n9613 & n9617 ;
  assign n9620 = n9618 & ~n9619 ;
  buffer buf_n9621( .i (n9620), .o (n9621) );
  assign n9622 = ~n9608 & n9621 ;
  assign n9623 = n9608 & ~n9621 ;
  assign n9624 = n9622 | n9623 ;
  buffer buf_n9625( .i (n9624), .o (n9625) );
  buffer buf_n9626( .i (n9625), .o (n9626) );
  buffer buf_n9627( .i (n9626), .o (n9627) );
  buffer buf_n9628( .i (n9627), .o (n9628) );
  buffer buf_n9629( .i (n9628), .o (n9629) );
  buffer buf_n9630( .i (n9629), .o (n9630) );
  buffer buf_n9631( .i (n9630), .o (n9631) );
  buffer buf_n9632( .i (n9631), .o (n9632) );
  buffer buf_n9633( .i (n9632), .o (n9633) );
  buffer buf_n9634( .i (n9633), .o (n9634) );
  buffer buf_n9635( .i (n9634), .o (n9635) );
  buffer buf_n9636( .i (n9635), .o (n9636) );
  buffer buf_n9637( .i (n9636), .o (n9637) );
  buffer buf_n9638( .i (n9637), .o (n9638) );
  buffer buf_n9639( .i (n9638), .o (n9639) );
  buffer buf_n9640( .i (n9639), .o (n9640) );
  buffer buf_n9641( .i (n9640), .o (n9641) );
  buffer buf_n9642( .i (n9641), .o (n9642) );
  buffer buf_n9643( .i (n9642), .o (n9643) );
  buffer buf_n9644( .i (n9643), .o (n9644) );
  buffer buf_n9645( .i (n9644), .o (n9645) );
  buffer buf_n9646( .i (n9645), .o (n9646) );
  buffer buf_n9647( .i (n9646), .o (n9647) );
  buffer buf_n9648( .i (n9647), .o (n9648) );
  buffer buf_n9649( .i (n9648), .o (n9649) );
  buffer buf_n9650( .i (n9649), .o (n9650) );
  assign n9651 = n5961 & ~n9650 ;
  assign n9652 = n4324 & n4432 ;
  assign n9653 = n4464 & ~n9652 ;
  buffer buf_n9654( .i (n9653), .o (n9654) );
  assign n9655 = ~n4497 & n9654 ;
  assign n9656 = n4497 & ~n9654 ;
  assign n9657 = n9655 | n9656 ;
  buffer buf_n9658( .i (n9657), .o (n9658) );
  buffer buf_n9659( .i (n9658), .o (n9659) );
  buffer buf_n9660( .i (n9659), .o (n9660) );
  buffer buf_n9661( .i (n9660), .o (n9661) );
  buffer buf_n9662( .i (n9661), .o (n9662) );
  buffer buf_n9663( .i (n9662), .o (n9663) );
  assign n9664 = n8810 | n8868 ;
  assign n9665 = ~n4466 & n9664 ;
  buffer buf_n9666( .i (n9665), .o (n9666) );
  assign n9667 = n8731 & n9666 ;
  assign n9668 = n8731 | n9666 ;
  assign n9669 = ~n9667 & n9668 ;
  buffer buf_n9670( .i (n9669), .o (n9670) );
  assign n9671 = n4532 | n9670 ;
  assign n9672 = n4532 & n9670 ;
  assign n9673 = n9671 & ~n9672 ;
  buffer buf_n9674( .i (n9673), .o (n9674) );
  assign n9675 = n9663 & n9674 ;
  assign n9676 = n9663 | n9674 ;
  assign n9677 = ~n9675 & n9676 ;
  buffer buf_n9678( .i (n9677), .o (n9678) );
  buffer buf_n9679( .i (n9678), .o (n9679) );
  buffer buf_n9680( .i (n9679), .o (n9680) );
  buffer buf_n9681( .i (n9680), .o (n9681) );
  buffer buf_n9682( .i (n9681), .o (n9682) );
  buffer buf_n9683( .i (n9682), .o (n9683) );
  buffer buf_n9684( .i (n9683), .o (n9684) );
  buffer buf_n9685( .i (n9684), .o (n9685) );
  buffer buf_n9686( .i (n9685), .o (n9686) );
  buffer buf_n9687( .i (n9686), .o (n9687) );
  buffer buf_n9688( .i (n9687), .o (n9688) );
  buffer buf_n9689( .i (n9688), .o (n9689) );
  buffer buf_n9690( .i (n9689), .o (n9690) );
  buffer buf_n9691( .i (n9690), .o (n9691) );
  buffer buf_n9692( .i (n9691), .o (n9692) );
  buffer buf_n9693( .i (n9692), .o (n9693) );
  buffer buf_n9694( .i (n9693), .o (n9694) );
  buffer buf_n9695( .i (n9694), .o (n9695) );
  buffer buf_n9696( .i (n9695), .o (n9696) );
  buffer buf_n9697( .i (n9696), .o (n9697) );
  buffer buf_n9698( .i (n9697), .o (n9698) );
  buffer buf_n9699( .i (n9698), .o (n9699) );
  assign n9700 = ~n5961 & n9699 ;
  assign n9701 = n9651 | n9700 ;
  buffer buf_n9702( .i (n9701), .o (n9702) );
  assign n9703 = n9603 & ~n9702 ;
  assign n9704 = ~n9603 & n9702 ;
  assign n9705 = n9703 | n9704 ;
  buffer buf_n9706( .i (n9705), .o (n9706) );
  buffer buf_n9707( .i (n9706), .o (n9707) );
  buffer buf_n9708( .i (n9707), .o (n9708) );
  buffer buf_n9709( .i (n9708), .o (n9709) );
  buffer buf_n9710( .i (n9709), .o (n9710) );
  buffer buf_n9711( .i (n9710), .o (n9711) );
  buffer buf_n9712( .i (n9711), .o (n9712) );
  buffer buf_n9713( .i (n9712), .o (n9713) );
  buffer buf_n9714( .i (n9713), .o (n9714) );
  buffer buf_n9715( .i (n9714), .o (n9715) );
  buffer buf_n9716( .i (n9715), .o (n9716) );
  buffer buf_n9717( .i (n9716), .o (n9717) );
  buffer buf_n9718( .i (n9717), .o (n9718) );
  buffer buf_n9719( .i (n9718), .o (n9719) );
  buffer buf_n3871( .i (n3870), .o (n3871) );
  buffer buf_n9720( .i (n6189), .o (n9720) );
  assign n9721 = n3875 & n9720 ;
  assign n9722 = n3871 | n9721 ;
  buffer buf_n9723( .i (n9722), .o (n9723) );
  assign n9724 = ~n4163 & n6014 ;
  assign n9725 = n4163 & ~n6014 ;
  assign n9726 = n9724 | n9725 ;
  buffer buf_n9727( .i (n9726), .o (n9727) );
  assign n9728 = ~n3738 & n9727 ;
  assign n9729 = n3738 & ~n9727 ;
  assign n9730 = n9728 | n9729 ;
  buffer buf_n9731( .i (n9730), .o (n9731) );
  assign n9732 = n6018 | n6062 ;
  buffer buf_n9733( .i (n9732), .o (n9733) );
  assign n9734 = ~n6110 & n9733 ;
  buffer buf_n9735( .i (n9734), .o (n9735) );
  buffer buf_n9736( .i (n9735), .o (n9736) );
  buffer buf_n9737( .i (n9736), .o (n9737) );
  buffer buf_n9738( .i (n9737), .o (n9738) );
  buffer buf_n9739( .i (n9738), .o (n9739) );
  buffer buf_n9740( .i (n9739), .o (n9740) );
  assign n9741 = n8298 & ~n9740 ;
  assign n9742 = ~n8298 & n9740 ;
  assign n9743 = n9741 | n9742 ;
  buffer buf_n9744( .i (n9743), .o (n9744) );
  assign n9745 = n4128 & n6146 ;
  buffer buf_n9746( .i (n9745), .o (n9746) );
  buffer buf_n9747( .i (n9746), .o (n9747) );
  buffer buf_n9748( .i (n9747), .o (n9748) );
  buffer buf_n9749( .i (n9748), .o (n9749) );
  buffer buf_n9750( .i (n9749), .o (n9750) );
  buffer buf_n9751( .i (n9750), .o (n9751) );
  buffer buf_n9752( .i (n9751), .o (n9752) );
  assign n9753 = n9744 & ~n9752 ;
  buffer buf_n9754( .i (n9753), .o (n9754) );
  assign n9755 = n4080 & ~n6148 ;
  buffer buf_n9756( .i (n9755), .o (n9756) );
  assign n9757 = n3981 | n6016 ;
  assign n9758 = n4037 & n6016 ;
  assign n9759 = n9757 & ~n9758 ;
  buffer buf_n9760( .i (n9759), .o (n9760) );
  assign n9761 = n4167 & n9760 ;
  assign n9762 = n4167 | n9760 ;
  assign n9763 = ~n9761 & n9762 ;
  buffer buf_n9764( .i (n9763), .o (n9764) );
  buffer buf_n9765( .i (n9764), .o (n9765) );
  buffer buf_n9766( .i (n9765), .o (n9766) );
  buffer buf_n9767( .i (n9766), .o (n9767) );
  buffer buf_n9768( .i (n9767), .o (n9768) );
  assign n9769 = ~n9756 & n9768 ;
  assign n9770 = n9756 & ~n9768 ;
  assign n9771 = n9769 | n9770 ;
  buffer buf_n9772( .i (n9771), .o (n9772) );
  buffer buf_n9773( .i (n9772), .o (n9773) );
  buffer buf_n9774( .i (n9773), .o (n9774) );
  buffer buf_n9775( .i (n9774), .o (n9775) );
  assign n9776 = n9754 & ~n9775 ;
  assign n9777 = ~n9754 & n9775 ;
  assign n9778 = n9776 | n9777 ;
  buffer buf_n9779( .i (n9778), .o (n9779) );
  buffer buf_n9780( .i (n9779), .o (n9780) );
  buffer buf_n9781( .i (n9780), .o (n9781) );
  buffer buf_n9782( .i (n9781), .o (n9782) );
  buffer buf_n9783( .i (n9782), .o (n9783) );
  buffer buf_n9784( .i (n9783), .o (n9784) );
  buffer buf_n9785( .i (n9784), .o (n9785) );
  buffer buf_n9786( .i (n9785), .o (n9786) );
  buffer buf_n9787( .i (n9786), .o (n9787) );
  buffer buf_n9788( .i (n9787), .o (n9788) );
  buffer buf_n9789( .i (n9788), .o (n9789) );
  buffer buf_n9790( .i (n9789), .o (n9790) );
  buffer buf_n9791( .i (n9790), .o (n9791) );
  buffer buf_n9792( .i (n9791), .o (n9792) );
  buffer buf_n9793( .i (n9792), .o (n9793) );
  buffer buf_n9794( .i (n9793), .o (n9794) );
  buffer buf_n9795( .i (n9794), .o (n9795) );
  buffer buf_n9796( .i (n9795), .o (n9796) );
  buffer buf_n9797( .i (n9796), .o (n9797) );
  buffer buf_n9798( .i (n9797), .o (n9798) );
  buffer buf_n9799( .i (n9798), .o (n9799) );
  buffer buf_n9800( .i (n9799), .o (n9800) );
  buffer buf_n9801( .i (n9800), .o (n9801) );
  buffer buf_n9802( .i (n9801), .o (n9802) );
  buffer buf_n9803( .i (n9802), .o (n9803) );
  buffer buf_n9804( .i (n9803), .o (n9804) );
  assign n9805 = n5973 | n9804 ;
  assign n9806 = n3981 | n3989 ;
  buffer buf_n9807( .i (n9806), .o (n9807) );
  assign n9808 = ~n4039 & n9807 ;
  buffer buf_n9809( .i (n9808), .o (n9809) );
  assign n9810 = ~n4168 & n9809 ;
  assign n9811 = n4168 & ~n9809 ;
  assign n9812 = n9810 | n9811 ;
  buffer buf_n9813( .i (n9812), .o (n9813) );
  buffer buf_n9814( .i (n9813), .o (n9814) );
  assign n9815 = n4080 | n9814 ;
  buffer buf_n9816( .i (n4079), .o (n9816) );
  assign n9817 = n9814 & n9816 ;
  assign n9818 = n9815 & ~n9817 ;
  buffer buf_n9819( .i (n9818), .o (n9819) );
  buffer buf_n9820( .i (n9819), .o (n9820) );
  buffer buf_n9821( .i (n9820), .o (n9821) );
  buffer buf_n9822( .i (n9821), .o (n9822) );
  assign n9823 = n9744 & n9822 ;
  assign n9824 = n9744 | n9822 ;
  assign n9825 = ~n9823 & n9824 ;
  buffer buf_n9826( .i (n9825), .o (n9826) );
  buffer buf_n9827( .i (n9826), .o (n9827) );
  buffer buf_n9828( .i (n9827), .o (n9828) );
  buffer buf_n9829( .i (n9828), .o (n9829) );
  buffer buf_n9830( .i (n9829), .o (n9830) );
  buffer buf_n9831( .i (n9830), .o (n9831) );
  buffer buf_n9832( .i (n9831), .o (n9832) );
  buffer buf_n9833( .i (n9832), .o (n9833) );
  buffer buf_n9834( .i (n9833), .o (n9834) );
  buffer buf_n9835( .i (n9834), .o (n9835) );
  buffer buf_n9836( .i (n9835), .o (n9836) );
  buffer buf_n9837( .i (n9836), .o (n9837) );
  buffer buf_n9838( .i (n9837), .o (n9838) );
  buffer buf_n9839( .i (n9838), .o (n9839) );
  buffer buf_n9840( .i (n9839), .o (n9840) );
  buffer buf_n9841( .i (n9840), .o (n9841) );
  buffer buf_n9842( .i (n9841), .o (n9842) );
  buffer buf_n9843( .i (n9842), .o (n9843) );
  buffer buf_n9844( .i (n9843), .o (n9844) );
  buffer buf_n9845( .i (n9844), .o (n9845) );
  buffer buf_n9846( .i (n9845), .o (n9846) );
  buffer buf_n9847( .i (n9846), .o (n9847) );
  buffer buf_n9848( .i (n9847), .o (n9848) );
  buffer buf_n9849( .i (n9848), .o (n9849) );
  buffer buf_n9850( .i (n9849), .o (n9850) );
  buffer buf_n9851( .i (n9850), .o (n9851) );
  buffer buf_n9852( .i (n9851), .o (n9852) );
  buffer buf_n9853( .i (n9852), .o (n9853) );
  assign n9854 = n5973 & n9853 ;
  assign n9855 = n9805 & ~n9854 ;
  buffer buf_n9856( .i (n9855), .o (n9856) );
  assign n9857 = ~n9731 & n9856 ;
  assign n9858 = n9731 & ~n9856 ;
  assign n9859 = n9857 | n9858 ;
  buffer buf_n9860( .i (n9859), .o (n9860) );
  buffer buf_n9861( .i (n9860), .o (n9861) );
  buffer buf_n9862( .i (n9861), .o (n9862) );
  buffer buf_n9863( .i (n9862), .o (n9863) );
  assign n9864 = n9723 | n9863 ;
  assign n9865 = n9723 & n9863 ;
  assign n9866 = n9864 & ~n9865 ;
  buffer buf_n9867( .i (n9866), .o (n9867) );
  assign n9868 = n5074 & n5084 ;
  buffer buf_n9869( .i (n9868), .o (n9869) );
  assign n9870 = n5109 & ~n9869 ;
  buffer buf_n9871( .i (n9870), .o (n9871) );
  assign n9872 = ~n5153 & n5181 ;
  assign n9873 = n9871 | n9872 ;
  buffer buf_n9874( .i (n9873), .o (n9874) );
  assign n9875 = ~n9168 & n9225 ;
  assign n9876 = n9168 & ~n9225 ;
  assign n9877 = n9875 | n9876 ;
  buffer buf_n9878( .i (n9877), .o (n9878) );
  assign n9879 = n9874 & ~n9878 ;
  assign n9880 = ~n9874 & n9878 ;
  assign n9881 = n9879 | n9880 ;
  buffer buf_n9882( .i (n9881), .o (n9882) );
  assign n9883 = n5248 & n9882 ;
  assign n9884 = n5248 | n9882 ;
  assign n9885 = ~n9883 & n9884 ;
  buffer buf_n9886( .i (n9885), .o (n9886) );
  buffer buf_n9887( .i (n9886), .o (n9887) );
  buffer buf_n9888( .i (n9887), .o (n9888) );
  buffer buf_n9889( .i (n9888), .o (n9889) );
  buffer buf_n9890( .i (n9889), .o (n9890) );
  buffer buf_n9891( .i (n9890), .o (n9891) );
  buffer buf_n9892( .i (n9891), .o (n9892) );
  buffer buf_n9893( .i (n9892), .o (n9893) );
  buffer buf_n9894( .i (n9893), .o (n9894) );
  buffer buf_n9895( .i (n9894), .o (n9895) );
  buffer buf_n9896( .i (n9895), .o (n9896) );
  buffer buf_n9897( .i (n9896), .o (n9897) );
  buffer buf_n9898( .i (n9897), .o (n9898) );
  buffer buf_n9899( .i (n9898), .o (n9899) );
  buffer buf_n9900( .i (n9899), .o (n9900) );
  assign n9901 = n5943 & ~n9900 ;
  buffer buf_n5062( .i (n5061), .o (n5062) );
  assign n9902 = n5053 | n5111 ;
  assign n9903 = ~n5062 & n9902 ;
  buffer buf_n9904( .i (n9903), .o (n9904) );
  assign n9905 = n5157 & ~n9904 ;
  assign n9906 = ~n5157 & n9904 ;
  assign n9907 = n9905 | n9906 ;
  buffer buf_n9908( .i (n9907), .o (n9908) );
  assign n9909 = n5111 & ~n5182 ;
  buffer buf_n5075( .i (n5074), .o (n5075) );
  assign n9910 = ~n5075 & n5179 ;
  buffer buf_n9911( .i (n9910), .o (n9911) );
  buffer buf_n9912( .i (n9911), .o (n9912) );
  buffer buf_n9913( .i (n9912), .o (n9913) );
  assign n9914 = n9909 | n9913 ;
  buffer buf_n9915( .i (n9914), .o (n9915) );
  assign n9916 = n9172 & ~n9915 ;
  assign n9917 = ~n9172 & n9915 ;
  assign n9918 = n9916 | n9917 ;
  buffer buf_n9919( .i (n9918), .o (n9919) );
  assign n9920 = n9908 | n9919 ;
  assign n9921 = n9908 & n9919 ;
  assign n9922 = n9920 & ~n9921 ;
  buffer buf_n9923( .i (n9922), .o (n9923) );
  buffer buf_n9924( .i (n9923), .o (n9924) );
  buffer buf_n9925( .i (n9924), .o (n9925) );
  buffer buf_n9926( .i (n9925), .o (n9926) );
  buffer buf_n9927( .i (n9926), .o (n9927) );
  buffer buf_n9928( .i (n9927), .o (n9928) );
  buffer buf_n9929( .i (n9928), .o (n9929) );
  buffer buf_n9930( .i (n9929), .o (n9930) );
  buffer buf_n9931( .i (n9930), .o (n9931) );
  buffer buf_n9932( .i (n9931), .o (n9932) );
  buffer buf_n9933( .i (n9932), .o (n9933) );
  buffer buf_n9934( .i (n9933), .o (n9934) );
  buffer buf_n9935( .i (n9934), .o (n9935) );
  buffer buf_n9936( .i (n9935), .o (n9936) );
  assign n9937 = n5943 | n9936 ;
  assign n9938 = ~n9901 & n9937 ;
  buffer buf_n9939( .i (n9938), .o (n9939) );
  assign n9940 = n5406 | n5889 ;
  buffer buf_n9941( .i (n9940), .o (n9941) );
  assign n9942 = ~n5911 & n9941 ;
  buffer buf_n9943( .i (n9942), .o (n9943) );
  assign n9944 = n5314 | n9077 ;
  assign n9945 = n5314 & n9077 ;
  assign n9946 = n9944 & ~n9945 ;
  buffer buf_n9947( .i (n9946), .o (n9947) );
  assign n9948 = n9943 & n9947 ;
  assign n9949 = n9943 | n9947 ;
  assign n9950 = ~n9948 & n9949 ;
  buffer buf_n9951( .i (n9950), .o (n9951) );
  buffer buf_n9952( .i (n9951), .o (n9952) );
  buffer buf_n9953( .i (n9952), .o (n9953) );
  buffer buf_n9954( .i (n9953), .o (n9954) );
  assign n9955 = n8979 | n9954 ;
  assign n9956 = n8979 & n9954 ;
  assign n9957 = n9955 & ~n9956 ;
  buffer buf_n9958( .i (n9957), .o (n9958) );
  buffer buf_n9959( .i (n9958), .o (n9959) );
  buffer buf_n9960( .i (n9959), .o (n9960) );
  buffer buf_n9961( .i (n9960), .o (n9961) );
  buffer buf_n9962( .i (n9961), .o (n9962) );
  assign n9963 = n5884 | n9962 ;
  assign n9964 = n5444 & n8979 ;
  assign n9965 = n5500 & ~n9964 ;
  buffer buf_n9966( .i (n9965), .o (n9966) );
  assign n9967 = ~n5913 & n9023 ;
  buffer buf_n9968( .i (n9967), .o (n9968) );
  assign n9969 = n5272 & ~n5331 ;
  buffer buf_n9970( .i (n9969), .o (n9970) );
  buffer buf_n9971( .i (n9970), .o (n9971) );
  buffer buf_n9972( .i (n9971), .o (n9972) );
  assign n9973 = ~n5307 & n5335 ;
  assign n9974 = n9972 | n9973 ;
  buffer buf_n9975( .i (n9974), .o (n9975) );
  buffer buf_n9976( .i (n9975), .o (n9976) );
  buffer buf_n9977( .i (n9976), .o (n9977) );
  buffer buf_n9978( .i (n9977), .o (n9978) );
  assign n9979 = n9968 | n9978 ;
  assign n9980 = n9968 & n9978 ;
  assign n9981 = n9979 & ~n9980 ;
  buffer buf_n9982( .i (n9981), .o (n9982) );
  buffer buf_n9983( .i (n9982), .o (n9983) );
  buffer buf_n9984( .i (n9983), .o (n9984) );
  buffer buf_n9985( .i (n9984), .o (n9985) );
  buffer buf_n9986( .i (n9985), .o (n9986) );
  assign n9987 = n9966 & ~n9986 ;
  assign n9988 = ~n9966 & n9986 ;
  assign n9989 = n9987 | n9988 ;
  buffer buf_n9990( .i (n9989), .o (n9990) );
  buffer buf_n9991( .i (n9990), .o (n9991) );
  assign n9992 = n5884 & n9991 ;
  assign n9993 = n9963 & ~n9992 ;
  buffer buf_n9994( .i (n9993), .o (n9994) );
  assign n9995 = n5369 & n5413 ;
  assign n9996 = n5436 & ~n9995 ;
  buffer buf_n9997( .i (n9996), .o (n9997) );
  buffer buf_n9998( .i (n9997), .o (n9998) );
  buffer buf_n9999( .i (n9998), .o (n9999) );
  buffer buf_n10000( .i (n9999), .o (n10000) );
  buffer buf_n10001( .i (n10000), .o (n10001) );
  buffer buf_n10002( .i (n10001), .o (n10002) );
  buffer buf_n10003( .i (n10002), .o (n10003) );
  buffer buf_n10004( .i (n10003), .o (n10004) );
  buffer buf_n10005( .i (n10004), .o (n10005) );
  buffer buf_n10006( .i (n10005), .o (n10006) );
  buffer buf_n10007( .i (n10006), .o (n10007) );
  buffer buf_n10008( .i (n10007), .o (n10008) );
  buffer buf_n10009( .i (n10008), .o (n10009) );
  buffer buf_n10010( .i (n10009), .o (n10010) );
  buffer buf_n10011( .i (n10010), .o (n10011) );
  buffer buf_n10012( .i (n10011), .o (n10012) );
  buffer buf_n10013( .i (n10012), .o (n10013) );
  assign n10014 = n9994 & ~n10013 ;
  assign n10015 = ~n9994 & n10013 ;
  assign n10016 = n10014 | n10015 ;
  buffer buf_n10017( .i (n10016), .o (n10017) );
  buffer buf_n10018( .i (n10017), .o (n10018) );
  buffer buf_n10019( .i (n10018), .o (n10019) );
  assign n10020 = ~n9939 & n10019 ;
  assign n10021 = n9939 & ~n10019 ;
  assign n10022 = n10020 | n10021 ;
  buffer buf_n10023( .i (n10022), .o (n10023) );
  buffer buf_n10024( .i (n10023), .o (n10024) );
  buffer buf_n10025( .i (n10024), .o (n10025) );
  buffer buf_n10026( .i (n10025), .o (n10026) );
  buffer buf_n10027( .i (n10026), .o (n10027) );
  buffer buf_n10028( .i (n10027), .o (n10028) );
  buffer buf_n10029( .i (n10028), .o (n10029) );
  buffer buf_n10030( .i (n10029), .o (n10030) );
  buffer buf_n10031( .i (n10030), .o (n10031) );
  buffer buf_n10032( .i (n10031), .o (n10032) );
  buffer buf_n10033( .i (n10032), .o (n10033) );
  buffer buf_n10034( .i (n10033), .o (n10034) );
  buffer buf_n10035( .i (n10034), .o (n10035) );
  buffer buf_n10036( .i (n10035), .o (n10036) );
  buffer buf_n10037( .i (n10036), .o (n10037) );
  buffer buf_n10038( .i (n10037), .o (n10038) );
  buffer buf_n10039( .i (n10038), .o (n10039) );
  buffer buf_n10040( .i (n10039), .o (n10040) );
  buffer buf_n10041( .i (n10040), .o (n10041) );
  buffer buf_n10042( .i (n10041), .o (n10042) );
  buffer buf_n10043( .i (n10042), .o (n10043) );
  buffer buf_n10044( .i (n10043), .o (n10044) );
  buffer buf_n10045( .i (n10044), .o (n10045) );
  buffer buf_n10046( .i (n10045), .o (n10046) );
  buffer buf_n10047( .i (n10046), .o (n10047) );
  assign n10048 = n5587 | n5795 ;
  assign n10049 = n5557 & n5792 ;
  buffer buf_n10050( .i (n10049), .o (n10050) );
  buffer buf_n10051( .i (n10050), .o (n10051) );
  buffer buf_n10052( .i (n10051), .o (n10052) );
  assign n10053 = n10048 & ~n10052 ;
  buffer buf_n10054( .i (n10053), .o (n10054) );
  buffer buf_n10055( .i (n10054), .o (n10055) );
  buffer buf_n10056( .i (n10055), .o (n10056) );
  assign n10057 = n5608 | n10056 ;
  assign n10058 = n5608 & n10056 ;
  assign n10059 = n10057 & ~n10058 ;
  buffer buf_n10060( .i (n10059), .o (n10060) );
  assign n10061 = n5830 & n5851 ;
  assign n10062 = n5868 & ~n10061 ;
  buffer buf_n10063( .i (n10062), .o (n10063) );
  assign n10068 = n5777 & ~n10063 ;
  assign n10069 = ~n5777 & n10063 ;
  assign n10070 = n10068 | n10069 ;
  buffer buf_n10071( .i (n10070), .o (n10071) );
  buffer buf_n10072( .i (n10071), .o (n10072) );
  assign n10073 = n10060 & n10072 ;
  assign n10074 = n10060 | n10072 ;
  assign n10075 = ~n10073 & n10074 ;
  buffer buf_n10076( .i (n10075), .o (n10076) );
  assign n10077 = n5767 & ~n10076 ;
  buffer buf_n10078( .i (n10077), .o (n10078) );
  buffer buf_n3334( .i (n3333), .o (n3334) );
  buffer buf_n3335( .i (n3334), .o (n3335) );
  buffer buf_n3336( .i (n3335), .o (n3336) );
  buffer buf_n10064( .i (n10063), .o (n10064) );
  buffer buf_n10065( .i (n10064), .o (n10065) );
  buffer buf_n10066( .i (n10065), .o (n10066) );
  buffer buf_n10067( .i (n10066), .o (n10067) );
  assign n10079 = n5555 & ~n5567 ;
  buffer buf_n5558( .i (n5557), .o (n5558) );
  assign n10080 = n5558 & n5567 ;
  assign n10081 = n10079 | n10080 ;
  buffer buf_n10082( .i (n10081), .o (n10082) );
  buffer buf_n10083( .i (n10082), .o (n10083) );
  assign n10084 = n5826 & ~n10083 ;
  buffer buf_n10085( .i (n10084), .o (n10085) );
  buffer buf_n10086( .i (n10085), .o (n10086) );
  assign n10087 = n5608 & n10086 ;
  assign n10088 = n7238 & ~n10085 ;
  buffer buf_n10089( .i (n5607), .o (n10089) );
  assign n10090 = n10088 & ~n10089 ;
  assign n10091 = n10087 | n10090 ;
  buffer buf_n10092( .i (n10091), .o (n10092) );
  assign n10093 = ~n10067 & n10092 ;
  assign n10094 = n10067 & ~n10092 ;
  assign n10095 = n10093 | n10094 ;
  buffer buf_n10096( .i (n10095), .o (n10096) );
  assign n10097 = n5767 | n10096 ;
  assign n10098 = n3336 & n10097 ;
  assign n10099 = ~n10078 & n10098 ;
  assign n10100 = ~n5736 & n10076 ;
  assign n10101 = ~n3333 & n5734 ;
  buffer buf_n10102( .i (n10101), .o (n10102) );
  assign n10103 = n10096 & n10102 ;
  assign n10104 = n10100 | n10103 ;
  buffer buf_n10105( .i (n10104), .o (n10105) );
  assign n10106 = n10099 | n10105 ;
  buffer buf_n10107( .i (n10106), .o (n10107) );
  buffer buf_n10108( .i (n10107), .o (n10108) );
  buffer buf_n10109( .i (n10108), .o (n10109) );
  buffer buf_n10110( .i (n10109), .o (n10110) );
  assign n10111 = ~n5675 & n5723 ;
  buffer buf_n10112( .i (n10111), .o (n10112) );
  assign n10113 = n5728 & ~n10112 ;
  buffer buf_n10114( .i (n10113), .o (n10114) );
  buffer buf_n10115( .i (n10114), .o (n10115) );
  buffer buf_n10116( .i (n10115), .o (n10116) );
  buffer buf_n10117( .i (n10116), .o (n10117) );
  assign n10118 = ~n5712 & n7126 ;
  buffer buf_n10119( .i (n10118), .o (n10119) );
  buffer buf_n10120( .i (n10119), .o (n10120) );
  buffer buf_n10121( .i (n10120), .o (n10121) );
  buffer buf_n10122( .i (n10121), .o (n10122) );
  buffer buf_n10123( .i (n10122), .o (n10123) );
  buffer buf_n10124( .i (n10123), .o (n10124) );
  assign n10125 = n3628 & n5743 ;
  buffer buf_n10126( .i (n10125), .o (n10126) );
  assign n10127 = n5747 & ~n10126 ;
  buffer buf_n10128( .i (n10127), .o (n10128) );
  assign n10129 = n7019 & n10128 ;
  assign n10130 = n7019 | n10128 ;
  assign n10131 = ~n10129 & n10130 ;
  buffer buf_n10132( .i (n10131), .o (n10132) );
  assign n10135 = ~n10124 & n10132 ;
  assign n10136 = n10124 & ~n10132 ;
  assign n10137 = n10135 | n10136 ;
  buffer buf_n10138( .i (n10137), .o (n10138) );
  assign n10139 = n10117 & ~n10138 ;
  buffer buf_n10140( .i (n10139), .o (n10140) );
  assign n10141 = ~n10117 & n10138 ;
  assign n10142 = n3334 | n10141 ;
  assign n10143 = n10140 | n10142 ;
  buffer buf_n10144( .i (n10143), .o (n10144) );
  buffer buf_n10145( .i (n10144), .o (n10145) );
  assign n10146 = ~n5724 & n5749 ;
  buffer buf_n10147( .i (n10146), .o (n10147) );
  buffer buf_n3620( .i (n3619), .o (n3620) );
  buffer buf_n3621( .i (n3620), .o (n3621) );
  assign n10148 = n3621 | n5707 ;
  buffer buf_n10149( .i (n10148), .o (n10149) );
  buffer buf_n10150( .i (n10149), .o (n10150) );
  buffer buf_n10151( .i (n10150), .o (n10151) );
  buffer buf_n3622( .i (n3621), .o (n3622) );
  buffer buf_n3623( .i (n3622), .o (n3623) );
  buffer buf_n3624( .i (n3623), .o (n3624) );
  buffer buf_n5717( .i (n5716), .o (n5717) );
  buffer buf_n5718( .i (n5717), .o (n5718) );
  assign n10152 = n5712 | n5718 ;
  assign n10153 = n3624 & ~n10152 ;
  assign n10154 = n10151 & ~n10153 ;
  buffer buf_n10155( .i (n10154), .o (n10155) );
  buffer buf_n10156( .i (n10155), .o (n10156) );
  buffer buf_n10157( .i (n10156), .o (n10157) );
  assign n10158 = ~n10147 & n10157 ;
  assign n10159 = n10147 & ~n10157 ;
  assign n10160 = n10158 | n10159 ;
  buffer buf_n10161( .i (n10160), .o (n10161) );
  buffer buf_n10162( .i (n10161), .o (n10162) );
  buffer buf_n10163( .i (n10162), .o (n10163) );
  buffer buf_n10164( .i (n10163), .o (n10164) );
  buffer buf_n10133( .i (n10132), .o (n10133) );
  buffer buf_n10134( .i (n10133), .o (n10134) );
  assign n10165 = n5764 & ~n10134 ;
  assign n10166 = ~n5764 & n10134 ;
  assign n10167 = n10165 | n10166 ;
  buffer buf_n10168( .i (n10167), .o (n10168) );
  assign n10169 = n10164 & n10168 ;
  buffer buf_n10170( .i (n10169), .o (n10170) );
  assign n10171 = n10164 | n10168 ;
  assign n10172 = n3336 & n10171 ;
  assign n10173 = ~n10170 & n10172 ;
  assign n10174 = n10145 & ~n10173 ;
  buffer buf_n10175( .i (n10174), .o (n10175) );
  assign n10176 = n5739 & n5752 ;
  assign n10177 = n5739 | n5752 ;
  assign n10178 = ~n10176 & n10177 ;
  buffer buf_n10179( .i (n10178), .o (n10179) );
  buffer buf_n10180( .i (n10179), .o (n10180) );
  buffer buf_n10181( .i (n10180), .o (n10181) );
  buffer buf_n10182( .i (n10181), .o (n10182) );
  buffer buf_n10183( .i (n10182), .o (n10183) );
  buffer buf_n10184( .i (n10183), .o (n10184) );
  buffer buf_n10185( .i (n10184), .o (n10185) );
  buffer buf_n10186( .i (n10185), .o (n10186) );
  buffer buf_n10187( .i (n10186), .o (n10187) );
  buffer buf_n10188( .i (n10187), .o (n10188) );
  buffer buf_n10189( .i (n10188), .o (n10189) );
  buffer buf_n10190( .i (n10189), .o (n10190) );
  buffer buf_n10191( .i (n10190), .o (n10191) );
  buffer buf_n10192( .i (n10191), .o (n10192) );
  assign n10193 = n10175 | n10192 ;
  assign n10194 = n10175 & n10192 ;
  assign n10195 = n10193 & ~n10194 ;
  buffer buf_n10196( .i (n10195), .o (n10196) );
  assign n10197 = n10110 | n10196 ;
  assign n10198 = n10110 & n10196 ;
  assign n10199 = n10197 & ~n10198 ;
  buffer buf_n10200( .i (n10199), .o (n10200) );
  buffer buf_n10201( .i (n10200), .o (n10201) );
  buffer buf_n10202( .i (n10201), .o (n10202) );
  buffer buf_n10203( .i (n10202), .o (n10203) );
  buffer buf_n10204( .i (n10203), .o (n10204) );
  buffer buf_n10205( .i (n10204), .o (n10205) );
  buffer buf_n10206( .i (n10205), .o (n10206) );
  buffer buf_n10207( .i (n10206), .o (n10207) );
  buffer buf_n10208( .i (n10207), .o (n10208) );
  buffer buf_n10209( .i (n10208), .o (n10209) );
  buffer buf_n10210( .i (n10209), .o (n10210) );
  buffer buf_n10211( .i (n10210), .o (n10211) );
  buffer buf_n10212( .i (n10211), .o (n10212) );
  buffer buf_n10213( .i (n10212), .o (n10213) );
  buffer buf_n10214( .i (n10213), .o (n10214) );
  buffer buf_n10215( .i (n10214), .o (n10215) );
  buffer buf_n10216( .i (n10215), .o (n10216) );
  buffer buf_n10217( .i (n10216), .o (n10217) );
  buffer buf_n10218( .i (n10217), .o (n10218) );
  buffer buf_n10219( .i (n10218), .o (n10219) );
  buffer buf_n10220( .i (n10219), .o (n10220) );
  buffer buf_n10221( .i (n10220), .o (n10221) );
  buffer buf_n10222( .i (n10221), .o (n10222) );
  buffer buf_n10223( .i (n10222), .o (n10223) );
  buffer buf_n10224( .i (n10223), .o (n10224) );
  buffer buf_n10225( .i (n10224), .o (n10225) );
  buffer buf_n10226( .i (n10225), .o (n10226) );
  buffer buf_n10227( .i (n10226), .o (n10227) );
  buffer buf_n10228( .i (n10227), .o (n10228) );
  buffer buf_n10229( .i (n10228), .o (n10229) );
  buffer buf_n10230( .i (n10229), .o (n10230) );
  buffer buf_n10231( .i (n10230), .o (n10231) );
  buffer buf_n208( .i (N1), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n528( .i (N163), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  assign n10232 = n209 & n529 ;
  buffer buf_n10233( .i (n10232), .o (n10233) );
  buffer buf_n10234( .i (n10233), .o (n10234) );
  buffer buf_n10235( .i (n10234), .o (n10235) );
  buffer buf_n10236( .i (n10235), .o (n10236) );
  buffer buf_n10237( .i (n10236), .o (n10237) );
  buffer buf_n10238( .i (n10237), .o (n10238) );
  buffer buf_n10239( .i (n10238), .o (n10239) );
  buffer buf_n10240( .i (n10239), .o (n10240) );
  buffer buf_n10241( .i (n10240), .o (n10241) );
  buffer buf_n10242( .i (n10241), .o (n10242) );
  buffer buf_n10243( .i (n10242), .o (n10243) );
  buffer buf_n10244( .i (n10243), .o (n10244) );
  buffer buf_n10245( .i (n10244), .o (n10245) );
  buffer buf_n10246( .i (n10245), .o (n10246) );
  buffer buf_n10247( .i (n10246), .o (n10247) );
  buffer buf_n10248( .i (n10247), .o (n10248) );
  buffer buf_n10249( .i (n10248), .o (n10249) );
  buffer buf_n10250( .i (n10249), .o (n10250) );
  buffer buf_n10251( .i (n10250), .o (n10251) );
  buffer buf_n10252( .i (n10251), .o (n10252) );
  buffer buf_n10253( .i (n10252), .o (n10253) );
  buffer buf_n10254( .i (n10253), .o (n10254) );
  buffer buf_n10255( .i (n10254), .o (n10255) );
  buffer buf_n10256( .i (n10255), .o (n10256) );
  buffer buf_n10257( .i (n10256), .o (n10257) );
  buffer buf_n10258( .i (n10257), .o (n10258) );
  buffer buf_n10259( .i (n10258), .o (n10259) );
  buffer buf_n10260( .i (n10259), .o (n10260) );
  buffer buf_n10261( .i (n10260), .o (n10261) );
  buffer buf_n10262( .i (n10261), .o (n10262) );
  buffer buf_n10263( .i (n10262), .o (n10263) );
  buffer buf_n10264( .i (n10263), .o (n10264) );
  buffer buf_n10265( .i (n10264), .o (n10265) );
  buffer buf_n10266( .i (n10265), .o (n10266) );
  buffer buf_n10267( .i (n10266), .o (n10267) );
  buffer buf_n10268( .i (n10267), .o (n10268) );
  buffer buf_n10269( .i (n10268), .o (n10269) );
  buffer buf_n10270( .i (n10269), .o (n10270) );
  buffer buf_n10271( .i (n10270), .o (n10271) );
  buffer buf_n10272( .i (n10271), .o (n10272) );
  buffer buf_n10273( .i (n10272), .o (n10273) );
  buffer buf_n10274( .i (n10273), .o (n10274) );
  buffer buf_n10275( .i (n10274), .o (n10275) );
  buffer buf_n10276( .i (n10275), .o (n10276) );
  buffer buf_n10277( .i (n10276), .o (n10277) );
  buffer buf_n10278( .i (n10277), .o (n10278) );
  buffer buf_n10279( .i (n10278), .o (n10279) );
  buffer buf_n10280( .i (n10279), .o (n10280) );
  buffer buf_n10281( .i (n10280), .o (n10281) );
  buffer buf_n10282( .i (n10281), .o (n10282) );
  buffer buf_n10283( .i (n10282), .o (n10283) );
  buffer buf_n10284( .i (n10283), .o (n10284) );
  buffer buf_n10285( .i (n10284), .o (n10285) );
  buffer buf_n10286( .i (n10285), .o (n10286) );
  buffer buf_n10287( .i (n10286), .o (n10287) );
  buffer buf_n10288( .i (n10287), .o (n10288) );
  buffer buf_n10289( .i (n10288), .o (n10289) );
  buffer buf_n10290( .i (n10289), .o (n10290) );
  buffer buf_n10291( .i (n10290), .o (n10291) );
  buffer buf_n10292( .i (n10291), .o (n10292) );
  buffer buf_n10293( .i (n10292), .o (n10293) );
  buffer buf_n10294( .i (n10293), .o (n10294) );
  buffer buf_n10295( .i (n10294), .o (n10295) );
  buffer buf_n785( .i (N241_I), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n1247( .i (n1246), .o (n1247) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n1488( .i (n1487), .o (n1488) );
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  buffer buf_n1534( .i (n1533), .o (n1534) );
  buffer buf_n1535( .i (n1534), .o (n1535) );
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n1556( .i (n1555), .o (n1556) );
  buffer buf_n1557( .i (n1556), .o (n1557) );
  buffer buf_n1558( .i (n1557), .o (n1558) );
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n1633( .i (n1632), .o (n1633) );
  buffer buf_n1634( .i (n1633), .o (n1634) );
  buffer buf_n1635( .i (n1634), .o (n1635) );
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n1637( .i (n1636), .o (n1637) );
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1658( .i (n1657), .o (n1658) );
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  buffer buf_n1813( .i (n1812), .o (n1813) );
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  buffer buf_n1821( .i (n1820), .o (n1821) );
  buffer buf_n1822( .i (n1821), .o (n1822) );
  buffer buf_n1823( .i (n1822), .o (n1823) );
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1825( .i (n1824), .o (n1825) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  buffer buf_n1846( .i (n1845), .o (n1846) );
  buffer buf_n1847( .i (n1846), .o (n1847) );
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  buffer buf_n1872( .i (n1871), .o (n1872) );
  buffer buf_n1873( .i (n1872), .o (n1873) );
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  buffer buf_n1879( .i (n1878), .o (n1879) );
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n1888( .i (n1887), .o (n1888) );
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1907( .i (n1906), .o (n1907) );
  buffer buf_n1908( .i (n1907), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n1915( .i (n1914), .o (n1915) );
  buffer buf_n1916( .i (n1915), .o (n1916) );
  buffer buf_n1917( .i (n1916), .o (n1917) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  buffer buf_n1930( .i (n1929), .o (n1930) );
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n1934( .i (n1933), .o (n1934) );
  buffer buf_n1935( .i (n1934), .o (n1935) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  buffer buf_n1954( .i (n1953), .o (n1954) );
  buffer buf_n1955( .i (n1954), .o (n1955) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  buffer buf_n1960( .i (n1959), .o (n1960) );
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n1967( .i (n1966), .o (n1967) );
  buffer buf_n1968( .i (n1967), .o (n1968) );
  buffer buf_n1969( .i (n1968), .o (n1969) );
  buffer buf_n1970( .i (n1969), .o (n1970) );
  buffer buf_n1971( .i (n1970), .o (n1971) );
  buffer buf_n1972( .i (n1971), .o (n1972) );
  buffer buf_n1973( .i (n1972), .o (n1973) );
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  buffer buf_n1983( .i (n1982), .o (n1983) );
  buffer buf_n1988( .i (n1987), .o (n1988) );
  buffer buf_n1989( .i (n1988), .o (n1989) );
  buffer buf_n1990( .i (n1989), .o (n1990) );
  buffer buf_n1991( .i (n1990), .o (n1991) );
  buffer buf_n1992( .i (n1991), .o (n1992) );
  buffer buf_n1993( .i (n1992), .o (n1993) );
  buffer buf_n1994( .i (n1993), .o (n1994) );
  buffer buf_n1995( .i (n1994), .o (n1995) );
  buffer buf_n1996( .i (n1995), .o (n1996) );
  buffer buf_n1997( .i (n1996), .o (n1997) );
  buffer buf_n1998( .i (n1997), .o (n1998) );
  buffer buf_n1999( .i (n1998), .o (n1999) );
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n2001( .i (n2000), .o (n2001) );
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n2003), .o (n2004) );
  buffer buf_n2005( .i (n2004), .o (n2005) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n2007( .i (n2006), .o (n2007) );
  buffer buf_n2008( .i (n2007), .o (n2008) );
  buffer buf_n2009( .i (n2008), .o (n2009) );
  buffer buf_n2010( .i (n2009), .o (n2010) );
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n2012( .i (n2011), .o (n2012) );
  buffer buf_n2013( .i (n2012), .o (n2013) );
  buffer buf_n2014( .i (n2013), .o (n2014) );
  buffer buf_n2015( .i (n2014), .o (n2015) );
  buffer buf_n2016( .i (n2015), .o (n2016) );
  buffer buf_n2017( .i (n2016), .o (n2017) );
  buffer buf_n2018( .i (n2017), .o (n2018) );
  buffer buf_n2019( .i (n2018), .o (n2019) );
  buffer buf_n2020( .i (n2019), .o (n2020) );
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2028( .i (n2027), .o (n2028) );
  buffer buf_n2029( .i (n2028), .o (n2029) );
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n2031( .i (n2030), .o (n2031) );
  buffer buf_n2032( .i (n2031), .o (n2032) );
  buffer buf_n2033( .i (n2032), .o (n2033) );
  buffer buf_n2034( .i (n2033), .o (n2034) );
  buffer buf_n2035( .i (n2034), .o (n2035) );
  buffer buf_n2036( .i (n2035), .o (n2036) );
  buffer buf_n2037( .i (n2036), .o (n2037) );
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2056( .i (n2055), .o (n2056) );
  buffer buf_n2057( .i (n2056), .o (n2057) );
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  buffer buf_n2064( .i (n2063), .o (n2064) );
  buffer buf_n2065( .i (n2064), .o (n2065) );
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n2073( .i (n2072), .o (n2073) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n2075( .i (n2074), .o (n2075) );
  buffer buf_n2076( .i (n2075), .o (n2076) );
  buffer buf_n2077( .i (n2076), .o (n2077) );
  buffer buf_n2078( .i (n2077), .o (n2078) );
  buffer buf_n2079( .i (n2078), .o (n2079) );
  buffer buf_n2080( .i (n2079), .o (n2080) );
  buffer buf_n2081( .i (n2080), .o (n2081) );
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2089( .i (n2088), .o (n2089) );
  buffer buf_n2090( .i (n2089), .o (n2090) );
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n2099( .i (n2098), .o (n2099) );
  buffer buf_n2100( .i (n2099), .o (n2100) );
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n2102( .i (n2101), .o (n2102) );
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n2111( .i (n2110), .o (n2111) );
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  buffer buf_n2129( .i (n2128), .o (n2129) );
  buffer buf_n2130( .i (n2129), .o (n2130) );
  buffer buf_n2131( .i (n2130), .o (n2131) );
  buffer buf_n2132( .i (n2131), .o (n2132) );
  buffer buf_n2133( .i (n2132), .o (n2133) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  buffer buf_n2137( .i (n2136), .o (n2137) );
  buffer buf_n2138( .i (n2137), .o (n2138) );
  buffer buf_n2139( .i (n2138), .o (n2139) );
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n2143( .i (n2142), .o (n2143) );
  buffer buf_n2144( .i (n2143), .o (n2144) );
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  buffer buf_n2152( .i (n2151), .o (n2152) );
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n2155( .i (n2154), .o (n2155) );
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n2158( .i (n2157), .o (n2158) );
  buffer buf_n2159( .i (n2158), .o (n2159) );
  buffer buf_n2160( .i (n2159), .o (n2160) );
  buffer buf_n2161( .i (n2160), .o (n2161) );
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n2163( .i (n2162), .o (n2163) );
  buffer buf_n2164( .i (n2163), .o (n2164) );
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n2166( .i (n2165), .o (n2166) );
  buffer buf_n2167( .i (n2166), .o (n2167) );
  buffer buf_n2168( .i (n2167), .o (n2168) );
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  buffer buf_n2171( .i (n2170), .o (n2171) );
  buffer buf_n2172( .i (n2171), .o (n2172) );
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n2175( .i (n2174), .o (n2175) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n2177), .o (n2178) );
  buffer buf_n2179( .i (n2178), .o (n2179) );
  buffer buf_n2180( .i (n2179), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  buffer buf_n2190( .i (n2189), .o (n2190) );
  buffer buf_n2191( .i (n2190), .o (n2191) );
  buffer buf_n2192( .i (n2191), .o (n2192) );
  buffer buf_n2193( .i (n2192), .o (n2193) );
  buffer buf_n2194( .i (n2193), .o (n2194) );
  buffer buf_n2195( .i (n2194), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  buffer buf_n2197( .i (n2196), .o (n2197) );
  buffer buf_n2198( .i (n2197), .o (n2198) );
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n2200( .i (n2199), .o (n2200) );
  buffer buf_n2201( .i (n2200), .o (n2201) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  buffer buf_n2203( .i (n2202), .o (n2203) );
  buffer buf_n2204( .i (n2203), .o (n2204) );
  buffer buf_n2205( .i (n2204), .o (n2205) );
  buffer buf_n2206( .i (n2205), .o (n2206) );
  buffer buf_n2207( .i (n2206), .o (n2207) );
  buffer buf_n2208( .i (n2207), .o (n2208) );
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n2211( .i (n2210), .o (n2211) );
  buffer buf_n2212( .i (n2211), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  buffer buf_n2214( .i (n2213), .o (n2214) );
  buffer buf_n2215( .i (n2214), .o (n2215) );
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n2221( .i (n2220), .o (n2221) );
  buffer buf_n2222( .i (n2221), .o (n2222) );
  buffer buf_n2223( .i (n2222), .o (n2223) );
  buffer buf_n2224( .i (n2223), .o (n2224) );
  buffer buf_n2225( .i (n2224), .o (n2225) );
  buffer buf_n2226( .i (n2225), .o (n2226) );
  buffer buf_n2227( .i (n2226), .o (n2227) );
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  buffer buf_n2231( .i (n2230), .o (n2231) );
  buffer buf_n2232( .i (n2231), .o (n2232) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  buffer buf_n2235( .i (n2234), .o (n2235) );
  buffer buf_n2236( .i (n2235), .o (n2236) );
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  buffer buf_n2265( .i (n2264), .o (n2265) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  buffer buf_n2269( .i (n2268), .o (n2269) );
  buffer buf_n2270( .i (n2269), .o (n2270) );
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2273( .i (n2272), .o (n2273) );
  buffer buf_n2274( .i (n2273), .o (n2274) );
  buffer buf_n2275( .i (n2274), .o (n2275) );
  buffer buf_n2276( .i (n2275), .o (n2276) );
  buffer buf_n2277( .i (n2276), .o (n2277) );
  buffer buf_n2278( .i (n2277), .o (n2278) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  buffer buf_n2280( .i (n2279), .o (n2280) );
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n2289( .i (n2288), .o (n2289) );
  buffer buf_n2290( .i (n2289), .o (n2290) );
  buffer buf_n2291( .i (n2290), .o (n2291) );
  buffer buf_n2292( .i (n2291), .o (n2292) );
  buffer buf_n2293( .i (n2292), .o (n2293) );
  buffer buf_n2294( .i (n2293), .o (n2294) );
  buffer buf_n2295( .i (n2294), .o (n2295) );
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n2297( .i (n2296), .o (n2297) );
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  buffer buf_n2307( .i (n2306), .o (n2307) );
  buffer buf_n2308( .i (n2307), .o (n2308) );
  buffer buf_n2309( .i (n2308), .o (n2309) );
  buffer buf_n2310( .i (n2309), .o (n2310) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  buffer buf_n2326( .i (n2325), .o (n2326) );
  buffer buf_n2327( .i (n2326), .o (n2327) );
  buffer buf_n2328( .i (n2327), .o (n2328) );
  buffer buf_n2329( .i (n2328), .o (n2329) );
  buffer buf_n2330( .i (n2329), .o (n2330) );
  buffer buf_n2331( .i (n2330), .o (n2331) );
  buffer buf_n2332( .i (n2331), .o (n2332) );
  buffer buf_n2333( .i (n2332), .o (n2333) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n2335( .i (n2334), .o (n2335) );
  buffer buf_n2336( .i (n2335), .o (n2336) );
  buffer buf_n2337( .i (n2336), .o (n2337) );
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  buffer buf_n2340( .i (n2339), .o (n2340) );
  buffer buf_n2341( .i (n2340), .o (n2341) );
  buffer buf_n2342( .i (n2341), .o (n2342) );
  buffer buf_n2343( .i (n2342), .o (n2343) );
  buffer buf_n2344( .i (n2343), .o (n2344) );
  buffer buf_n2345( .i (n2344), .o (n2345) );
  buffer buf_n2346( .i (n2345), .o (n2346) );
  buffer buf_n2347( .i (n2346), .o (n2347) );
  buffer buf_n2348( .i (n2347), .o (n2348) );
  buffer buf_n2349( .i (n2348), .o (n2349) );
  buffer buf_n2350( .i (n2349), .o (n2350) );
  buffer buf_n2351( .i (n2350), .o (n2351) );
  buffer buf_n2352( .i (n2351), .o (n2352) );
  buffer buf_n2353( .i (n2352), .o (n2353) );
  buffer buf_n2354( .i (n2353), .o (n2354) );
  buffer buf_n2355( .i (n2354), .o (n2355) );
  buffer buf_n2356( .i (n2355), .o (n2356) );
  buffer buf_n2357( .i (n2356), .o (n2357) );
  buffer buf_n2358( .i (n2357), .o (n2358) );
  buffer buf_n2359( .i (n2358), .o (n2359) );
  buffer buf_n2360( .i (n2359), .o (n2360) );
  buffer buf_n2361( .i (n2360), .o (n2361) );
  buffer buf_n2362( .i (n2361), .o (n2362) );
  buffer buf_n2363( .i (n2362), .o (n2363) );
  buffer buf_n2364( .i (n2363), .o (n2364) );
  buffer buf_n2365( .i (n2364), .o (n2365) );
  buffer buf_n2366( .i (n2365), .o (n2366) );
  buffer buf_n2367( .i (n2366), .o (n2367) );
  buffer buf_n2368( .i (n2367), .o (n2368) );
  buffer buf_n2369( .i (n2368), .o (n2369) );
  buffer buf_n2370( .i (n2369), .o (n2370) );
  buffer buf_n2371( .i (n2370), .o (n2371) );
  buffer buf_n2372( .i (n2371), .o (n2372) );
  buffer buf_n2373( .i (n2372), .o (n2373) );
  buffer buf_n2374( .i (n2373), .o (n2374) );
  buffer buf_n2375( .i (n2374), .o (n2375) );
  buffer buf_n2376( .i (n2375), .o (n2376) );
  buffer buf_n2377( .i (n2376), .o (n2377) );
  buffer buf_n2378( .i (n2377), .o (n2378) );
  buffer buf_n2379( .i (n2378), .o (n2379) );
  buffer buf_n2380( .i (n2379), .o (n2380) );
  buffer buf_n2381( .i (n2380), .o (n2381) );
  buffer buf_n2382( .i (n2381), .o (n2382) );
  buffer buf_n2383( .i (n2382), .o (n2383) );
  buffer buf_n2392( .i (n2391), .o (n2392) );
  buffer buf_n2393( .i (n2392), .o (n2393) );
  buffer buf_n2394( .i (n2393), .o (n2394) );
  buffer buf_n2395( .i (n2394), .o (n2395) );
  buffer buf_n2396( .i (n2395), .o (n2396) );
  buffer buf_n2397( .i (n2396), .o (n2397) );
  buffer buf_n2398( .i (n2397), .o (n2398) );
  buffer buf_n2399( .i (n2398), .o (n2399) );
  buffer buf_n2400( .i (n2399), .o (n2400) );
  buffer buf_n2401( .i (n2400), .o (n2401) );
  buffer buf_n2402( .i (n2401), .o (n2402) );
  buffer buf_n2403( .i (n2402), .o (n2403) );
  buffer buf_n2404( .i (n2403), .o (n2404) );
  buffer buf_n2405( .i (n2404), .o (n2405) );
  buffer buf_n2406( .i (n2405), .o (n2406) );
  buffer buf_n2407( .i (n2406), .o (n2407) );
  buffer buf_n2408( .i (n2407), .o (n2408) );
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  buffer buf_n2411( .i (n2410), .o (n2411) );
  buffer buf_n2412( .i (n2411), .o (n2412) );
  buffer buf_n2413( .i (n2412), .o (n2413) );
  buffer buf_n2414( .i (n2413), .o (n2414) );
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n2416( .i (n2415), .o (n2416) );
  buffer buf_n2417( .i (n2416), .o (n2417) );
  buffer buf_n2418( .i (n2417), .o (n2418) );
  buffer buf_n2419( .i (n2418), .o (n2419) );
  buffer buf_n2420( .i (n2419), .o (n2420) );
  buffer buf_n2421( .i (n2420), .o (n2421) );
  buffer buf_n2422( .i (n2421), .o (n2422) );
  buffer buf_n2423( .i (n2422), .o (n2423) );
  buffer buf_n2424( .i (n2423), .o (n2424) );
  buffer buf_n2425( .i (n2424), .o (n2425) );
  buffer buf_n2426( .i (n2425), .o (n2426) );
  buffer buf_n2427( .i (n2426), .o (n2427) );
  buffer buf_n2428( .i (n2427), .o (n2428) );
  buffer buf_n2429( .i (n2428), .o (n2429) );
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  buffer buf_n2432( .i (n2431), .o (n2432) );
  buffer buf_n2433( .i (n2432), .o (n2433) );
  buffer buf_n2434( .i (n2433), .o (n2434) );
  buffer buf_n2435( .i (n2434), .o (n2435) );
  buffer buf_n2436( .i (n2435), .o (n2436) );
  buffer buf_n2437( .i (n2436), .o (n2437) );
  buffer buf_n2438( .i (n2437), .o (n2438) );
  buffer buf_n2439( .i (n2438), .o (n2439) );
  buffer buf_n2440( .i (n2439), .o (n2440) );
  buffer buf_n2441( .i (n2440), .o (n2441) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  buffer buf_n2443( .i (n2442), .o (n2443) );
  buffer buf_n2444( .i (n2443), .o (n2444) );
  buffer buf_n2445( .i (n2444), .o (n2445) );
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n2448( .i (n2447), .o (n2448) );
  buffer buf_n2449( .i (n2448), .o (n2449) );
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n2460( .i (n2459), .o (n2460) );
  buffer buf_n2461( .i (n2460), .o (n2461) );
  buffer buf_n2462( .i (n2461), .o (n2462) );
  buffer buf_n2463( .i (n2462), .o (n2463) );
  buffer buf_n2464( .i (n2463), .o (n2464) );
  buffer buf_n2465( .i (n2464), .o (n2465) );
  buffer buf_n2466( .i (n2465), .o (n2466) );
  buffer buf_n2467( .i (n2466), .o (n2467) );
  buffer buf_n2468( .i (n2467), .o (n2468) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  buffer buf_n2470( .i (n2469), .o (n2470) );
  buffer buf_n2471( .i (n2470), .o (n2471) );
  buffer buf_n2472( .i (n2471), .o (n2472) );
  buffer buf_n2473( .i (n2472), .o (n2473) );
  buffer buf_n2474( .i (n2473), .o (n2474) );
  buffer buf_n2475( .i (n2474), .o (n2475) );
  buffer buf_n2476( .i (n2475), .o (n2476) );
  buffer buf_n2477( .i (n2476), .o (n2477) );
  buffer buf_n2478( .i (n2477), .o (n2478) );
  buffer buf_n2479( .i (n2478), .o (n2479) );
  buffer buf_n2480( .i (n2479), .o (n2480) );
  buffer buf_n2481( .i (n2480), .o (n2481) );
  buffer buf_n2482( .i (n2481), .o (n2482) );
  buffer buf_n2483( .i (n2482), .o (n2483) );
  buffer buf_n2484( .i (n2483), .o (n2484) );
  buffer buf_n2485( .i (n2484), .o (n2485) );
  buffer buf_n2486( .i (n2485), .o (n2486) );
  buffer buf_n2487( .i (n2486), .o (n2487) );
  buffer buf_n2488( .i (n2487), .o (n2488) );
  buffer buf_n2489( .i (n2488), .o (n2489) );
  buffer buf_n2490( .i (n2489), .o (n2490) );
  buffer buf_n2491( .i (n2490), .o (n2491) );
  buffer buf_n2492( .i (n2491), .o (n2492) );
  buffer buf_n2493( .i (n2492), .o (n2493) );
  buffer buf_n2494( .i (n2493), .o (n2494) );
  buffer buf_n2495( .i (n2494), .o (n2495) );
  buffer buf_n2496( .i (n2495), .o (n2496) );
  buffer buf_n2497( .i (n2496), .o (n2497) );
  buffer buf_n2498( .i (n2497), .o (n2498) );
  buffer buf_n2499( .i (n2498), .o (n2499) );
  buffer buf_n2500( .i (n2499), .o (n2500) );
  buffer buf_n2501( .i (n2500), .o (n2501) );
  buffer buf_n2502( .i (n2501), .o (n2502) );
  buffer buf_n2503( .i (n2502), .o (n2503) );
  buffer buf_n2504( .i (n2503), .o (n2504) );
  buffer buf_n2505( .i (n2504), .o (n2505) );
  buffer buf_n2506( .i (n2505), .o (n2506) );
  buffer buf_n2507( .i (n2506), .o (n2507) );
  buffer buf_n2508( .i (n2507), .o (n2508) );
  buffer buf_n2509( .i (n2508), .o (n2509) );
  buffer buf_n2510( .i (n2509), .o (n2510) );
  buffer buf_n2511( .i (n2510), .o (n2511) );
  buffer buf_n2512( .i (n2511), .o (n2512) );
  buffer buf_n2513( .i (n2512), .o (n2513) );
  buffer buf_n2514( .i (n2513), .o (n2514) );
  buffer buf_n2515( .i (n2514), .o (n2515) );
  buffer buf_n2524( .i (n2523), .o (n2524) );
  buffer buf_n2525( .i (n2524), .o (n2525) );
  buffer buf_n2526( .i (n2525), .o (n2526) );
  buffer buf_n2527( .i (n2526), .o (n2527) );
  buffer buf_n2528( .i (n2527), .o (n2528) );
  buffer buf_n2529( .i (n2528), .o (n2529) );
  buffer buf_n2530( .i (n2529), .o (n2530) );
  buffer buf_n2531( .i (n2530), .o (n2531) );
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n2532), .o (n2533) );
  buffer buf_n2534( .i (n2533), .o (n2534) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  buffer buf_n2536( .i (n2535), .o (n2536) );
  buffer buf_n2537( .i (n2536), .o (n2537) );
  buffer buf_n2538( .i (n2537), .o (n2538) );
  buffer buf_n2539( .i (n2538), .o (n2539) );
  buffer buf_n2540( .i (n2539), .o (n2540) );
  buffer buf_n2541( .i (n2540), .o (n2541) );
  buffer buf_n2542( .i (n2541), .o (n2542) );
  buffer buf_n2543( .i (n2542), .o (n2543) );
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  buffer buf_n2551( .i (n2550), .o (n2551) );
  buffer buf_n2552( .i (n2551), .o (n2552) );
  buffer buf_n2553( .i (n2552), .o (n2553) );
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2555( .i (n2554), .o (n2555) );
  buffer buf_n2556( .i (n2555), .o (n2556) );
  buffer buf_n2557( .i (n2556), .o (n2557) );
  buffer buf_n2558( .i (n2557), .o (n2558) );
  buffer buf_n2559( .i (n2558), .o (n2559) );
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  buffer buf_n2563( .i (n2562), .o (n2563) );
  buffer buf_n2564( .i (n2563), .o (n2564) );
  buffer buf_n2565( .i (n2564), .o (n2565) );
  buffer buf_n2566( .i (n2565), .o (n2566) );
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n2568( .i (n2567), .o (n2568) );
  buffer buf_n2569( .i (n2568), .o (n2569) );
  buffer buf_n2570( .i (n2569), .o (n2570) );
  buffer buf_n2571( .i (n2570), .o (n2571) );
  buffer buf_n2572( .i (n2571), .o (n2572) );
  buffer buf_n2573( .i (n2572), .o (n2573) );
  buffer buf_n2574( .i (n2573), .o (n2574) );
  buffer buf_n2575( .i (n2574), .o (n2575) );
  buffer buf_n2576( .i (n2575), .o (n2576) );
  buffer buf_n2577( .i (n2576), .o (n2577) );
  buffer buf_n2578( .i (n2577), .o (n2578) );
  buffer buf_n2579( .i (n2578), .o (n2579) );
  buffer buf_n2580( .i (n2579), .o (n2580) );
  buffer buf_n2581( .i (n2580), .o (n2581) );
  buffer buf_n2590( .i (n2589), .o (n2590) );
  buffer buf_n2591( .i (n2590), .o (n2591) );
  buffer buf_n2592( .i (n2591), .o (n2592) );
  buffer buf_n2593( .i (n2592), .o (n2593) );
  buffer buf_n2594( .i (n2593), .o (n2594) );
  buffer buf_n2595( .i (n2594), .o (n2595) );
  buffer buf_n2596( .i (n2595), .o (n2596) );
  buffer buf_n2597( .i (n2596), .o (n2597) );
  buffer buf_n2598( .i (n2597), .o (n2598) );
  buffer buf_n2599( .i (n2598), .o (n2599) );
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  buffer buf_n2602( .i (n2601), .o (n2602) );
  buffer buf_n2603( .i (n2602), .o (n2603) );
  buffer buf_n2604( .i (n2603), .o (n2604) );
  buffer buf_n2605( .i (n2604), .o (n2605) );
  buffer buf_n2606( .i (n2605), .o (n2606) );
  buffer buf_n2607( .i (n2606), .o (n2607) );
  buffer buf_n2608( .i (n2607), .o (n2608) );
  buffer buf_n2609( .i (n2608), .o (n2609) );
  buffer buf_n2610( .i (n2609), .o (n2610) );
  buffer buf_n2611( .i (n2610), .o (n2611) );
  buffer buf_n2612( .i (n2611), .o (n2612) );
  buffer buf_n2613( .i (n2612), .o (n2613) );
  buffer buf_n2614( .i (n2613), .o (n2614) );
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  buffer buf_n2617( .i (n2616), .o (n2617) );
  buffer buf_n2618( .i (n2617), .o (n2618) );
  buffer buf_n2619( .i (n2618), .o (n2619) );
  buffer buf_n2620( .i (n2619), .o (n2620) );
  buffer buf_n2621( .i (n2620), .o (n2621) );
  buffer buf_n2622( .i (n2621), .o (n2622) );
  buffer buf_n2623( .i (n2622), .o (n2623) );
  buffer buf_n2624( .i (n2623), .o (n2624) );
  buffer buf_n2625( .i (n2624), .o (n2625) );
  buffer buf_n2626( .i (n2625), .o (n2626) );
  buffer buf_n2627( .i (n2626), .o (n2627) );
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  buffer buf_n2631( .i (n2630), .o (n2631) );
  buffer buf_n2632( .i (n2631), .o (n2632) );
  buffer buf_n2633( .i (n2632), .o (n2633) );
  buffer buf_n2634( .i (n2633), .o (n2634) );
  buffer buf_n2635( .i (n2634), .o (n2635) );
  buffer buf_n2636( .i (n2635), .o (n2636) );
  buffer buf_n2637( .i (n2636), .o (n2637) );
  buffer buf_n2638( .i (n2637), .o (n2638) );
  buffer buf_n2639( .i (n2638), .o (n2639) );
  buffer buf_n2640( .i (n2639), .o (n2640) );
  buffer buf_n2641( .i (n2640), .o (n2641) );
  buffer buf_n2642( .i (n2641), .o (n2642) );
  buffer buf_n2643( .i (n2642), .o (n2643) );
  buffer buf_n2644( .i (n2643), .o (n2644) );
  buffer buf_n2645( .i (n2644), .o (n2645) );
  buffer buf_n2646( .i (n2645), .o (n2646) );
  buffer buf_n2647( .i (n2646), .o (n2647) );
  buffer buf_n2652( .i (n2651), .o (n2652) );
  buffer buf_n2653( .i (n2652), .o (n2653) );
  buffer buf_n2654( .i (n2653), .o (n2654) );
  buffer buf_n2655( .i (n2654), .o (n2655) );
  buffer buf_n2656( .i (n2655), .o (n2656) );
  buffer buf_n2657( .i (n2656), .o (n2657) );
  buffer buf_n2658( .i (n2657), .o (n2658) );
  buffer buf_n2659( .i (n2658), .o (n2659) );
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2660), .o (n2661) );
  buffer buf_n2662( .i (n2661), .o (n2662) );
  buffer buf_n2663( .i (n2662), .o (n2663) );
  buffer buf_n2664( .i (n2663), .o (n2664) );
  buffer buf_n2665( .i (n2664), .o (n2665) );
  buffer buf_n2666( .i (n2665), .o (n2666) );
  buffer buf_n2667( .i (n2666), .o (n2667) );
  buffer buf_n2668( .i (n2667), .o (n2668) );
  buffer buf_n2669( .i (n2668), .o (n2669) );
  buffer buf_n2670( .i (n2669), .o (n2670) );
  buffer buf_n2671( .i (n2670), .o (n2671) );
  buffer buf_n2672( .i (n2671), .o (n2672) );
  buffer buf_n2673( .i (n2672), .o (n2673) );
  buffer buf_n2674( .i (n2673), .o (n2674) );
  buffer buf_n2675( .i (n2674), .o (n2675) );
  buffer buf_n2676( .i (n2675), .o (n2676) );
  buffer buf_n2677( .i (n2676), .o (n2677) );
  buffer buf_n2678( .i (n2677), .o (n2678) );
  buffer buf_n2679( .i (n2678), .o (n2679) );
  buffer buf_n2680( .i (n2679), .o (n2680) );
  buffer buf_n2681( .i (n2680), .o (n2681) );
  buffer buf_n2682( .i (n2681), .o (n2682) );
  buffer buf_n2683( .i (n2682), .o (n2683) );
  buffer buf_n2684( .i (n2683), .o (n2684) );
  buffer buf_n2685( .i (n2684), .o (n2685) );
  buffer buf_n2686( .i (n2685), .o (n2686) );
  buffer buf_n2687( .i (n2686), .o (n2687) );
  buffer buf_n2688( .i (n2687), .o (n2688) );
  buffer buf_n2689( .i (n2688), .o (n2689) );
  buffer buf_n2690( .i (n2689), .o (n2690) );
  buffer buf_n2691( .i (n2690), .o (n2691) );
  buffer buf_n2692( .i (n2691), .o (n2692) );
  buffer buf_n2693( .i (n2692), .o (n2693) );
  buffer buf_n2694( .i (n2693), .o (n2694) );
  buffer buf_n2695( .i (n2694), .o (n2695) );
  buffer buf_n2696( .i (n2695), .o (n2696) );
  buffer buf_n2697( .i (n2696), .o (n2697) );
  buffer buf_n2698( .i (n2697), .o (n2698) );
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n2700( .i (n2699), .o (n2700) );
  buffer buf_n2701( .i (n2700), .o (n2701) );
  buffer buf_n2702( .i (n2701), .o (n2702) );
  buffer buf_n2703( .i (n2702), .o (n2703) );
  buffer buf_n2704( .i (n2703), .o (n2704) );
  buffer buf_n2705( .i (n2704), .o (n2705) );
  buffer buf_n2706( .i (n2705), .o (n2706) );
  buffer buf_n2707( .i (n2706), .o (n2707) );
  buffer buf_n2708( .i (n2707), .o (n2708) );
  buffer buf_n2709( .i (n2708), .o (n2709) );
  buffer buf_n2710( .i (n2709), .o (n2710) );
  buffer buf_n2711( .i (n2710), .o (n2711) );
  buffer buf_n2712( .i (n2711), .o (n2712) );
  buffer buf_n2713( .i (n2712), .o (n2713) );
  buffer buf_n2788( .i (n2787), .o (n2788) );
  buffer buf_n2789( .i (n2788), .o (n2789) );
  buffer buf_n2790( .i (n2789), .o (n2790) );
  buffer buf_n2791( .i (n2790), .o (n2791) );
  buffer buf_n2792( .i (n2791), .o (n2792) );
  buffer buf_n2793( .i (n2792), .o (n2793) );
  buffer buf_n2794( .i (n2793), .o (n2794) );
  buffer buf_n2795( .i (n2794), .o (n2795) );
  buffer buf_n2796( .i (n2795), .o (n2796) );
  buffer buf_n2797( .i (n2796), .o (n2797) );
  buffer buf_n2798( .i (n2797), .o (n2798) );
  buffer buf_n2799( .i (n2798), .o (n2799) );
  buffer buf_n2800( .i (n2799), .o (n2800) );
  buffer buf_n2801( .i (n2800), .o (n2801) );
  buffer buf_n2802( .i (n2801), .o (n2802) );
  buffer buf_n2803( .i (n2802), .o (n2803) );
  buffer buf_n2804( .i (n2803), .o (n2804) );
  buffer buf_n2805( .i (n2804), .o (n2805) );
  buffer buf_n2806( .i (n2805), .o (n2806) );
  buffer buf_n2807( .i (n2806), .o (n2807) );
  buffer buf_n2808( .i (n2807), .o (n2808) );
  buffer buf_n2809( .i (n2808), .o (n2809) );
  buffer buf_n2810( .i (n2809), .o (n2810) );
  buffer buf_n2811( .i (n2810), .o (n2811) );
  buffer buf_n2812( .i (n2811), .o (n2812) );
  buffer buf_n2813( .i (n2812), .o (n2813) );
  buffer buf_n2814( .i (n2813), .o (n2814) );
  buffer buf_n2815( .i (n2814), .o (n2815) );
  buffer buf_n2816( .i (n2815), .o (n2816) );
  buffer buf_n2817( .i (n2816), .o (n2817) );
  buffer buf_n2818( .i (n2817), .o (n2818) );
  buffer buf_n2819( .i (n2818), .o (n2819) );
  buffer buf_n2820( .i (n2819), .o (n2820) );
  buffer buf_n2821( .i (n2820), .o (n2821) );
  buffer buf_n2822( .i (n2821), .o (n2822) );
  buffer buf_n2823( .i (n2822), .o (n2823) );
  buffer buf_n2824( .i (n2823), .o (n2824) );
  buffer buf_n2825( .i (n2824), .o (n2825) );
  buffer buf_n2826( .i (n2825), .o (n2826) );
  buffer buf_n2827( .i (n2826), .o (n2827) );
  buffer buf_n2828( .i (n2827), .o (n2828) );
  buffer buf_n2829( .i (n2828), .o (n2829) );
  buffer buf_n2830( .i (n2829), .o (n2830) );
  buffer buf_n2831( .i (n2830), .o (n2831) );
  buffer buf_n2832( .i (n2831), .o (n2832) );
  buffer buf_n2833( .i (n2832), .o (n2833) );
  buffer buf_n2834( .i (n2833), .o (n2834) );
  buffer buf_n2835( .i (n2834), .o (n2835) );
  buffer buf_n2836( .i (n2835), .o (n2836) );
  buffer buf_n2837( .i (n2836), .o (n2837) );
  buffer buf_n2838( .i (n2837), .o (n2838) );
  buffer buf_n2839( .i (n2838), .o (n2839) );
  buffer buf_n2840( .i (n2839), .o (n2840) );
  buffer buf_n2841( .i (n2840), .o (n2841) );
  buffer buf_n2842( .i (n2841), .o (n2842) );
  buffer buf_n2843( .i (n2842), .o (n2843) );
  buffer buf_n2844( .i (n2843), .o (n2844) );
  buffer buf_n2845( .i (n2844), .o (n2845) );
  buffer buf_n2854( .i (n2853), .o (n2854) );
  buffer buf_n2855( .i (n2854), .o (n2855) );
  buffer buf_n2856( .i (n2855), .o (n2856) );
  buffer buf_n2857( .i (n2856), .o (n2857) );
  buffer buf_n2858( .i (n2857), .o (n2858) );
  buffer buf_n2859( .i (n2858), .o (n2859) );
  buffer buf_n2860( .i (n2859), .o (n2860) );
  buffer buf_n2861( .i (n2860), .o (n2861) );
  buffer buf_n2862( .i (n2861), .o (n2862) );
  buffer buf_n2863( .i (n2862), .o (n2863) );
  buffer buf_n2864( .i (n2863), .o (n2864) );
  buffer buf_n2865( .i (n2864), .o (n2865) );
  buffer buf_n2866( .i (n2865), .o (n2866) );
  buffer buf_n2867( .i (n2866), .o (n2867) );
  buffer buf_n2868( .i (n2867), .o (n2868) );
  buffer buf_n2869( .i (n2868), .o (n2869) );
  buffer buf_n2870( .i (n2869), .o (n2870) );
  buffer buf_n2871( .i (n2870), .o (n2871) );
  buffer buf_n2872( .i (n2871), .o (n2872) );
  buffer buf_n2873( .i (n2872), .o (n2873) );
  buffer buf_n2874( .i (n2873), .o (n2874) );
  buffer buf_n2875( .i (n2874), .o (n2875) );
  buffer buf_n2876( .i (n2875), .o (n2876) );
  buffer buf_n2877( .i (n2876), .o (n2877) );
  buffer buf_n2878( .i (n2877), .o (n2878) );
  buffer buf_n2879( .i (n2878), .o (n2879) );
  buffer buf_n2880( .i (n2879), .o (n2880) );
  buffer buf_n2881( .i (n2880), .o (n2881) );
  buffer buf_n2882( .i (n2881), .o (n2882) );
  buffer buf_n2883( .i (n2882), .o (n2883) );
  buffer buf_n2884( .i (n2883), .o (n2884) );
  buffer buf_n2885( .i (n2884), .o (n2885) );
  buffer buf_n2886( .i (n2885), .o (n2886) );
  buffer buf_n2887( .i (n2886), .o (n2887) );
  buffer buf_n2888( .i (n2887), .o (n2888) );
  buffer buf_n2889( .i (n2888), .o (n2889) );
  buffer buf_n2890( .i (n2889), .o (n2890) );
  buffer buf_n2891( .i (n2890), .o (n2891) );
  buffer buf_n2892( .i (n2891), .o (n2892) );
  buffer buf_n2893( .i (n2892), .o (n2893) );
  buffer buf_n2894( .i (n2893), .o (n2894) );
  buffer buf_n2895( .i (n2894), .o (n2895) );
  buffer buf_n2896( .i (n2895), .o (n2896) );
  buffer buf_n2897( .i (n2896), .o (n2897) );
  buffer buf_n2898( .i (n2897), .o (n2898) );
  buffer buf_n2899( .i (n2898), .o (n2899) );
  buffer buf_n2900( .i (n2899), .o (n2900) );
  buffer buf_n2901( .i (n2900), .o (n2901) );
  buffer buf_n2902( .i (n2901), .o (n2902) );
  buffer buf_n2903( .i (n2902), .o (n2903) );
  buffer buf_n2904( .i (n2903), .o (n2904) );
  buffer buf_n2905( .i (n2904), .o (n2905) );
  buffer buf_n2906( .i (n2905), .o (n2906) );
  buffer buf_n2907( .i (n2906), .o (n2907) );
  buffer buf_n2908( .i (n2907), .o (n2908) );
  buffer buf_n2909( .i (n2908), .o (n2909) );
  buffer buf_n2910( .i (n2909), .o (n2910) );
  buffer buf_n2911( .i (n2910), .o (n2911) );
  buffer buf_n2920( .i (n2919), .o (n2920) );
  buffer buf_n2921( .i (n2920), .o (n2921) );
  buffer buf_n2922( .i (n2921), .o (n2922) );
  buffer buf_n2923( .i (n2922), .o (n2923) );
  buffer buf_n2924( .i (n2923), .o (n2924) );
  buffer buf_n2925( .i (n2924), .o (n2925) );
  buffer buf_n2926( .i (n2925), .o (n2926) );
  buffer buf_n2927( .i (n2926), .o (n2927) );
  buffer buf_n2928( .i (n2927), .o (n2928) );
  buffer buf_n2929( .i (n2928), .o (n2929) );
  buffer buf_n2930( .i (n2929), .o (n2930) );
  buffer buf_n2931( .i (n2930), .o (n2931) );
  buffer buf_n2932( .i (n2931), .o (n2932) );
  buffer buf_n2933( .i (n2932), .o (n2933) );
  buffer buf_n2934( .i (n2933), .o (n2934) );
  buffer buf_n2935( .i (n2934), .o (n2935) );
  buffer buf_n2936( .i (n2935), .o (n2936) );
  buffer buf_n2937( .i (n2936), .o (n2937) );
  buffer buf_n2938( .i (n2937), .o (n2938) );
  buffer buf_n2939( .i (n2938), .o (n2939) );
  buffer buf_n2940( .i (n2939), .o (n2940) );
  buffer buf_n2941( .i (n2940), .o (n2941) );
  buffer buf_n2942( .i (n2941), .o (n2942) );
  buffer buf_n2943( .i (n2942), .o (n2943) );
  buffer buf_n2944( .i (n2943), .o (n2944) );
  buffer buf_n2945( .i (n2944), .o (n2945) );
  buffer buf_n2946( .i (n2945), .o (n2946) );
  buffer buf_n2947( .i (n2946), .o (n2947) );
  buffer buf_n2948( .i (n2947), .o (n2948) );
  buffer buf_n2949( .i (n2948), .o (n2949) );
  buffer buf_n2950( .i (n2949), .o (n2950) );
  buffer buf_n2951( .i (n2950), .o (n2951) );
  buffer buf_n2952( .i (n2951), .o (n2952) );
  buffer buf_n2953( .i (n2952), .o (n2953) );
  buffer buf_n2954( .i (n2953), .o (n2954) );
  buffer buf_n2955( .i (n2954), .o (n2955) );
  buffer buf_n2956( .i (n2955), .o (n2956) );
  buffer buf_n2957( .i (n2956), .o (n2957) );
  buffer buf_n2958( .i (n2957), .o (n2958) );
  buffer buf_n2959( .i (n2958), .o (n2959) );
  buffer buf_n2960( .i (n2959), .o (n2960) );
  buffer buf_n2961( .i (n2960), .o (n2961) );
  buffer buf_n2962( .i (n2961), .o (n2962) );
  buffer buf_n2963( .i (n2962), .o (n2963) );
  buffer buf_n2964( .i (n2963), .o (n2964) );
  buffer buf_n2965( .i (n2964), .o (n2965) );
  buffer buf_n2966( .i (n2965), .o (n2966) );
  buffer buf_n2967( .i (n2966), .o (n2967) );
  buffer buf_n2968( .i (n2967), .o (n2968) );
  buffer buf_n2969( .i (n2968), .o (n2969) );
  buffer buf_n2970( .i (n2969), .o (n2970) );
  buffer buf_n2971( .i (n2970), .o (n2971) );
  buffer buf_n2972( .i (n2971), .o (n2972) );
  buffer buf_n2973( .i (n2972), .o (n2973) );
  buffer buf_n2974( .i (n2973), .o (n2974) );
  buffer buf_n2975( .i (n2974), .o (n2975) );
  buffer buf_n2976( .i (n2975), .o (n2976) );
  buffer buf_n2977( .i (n2976), .o (n2977) );
  buffer buf_n2990( .i (n2989), .o (n2990) );
  buffer buf_n2991( .i (n2990), .o (n2991) );
  buffer buf_n2992( .i (n2991), .o (n2992) );
  buffer buf_n2993( .i (n2992), .o (n2993) );
  buffer buf_n2994( .i (n2993), .o (n2994) );
  buffer buf_n2995( .i (n2994), .o (n2995) );
  buffer buf_n2996( .i (n2995), .o (n2996) );
  buffer buf_n2997( .i (n2996), .o (n2997) );
  buffer buf_n2998( .i (n2997), .o (n2998) );
  buffer buf_n2999( .i (n2998), .o (n2999) );
  buffer buf_n3000( .i (n2999), .o (n3000) );
  buffer buf_n3001( .i (n3000), .o (n3001) );
  buffer buf_n3002( .i (n3001), .o (n3002) );
  buffer buf_n3003( .i (n3002), .o (n3003) );
  buffer buf_n3004( .i (n3003), .o (n3004) );
  buffer buf_n3005( .i (n3004), .o (n3005) );
  buffer buf_n3006( .i (n3005), .o (n3006) );
  buffer buf_n3007( .i (n3006), .o (n3007) );
  buffer buf_n3008( .i (n3007), .o (n3008) );
  buffer buf_n3009( .i (n3008), .o (n3009) );
  buffer buf_n3010( .i (n3009), .o (n3010) );
  buffer buf_n3011( .i (n3010), .o (n3011) );
  buffer buf_n3012( .i (n3011), .o (n3012) );
  buffer buf_n3013( .i (n3012), .o (n3013) );
  buffer buf_n3014( .i (n3013), .o (n3014) );
  buffer buf_n3015( .i (n3014), .o (n3015) );
  buffer buf_n3016( .i (n3015), .o (n3016) );
  buffer buf_n3017( .i (n3016), .o (n3017) );
  buffer buf_n3018( .i (n3017), .o (n3018) );
  buffer buf_n3019( .i (n3018), .o (n3019) );
  buffer buf_n3020( .i (n3019), .o (n3020) );
  buffer buf_n3021( .i (n3020), .o (n3021) );
  buffer buf_n3022( .i (n3021), .o (n3022) );
  buffer buf_n3023( .i (n3022), .o (n3023) );
  buffer buf_n3024( .i (n3023), .o (n3024) );
  buffer buf_n3025( .i (n3024), .o (n3025) );
  buffer buf_n3026( .i (n3025), .o (n3026) );
  buffer buf_n3027( .i (n3026), .o (n3027) );
  buffer buf_n3028( .i (n3027), .o (n3028) );
  buffer buf_n3029( .i (n3028), .o (n3029) );
  buffer buf_n3030( .i (n3029), .o (n3030) );
  buffer buf_n3031( .i (n3030), .o (n3031) );
  buffer buf_n3032( .i (n3031), .o (n3032) );
  buffer buf_n3033( .i (n3032), .o (n3033) );
  buffer buf_n3034( .i (n3033), .o (n3034) );
  buffer buf_n3035( .i (n3034), .o (n3035) );
  buffer buf_n3036( .i (n3035), .o (n3036) );
  buffer buf_n3037( .i (n3036), .o (n3037) );
  buffer buf_n3038( .i (n3037), .o (n3038) );
  buffer buf_n3039( .i (n3038), .o (n3039) );
  buffer buf_n3040( .i (n3039), .o (n3040) );
  buffer buf_n3041( .i (n3040), .o (n3041) );
  buffer buf_n3042( .i (n3041), .o (n3042) );
  buffer buf_n3043( .i (n3042), .o (n3043) );
  buffer buf_n3044( .i (n3043), .o (n3044) );
  buffer buf_n3045( .i (n3044), .o (n3045) );
  buffer buf_n3046( .i (n3045), .o (n3046) );
  buffer buf_n3047( .i (n3046), .o (n3047) );
  buffer buf_n3056( .i (n3055), .o (n3056) );
  buffer buf_n3057( .i (n3056), .o (n3057) );
  buffer buf_n3058( .i (n3057), .o (n3058) );
  buffer buf_n3059( .i (n3058), .o (n3059) );
  buffer buf_n3060( .i (n3059), .o (n3060) );
  buffer buf_n3061( .i (n3060), .o (n3061) );
  buffer buf_n3062( .i (n3061), .o (n3062) );
  buffer buf_n3063( .i (n3062), .o (n3063) );
  buffer buf_n3064( .i (n3063), .o (n3064) );
  buffer buf_n3065( .i (n3064), .o (n3065) );
  buffer buf_n3066( .i (n3065), .o (n3066) );
  buffer buf_n3067( .i (n3066), .o (n3067) );
  buffer buf_n3068( .i (n3067), .o (n3068) );
  buffer buf_n3069( .i (n3068), .o (n3069) );
  buffer buf_n3070( .i (n3069), .o (n3070) );
  buffer buf_n3071( .i (n3070), .o (n3071) );
  buffer buf_n3072( .i (n3071), .o (n3072) );
  buffer buf_n3073( .i (n3072), .o (n3073) );
  buffer buf_n3074( .i (n3073), .o (n3074) );
  buffer buf_n3075( .i (n3074), .o (n3075) );
  buffer buf_n3076( .i (n3075), .o (n3076) );
  buffer buf_n3077( .i (n3076), .o (n3077) );
  buffer buf_n3078( .i (n3077), .o (n3078) );
  buffer buf_n3079( .i (n3078), .o (n3079) );
  buffer buf_n3080( .i (n3079), .o (n3080) );
  buffer buf_n3081( .i (n3080), .o (n3081) );
  buffer buf_n3082( .i (n3081), .o (n3082) );
  buffer buf_n3083( .i (n3082), .o (n3083) );
  buffer buf_n3084( .i (n3083), .o (n3084) );
  buffer buf_n3085( .i (n3084), .o (n3085) );
  buffer buf_n3086( .i (n3085), .o (n3086) );
  buffer buf_n3087( .i (n3086), .o (n3087) );
  buffer buf_n3088( .i (n3087), .o (n3088) );
  buffer buf_n3089( .i (n3088), .o (n3089) );
  buffer buf_n3090( .i (n3089), .o (n3090) );
  buffer buf_n3091( .i (n3090), .o (n3091) );
  buffer buf_n3092( .i (n3091), .o (n3092) );
  buffer buf_n3093( .i (n3092), .o (n3093) );
  buffer buf_n3094( .i (n3093), .o (n3094) );
  buffer buf_n3095( .i (n3094), .o (n3095) );
  buffer buf_n3096( .i (n3095), .o (n3096) );
  buffer buf_n3097( .i (n3096), .o (n3097) );
  buffer buf_n3098( .i (n3097), .o (n3098) );
  buffer buf_n3099( .i (n3098), .o (n3099) );
  buffer buf_n3100( .i (n3099), .o (n3100) );
  buffer buf_n3101( .i (n3100), .o (n3101) );
  buffer buf_n3102( .i (n3101), .o (n3102) );
  buffer buf_n3103( .i (n3102), .o (n3103) );
  buffer buf_n3104( .i (n3103), .o (n3104) );
  buffer buf_n3105( .i (n3104), .o (n3105) );
  buffer buf_n3106( .i (n3105), .o (n3106) );
  buffer buf_n3107( .i (n3106), .o (n3107) );
  buffer buf_n3108( .i (n3107), .o (n3108) );
  buffer buf_n3109( .i (n3108), .o (n3109) );
  buffer buf_n3110( .i (n3109), .o (n3110) );
  buffer buf_n3111( .i (n3110), .o (n3111) );
  buffer buf_n3112( .i (n3111), .o (n3112) );
  buffer buf_n3113( .i (n3112), .o (n3113) );
  buffer buf_n3122( .i (n3121), .o (n3122) );
  buffer buf_n3123( .i (n3122), .o (n3123) );
  buffer buf_n3124( .i (n3123), .o (n3124) );
  buffer buf_n3125( .i (n3124), .o (n3125) );
  buffer buf_n3126( .i (n3125), .o (n3126) );
  buffer buf_n3127( .i (n3126), .o (n3127) );
  buffer buf_n3128( .i (n3127), .o (n3128) );
  buffer buf_n3129( .i (n3128), .o (n3129) );
  buffer buf_n3130( .i (n3129), .o (n3130) );
  buffer buf_n3131( .i (n3130), .o (n3131) );
  buffer buf_n3132( .i (n3131), .o (n3132) );
  buffer buf_n3133( .i (n3132), .o (n3133) );
  buffer buf_n3134( .i (n3133), .o (n3134) );
  buffer buf_n3135( .i (n3134), .o (n3135) );
  buffer buf_n3136( .i (n3135), .o (n3136) );
  buffer buf_n3137( .i (n3136), .o (n3137) );
  buffer buf_n3138( .i (n3137), .o (n3138) );
  buffer buf_n3139( .i (n3138), .o (n3139) );
  buffer buf_n3140( .i (n3139), .o (n3140) );
  buffer buf_n3141( .i (n3140), .o (n3141) );
  buffer buf_n3142( .i (n3141), .o (n3142) );
  buffer buf_n3143( .i (n3142), .o (n3143) );
  buffer buf_n3144( .i (n3143), .o (n3144) );
  buffer buf_n3145( .i (n3144), .o (n3145) );
  buffer buf_n3146( .i (n3145), .o (n3146) );
  buffer buf_n3147( .i (n3146), .o (n3147) );
  buffer buf_n3148( .i (n3147), .o (n3148) );
  buffer buf_n3149( .i (n3148), .o (n3149) );
  buffer buf_n3150( .i (n3149), .o (n3150) );
  buffer buf_n3151( .i (n3150), .o (n3151) );
  buffer buf_n3152( .i (n3151), .o (n3152) );
  buffer buf_n3153( .i (n3152), .o (n3153) );
  buffer buf_n3154( .i (n3153), .o (n3154) );
  buffer buf_n3155( .i (n3154), .o (n3155) );
  buffer buf_n3156( .i (n3155), .o (n3156) );
  buffer buf_n3157( .i (n3156), .o (n3157) );
  buffer buf_n3158( .i (n3157), .o (n3158) );
  buffer buf_n3159( .i (n3158), .o (n3159) );
  buffer buf_n3160( .i (n3159), .o (n3160) );
  buffer buf_n3161( .i (n3160), .o (n3161) );
  buffer buf_n3162( .i (n3161), .o (n3162) );
  buffer buf_n3163( .i (n3162), .o (n3163) );
  buffer buf_n3164( .i (n3163), .o (n3164) );
  buffer buf_n3165( .i (n3164), .o (n3165) );
  buffer buf_n3166( .i (n3165), .o (n3166) );
  buffer buf_n3167( .i (n3166), .o (n3167) );
  buffer buf_n3168( .i (n3167), .o (n3168) );
  buffer buf_n3169( .i (n3168), .o (n3169) );
  buffer buf_n3170( .i (n3169), .o (n3170) );
  buffer buf_n3171( .i (n3170), .o (n3171) );
  buffer buf_n3172( .i (n3171), .o (n3172) );
  buffer buf_n3173( .i (n3172), .o (n3173) );
  buffer buf_n3174( .i (n3173), .o (n3174) );
  buffer buf_n3175( .i (n3174), .o (n3175) );
  buffer buf_n3176( .i (n3175), .o (n3176) );
  buffer buf_n3177( .i (n3176), .o (n3177) );
  buffer buf_n3178( .i (n3177), .o (n3178) );
  buffer buf_n3179( .i (n3178), .o (n3179) );
  buffer buf_n3188( .i (n3187), .o (n3188) );
  buffer buf_n3189( .i (n3188), .o (n3189) );
  buffer buf_n3190( .i (n3189), .o (n3190) );
  buffer buf_n3191( .i (n3190), .o (n3191) );
  buffer buf_n3192( .i (n3191), .o (n3192) );
  buffer buf_n3193( .i (n3192), .o (n3193) );
  buffer buf_n3194( .i (n3193), .o (n3194) );
  buffer buf_n3195( .i (n3194), .o (n3195) );
  buffer buf_n3196( .i (n3195), .o (n3196) );
  buffer buf_n3197( .i (n3196), .o (n3197) );
  buffer buf_n3198( .i (n3197), .o (n3198) );
  buffer buf_n3199( .i (n3198), .o (n3199) );
  buffer buf_n3200( .i (n3199), .o (n3200) );
  buffer buf_n3201( .i (n3200), .o (n3201) );
  buffer buf_n3202( .i (n3201), .o (n3202) );
  buffer buf_n3203( .i (n3202), .o (n3203) );
  buffer buf_n3204( .i (n3203), .o (n3204) );
  buffer buf_n3205( .i (n3204), .o (n3205) );
  buffer buf_n3206( .i (n3205), .o (n3206) );
  buffer buf_n3207( .i (n3206), .o (n3207) );
  buffer buf_n3208( .i (n3207), .o (n3208) );
  buffer buf_n3209( .i (n3208), .o (n3209) );
  buffer buf_n3210( .i (n3209), .o (n3210) );
  buffer buf_n3211( .i (n3210), .o (n3211) );
  buffer buf_n3212( .i (n3211), .o (n3212) );
  buffer buf_n3213( .i (n3212), .o (n3213) );
  buffer buf_n3214( .i (n3213), .o (n3214) );
  buffer buf_n3215( .i (n3214), .o (n3215) );
  buffer buf_n3216( .i (n3215), .o (n3216) );
  buffer buf_n3217( .i (n3216), .o (n3217) );
  buffer buf_n3218( .i (n3217), .o (n3218) );
  buffer buf_n3219( .i (n3218), .o (n3219) );
  buffer buf_n3220( .i (n3219), .o (n3220) );
  buffer buf_n3221( .i (n3220), .o (n3221) );
  buffer buf_n3222( .i (n3221), .o (n3222) );
  buffer buf_n3223( .i (n3222), .o (n3223) );
  buffer buf_n3224( .i (n3223), .o (n3224) );
  buffer buf_n3225( .i (n3224), .o (n3225) );
  buffer buf_n3226( .i (n3225), .o (n3226) );
  buffer buf_n3227( .i (n3226), .o (n3227) );
  buffer buf_n3228( .i (n3227), .o (n3228) );
  buffer buf_n3229( .i (n3228), .o (n3229) );
  buffer buf_n3230( .i (n3229), .o (n3230) );
  buffer buf_n3231( .i (n3230), .o (n3231) );
  buffer buf_n3232( .i (n3231), .o (n3232) );
  buffer buf_n3233( .i (n3232), .o (n3233) );
  buffer buf_n3234( .i (n3233), .o (n3234) );
  buffer buf_n3235( .i (n3234), .o (n3235) );
  buffer buf_n3236( .i (n3235), .o (n3236) );
  buffer buf_n3237( .i (n3236), .o (n3237) );
  buffer buf_n3238( .i (n3237), .o (n3238) );
  buffer buf_n3239( .i (n3238), .o (n3239) );
  buffer buf_n3240( .i (n3239), .o (n3240) );
  buffer buf_n3241( .i (n3240), .o (n3241) );
  buffer buf_n3242( .i (n3241), .o (n3242) );
  buffer buf_n3243( .i (n3242), .o (n3243) );
  buffer buf_n3244( .i (n3243), .o (n3244) );
  buffer buf_n3245( .i (n3244), .o (n3245) );
  buffer buf_n3254( .i (n3253), .o (n3254) );
  buffer buf_n3255( .i (n3254), .o (n3255) );
  buffer buf_n3256( .i (n3255), .o (n3256) );
  buffer buf_n3257( .i (n3256), .o (n3257) );
  buffer buf_n3258( .i (n3257), .o (n3258) );
  buffer buf_n3259( .i (n3258), .o (n3259) );
  buffer buf_n3260( .i (n3259), .o (n3260) );
  buffer buf_n3261( .i (n3260), .o (n3261) );
  buffer buf_n3262( .i (n3261), .o (n3262) );
  buffer buf_n3263( .i (n3262), .o (n3263) );
  buffer buf_n3264( .i (n3263), .o (n3264) );
  buffer buf_n3265( .i (n3264), .o (n3265) );
  buffer buf_n3266( .i (n3265), .o (n3266) );
  buffer buf_n3267( .i (n3266), .o (n3267) );
  buffer buf_n3268( .i (n3267), .o (n3268) );
  buffer buf_n3269( .i (n3268), .o (n3269) );
  buffer buf_n3270( .i (n3269), .o (n3270) );
  buffer buf_n3271( .i (n3270), .o (n3271) );
  buffer buf_n3272( .i (n3271), .o (n3272) );
  buffer buf_n3273( .i (n3272), .o (n3273) );
  buffer buf_n3274( .i (n3273), .o (n3274) );
  buffer buf_n3275( .i (n3274), .o (n3275) );
  buffer buf_n3276( .i (n3275), .o (n3276) );
  buffer buf_n3277( .i (n3276), .o (n3277) );
  buffer buf_n3278( .i (n3277), .o (n3278) );
  buffer buf_n3279( .i (n3278), .o (n3279) );
  buffer buf_n3280( .i (n3279), .o (n3280) );
  buffer buf_n3281( .i (n3280), .o (n3281) );
  buffer buf_n3282( .i (n3281), .o (n3282) );
  buffer buf_n3283( .i (n3282), .o (n3283) );
  buffer buf_n3284( .i (n3283), .o (n3284) );
  buffer buf_n3285( .i (n3284), .o (n3285) );
  buffer buf_n3286( .i (n3285), .o (n3286) );
  buffer buf_n3287( .i (n3286), .o (n3287) );
  buffer buf_n3288( .i (n3287), .o (n3288) );
  buffer buf_n3289( .i (n3288), .o (n3289) );
  buffer buf_n3290( .i (n3289), .o (n3290) );
  buffer buf_n3291( .i (n3290), .o (n3291) );
  buffer buf_n3292( .i (n3291), .o (n3292) );
  buffer buf_n3293( .i (n3292), .o (n3293) );
  buffer buf_n3294( .i (n3293), .o (n3294) );
  buffer buf_n3295( .i (n3294), .o (n3295) );
  buffer buf_n3296( .i (n3295), .o (n3296) );
  buffer buf_n3297( .i (n3296), .o (n3297) );
  buffer buf_n3298( .i (n3297), .o (n3298) );
  buffer buf_n3299( .i (n3298), .o (n3299) );
  buffer buf_n3300( .i (n3299), .o (n3300) );
  buffer buf_n3301( .i (n3300), .o (n3301) );
  buffer buf_n3302( .i (n3301), .o (n3302) );
  buffer buf_n3303( .i (n3302), .o (n3303) );
  buffer buf_n3304( .i (n3303), .o (n3304) );
  buffer buf_n3305( .i (n3304), .o (n3305) );
  buffer buf_n3306( .i (n3305), .o (n3306) );
  buffer buf_n3307( .i (n3306), .o (n3307) );
  buffer buf_n3308( .i (n3307), .o (n3308) );
  buffer buf_n3309( .i (n3308), .o (n3309) );
  buffer buf_n3310( .i (n3309), .o (n3310) );
  buffer buf_n3311( .i (n3310), .o (n3311) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n2722( .i (n2721), .o (n2722) );
  buffer buf_n2723( .i (n2722), .o (n2723) );
  buffer buf_n2724( .i (n2723), .o (n2724) );
  buffer buf_n2725( .i (n2724), .o (n2725) );
  buffer buf_n2726( .i (n2725), .o (n2726) );
  buffer buf_n2727( .i (n2726), .o (n2727) );
  buffer buf_n2728( .i (n2727), .o (n2728) );
  buffer buf_n2729( .i (n2728), .o (n2729) );
  buffer buf_n2730( .i (n2729), .o (n2730) );
  buffer buf_n2731( .i (n2730), .o (n2731) );
  buffer buf_n2732( .i (n2731), .o (n2732) );
  buffer buf_n2733( .i (n2732), .o (n2733) );
  buffer buf_n2734( .i (n2733), .o (n2734) );
  buffer buf_n2735( .i (n2734), .o (n2735) );
  buffer buf_n2736( .i (n2735), .o (n2736) );
  buffer buf_n2737( .i (n2736), .o (n2737) );
  buffer buf_n2738( .i (n2737), .o (n2738) );
  buffer buf_n2739( .i (n2738), .o (n2739) );
  buffer buf_n2740( .i (n2739), .o (n2740) );
  buffer buf_n2741( .i (n2740), .o (n2741) );
  buffer buf_n2742( .i (n2741), .o (n2742) );
  buffer buf_n2743( .i (n2742), .o (n2743) );
  buffer buf_n2744( .i (n2743), .o (n2744) );
  buffer buf_n2745( .i (n2744), .o (n2745) );
  buffer buf_n2746( .i (n2745), .o (n2746) );
  buffer buf_n2747( .i (n2746), .o (n2747) );
  buffer buf_n2748( .i (n2747), .o (n2748) );
  buffer buf_n2749( .i (n2748), .o (n2749) );
  buffer buf_n2750( .i (n2749), .o (n2750) );
  buffer buf_n2751( .i (n2750), .o (n2751) );
  buffer buf_n2752( .i (n2751), .o (n2752) );
  buffer buf_n2753( .i (n2752), .o (n2753) );
  buffer buf_n2754( .i (n2753), .o (n2754) );
  buffer buf_n2755( .i (n2754), .o (n2755) );
  buffer buf_n2756( .i (n2755), .o (n2756) );
  buffer buf_n2757( .i (n2756), .o (n2757) );
  buffer buf_n2758( .i (n2757), .o (n2758) );
  buffer buf_n2759( .i (n2758), .o (n2759) );
  buffer buf_n2760( .i (n2759), .o (n2760) );
  buffer buf_n2761( .i (n2760), .o (n2761) );
  buffer buf_n2762( .i (n2761), .o (n2762) );
  buffer buf_n2763( .i (n2762), .o (n2763) );
  buffer buf_n2764( .i (n2763), .o (n2764) );
  buffer buf_n2765( .i (n2764), .o (n2765) );
  buffer buf_n2766( .i (n2765), .o (n2766) );
  buffer buf_n2767( .i (n2766), .o (n2767) );
  buffer buf_n2768( .i (n2767), .o (n2768) );
  buffer buf_n2769( .i (n2768), .o (n2769) );
  buffer buf_n2770( .i (n2769), .o (n2770) );
  buffer buf_n2771( .i (n2770), .o (n2771) );
  buffer buf_n2772( .i (n2771), .o (n2772) );
  buffer buf_n2773( .i (n2772), .o (n2773) );
  buffer buf_n2774( .i (n2773), .o (n2774) );
  buffer buf_n2775( .i (n2774), .o (n2775) );
  buffer buf_n2776( .i (n2775), .o (n2776) );
  buffer buf_n2777( .i (n2776), .o (n2777) );
  buffer buf_n2778( .i (n2777), .o (n2778) );
  buffer buf_n2779( .i (n2778), .o (n2779) );
  buffer buf_n3480( .i (N57), .o (n3480) );
  assign n10296 = n3459 | n3480 ;
  buffer buf_n10297( .i (n10296), .o (n10297) );
  buffer buf_n10298( .i (n10297), .o (n10298) );
  buffer buf_n10299( .i (n10298), .o (n10299) );
  buffer buf_n10300( .i (n10299), .o (n10300) );
  buffer buf_n10301( .i (n10300), .o (n10301) );
  buffer buf_n10302( .i (n10301), .o (n10302) );
  buffer buf_n10303( .i (n10302), .o (n10303) );
  buffer buf_n10304( .i (n10303), .o (n10304) );
  buffer buf_n10305( .i (n10304), .o (n10305) );
  buffer buf_n10306( .i (n10305), .o (n10306) );
  buffer buf_n10307( .i (n10306), .o (n10307) );
  buffer buf_n10308( .i (n10307), .o (n10308) );
  buffer buf_n10309( .i (n10308), .o (n10309) );
  buffer buf_n10310( .i (n10309), .o (n10310) );
  buffer buf_n10311( .i (n10310), .o (n10311) );
  buffer buf_n10312( .i (n10311), .o (n10312) );
  buffer buf_n10313( .i (n10312), .o (n10313) );
  buffer buf_n10314( .i (n10313), .o (n10314) );
  buffer buf_n10315( .i (n10314), .o (n10315) );
  buffer buf_n10316( .i (n10315), .o (n10316) );
  buffer buf_n10317( .i (n10316), .o (n10317) );
  buffer buf_n10318( .i (n10317), .o (n10318) );
  buffer buf_n10319( .i (n10318), .o (n10319) );
  buffer buf_n10320( .i (n10319), .o (n10320) );
  buffer buf_n10321( .i (n10320), .o (n10321) );
  buffer buf_n10322( .i (n10321), .o (n10322) );
  buffer buf_n10323( .i (n10322), .o (n10323) );
  buffer buf_n10324( .i (n10323), .o (n10324) );
  buffer buf_n10325( .i (n10324), .o (n10325) );
  buffer buf_n10326( .i (n10325), .o (n10326) );
  buffer buf_n10327( .i (n10326), .o (n10327) );
  buffer buf_n10328( .i (n10327), .o (n10328) );
  buffer buf_n10329( .i (n10328), .o (n10329) );
  buffer buf_n10330( .i (n10329), .o (n10330) );
  buffer buf_n10331( .i (n10330), .o (n10331) );
  buffer buf_n10332( .i (n10331), .o (n10332) );
  buffer buf_n10333( .i (n10332), .o (n10333) );
  buffer buf_n10334( .i (n10333), .o (n10334) );
  buffer buf_n10335( .i (n10334), .o (n10335) );
  buffer buf_n10336( .i (n10335), .o (n10336) );
  buffer buf_n10337( .i (n10336), .o (n10337) );
  buffer buf_n10338( .i (n10337), .o (n10338) );
  buffer buf_n10339( .i (n10338), .o (n10339) );
  buffer buf_n10340( .i (n10339), .o (n10340) );
  buffer buf_n10341( .i (n10340), .o (n10341) );
  buffer buf_n10342( .i (n10341), .o (n10342) );
  buffer buf_n10343( .i (n10342), .o (n10343) );
  buffer buf_n10344( .i (n10343), .o (n10344) );
  buffer buf_n10345( .i (n10344), .o (n10345) );
  buffer buf_n10346( .i (n10345), .o (n10346) );
  buffer buf_n10347( .i (n10346), .o (n10347) );
  buffer buf_n10348( .i (n10347), .o (n10348) );
  buffer buf_n10349( .i (n10348), .o (n10349) );
  buffer buf_n10350( .i (n10349), .o (n10350) );
  buffer buf_n10351( .i (n10350), .o (n10351) );
  buffer buf_n10352( .i (n10351), .o (n10352) );
  buffer buf_n10353( .i (n10352), .o (n10353) );
  buffer buf_n10354( .i (n10353), .o (n10354) );
  buffer buf_n10355( .i (n10354), .o (n10355) );
  buffer buf_n10356( .i (n10355), .o (n10356) );
  buffer buf_n10357( .i (n10356), .o (n10357) );
  buffer buf_n10358( .i (n10357), .o (n10358) );
  buffer buf_n10359( .i (n10358), .o (n10359) );
  buffer buf_n10360( .i (n10359), .o (n10360) );
  buffer buf_n8397( .i (n8396), .o (n8397) );
  buffer buf_n8398( .i (n8397), .o (n8398) );
  buffer buf_n8399( .i (n8398), .o (n8399) );
  buffer buf_n8400( .i (n8399), .o (n8400) );
  buffer buf_n8401( .i (n8400), .o (n8401) );
  buffer buf_n8402( .i (n8401), .o (n8402) );
  buffer buf_n8403( .i (n8402), .o (n8403) );
  buffer buf_n8404( .i (n8403), .o (n8404) );
  buffer buf_n8405( .i (n8404), .o (n8405) );
  buffer buf_n8406( .i (n8405), .o (n8406) );
  buffer buf_n8407( .i (n8406), .o (n8407) );
  buffer buf_n8408( .i (n8407), .o (n8408) );
  buffer buf_n8409( .i (n8408), .o (n8409) );
  buffer buf_n8410( .i (n8409), .o (n8410) );
  buffer buf_n8411( .i (n8410), .o (n8411) );
  buffer buf_n8412( .i (n8411), .o (n8412) );
  buffer buf_n8413( .i (n8412), .o (n8413) );
  buffer buf_n8414( .i (n8413), .o (n8414) );
  buffer buf_n8415( .i (n8414), .o (n8415) );
  buffer buf_n8416( .i (n8415), .o (n8416) );
  buffer buf_n8417( .i (n8416), .o (n8417) );
  buffer buf_n8418( .i (n8417), .o (n8418) );
  buffer buf_n8419( .i (n8418), .o (n8419) );
  buffer buf_n8420( .i (n8419), .o (n8420) );
  buffer buf_n8421( .i (n8420), .o (n8421) );
  buffer buf_n8422( .i (n8421), .o (n8422) );
  buffer buf_n8423( .i (n8422), .o (n8423) );
  buffer buf_n8424( .i (n8423), .o (n8424) );
  buffer buf_n8425( .i (n8424), .o (n8425) );
  buffer buf_n8426( .i (n8425), .o (n8426) );
  buffer buf_n8427( .i (n8426), .o (n8427) );
  buffer buf_n8428( .i (n8427), .o (n8428) );
  buffer buf_n8429( .i (n8428), .o (n8429) );
  buffer buf_n8430( .i (n8429), .o (n8430) );
  buffer buf_n8431( .i (n8430), .o (n8431) );
  buffer buf_n8432( .i (n8431), .o (n8432) );
  buffer buf_n8433( .i (n8432), .o (n8433) );
  buffer buf_n8434( .i (n8433), .o (n8434) );
  buffer buf_n8435( .i (n8434), .o (n8435) );
  buffer buf_n8436( .i (n8435), .o (n8436) );
  buffer buf_n8437( .i (n8436), .o (n8437) );
  buffer buf_n8438( .i (n8437), .o (n8438) );
  buffer buf_n8439( .i (n8438), .o (n8439) );
  buffer buf_n8440( .i (n8439), .o (n8440) );
  buffer buf_n8441( .i (n8440), .o (n8441) );
  buffer buf_n8442( .i (n8441), .o (n8442) );
  buffer buf_n8443( .i (n8442), .o (n8443) );
  buffer buf_n8444( .i (n8443), .o (n8444) );
  buffer buf_n8445( .i (n8444), .o (n8445) );
  buffer buf_n8446( .i (n8445), .o (n8446) );
  buffer buf_n8447( .i (n8446), .o (n8447) );
  buffer buf_n8448( .i (n8447), .o (n8448) );
  buffer buf_n8449( .i (n8448), .o (n8449) );
  buffer buf_n8450( .i (n8449), .o (n8450) );
  buffer buf_n8451( .i (n8450), .o (n8451) );
  buffer buf_n8452( .i (n8451), .o (n8452) );
  buffer buf_n8453( .i (n8452), .o (n8453) );
  buffer buf_n8454( .i (n8453), .o (n8454) );
  buffer buf_n8455( .i (n8454), .o (n8455) );
  buffer buf_n8456( .i (n8455), .o (n8456) );
  buffer buf_n8457( .i (n8456), .o (n8457) );
  buffer buf_n8458( .i (n8457), .o (n8458) );
  buffer buf_n8459( .i (n8458), .o (n8459) );
  buffer buf_n8464( .i (n8463), .o (n8464) );
  buffer buf_n8465( .i (n8464), .o (n8465) );
  buffer buf_n8466( .i (n8465), .o (n8466) );
  buffer buf_n8467( .i (n8466), .o (n8467) );
  buffer buf_n8468( .i (n8467), .o (n8468) );
  buffer buf_n8469( .i (n8468), .o (n8469) );
  buffer buf_n8470( .i (n8469), .o (n8470) );
  buffer buf_n8471( .i (n8470), .o (n8471) );
  buffer buf_n8472( .i (n8471), .o (n8472) );
  buffer buf_n8473( .i (n8472), .o (n8473) );
  buffer buf_n8474( .i (n8473), .o (n8474) );
  buffer buf_n8475( .i (n8474), .o (n8475) );
  buffer buf_n8476( .i (n8475), .o (n8476) );
  buffer buf_n8477( .i (n8476), .o (n8477) );
  buffer buf_n8478( .i (n8477), .o (n8478) );
  buffer buf_n8479( .i (n8478), .o (n8479) );
  buffer buf_n8480( .i (n8479), .o (n8480) );
  buffer buf_n8481( .i (n8480), .o (n8481) );
  buffer buf_n8482( .i (n8481), .o (n8482) );
  buffer buf_n8483( .i (n8482), .o (n8483) );
  buffer buf_n8484( .i (n8483), .o (n8484) );
  buffer buf_n8485( .i (n8484), .o (n8485) );
  buffer buf_n8486( .i (n8485), .o (n8486) );
  buffer buf_n8487( .i (n8486), .o (n8487) );
  buffer buf_n8488( .i (n8487), .o (n8488) );
  buffer buf_n8489( .i (n8488), .o (n8489) );
  buffer buf_n8490( .i (n8489), .o (n8490) );
  buffer buf_n8491( .i (n8490), .o (n8491) );
  buffer buf_n8492( .i (n8491), .o (n8492) );
  buffer buf_n8493( .i (n8492), .o (n8493) );
  buffer buf_n8494( .i (n8493), .o (n8494) );
  buffer buf_n8495( .i (n8494), .o (n8495) );
  buffer buf_n8496( .i (n8495), .o (n8496) );
  buffer buf_n8497( .i (n8496), .o (n8497) );
  buffer buf_n8498( .i (n8497), .o (n8498) );
  buffer buf_n8499( .i (n8498), .o (n8499) );
  buffer buf_n8500( .i (n8499), .o (n8500) );
  buffer buf_n8501( .i (n8500), .o (n8501) );
  buffer buf_n8502( .i (n8501), .o (n8502) );
  buffer buf_n8503( .i (n8502), .o (n8503) );
  buffer buf_n8504( .i (n8503), .o (n8504) );
  buffer buf_n8505( .i (n8504), .o (n8505) );
  buffer buf_n8506( .i (n8505), .o (n8506) );
  buffer buf_n8507( .i (n8506), .o (n8507) );
  buffer buf_n8508( .i (n8507), .o (n8508) );
  buffer buf_n8509( .i (n8508), .o (n8509) );
  buffer buf_n8510( .i (n8509), .o (n8510) );
  buffer buf_n8511( .i (n8510), .o (n8511) );
  buffer buf_n8512( .i (n8511), .o (n8512) );
  buffer buf_n8513( .i (n8512), .o (n8513) );
  buffer buf_n8514( .i (n8513), .o (n8514) );
  buffer buf_n8515( .i (n8514), .o (n8515) );
  buffer buf_n8516( .i (n8515), .o (n8516) );
  buffer buf_n8517( .i (n8516), .o (n8517) );
  buffer buf_n8518( .i (n8517), .o (n8518) );
  buffer buf_n8519( .i (n8518), .o (n8519) );
  buffer buf_n8520( .i (n8519), .o (n8520) );
  buffer buf_n8521( .i (n8520), .o (n8521) );
  buffer buf_n8522( .i (n8521), .o (n8522) );
  buffer buf_n8523( .i (n8522), .o (n8523) );
  buffer buf_n8524( .i (n8523), .o (n8524) );
  buffer buf_n8525( .i (n8524), .o (n8525) );
  buffer buf_n8526( .i (n8525), .o (n8526) );
  buffer buf_n8532( .i (n8531), .o (n8532) );
  buffer buf_n8533( .i (n8532), .o (n8533) );
  buffer buf_n8534( .i (n8533), .o (n8534) );
  buffer buf_n8535( .i (n8534), .o (n8535) );
  buffer buf_n8536( .i (n8535), .o (n8536) );
  buffer buf_n8537( .i (n8536), .o (n8537) );
  buffer buf_n8538( .i (n8537), .o (n8538) );
  buffer buf_n8539( .i (n8538), .o (n8539) );
  buffer buf_n8540( .i (n8539), .o (n8540) );
  buffer buf_n8541( .i (n8540), .o (n8541) );
  buffer buf_n8542( .i (n8541), .o (n8542) );
  buffer buf_n8543( .i (n8542), .o (n8543) );
  buffer buf_n8544( .i (n8543), .o (n8544) );
  buffer buf_n8545( .i (n8544), .o (n8545) );
  buffer buf_n8546( .i (n8545), .o (n8546) );
  buffer buf_n8547( .i (n8546), .o (n8547) );
  buffer buf_n8548( .i (n8547), .o (n8548) );
  buffer buf_n8549( .i (n8548), .o (n8549) );
  buffer buf_n8550( .i (n8549), .o (n8550) );
  buffer buf_n8551( .i (n8550), .o (n8551) );
  buffer buf_n8552( .i (n8551), .o (n8552) );
  buffer buf_n8553( .i (n8552), .o (n8553) );
  buffer buf_n8554( .i (n8553), .o (n8554) );
  buffer buf_n8555( .i (n8554), .o (n8555) );
  buffer buf_n8556( .i (n8555), .o (n8556) );
  buffer buf_n8557( .i (n8556), .o (n8557) );
  buffer buf_n8558( .i (n8557), .o (n8558) );
  buffer buf_n8559( .i (n8558), .o (n8559) );
  buffer buf_n8560( .i (n8559), .o (n8560) );
  buffer buf_n8561( .i (n8560), .o (n8561) );
  buffer buf_n8562( .i (n8561), .o (n8562) );
  buffer buf_n8563( .i (n8562), .o (n8563) );
  buffer buf_n8564( .i (n8563), .o (n8564) );
  buffer buf_n8565( .i (n8564), .o (n8565) );
  buffer buf_n8566( .i (n8565), .o (n8566) );
  buffer buf_n8567( .i (n8566), .o (n8567) );
  buffer buf_n8568( .i (n8567), .o (n8568) );
  buffer buf_n8569( .i (n8568), .o (n8569) );
  buffer buf_n8570( .i (n8569), .o (n8570) );
  buffer buf_n8571( .i (n8570), .o (n8571) );
  buffer buf_n8572( .i (n8571), .o (n8572) );
  buffer buf_n8573( .i (n8572), .o (n8573) );
  buffer buf_n8574( .i (n8573), .o (n8574) );
  buffer buf_n8575( .i (n8574), .o (n8575) );
  buffer buf_n8576( .i (n8575), .o (n8576) );
  buffer buf_n8577( .i (n8576), .o (n8577) );
  buffer buf_n8578( .i (n8577), .o (n8578) );
  buffer buf_n8579( .i (n8578), .o (n8579) );
  buffer buf_n8580( .i (n8579), .o (n8580) );
  buffer buf_n8581( .i (n8580), .o (n8581) );
  buffer buf_n8582( .i (n8581), .o (n8582) );
  buffer buf_n8583( .i (n8582), .o (n8583) );
  buffer buf_n8584( .i (n8583), .o (n8584) );
  buffer buf_n8585( .i (n8584), .o (n8585) );
  buffer buf_n8586( .i (n8585), .o (n8586) );
  buffer buf_n8587( .i (n8586), .o (n8587) );
  buffer buf_n8588( .i (n8587), .o (n8588) );
  buffer buf_n8589( .i (n8588), .o (n8589) );
  buffer buf_n8590( .i (n8589), .o (n8590) );
  buffer buf_n8591( .i (n8590), .o (n8591) );
  buffer buf_n8592( .i (n8591), .o (n8592) );
  buffer buf_n8593( .i (n8592), .o (n8593) );
  buffer buf_n8594( .i (n8593), .o (n8594) );
  buffer buf_n8599( .i (n8598), .o (n8599) );
  buffer buf_n8600( .i (n8599), .o (n8600) );
  buffer buf_n8601( .i (n8600), .o (n8601) );
  buffer buf_n8602( .i (n8601), .o (n8602) );
  buffer buf_n8603( .i (n8602), .o (n8603) );
  buffer buf_n8604( .i (n8603), .o (n8604) );
  buffer buf_n8605( .i (n8604), .o (n8605) );
  buffer buf_n8606( .i (n8605), .o (n8606) );
  buffer buf_n8607( .i (n8606), .o (n8607) );
  buffer buf_n8608( .i (n8607), .o (n8608) );
  buffer buf_n8609( .i (n8608), .o (n8609) );
  buffer buf_n8610( .i (n8609), .o (n8610) );
  buffer buf_n8611( .i (n8610), .o (n8611) );
  buffer buf_n8612( .i (n8611), .o (n8612) );
  buffer buf_n8613( .i (n8612), .o (n8613) );
  buffer buf_n8614( .i (n8613), .o (n8614) );
  buffer buf_n8615( .i (n8614), .o (n8615) );
  buffer buf_n8616( .i (n8615), .o (n8616) );
  buffer buf_n8617( .i (n8616), .o (n8617) );
  buffer buf_n8618( .i (n8617), .o (n8618) );
  buffer buf_n8619( .i (n8618), .o (n8619) );
  buffer buf_n8620( .i (n8619), .o (n8620) );
  buffer buf_n8621( .i (n8620), .o (n8621) );
  buffer buf_n8622( .i (n8621), .o (n8622) );
  buffer buf_n8623( .i (n8622), .o (n8623) );
  buffer buf_n8624( .i (n8623), .o (n8624) );
  buffer buf_n8625( .i (n8624), .o (n8625) );
  buffer buf_n8626( .i (n8625), .o (n8626) );
  buffer buf_n8627( .i (n8626), .o (n8627) );
  buffer buf_n8628( .i (n8627), .o (n8628) );
  buffer buf_n8629( .i (n8628), .o (n8629) );
  buffer buf_n8630( .i (n8629), .o (n8630) );
  buffer buf_n8631( .i (n8630), .o (n8631) );
  buffer buf_n8632( .i (n8631), .o (n8632) );
  buffer buf_n8633( .i (n8632), .o (n8633) );
  buffer buf_n8634( .i (n8633), .o (n8634) );
  buffer buf_n8635( .i (n8634), .o (n8635) );
  buffer buf_n8636( .i (n8635), .o (n8636) );
  buffer buf_n8637( .i (n8636), .o (n8637) );
  buffer buf_n8638( .i (n8637), .o (n8638) );
  buffer buf_n8639( .i (n8638), .o (n8639) );
  buffer buf_n8640( .i (n8639), .o (n8640) );
  buffer buf_n8641( .i (n8640), .o (n8641) );
  buffer buf_n8642( .i (n8641), .o (n8642) );
  buffer buf_n8643( .i (n8642), .o (n8643) );
  buffer buf_n8644( .i (n8643), .o (n8644) );
  buffer buf_n8645( .i (n8644), .o (n8645) );
  buffer buf_n8646( .i (n8645), .o (n8646) );
  buffer buf_n8647( .i (n8646), .o (n8647) );
  buffer buf_n8648( .i (n8647), .o (n8648) );
  buffer buf_n8649( .i (n8648), .o (n8649) );
  buffer buf_n8650( .i (n8649), .o (n8650) );
  buffer buf_n8651( .i (n8650), .o (n8651) );
  buffer buf_n8652( .i (n8651), .o (n8652) );
  buffer buf_n8653( .i (n8652), .o (n8653) );
  buffer buf_n8654( .i (n8653), .o (n8654) );
  buffer buf_n8655( .i (n8654), .o (n8655) );
  buffer buf_n8656( .i (n8655), .o (n8656) );
  buffer buf_n8657( .i (n8656), .o (n8657) );
  buffer buf_n8658( .i (n8657), .o (n8658) );
  buffer buf_n8659( .i (n8658), .o (n8659) );
  buffer buf_n8660( .i (n8659), .o (n8660) );
  buffer buf_n8661( .i (n8660), .o (n8661) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  assign N10025 = ~n3686 ;
  assign N10101 = ~n6196 ;
  assign N10102 = n7013 ;
  assign N10103 = n7013 ;
  assign N10104 = ~n6196 ;
  assign N10109 = ~n7075 ;
  assign N10110 = ~n7124 ;
  assign N10111 = ~n7181 ;
  assign N10112 = ~n7236 ;
  assign N10350 = ~n7288 ;
  assign N10351 = ~n7329 ;
  assign N10352 = ~n7368 ;
  assign N10353 = ~n7408 ;
  assign N10574 = ~n7643 ;
  assign N10575 = ~n7866 ;
  assign N10576 = ~n8093 ;
  assign N10628 = n7013 ;
  assign N10632 = ~n8118 ;
  assign N10641 = ~n8132 ;
  assign N10704 = n6607 ;
  assign N10706 = ~n6196 ;
  assign N10711 = n8219 ;
  assign N10712 = ~n8245 ;
  assign N10713 = ~n8273 ;
  assign N10714 = ~n8295 ;
  assign N10715 = ~n8345 ;
  assign N10716 = ~n8362 ;
  assign N10717 = ~n8381 ;
  assign N10718 = ~n8392 ;
  assign N10729 = ~n8725 ;
  assign N10759 = ~n6196 ;
  assign N10760 = ~n8781 ;
  assign N10761 = ~n8806 ;
  assign N10762 = ~n8866 ;
  assign N10763 = ~n8921 ;
  assign N10827 = ~n8960 ;
  assign N10837 = n8968 ;
  assign N10838 = n8968 ;
  assign N10839 = n8974 ;
  assign N10840 = n8974 ;
  assign N10868 = ~n9021 ;
  assign N10869 = ~n9072 ;
  assign N10870 = ~n9131 ;
  assign N10871 = ~n9165 ;
  assign N10905 = ~n9222 ;
  assign N10906 = ~n9282 ;
  assign N10907 = ~n9316 ;
  assign N10908 = ~n9347 ;
  assign N1110 = ~n9412 ;
  assign N1111 = ~n484 ;
  assign N1112 = ~n9412 ;
  assign N1113 = ~n9477 ;
  assign N1114 = ~n484 ;
  assign N11333 = ~n9719 ;
  assign N11334 = n9867 ;
  assign N11340 = n10047 ;
  assign N11342 = n10231 ;
  assign N1489 = ~n9477 ;
  assign N1490 = n273 ;
  assign N1781 = n10295 ;
  assign N241_O = n850 ;
  assign N387 = n273 ;
  assign N388 = n273 ;
  assign N478 = n918 ;
  assign N482 = n1050 ;
  assign N484 = n1116 ;
  assign N486 = n1186 ;
  assign N489 = n1252 ;
  assign N492 = n1318 ;
  assign N501 = n1385 ;
  assign N505 = n1517 ;
  assign N507 = n1583 ;
  assign N509 = n1649 ;
  assign N511 = n1715 ;
  assign N513 = n1785 ;
  assign N515 = n1851 ;
  assign N517 = n1917 ;
  assign N519 = n1983 ;
  assign N535 = n2049 ;
  assign N537 = n2115 ;
  assign N539 = n2181 ;
  assign N541 = n2247 ;
  assign N543 = n2313 ;
  assign N545 = n2383 ;
  assign N547 = n2449 ;
  assign N549 = n2515 ;
  assign N551 = n2581 ;
  assign N553 = n2647 ;
  assign N556 = n2713 ;
  assign N559 = n2845 ;
  assign N561 = n2911 ;
  assign N563 = n2977 ;
  assign N565 = n3047 ;
  assign N567 = n3113 ;
  assign N569 = n3179 ;
  assign N571 = n3245 ;
  assign N573 = n3311 ;
  assign N582 = ~n484 ;
  assign N643 = n984 ;
  assign N707 = n1451 ;
  assign N813 = n2779 ;
  assign N881 = n10360 ;
  assign N882 = ~n8459 ;
  assign N883 = ~n8526 ;
  assign N884 = ~n8594 ;
  assign N885 = ~n8661 ;
  assign N889 = n273 ;
  assign N945 = n347 ;
endmodule
