module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( N1 , N103 , N120 , N137 , N154 , N171 , N18 , N188 , N205 , N222 , N239 , N256 , N273 , N290 , N307 , N324 , N341 , N35 , N358 , N375 , N392 , N409 , N426 , N443 , N460 , N477 , N494 , N511 , N52 , N528 , N69 , N86 , N1581 , N1901 , N2223 , N2548 , N2877 , N3211 , N3552 , N3895 , N4241 , N4591 , N4946 , N5308 , N545 , N5672 , N5971 , N6123 , N6150 , N6160 , N6170 , N6180 , N6190 , N6200 , N6210 , N6220 , N6230 , N6240 , N6250 , N6260 , N6270 , N6280 , N6287 , N6288 );
  input N1 , N103 , N120 , N137 , N154 , N171 , N18 , N188 , N205 , N222 , N239 , N256 , N273 , N290 , N307 , N324 , N341 , N35 , N358 , N375 , N392 , N409 , N426 , N443 , N460 , N477 , N494 , N511 , N52 , N528 , N69 , N86 ;
  output N1581 , N1901 , N2223 , N2548 , N2877 , N3211 , N3552 , N3895 , N4241 , N4591 , N4946 , N5308 , N545 , N5672 , N5971 , N6123 , N6150 , N6160 , N6170 , N6180 , N6190 , N6200 , N6210 , N6220 , N6230 , N6240 , N6250 , N6260 , N6270 , N6280 , N6287 , N6288 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 ;
  assign n33 = N18 & N290 ;
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  assign n36 = N1 & N273 ;
  buffer buf_n37( .i (n36), .o (n37) );
  assign n38 = n35 & n37 ;
  buffer buf_n39( .i (n38), .o (n39) );
  assign n41 = N18 & N273 ;
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  assign n46 = N1 & N290 ;
  assign n47 = n45 | n46 ;
  assign n48 = ~n39 & n47 ;
  assign n49 = N1 & N307 ;
  buffer buf_n50( .i (n49), .o (n50) );
  assign n52 = N290 & N35 ;
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  assign n55 = n42 & n54 ;
  buffer buf_n56( .i (n55), .o (n56) );
  assign n58 = N273 & N35 ;
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  assign n63 = n34 | n62 ;
  assign n64 = ~n56 & n63 ;
  buffer buf_n65( .i (n64), .o (n65) );
  assign n67 = n39 | n65 ;
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n66( .i (n65), .o (n66) );
  assign n73 = n40 & n66 ;
  assign n74 = n68 & ~n73 ;
  buffer buf_n75( .i (n74), .o (n75) );
  assign n77 = ~n50 & n75 ;
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n76( .i (n75), .o (n76) );
  assign n79 = n51 & ~n76 ;
  assign n80 = n78 | n79 ;
  assign n81 = N1 & N324 ;
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  assign n84 = n72 & ~n78 ;
  buffer buf_n85( .i (n84), .o (n85) );
  assign n87 = N18 & N307 ;
  buffer buf_n88( .i (n87), .o (n88) );
  assign n92 = N290 & N52 ;
  buffer buf_n93( .i (n92), .o (n93) );
  assign n95 = n59 & n93 ;
  buffer buf_n96( .i (n95), .o (n96) );
  assign n100 = N273 & N52 ;
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  assign n103 = n53 | n102 ;
  assign n104 = ~n96 & n103 ;
  buffer buf_n105( .i (n104), .o (n105) );
  assign n107 = n56 | n105 ;
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n106( .i (n105), .o (n106) );
  assign n113 = n57 & n106 ;
  assign n114 = n108 & ~n113 ;
  buffer buf_n115( .i (n114), .o (n115) );
  assign n119 = ~n88 & n115 ;
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  assign n123 = n91 & ~n118 ;
  assign n124 = n122 | n123 ;
  buffer buf_n125( .i (n124), .o (n125) );
  assign n127 = n85 | n125 ;
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n126( .i (n125), .o (n126) );
  assign n133 = n86 & n126 ;
  assign n134 = n128 & ~n133 ;
  buffer buf_n135( .i (n134), .o (n135) );
  assign n137 = ~n82 & n135 ;
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n136( .i (n135), .o (n136) );
  assign n139 = n83 & ~n136 ;
  assign n140 = n138 | n139 ;
  assign n141 = N1 & N341 ;
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  assign n144 = n132 & ~n138 ;
  buffer buf_n145( .i (n144), .o (n145) );
  assign n147 = N18 & N324 ;
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  assign n152 = n112 & ~n120 ;
  buffer buf_n153( .i (n152), .o (n153) );
  assign n155 = N307 & N35 ;
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  assign n158 = N290 & N69 ;
  buffer buf_n159( .i (n158), .o (n159) );
  assign n161 = n101 & n159 ;
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n94( .i (n93), .o (n94) );
  assign n166 = N273 & N69 ;
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = n94 | n168 ;
  assign n170 = ~n162 & n169 ;
  buffer buf_n171( .i (n170), .o (n171) );
  assign n173 = n98 | n171 ;
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n172( .i (n171), .o (n172) );
  assign n179 = n99 & n172 ;
  assign n180 = n174 & ~n179 ;
  buffer buf_n181( .i (n180), .o (n181) );
  assign n183 = ~n156 & n181 ;
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n182( .i (n181), .o (n182) );
  assign n185 = n157 & ~n182 ;
  assign n186 = n184 | n185 ;
  buffer buf_n187( .i (n186), .o (n187) );
  assign n189 = n153 | n187 ;
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n188( .i (n187), .o (n188) );
  assign n195 = n154 & n188 ;
  assign n196 = n190 & ~n195 ;
  buffer buf_n197( .i (n196), .o (n197) );
  assign n201 = ~n148 & n197 ;
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  assign n205 = n151 & ~n200 ;
  assign n206 = n204 | n205 ;
  buffer buf_n207( .i (n206), .o (n207) );
  assign n209 = n145 | n207 ;
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n208( .i (n207), .o (n208) );
  assign n215 = n146 & n208 ;
  assign n216 = n210 & ~n215 ;
  buffer buf_n217( .i (n216), .o (n217) );
  assign n219 = ~n142 & n217 ;
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n218( .i (n217), .o (n218) );
  assign n221 = n143 & ~n218 ;
  assign n222 = n220 | n221 ;
  assign n223 = N1 & N358 ;
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n226 = n214 & ~n220 ;
  buffer buf_n227( .i (n226), .o (n227) );
  assign n229 = N18 & N341 ;
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  assign n234 = n194 & ~n202 ;
  buffer buf_n235( .i (n234), .o (n235) );
  assign n237 = N324 & N35 ;
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  assign n240 = n178 & ~n184 ;
  buffer buf_n241( .i (n240), .o (n241) );
  assign n243 = N307 & N52 ;
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  assign n246 = N290 & N86 ;
  buffer buf_n247( .i (n246), .o (n247) );
  assign n249 = n167 & n247 ;
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n160( .i (n159), .o (n160) );
  assign n254 = N273 & N86 ;
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  assign n257 = n160 | n256 ;
  assign n258 = ~n250 & n257 ;
  buffer buf_n259( .i (n258), .o (n259) );
  assign n261 = n164 | n259 ;
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n260( .i (n259), .o (n260) );
  assign n267 = n165 & n260 ;
  assign n268 = n262 & ~n267 ;
  buffer buf_n269( .i (n268), .o (n269) );
  assign n271 = ~n244 & n269 ;
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n270( .i (n269), .o (n270) );
  assign n273 = n245 & ~n270 ;
  assign n274 = n272 | n273 ;
  buffer buf_n275( .i (n274), .o (n275) );
  assign n277 = n241 | n275 ;
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n276( .i (n275), .o (n276) );
  assign n283 = n242 & n276 ;
  assign n284 = n278 & ~n283 ;
  buffer buf_n285( .i (n284), .o (n285) );
  assign n287 = ~n238 & n285 ;
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n286( .i (n285), .o (n286) );
  assign n289 = n239 & ~n286 ;
  assign n290 = n288 | n289 ;
  buffer buf_n291( .i (n290), .o (n291) );
  assign n293 = n235 | n291 ;
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n292( .i (n291), .o (n292) );
  assign n299 = n236 & n292 ;
  assign n300 = n294 & ~n299 ;
  buffer buf_n301( .i (n300), .o (n301) );
  assign n305 = ~n230 & n301 ;
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  assign n309 = n233 & ~n304 ;
  assign n310 = n308 | n309 ;
  buffer buf_n311( .i (n310), .o (n311) );
  assign n313 = n227 | n311 ;
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n312( .i (n311), .o (n312) );
  assign n319 = n228 & n312 ;
  assign n320 = n314 & ~n319 ;
  buffer buf_n321( .i (n320), .o (n321) );
  assign n323 = ~n224 & n321 ;
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n322( .i (n321), .o (n322) );
  assign n325 = n225 & ~n322 ;
  assign n326 = n324 | n325 ;
  assign n327 = N1 & N375 ;
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  assign n330 = n318 & ~n324 ;
  buffer buf_n331( .i (n330), .o (n331) );
  assign n333 = N18 & N358 ;
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  assign n338 = n298 & ~n306 ;
  buffer buf_n339( .i (n338), .o (n339) );
  assign n341 = N341 & N35 ;
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  assign n344 = n282 & ~n288 ;
  buffer buf_n345( .i (n344), .o (n345) );
  assign n347 = N324 & N52 ;
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  assign n350 = n266 & ~n272 ;
  buffer buf_n351( .i (n350), .o (n351) );
  assign n353 = N307 & N69 ;
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  assign n356 = N103 & N290 ;
  buffer buf_n357( .i (n356), .o (n357) );
  assign n359 = n255 & n357 ;
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n248( .i (n247), .o (n248) );
  assign n364 = N103 & N273 ;
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  assign n367 = n248 | n366 ;
  assign n368 = ~n360 & n367 ;
  buffer buf_n369( .i (n368), .o (n369) );
  assign n371 = n252 | n369 ;
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n370( .i (n369), .o (n370) );
  assign n377 = n253 & n370 ;
  assign n378 = n372 & ~n377 ;
  buffer buf_n379( .i (n378), .o (n379) );
  assign n381 = ~n354 & n379 ;
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n380( .i (n379), .o (n380) );
  assign n383 = n355 & ~n380 ;
  assign n384 = n382 | n383 ;
  buffer buf_n385( .i (n384), .o (n385) );
  assign n387 = n351 | n385 ;
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n386( .i (n385), .o (n386) );
  assign n393 = n352 & n386 ;
  assign n394 = n388 & ~n393 ;
  buffer buf_n395( .i (n394), .o (n395) );
  assign n397 = ~n348 & n395 ;
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n396( .i (n395), .o (n396) );
  assign n399 = n349 & ~n396 ;
  assign n400 = n398 | n399 ;
  buffer buf_n401( .i (n400), .o (n401) );
  assign n403 = n345 | n401 ;
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n402( .i (n401), .o (n402) );
  assign n409 = n346 & n402 ;
  assign n410 = n404 & ~n409 ;
  buffer buf_n411( .i (n410), .o (n411) );
  assign n413 = ~n342 & n411 ;
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n412( .i (n411), .o (n412) );
  assign n415 = n343 & ~n412 ;
  assign n416 = n414 | n415 ;
  buffer buf_n417( .i (n416), .o (n417) );
  assign n419 = n339 | n417 ;
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n418( .i (n417), .o (n418) );
  assign n425 = n340 & n418 ;
  assign n426 = n420 & ~n425 ;
  buffer buf_n427( .i (n426), .o (n427) );
  assign n431 = ~n334 & n427 ;
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  assign n435 = n337 & ~n430 ;
  assign n436 = n434 | n435 ;
  buffer buf_n437( .i (n436), .o (n437) );
  assign n439 = n331 | n437 ;
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n438( .i (n437), .o (n438) );
  assign n445 = n332 & n438 ;
  assign n446 = n440 & ~n445 ;
  buffer buf_n447( .i (n446), .o (n447) );
  assign n449 = ~n328 & n447 ;
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n448( .i (n447), .o (n448) );
  assign n451 = n329 & ~n448 ;
  assign n452 = n450 | n451 ;
  assign n453 = N1 & N392 ;
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  assign n456 = n444 & ~n450 ;
  buffer buf_n457( .i (n456), .o (n457) );
  assign n459 = N18 & N375 ;
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  assign n464 = n424 & ~n432 ;
  buffer buf_n465( .i (n464), .o (n465) );
  assign n467 = N35 & N358 ;
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  assign n470 = n408 & ~n414 ;
  buffer buf_n471( .i (n470), .o (n471) );
  assign n473 = N341 & N52 ;
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  assign n476 = n392 & ~n398 ;
  buffer buf_n477( .i (n476), .o (n477) );
  assign n479 = N324 & N69 ;
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  assign n482 = n376 & ~n382 ;
  buffer buf_n483( .i (n482), .o (n483) );
  assign n485 = N307 & N86 ;
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  assign n488 = N120 & N290 ;
  buffer buf_n489( .i (n488), .o (n489) );
  assign n491 = n365 & n489 ;
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n358( .i (n357), .o (n358) );
  assign n496 = N120 & N273 ;
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  assign n499 = n358 | n498 ;
  assign n500 = ~n492 & n499 ;
  buffer buf_n501( .i (n500), .o (n501) );
  assign n503 = n362 | n501 ;
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n502( .i (n501), .o (n502) );
  assign n509 = n363 & n502 ;
  assign n510 = n504 & ~n509 ;
  buffer buf_n511( .i (n510), .o (n511) );
  assign n513 = ~n486 & n511 ;
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n512( .i (n511), .o (n512) );
  assign n515 = n487 & ~n512 ;
  assign n516 = n514 | n515 ;
  buffer buf_n517( .i (n516), .o (n517) );
  assign n519 = n483 | n517 ;
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n518( .i (n517), .o (n518) );
  assign n525 = n484 & n518 ;
  assign n526 = n520 & ~n525 ;
  buffer buf_n527( .i (n526), .o (n527) );
  assign n529 = ~n480 & n527 ;
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n528( .i (n527), .o (n528) );
  assign n531 = n481 & ~n528 ;
  assign n532 = n530 | n531 ;
  buffer buf_n533( .i (n532), .o (n533) );
  assign n535 = n477 | n533 ;
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n534( .i (n533), .o (n534) );
  assign n541 = n478 & n534 ;
  assign n542 = n536 & ~n541 ;
  buffer buf_n543( .i (n542), .o (n543) );
  assign n545 = ~n474 & n543 ;
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n544( .i (n543), .o (n544) );
  assign n547 = n475 & ~n544 ;
  assign n548 = n546 | n547 ;
  buffer buf_n549( .i (n548), .o (n549) );
  assign n551 = n471 | n549 ;
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n550( .i (n549), .o (n550) );
  assign n557 = n472 & n550 ;
  assign n558 = n552 & ~n557 ;
  buffer buf_n559( .i (n558), .o (n559) );
  assign n561 = ~n468 & n559 ;
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n560( .i (n559), .o (n560) );
  assign n563 = n469 & ~n560 ;
  assign n564 = n562 | n563 ;
  buffer buf_n565( .i (n564), .o (n565) );
  assign n567 = n465 | n565 ;
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n566( .i (n565), .o (n566) );
  assign n573 = n466 & n566 ;
  assign n574 = n568 & ~n573 ;
  buffer buf_n575( .i (n574), .o (n575) );
  assign n579 = ~n460 & n575 ;
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  assign n583 = n463 & ~n578 ;
  assign n584 = n582 | n583 ;
  buffer buf_n585( .i (n584), .o (n585) );
  assign n587 = n457 | n585 ;
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n586( .i (n585), .o (n586) );
  assign n593 = n458 & n586 ;
  assign n594 = n588 & ~n593 ;
  buffer buf_n595( .i (n594), .o (n595) );
  assign n597 = ~n454 & n595 ;
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n596( .i (n595), .o (n596) );
  assign n599 = n455 & ~n596 ;
  assign n600 = n598 | n599 ;
  assign n601 = N1 & N409 ;
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  assign n604 = n592 & ~n598 ;
  buffer buf_n605( .i (n604), .o (n605) );
  assign n607 = N18 & N392 ;
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  assign n612 = n572 & ~n580 ;
  buffer buf_n613( .i (n612), .o (n613) );
  assign n615 = N35 & N375 ;
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  assign n618 = n556 & ~n562 ;
  buffer buf_n619( .i (n618), .o (n619) );
  assign n621 = N358 & N52 ;
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  assign n624 = n540 & ~n546 ;
  buffer buf_n625( .i (n624), .o (n625) );
  assign n627 = N341 & N69 ;
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  assign n630 = n524 & ~n530 ;
  buffer buf_n631( .i (n630), .o (n631) );
  assign n633 = N324 & N86 ;
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  assign n636 = n508 & ~n514 ;
  buffer buf_n637( .i (n636), .o (n637) );
  assign n639 = N103 & N307 ;
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  assign n642 = N137 & N290 ;
  buffer buf_n643( .i (n642), .o (n643) );
  assign n645 = n497 & n643 ;
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n490( .i (n489), .o (n490) );
  assign n650 = N137 & N273 ;
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  assign n653 = n490 | n652 ;
  assign n654 = ~n646 & n653 ;
  buffer buf_n655( .i (n654), .o (n655) );
  assign n657 = n494 | n655 ;
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n656( .i (n655), .o (n656) );
  assign n663 = n495 & n656 ;
  assign n664 = n658 & ~n663 ;
  buffer buf_n665( .i (n664), .o (n665) );
  assign n667 = ~n640 & n665 ;
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n666( .i (n665), .o (n666) );
  assign n669 = n641 & ~n666 ;
  assign n670 = n668 | n669 ;
  buffer buf_n671( .i (n670), .o (n671) );
  assign n673 = n637 | n671 ;
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n672( .i (n671), .o (n672) );
  assign n679 = n638 & n672 ;
  assign n680 = n674 & ~n679 ;
  buffer buf_n681( .i (n680), .o (n681) );
  assign n683 = ~n634 & n681 ;
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n682( .i (n681), .o (n682) );
  assign n685 = n635 & ~n682 ;
  assign n686 = n684 | n685 ;
  buffer buf_n687( .i (n686), .o (n687) );
  assign n689 = n631 | n687 ;
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n688( .i (n687), .o (n688) );
  assign n695 = n632 & n688 ;
  assign n696 = n690 & ~n695 ;
  buffer buf_n697( .i (n696), .o (n697) );
  assign n699 = ~n628 & n697 ;
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n698( .i (n697), .o (n698) );
  assign n701 = n629 & ~n698 ;
  assign n702 = n700 | n701 ;
  buffer buf_n703( .i (n702), .o (n703) );
  assign n705 = n625 | n703 ;
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n704( .i (n703), .o (n704) );
  assign n711 = n626 & n704 ;
  assign n712 = n706 & ~n711 ;
  buffer buf_n713( .i (n712), .o (n713) );
  assign n715 = ~n622 & n713 ;
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n714( .i (n713), .o (n714) );
  assign n717 = n623 & ~n714 ;
  assign n718 = n716 | n717 ;
  buffer buf_n719( .i (n718), .o (n719) );
  assign n721 = n619 | n719 ;
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n720( .i (n719), .o (n720) );
  assign n727 = n620 & n720 ;
  assign n728 = n722 & ~n727 ;
  buffer buf_n729( .i (n728), .o (n729) );
  assign n731 = ~n616 & n729 ;
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n730( .i (n729), .o (n730) );
  assign n733 = n617 & ~n730 ;
  assign n734 = n732 | n733 ;
  buffer buf_n735( .i (n734), .o (n735) );
  assign n737 = n613 | n735 ;
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n736( .i (n735), .o (n736) );
  assign n743 = n614 & n736 ;
  assign n744 = n738 & ~n743 ;
  buffer buf_n745( .i (n744), .o (n745) );
  assign n749 = ~n608 & n745 ;
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  assign n753 = n611 & ~n748 ;
  assign n754 = n752 | n753 ;
  buffer buf_n755( .i (n754), .o (n755) );
  assign n757 = n605 | n755 ;
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n756( .i (n755), .o (n756) );
  assign n763 = n606 & n756 ;
  assign n764 = n758 & ~n763 ;
  buffer buf_n765( .i (n764), .o (n765) );
  assign n767 = ~n602 & n765 ;
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n766( .i (n765), .o (n766) );
  assign n769 = n603 & ~n766 ;
  assign n770 = n768 | n769 ;
  assign n771 = N1 & N426 ;
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  assign n774 = n762 & ~n768 ;
  buffer buf_n775( .i (n774), .o (n775) );
  assign n777 = N18 & N409 ;
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  assign n782 = n742 & ~n750 ;
  buffer buf_n783( .i (n782), .o (n783) );
  assign n785 = N35 & N392 ;
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  assign n788 = n726 & ~n732 ;
  buffer buf_n789( .i (n788), .o (n789) );
  assign n791 = N375 & N52 ;
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  assign n794 = n710 & ~n716 ;
  buffer buf_n795( .i (n794), .o (n795) );
  assign n797 = N358 & N69 ;
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  assign n800 = n694 & ~n700 ;
  buffer buf_n801( .i (n800), .o (n801) );
  assign n803 = N341 & N86 ;
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  assign n806 = n678 & ~n684 ;
  buffer buf_n807( .i (n806), .o (n807) );
  assign n809 = N103 & N324 ;
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  assign n812 = n662 & ~n668 ;
  buffer buf_n813( .i (n812), .o (n813) );
  assign n815 = N120 & N307 ;
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  assign n818 = N154 & N290 ;
  buffer buf_n819( .i (n818), .o (n819) );
  assign n821 = n651 & n819 ;
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n644( .i (n643), .o (n644) );
  assign n826 = N154 & N273 ;
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  assign n829 = n644 | n828 ;
  assign n830 = ~n822 & n829 ;
  buffer buf_n831( .i (n830), .o (n831) );
  assign n833 = n648 | n831 ;
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n832( .i (n831), .o (n832) );
  assign n839 = n649 & n832 ;
  assign n840 = n834 & ~n839 ;
  buffer buf_n841( .i (n840), .o (n841) );
  assign n843 = ~n816 & n841 ;
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n842( .i (n841), .o (n842) );
  assign n845 = n817 & ~n842 ;
  assign n846 = n844 | n845 ;
  buffer buf_n847( .i (n846), .o (n847) );
  assign n849 = n813 | n847 ;
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n848( .i (n847), .o (n848) );
  assign n855 = n814 & n848 ;
  assign n856 = n850 & ~n855 ;
  buffer buf_n857( .i (n856), .o (n857) );
  assign n859 = ~n810 & n857 ;
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n858( .i (n857), .o (n858) );
  assign n861 = n811 & ~n858 ;
  assign n862 = n860 | n861 ;
  buffer buf_n863( .i (n862), .o (n863) );
  assign n865 = n807 | n863 ;
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n864( .i (n863), .o (n864) );
  assign n871 = n808 & n864 ;
  assign n872 = n866 & ~n871 ;
  buffer buf_n873( .i (n872), .o (n873) );
  assign n875 = ~n804 & n873 ;
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n874( .i (n873), .o (n874) );
  assign n877 = n805 & ~n874 ;
  assign n878 = n876 | n877 ;
  buffer buf_n879( .i (n878), .o (n879) );
  assign n881 = n801 | n879 ;
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n880( .i (n879), .o (n880) );
  assign n887 = n802 & n880 ;
  assign n888 = n882 & ~n887 ;
  buffer buf_n889( .i (n888), .o (n889) );
  assign n891 = ~n798 & n889 ;
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n890( .i (n889), .o (n890) );
  assign n893 = n799 & ~n890 ;
  assign n894 = n892 | n893 ;
  buffer buf_n895( .i (n894), .o (n895) );
  assign n897 = n795 | n895 ;
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n896( .i (n895), .o (n896) );
  assign n903 = n796 & n896 ;
  assign n904 = n898 & ~n903 ;
  buffer buf_n905( .i (n904), .o (n905) );
  assign n907 = ~n792 & n905 ;
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n906( .i (n905), .o (n906) );
  assign n909 = n793 & ~n906 ;
  assign n910 = n908 | n909 ;
  buffer buf_n911( .i (n910), .o (n911) );
  assign n913 = n789 | n911 ;
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n912( .i (n911), .o (n912) );
  assign n919 = n790 & n912 ;
  assign n920 = n914 & ~n919 ;
  buffer buf_n921( .i (n920), .o (n921) );
  assign n923 = ~n786 & n921 ;
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n922( .i (n921), .o (n922) );
  assign n925 = n787 & ~n922 ;
  assign n926 = n924 | n925 ;
  buffer buf_n927( .i (n926), .o (n927) );
  assign n929 = n783 | n927 ;
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n928( .i (n927), .o (n928) );
  assign n935 = n784 & n928 ;
  assign n936 = n930 & ~n935 ;
  buffer buf_n937( .i (n936), .o (n937) );
  assign n941 = ~n778 & n937 ;
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  assign n945 = n781 & ~n940 ;
  assign n946 = n944 | n945 ;
  buffer buf_n947( .i (n946), .o (n947) );
  assign n949 = n775 | n947 ;
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n948( .i (n947), .o (n948) );
  assign n955 = n776 & n948 ;
  assign n956 = n950 & ~n955 ;
  buffer buf_n957( .i (n956), .o (n957) );
  assign n959 = ~n772 & n957 ;
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n958( .i (n957), .o (n958) );
  assign n961 = n773 & ~n958 ;
  assign n962 = n960 | n961 ;
  assign n963 = N1 & N443 ;
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  assign n966 = n954 & ~n960 ;
  buffer buf_n967( .i (n966), .o (n967) );
  assign n969 = N18 & N426 ;
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  assign n974 = n934 & ~n942 ;
  buffer buf_n975( .i (n974), .o (n975) );
  assign n977 = N35 & N409 ;
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  assign n980 = n918 & ~n924 ;
  buffer buf_n981( .i (n980), .o (n981) );
  assign n983 = N392 & N52 ;
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  assign n986 = n902 & ~n908 ;
  buffer buf_n987( .i (n986), .o (n987) );
  assign n989 = N375 & N69 ;
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  assign n992 = n886 & ~n892 ;
  buffer buf_n993( .i (n992), .o (n993) );
  assign n995 = N358 & N86 ;
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  assign n998 = n870 & ~n876 ;
  buffer buf_n999( .i (n998), .o (n999) );
  assign n1001 = N103 & N341 ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  assign n1004 = n854 & ~n860 ;
  buffer buf_n1005( .i (n1004), .o (n1005) );
  assign n1007 = N120 & N324 ;
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  assign n1010 = n838 & ~n844 ;
  buffer buf_n1011( .i (n1010), .o (n1011) );
  assign n1013 = N137 & N307 ;
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  assign n1016 = N171 & N290 ;
  buffer buf_n1017( .i (n1016), .o (n1017) );
  assign n1019 = n827 & n1017 ;
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n820( .i (n819), .o (n820) );
  assign n1024 = N171 & N273 ;
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  assign n1027 = n820 | n1026 ;
  assign n1028 = ~n1020 & n1027 ;
  buffer buf_n1029( .i (n1028), .o (n1029) );
  assign n1031 = n824 | n1029 ;
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  assign n1037 = n825 & n1030 ;
  assign n1038 = n1032 & ~n1037 ;
  buffer buf_n1039( .i (n1038), .o (n1039) );
  assign n1041 = ~n1014 & n1039 ;
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  assign n1043 = n1015 & ~n1040 ;
  assign n1044 = n1042 | n1043 ;
  buffer buf_n1045( .i (n1044), .o (n1045) );
  assign n1047 = n1011 | n1045 ;
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  assign n1053 = n1012 & n1046 ;
  assign n1054 = n1048 & ~n1053 ;
  buffer buf_n1055( .i (n1054), .o (n1055) );
  assign n1057 = ~n1008 & n1055 ;
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  assign n1059 = n1009 & ~n1056 ;
  assign n1060 = n1058 | n1059 ;
  buffer buf_n1061( .i (n1060), .o (n1061) );
  assign n1063 = n1005 | n1061 ;
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  assign n1069 = n1006 & n1062 ;
  assign n1070 = n1064 & ~n1069 ;
  buffer buf_n1071( .i (n1070), .o (n1071) );
  assign n1073 = ~n1002 & n1071 ;
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  assign n1075 = n1003 & ~n1072 ;
  assign n1076 = n1074 | n1075 ;
  buffer buf_n1077( .i (n1076), .o (n1077) );
  assign n1079 = n999 | n1077 ;
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  assign n1085 = n1000 & n1078 ;
  assign n1086 = n1080 & ~n1085 ;
  buffer buf_n1087( .i (n1086), .o (n1087) );
  assign n1089 = ~n996 & n1087 ;
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  assign n1091 = n997 & ~n1088 ;
  assign n1092 = n1090 | n1091 ;
  buffer buf_n1093( .i (n1092), .o (n1093) );
  assign n1095 = n993 | n1093 ;
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  assign n1101 = n994 & n1094 ;
  assign n1102 = n1096 & ~n1101 ;
  buffer buf_n1103( .i (n1102), .o (n1103) );
  assign n1105 = ~n990 & n1103 ;
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  assign n1107 = n991 & ~n1104 ;
  assign n1108 = n1106 | n1107 ;
  buffer buf_n1109( .i (n1108), .o (n1109) );
  assign n1111 = n987 | n1109 ;
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  assign n1117 = n988 & n1110 ;
  assign n1118 = n1112 & ~n1117 ;
  buffer buf_n1119( .i (n1118), .o (n1119) );
  assign n1121 = ~n984 & n1119 ;
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  assign n1123 = n985 & ~n1120 ;
  assign n1124 = n1122 | n1123 ;
  buffer buf_n1125( .i (n1124), .o (n1125) );
  assign n1127 = n981 | n1125 ;
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  assign n1133 = n982 & n1126 ;
  assign n1134 = n1128 & ~n1133 ;
  buffer buf_n1135( .i (n1134), .o (n1135) );
  assign n1137 = ~n978 & n1135 ;
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  assign n1139 = n979 & ~n1136 ;
  assign n1140 = n1138 | n1139 ;
  buffer buf_n1141( .i (n1140), .o (n1141) );
  assign n1143 = n975 | n1141 ;
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  assign n1149 = n976 & n1142 ;
  assign n1150 = n1144 & ~n1149 ;
  buffer buf_n1151( .i (n1150), .o (n1151) );
  assign n1155 = ~n970 & n1151 ;
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  assign n1159 = n973 & ~n1154 ;
  assign n1160 = n1158 | n1159 ;
  buffer buf_n1161( .i (n1160), .o (n1161) );
  assign n1163 = n967 | n1161 ;
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  assign n1169 = n968 & n1162 ;
  assign n1170 = n1164 & ~n1169 ;
  buffer buf_n1171( .i (n1170), .o (n1171) );
  assign n1173 = ~n964 & n1171 ;
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  assign n1175 = n965 & ~n1172 ;
  assign n1176 = n1174 | n1175 ;
  assign n1177 = N1 & N460 ;
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  assign n1180 = n1168 & ~n1174 ;
  buffer buf_n1181( .i (n1180), .o (n1181) );
  assign n1183 = N18 & N443 ;
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  assign n1188 = n1148 & ~n1156 ;
  buffer buf_n1189( .i (n1188), .o (n1189) );
  assign n1191 = N35 & N426 ;
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  assign n1194 = n1132 & ~n1138 ;
  buffer buf_n1195( .i (n1194), .o (n1195) );
  assign n1197 = N409 & N52 ;
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  assign n1200 = n1116 & ~n1122 ;
  buffer buf_n1201( .i (n1200), .o (n1201) );
  assign n1203 = N392 & N69 ;
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  assign n1206 = n1100 & ~n1106 ;
  buffer buf_n1207( .i (n1206), .o (n1207) );
  assign n1209 = N375 & N86 ;
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  assign n1212 = n1084 & ~n1090 ;
  buffer buf_n1213( .i (n1212), .o (n1213) );
  assign n1215 = N103 & N358 ;
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  assign n1218 = n1068 & ~n1074 ;
  buffer buf_n1219( .i (n1218), .o (n1219) );
  assign n1221 = N120 & N341 ;
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  assign n1224 = n1052 & ~n1058 ;
  buffer buf_n1225( .i (n1224), .o (n1225) );
  assign n1227 = N137 & N324 ;
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  assign n1230 = n1036 & ~n1042 ;
  buffer buf_n1231( .i (n1230), .o (n1231) );
  assign n1233 = N154 & N307 ;
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  assign n1236 = N188 & N290 ;
  buffer buf_n1237( .i (n1236), .o (n1237) );
  assign n1239 = n1025 & n1237 ;
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  assign n1244 = N188 & N273 ;
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  assign n1247 = n1018 | n1246 ;
  assign n1248 = ~n1240 & n1247 ;
  buffer buf_n1249( .i (n1248), .o (n1249) );
  assign n1251 = n1022 | n1249 ;
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  assign n1257 = n1023 & n1250 ;
  assign n1258 = n1252 & ~n1257 ;
  buffer buf_n1259( .i (n1258), .o (n1259) );
  assign n1261 = ~n1234 & n1259 ;
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  assign n1263 = n1235 & ~n1260 ;
  assign n1264 = n1262 | n1263 ;
  buffer buf_n1265( .i (n1264), .o (n1265) );
  assign n1267 = n1231 | n1265 ;
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  assign n1273 = n1232 & n1266 ;
  assign n1274 = n1268 & ~n1273 ;
  buffer buf_n1275( .i (n1274), .o (n1275) );
  assign n1277 = ~n1228 & n1275 ;
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  assign n1279 = n1229 & ~n1276 ;
  assign n1280 = n1278 | n1279 ;
  buffer buf_n1281( .i (n1280), .o (n1281) );
  assign n1283 = n1225 | n1281 ;
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  assign n1289 = n1226 & n1282 ;
  assign n1290 = n1284 & ~n1289 ;
  buffer buf_n1291( .i (n1290), .o (n1291) );
  assign n1293 = ~n1222 & n1291 ;
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  assign n1295 = n1223 & ~n1292 ;
  assign n1296 = n1294 | n1295 ;
  buffer buf_n1297( .i (n1296), .o (n1297) );
  assign n1299 = n1219 | n1297 ;
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  assign n1305 = n1220 & n1298 ;
  assign n1306 = n1300 & ~n1305 ;
  buffer buf_n1307( .i (n1306), .o (n1307) );
  assign n1309 = ~n1216 & n1307 ;
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  assign n1311 = n1217 & ~n1308 ;
  assign n1312 = n1310 | n1311 ;
  buffer buf_n1313( .i (n1312), .o (n1313) );
  assign n1315 = n1213 | n1313 ;
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  assign n1321 = n1214 & n1314 ;
  assign n1322 = n1316 & ~n1321 ;
  buffer buf_n1323( .i (n1322), .o (n1323) );
  assign n1325 = ~n1210 & n1323 ;
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  assign n1327 = n1211 & ~n1324 ;
  assign n1328 = n1326 | n1327 ;
  buffer buf_n1329( .i (n1328), .o (n1329) );
  assign n1331 = n1207 | n1329 ;
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  assign n1337 = n1208 & n1330 ;
  assign n1338 = n1332 & ~n1337 ;
  buffer buf_n1339( .i (n1338), .o (n1339) );
  assign n1341 = ~n1204 & n1339 ;
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  assign n1343 = n1205 & ~n1340 ;
  assign n1344 = n1342 | n1343 ;
  buffer buf_n1345( .i (n1344), .o (n1345) );
  assign n1347 = n1201 | n1345 ;
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  assign n1353 = n1202 & n1346 ;
  assign n1354 = n1348 & ~n1353 ;
  buffer buf_n1355( .i (n1354), .o (n1355) );
  assign n1357 = ~n1198 & n1355 ;
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  assign n1359 = n1199 & ~n1356 ;
  assign n1360 = n1358 | n1359 ;
  buffer buf_n1361( .i (n1360), .o (n1361) );
  assign n1363 = n1195 | n1361 ;
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  assign n1369 = n1196 & n1362 ;
  assign n1370 = n1364 & ~n1369 ;
  buffer buf_n1371( .i (n1370), .o (n1371) );
  assign n1373 = ~n1192 & n1371 ;
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  assign n1375 = n1193 & ~n1372 ;
  assign n1376 = n1374 | n1375 ;
  buffer buf_n1377( .i (n1376), .o (n1377) );
  assign n1379 = n1189 | n1377 ;
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  assign n1385 = n1190 & n1378 ;
  assign n1386 = n1380 & ~n1385 ;
  buffer buf_n1387( .i (n1386), .o (n1387) );
  assign n1391 = ~n1184 & n1387 ;
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  assign n1395 = n1187 & ~n1390 ;
  assign n1396 = n1394 | n1395 ;
  buffer buf_n1397( .i (n1396), .o (n1397) );
  assign n1399 = n1181 | n1397 ;
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  assign n1405 = n1182 & n1398 ;
  assign n1406 = n1400 & ~n1405 ;
  buffer buf_n1407( .i (n1406), .o (n1407) );
  assign n1409 = ~n1178 & n1407 ;
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  assign n1411 = n1179 & ~n1408 ;
  assign n1412 = n1410 | n1411 ;
  assign n1413 = N1 & N477 ;
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  assign n1416 = n1404 & ~n1410 ;
  buffer buf_n1417( .i (n1416), .o (n1417) );
  assign n1419 = N18 & N460 ;
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  assign n1424 = n1384 & ~n1392 ;
  buffer buf_n1425( .i (n1424), .o (n1425) );
  assign n1427 = N35 & N443 ;
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  assign n1430 = n1368 & ~n1374 ;
  buffer buf_n1431( .i (n1430), .o (n1431) );
  assign n1433 = N426 & N52 ;
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  assign n1436 = n1352 & ~n1358 ;
  buffer buf_n1437( .i (n1436), .o (n1437) );
  assign n1439 = N409 & N69 ;
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  assign n1442 = n1336 & ~n1342 ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  assign n1445 = N392 & N86 ;
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  assign n1448 = n1320 & ~n1326 ;
  buffer buf_n1449( .i (n1448), .o (n1449) );
  assign n1451 = N103 & N375 ;
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  assign n1454 = n1304 & ~n1310 ;
  buffer buf_n1455( .i (n1454), .o (n1455) );
  assign n1457 = N120 & N358 ;
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  assign n1460 = n1288 & ~n1294 ;
  buffer buf_n1461( .i (n1460), .o (n1461) );
  assign n1463 = N137 & N341 ;
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  assign n1466 = n1272 & ~n1278 ;
  buffer buf_n1467( .i (n1466), .o (n1467) );
  assign n1469 = N154 & N324 ;
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  assign n1472 = n1256 & ~n1262 ;
  buffer buf_n1473( .i (n1472), .o (n1473) );
  assign n1475 = N171 & N307 ;
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  assign n1478 = N205 & N290 ;
  buffer buf_n1479( .i (n1478), .o (n1479) );
  assign n1481 = n1245 & n1479 ;
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  assign n1486 = N205 & N273 ;
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n1488( .i (n1487), .o (n1488) );
  assign n1489 = n1238 | n1488 ;
  assign n1490 = ~n1482 & n1489 ;
  buffer buf_n1491( .i (n1490), .o (n1491) );
  assign n1493 = n1242 | n1491 ;
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  assign n1499 = n1243 & n1492 ;
  assign n1500 = n1494 & ~n1499 ;
  buffer buf_n1501( .i (n1500), .o (n1501) );
  assign n1503 = ~n1476 & n1501 ;
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  assign n1505 = n1477 & ~n1502 ;
  assign n1506 = n1504 | n1505 ;
  buffer buf_n1507( .i (n1506), .o (n1507) );
  assign n1509 = n1473 | n1507 ;
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  assign n1515 = n1474 & n1508 ;
  assign n1516 = n1510 & ~n1515 ;
  buffer buf_n1517( .i (n1516), .o (n1517) );
  assign n1519 = ~n1470 & n1517 ;
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1518( .i (n1517), .o (n1518) );
  assign n1521 = n1471 & ~n1518 ;
  assign n1522 = n1520 | n1521 ;
  buffer buf_n1523( .i (n1522), .o (n1523) );
  assign n1525 = n1467 | n1523 ;
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  assign n1531 = n1468 & n1524 ;
  assign n1532 = n1526 & ~n1531 ;
  buffer buf_n1533( .i (n1532), .o (n1533) );
  assign n1535 = ~n1464 & n1533 ;
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1534( .i (n1533), .o (n1534) );
  assign n1537 = n1465 & ~n1534 ;
  assign n1538 = n1536 | n1537 ;
  buffer buf_n1539( .i (n1538), .o (n1539) );
  assign n1541 = n1461 | n1539 ;
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  assign n1547 = n1462 & n1540 ;
  assign n1548 = n1542 & ~n1547 ;
  buffer buf_n1549( .i (n1548), .o (n1549) );
  assign n1551 = ~n1458 & n1549 ;
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  assign n1553 = n1459 & ~n1550 ;
  assign n1554 = n1552 | n1553 ;
  buffer buf_n1555( .i (n1554), .o (n1555) );
  assign n1557 = n1455 | n1555 ;
  buffer buf_n1558( .i (n1557), .o (n1558) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  buffer buf_n1556( .i (n1555), .o (n1556) );
  assign n1563 = n1456 & n1556 ;
  assign n1564 = n1558 & ~n1563 ;
  buffer buf_n1565( .i (n1564), .o (n1565) );
  assign n1567 = ~n1452 & n1565 ;
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  assign n1569 = n1453 & ~n1566 ;
  assign n1570 = n1568 | n1569 ;
  buffer buf_n1571( .i (n1570), .o (n1571) );
  assign n1573 = n1449 | n1571 ;
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  assign n1579 = n1450 & n1572 ;
  assign n1580 = n1574 & ~n1579 ;
  buffer buf_n1581( .i (n1580), .o (n1581) );
  assign n1583 = ~n1446 & n1581 ;
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  assign n1585 = n1447 & ~n1582 ;
  assign n1586 = n1584 | n1585 ;
  buffer buf_n1587( .i (n1586), .o (n1587) );
  assign n1589 = n1443 | n1587 ;
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  assign n1595 = n1444 & n1588 ;
  assign n1596 = n1590 & ~n1595 ;
  buffer buf_n1597( .i (n1596), .o (n1597) );
  assign n1599 = ~n1440 & n1597 ;
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  assign n1601 = n1441 & ~n1598 ;
  assign n1602 = n1600 | n1601 ;
  buffer buf_n1603( .i (n1602), .o (n1603) );
  assign n1605 = n1437 | n1603 ;
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  assign n1611 = n1438 & n1604 ;
  assign n1612 = n1606 & ~n1611 ;
  buffer buf_n1613( .i (n1612), .o (n1613) );
  assign n1615 = ~n1434 & n1613 ;
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  assign n1617 = n1435 & ~n1614 ;
  assign n1618 = n1616 | n1617 ;
  buffer buf_n1619( .i (n1618), .o (n1619) );
  assign n1621 = n1431 | n1619 ;
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1620( .i (n1619), .o (n1620) );
  assign n1627 = n1432 & n1620 ;
  assign n1628 = n1622 & ~n1627 ;
  buffer buf_n1629( .i (n1628), .o (n1629) );
  assign n1631 = ~n1428 & n1629 ;
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  assign n1633 = n1429 & ~n1630 ;
  assign n1634 = n1632 | n1633 ;
  buffer buf_n1635( .i (n1634), .o (n1635) );
  assign n1637 = n1425 | n1635 ;
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1636( .i (n1635), .o (n1636) );
  assign n1643 = n1426 & n1636 ;
  assign n1644 = n1638 & ~n1643 ;
  buffer buf_n1645( .i (n1644), .o (n1645) );
  assign n1649 = ~n1420 & n1645 ;
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  assign n1653 = n1423 & ~n1648 ;
  assign n1654 = n1652 | n1653 ;
  buffer buf_n1655( .i (n1654), .o (n1655) );
  assign n1657 = n1417 | n1655 ;
  buffer buf_n1658( .i (n1657), .o (n1658) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  assign n1663 = n1418 & n1656 ;
  assign n1664 = n1658 & ~n1663 ;
  buffer buf_n1665( .i (n1664), .o (n1665) );
  assign n1667 = ~n1414 & n1665 ;
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  assign n1669 = n1415 & ~n1666 ;
  assign n1670 = n1668 | n1669 ;
  assign n1671 = N1 & N494 ;
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  assign n1674 = n1662 & ~n1668 ;
  buffer buf_n1675( .i (n1674), .o (n1675) );
  assign n1677 = N18 & N477 ;
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  assign n1682 = n1642 & ~n1650 ;
  buffer buf_n1683( .i (n1682), .o (n1683) );
  assign n1685 = N35 & N460 ;
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  assign n1688 = n1626 & ~n1632 ;
  buffer buf_n1689( .i (n1688), .o (n1689) );
  assign n1691 = N443 & N52 ;
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  assign n1694 = n1610 & ~n1616 ;
  buffer buf_n1695( .i (n1694), .o (n1695) );
  assign n1697 = N426 & N69 ;
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  assign n1700 = n1594 & ~n1600 ;
  buffer buf_n1701( .i (n1700), .o (n1701) );
  assign n1703 = N409 & N86 ;
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  assign n1706 = n1578 & ~n1584 ;
  buffer buf_n1707( .i (n1706), .o (n1707) );
  assign n1709 = N103 & N392 ;
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  assign n1712 = n1562 & ~n1568 ;
  buffer buf_n1713( .i (n1712), .o (n1713) );
  assign n1715 = N120 & N375 ;
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  assign n1718 = n1546 & ~n1552 ;
  buffer buf_n1719( .i (n1718), .o (n1719) );
  assign n1721 = N137 & N358 ;
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  assign n1724 = n1530 & ~n1536 ;
  buffer buf_n1725( .i (n1724), .o (n1725) );
  assign n1727 = N154 & N341 ;
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  assign n1730 = n1514 & ~n1520 ;
  buffer buf_n1731( .i (n1730), .o (n1731) );
  assign n1733 = N171 & N324 ;
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  assign n1736 = n1498 & ~n1504 ;
  buffer buf_n1737( .i (n1736), .o (n1737) );
  assign n1739 = N188 & N307 ;
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  assign n1742 = N222 & N290 ;
  buffer buf_n1743( .i (n1742), .o (n1743) );
  assign n1745 = n1487 & n1743 ;
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  assign n1750 = N222 & N273 ;
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  assign n1753 = n1480 | n1752 ;
  assign n1754 = ~n1746 & n1753 ;
  buffer buf_n1755( .i (n1754), .o (n1755) );
  assign n1757 = n1484 | n1755 ;
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  assign n1763 = n1485 & n1756 ;
  assign n1764 = n1758 & ~n1763 ;
  buffer buf_n1765( .i (n1764), .o (n1765) );
  assign n1767 = ~n1740 & n1765 ;
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  assign n1769 = n1741 & ~n1766 ;
  assign n1770 = n1768 | n1769 ;
  buffer buf_n1771( .i (n1770), .o (n1771) );
  assign n1773 = n1737 | n1771 ;
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  assign n1779 = n1738 & n1772 ;
  assign n1780 = n1774 & ~n1779 ;
  buffer buf_n1781( .i (n1780), .o (n1781) );
  assign n1783 = ~n1734 & n1781 ;
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  assign n1785 = n1735 & ~n1782 ;
  assign n1786 = n1784 | n1785 ;
  buffer buf_n1787( .i (n1786), .o (n1787) );
  assign n1789 = n1731 | n1787 ;
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  assign n1795 = n1732 & n1788 ;
  assign n1796 = n1790 & ~n1795 ;
  buffer buf_n1797( .i (n1796), .o (n1797) );
  assign n1799 = ~n1728 & n1797 ;
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  assign n1801 = n1729 & ~n1798 ;
  assign n1802 = n1800 | n1801 ;
  buffer buf_n1803( .i (n1802), .o (n1803) );
  assign n1805 = n1725 | n1803 ;
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  assign n1811 = n1726 & n1804 ;
  assign n1812 = n1806 & ~n1811 ;
  buffer buf_n1813( .i (n1812), .o (n1813) );
  assign n1815 = ~n1722 & n1813 ;
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1814( .i (n1813), .o (n1814) );
  assign n1817 = n1723 & ~n1814 ;
  assign n1818 = n1816 | n1817 ;
  buffer buf_n1819( .i (n1818), .o (n1819) );
  assign n1821 = n1719 | n1819 ;
  buffer buf_n1822( .i (n1821), .o (n1822) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  assign n1827 = n1720 & n1820 ;
  assign n1828 = n1822 & ~n1827 ;
  buffer buf_n1829( .i (n1828), .o (n1829) );
  assign n1831 = ~n1716 & n1829 ;
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  assign n1833 = n1717 & ~n1830 ;
  assign n1834 = n1832 | n1833 ;
  buffer buf_n1835( .i (n1834), .o (n1835) );
  assign n1837 = n1713 | n1835 ;
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  assign n1843 = n1714 & n1836 ;
  assign n1844 = n1838 & ~n1843 ;
  buffer buf_n1845( .i (n1844), .o (n1845) );
  assign n1847 = ~n1710 & n1845 ;
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1846( .i (n1845), .o (n1846) );
  assign n1849 = n1711 & ~n1846 ;
  assign n1850 = n1848 | n1849 ;
  buffer buf_n1851( .i (n1850), .o (n1851) );
  assign n1853 = n1707 | n1851 ;
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  assign n1859 = n1708 & n1852 ;
  assign n1860 = n1854 & ~n1859 ;
  buffer buf_n1861( .i (n1860), .o (n1861) );
  assign n1863 = ~n1704 & n1861 ;
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  assign n1865 = n1705 & ~n1862 ;
  assign n1866 = n1864 | n1865 ;
  buffer buf_n1867( .i (n1866), .o (n1867) );
  assign n1869 = n1701 | n1867 ;
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  assign n1875 = n1702 & n1868 ;
  assign n1876 = n1870 & ~n1875 ;
  buffer buf_n1877( .i (n1876), .o (n1877) );
  assign n1879 = ~n1698 & n1877 ;
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  assign n1881 = n1699 & ~n1878 ;
  assign n1882 = n1880 | n1881 ;
  buffer buf_n1883( .i (n1882), .o (n1883) );
  assign n1885 = n1695 | n1883 ;
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  assign n1891 = n1696 & n1884 ;
  assign n1892 = n1886 & ~n1891 ;
  buffer buf_n1893( .i (n1892), .o (n1893) );
  assign n1895 = ~n1692 & n1893 ;
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  assign n1897 = n1693 & ~n1894 ;
  assign n1898 = n1896 | n1897 ;
  buffer buf_n1899( .i (n1898), .o (n1899) );
  assign n1901 = n1689 | n1899 ;
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  assign n1907 = n1690 & n1900 ;
  assign n1908 = n1902 & ~n1907 ;
  buffer buf_n1909( .i (n1908), .o (n1909) );
  assign n1911 = ~n1686 & n1909 ;
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  assign n1913 = n1687 & ~n1910 ;
  assign n1914 = n1912 | n1913 ;
  buffer buf_n1915( .i (n1914), .o (n1915) );
  assign n1917 = n1683 | n1915 ;
  buffer buf_n1918( .i (n1917), .o (n1918) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1916( .i (n1915), .o (n1916) );
  assign n1923 = n1684 & n1916 ;
  assign n1924 = n1918 & ~n1923 ;
  buffer buf_n1925( .i (n1924), .o (n1925) );
  assign n1929 = ~n1678 & n1925 ;
  buffer buf_n1930( .i (n1929), .o (n1930) );
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  assign n1933 = n1681 & ~n1928 ;
  assign n1934 = n1932 | n1933 ;
  buffer buf_n1935( .i (n1934), .o (n1935) );
  assign n1937 = n1675 | n1935 ;
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  assign n1943 = n1676 & n1936 ;
  assign n1944 = n1938 & ~n1943 ;
  buffer buf_n1945( .i (n1944), .o (n1945) );
  assign n1947 = ~n1672 & n1945 ;
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  assign n1949 = n1673 & ~n1946 ;
  assign n1950 = n1948 | n1949 ;
  assign n1951 = N1 & N511 ;
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  assign n1954 = n1942 & ~n1948 ;
  buffer buf_n1955( .i (n1954), .o (n1955) );
  assign n1957 = N18 & N494 ;
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1919( .i (n1918), .o (n1919) );
  buffer buf_n1920( .i (n1919), .o (n1920) );
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  assign n1962 = n1922 & ~n1930 ;
  buffer buf_n1963( .i (n1962), .o (n1963) );
  assign n1965 = N35 & N477 ;
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  assign n1968 = n1906 & ~n1912 ;
  buffer buf_n1969( .i (n1968), .o (n1969) );
  assign n1971 = N460 & N52 ;
  buffer buf_n1972( .i (n1971), .o (n1972) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n1888( .i (n1887), .o (n1888) );
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  assign n1974 = n1890 & ~n1896 ;
  buffer buf_n1975( .i (n1974), .o (n1975) );
  assign n1977 = N443 & N69 ;
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  buffer buf_n1872( .i (n1871), .o (n1872) );
  buffer buf_n1873( .i (n1872), .o (n1873) );
  buffer buf_n1874( .i (n1873), .o (n1874) );
  assign n1980 = n1874 & ~n1880 ;
  buffer buf_n1981( .i (n1980), .o (n1981) );
  assign n1983 = N426 & N86 ;
  buffer buf_n1984( .i (n1983), .o (n1984) );
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  assign n1986 = n1858 & ~n1864 ;
  buffer buf_n1987( .i (n1986), .o (n1987) );
  assign n1989 = N103 & N409 ;
  buffer buf_n1990( .i (n1989), .o (n1990) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  assign n1992 = n1842 & ~n1848 ;
  buffer buf_n1993( .i (n1992), .o (n1993) );
  assign n1995 = N120 & N392 ;
  buffer buf_n1996( .i (n1995), .o (n1996) );
  buffer buf_n1823( .i (n1822), .o (n1823) );
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1825( .i (n1824), .o (n1825) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  assign n1998 = n1826 & ~n1832 ;
  buffer buf_n1999( .i (n1998), .o (n1999) );
  assign n2001 = N137 & N375 ;
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  assign n2004 = n1810 & ~n1816 ;
  buffer buf_n2005( .i (n2004), .o (n2005) );
  assign n2007 = N154 & N358 ;
  buffer buf_n2008( .i (n2007), .o (n2008) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  assign n2010 = n1794 & ~n1800 ;
  buffer buf_n2011( .i (n2010), .o (n2011) );
  assign n2013 = N171 & N341 ;
  buffer buf_n2014( .i (n2013), .o (n2014) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  assign n2016 = n1778 & ~n1784 ;
  buffer buf_n2017( .i (n2016), .o (n2017) );
  assign n2019 = N188 & N324 ;
  buffer buf_n2020( .i (n2019), .o (n2020) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  assign n2022 = n1762 & ~n1768 ;
  buffer buf_n2023( .i (n2022), .o (n2023) );
  assign n2025 = N205 & N307 ;
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  assign n2028 = N239 & N290 ;
  buffer buf_n2029( .i (n2028), .o (n2029) );
  assign n2033 = n1751 & n2029 ;
  buffer buf_n2034( .i (n2033), .o (n2034) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  assign n2038 = N239 & N273 ;
  buffer buf_n2039( .i (n2038), .o (n2039) );
  assign n2045 = n1744 | n2039 ;
  assign n2046 = ~n2034 & n2045 ;
  buffer buf_n2047( .i (n2046), .o (n2047) );
  assign n2049 = n1748 | n2047 ;
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  assign n2055 = n1749 & n2048 ;
  assign n2056 = n2050 & ~n2055 ;
  buffer buf_n2057( .i (n2056), .o (n2057) );
  assign n2059 = ~n2026 & n2057 ;
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2058( .i (n2057), .o (n2058) );
  assign n2061 = n2027 & ~n2058 ;
  assign n2062 = n2060 | n2061 ;
  buffer buf_n2063( .i (n2062), .o (n2063) );
  assign n2065 = n2023 | n2063 ;
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2064( .i (n2063), .o (n2064) );
  assign n2071 = n2024 & n2064 ;
  assign n2072 = n2066 & ~n2071 ;
  buffer buf_n2073( .i (n2072), .o (n2073) );
  assign n2075 = ~n2020 & n2073 ;
  buffer buf_n2076( .i (n2075), .o (n2076) );
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  assign n2077 = n2021 & ~n2074 ;
  assign n2078 = n2076 | n2077 ;
  buffer buf_n2079( .i (n2078), .o (n2079) );
  assign n2081 = n2017 | n2079 ;
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n2018( .i (n2017), .o (n2018) );
  buffer buf_n2080( .i (n2079), .o (n2080) );
  assign n2087 = n2018 & n2080 ;
  assign n2088 = n2082 & ~n2087 ;
  buffer buf_n2089( .i (n2088), .o (n2089) );
  assign n2091 = ~n2014 & n2089 ;
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n2015( .i (n2014), .o (n2015) );
  buffer buf_n2090( .i (n2089), .o (n2090) );
  assign n2093 = n2015 & ~n2090 ;
  assign n2094 = n2092 | n2093 ;
  buffer buf_n2095( .i (n2094), .o (n2095) );
  assign n2097 = n2011 | n2095 ;
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n2012( .i (n2011), .o (n2012) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  assign n2103 = n2012 & n2096 ;
  assign n2104 = n2098 & ~n2103 ;
  buffer buf_n2105( .i (n2104), .o (n2105) );
  assign n2107 = ~n2008 & n2105 ;
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2009( .i (n2008), .o (n2009) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  assign n2109 = n2009 & ~n2106 ;
  assign n2110 = n2108 | n2109 ;
  buffer buf_n2111( .i (n2110), .o (n2111) );
  assign n2113 = n2005 | n2111 ;
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n2112( .i (n2111), .o (n2112) );
  assign n2119 = n2006 & n2112 ;
  assign n2120 = n2114 & ~n2119 ;
  buffer buf_n2121( .i (n2120), .o (n2121) );
  assign n2123 = ~n2002 & n2121 ;
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2122( .i (n2121), .o (n2122) );
  assign n2125 = n2003 & ~n2122 ;
  assign n2126 = n2124 | n2125 ;
  buffer buf_n2127( .i (n2126), .o (n2127) );
  assign n2129 = n1999 | n2127 ;
  buffer buf_n2130( .i (n2129), .o (n2130) );
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  assign n2135 = n2000 & n2128 ;
  assign n2136 = n2130 & ~n2135 ;
  buffer buf_n2137( .i (n2136), .o (n2137) );
  assign n2139 = ~n1996 & n2137 ;
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n1997( .i (n1996), .o (n1997) );
  buffer buf_n2138( .i (n2137), .o (n2138) );
  assign n2141 = n1997 & ~n2138 ;
  assign n2142 = n2140 | n2141 ;
  buffer buf_n2143( .i (n2142), .o (n2143) );
  assign n2145 = n1993 | n2143 ;
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n1994( .i (n1993), .o (n1994) );
  buffer buf_n2144( .i (n2143), .o (n2144) );
  assign n2151 = n1994 & n2144 ;
  assign n2152 = n2146 & ~n2151 ;
  buffer buf_n2153( .i (n2152), .o (n2153) );
  assign n2155 = ~n1990 & n2153 ;
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n1991( .i (n1990), .o (n1991) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  assign n2157 = n1991 & ~n2154 ;
  assign n2158 = n2156 | n2157 ;
  buffer buf_n2159( .i (n2158), .o (n2159) );
  assign n2161 = n1987 | n2159 ;
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n1988( .i (n1987), .o (n1988) );
  buffer buf_n2160( .i (n2159), .o (n2160) );
  assign n2167 = n1988 & n2160 ;
  assign n2168 = n2162 & ~n2167 ;
  buffer buf_n2169( .i (n2168), .o (n2169) );
  assign n2171 = ~n1984 & n2169 ;
  buffer buf_n2172( .i (n2171), .o (n2172) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  assign n2173 = n1985 & ~n2170 ;
  assign n2174 = n2172 | n2173 ;
  buffer buf_n2175( .i (n2174), .o (n2175) );
  assign n2177 = n1981 | n2175 ;
  buffer buf_n2178( .i (n2177), .o (n2178) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  assign n2183 = n1982 & n2176 ;
  assign n2184 = n2178 & ~n2183 ;
  buffer buf_n2185( .i (n2184), .o (n2185) );
  assign n2187 = ~n1978 & n2185 ;
  buffer buf_n2188( .i (n2187), .o (n2188) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  assign n2189 = n1979 & ~n2186 ;
  assign n2190 = n2188 | n2189 ;
  buffer buf_n2191( .i (n2190), .o (n2191) );
  assign n2193 = n1975 | n2191 ;
  buffer buf_n2194( .i (n2193), .o (n2194) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n2192( .i (n2191), .o (n2192) );
  assign n2199 = n1976 & n2192 ;
  assign n2200 = n2194 & ~n2199 ;
  buffer buf_n2201( .i (n2200), .o (n2201) );
  assign n2203 = ~n1972 & n2201 ;
  buffer buf_n2204( .i (n2203), .o (n2204) );
  buffer buf_n1973( .i (n1972), .o (n1973) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  assign n2205 = n1973 & ~n2202 ;
  assign n2206 = n2204 | n2205 ;
  buffer buf_n2207( .i (n2206), .o (n2207) );
  assign n2209 = n1969 | n2207 ;
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n1970( .i (n1969), .o (n1970) );
  buffer buf_n2208( .i (n2207), .o (n2208) );
  assign n2215 = n1970 & n2208 ;
  assign n2216 = n2210 & ~n2215 ;
  buffer buf_n2217( .i (n2216), .o (n2217) );
  assign n2219 = ~n1966 & n2217 ;
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n1967( .i (n1966), .o (n1967) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  assign n2221 = n1967 & ~n2218 ;
  assign n2222 = n2220 | n2221 ;
  buffer buf_n2223( .i (n2222), .o (n2223) );
  assign n2225 = n1963 | n2223 ;
  buffer buf_n2226( .i (n2225), .o (n2226) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n2224( .i (n2223), .o (n2224) );
  assign n2231 = n1964 & n2224 ;
  assign n2232 = n2226 & ~n2231 ;
  buffer buf_n2233( .i (n2232), .o (n2233) );
  assign n2237 = ~n1958 & n2233 ;
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  buffer buf_n1960( .i (n1959), .o (n1960) );
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  buffer buf_n2235( .i (n2234), .o (n2235) );
  buffer buf_n2236( .i (n2235), .o (n2236) );
  assign n2241 = n1961 & ~n2236 ;
  assign n2242 = n2240 | n2241 ;
  buffer buf_n2243( .i (n2242), .o (n2243) );
  assign n2245 = n1955 | n2243 ;
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  assign n2251 = n1956 & n2244 ;
  assign n2252 = n2246 & ~n2251 ;
  buffer buf_n2253( .i (n2252), .o (n2253) );
  assign n2255 = ~n1952 & n2253 ;
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  assign n2257 = n1953 & ~n2254 ;
  assign n2258 = n2256 | n2257 ;
  assign n2259 = N1 & N528 ;
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  buffer buf_n2250( .i (n2249), .o (n2250) );
  assign n2262 = n2250 & ~n2256 ;
  buffer buf_n2263( .i (n2262), .o (n2263) );
  assign n2265 = N18 & N511 ;
  buffer buf_n2266( .i (n2265), .o (n2266) );
  buffer buf_n2227( .i (n2226), .o (n2227) );
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  assign n2270 = n2230 & ~n2238 ;
  buffer buf_n2271( .i (n2270), .o (n2271) );
  assign n2273 = N35 & N494 ;
  buffer buf_n2274( .i (n2273), .o (n2274) );
  buffer buf_n2211( .i (n2210), .o (n2211) );
  buffer buf_n2212( .i (n2211), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  buffer buf_n2214( .i (n2213), .o (n2214) );
  assign n2276 = n2214 & ~n2220 ;
  buffer buf_n2277( .i (n2276), .o (n2277) );
  assign n2279 = N477 & N52 ;
  buffer buf_n2280( .i (n2279), .o (n2280) );
  buffer buf_n2195( .i (n2194), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  buffer buf_n2197( .i (n2196), .o (n2197) );
  buffer buf_n2198( .i (n2197), .o (n2198) );
  assign n2282 = n2198 & ~n2204 ;
  buffer buf_n2283( .i (n2282), .o (n2283) );
  assign n2285 = N460 & N69 ;
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2179( .i (n2178), .o (n2179) );
  buffer buf_n2180( .i (n2179), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  buffer buf_n2182( .i (n2181), .o (n2182) );
  assign n2288 = n2182 & ~n2188 ;
  buffer buf_n2289( .i (n2288), .o (n2289) );
  assign n2291 = N443 & N86 ;
  buffer buf_n2292( .i (n2291), .o (n2292) );
  buffer buf_n2163( .i (n2162), .o (n2163) );
  buffer buf_n2164( .i (n2163), .o (n2164) );
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n2166( .i (n2165), .o (n2166) );
  assign n2294 = n2166 & ~n2172 ;
  buffer buf_n2295( .i (n2294), .o (n2295) );
  assign n2297 = N103 & N426 ;
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n2150( .i (n2149), .o (n2150) );
  assign n2300 = n2150 & ~n2156 ;
  buffer buf_n2301( .i (n2300), .o (n2301) );
  assign n2303 = N120 & N409 ;
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2131( .i (n2130), .o (n2131) );
  buffer buf_n2132( .i (n2131), .o (n2132) );
  buffer buf_n2133( .i (n2132), .o (n2133) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  assign n2306 = n2134 & ~n2140 ;
  buffer buf_n2307( .i (n2306), .o (n2307) );
  assign n2309 = N137 & N392 ;
  buffer buf_n2310( .i (n2309), .o (n2310) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  assign n2312 = n2118 & ~n2124 ;
  buffer buf_n2313( .i (n2312), .o (n2313) );
  assign n2315 = N154 & N375 ;
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2099( .i (n2098), .o (n2099) );
  buffer buf_n2100( .i (n2099), .o (n2100) );
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n2102( .i (n2101), .o (n2102) );
  assign n2318 = n2102 & ~n2108 ;
  buffer buf_n2319( .i (n2318), .o (n2319) );
  assign n2321 = N171 & N358 ;
  buffer buf_n2322( .i (n2321), .o (n2322) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  assign n2324 = n2086 & ~n2092 ;
  buffer buf_n2325( .i (n2324), .o (n2325) );
  assign n2327 = N188 & N341 ;
  buffer buf_n2328( .i (n2327), .o (n2328) );
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  assign n2330 = n2070 & ~n2076 ;
  buffer buf_n2331( .i (n2330), .o (n2331) );
  assign n2333 = N205 & N324 ;
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  assign n2336 = n2054 & ~n2060 ;
  buffer buf_n2337( .i (n2336), .o (n2337) );
  assign n2339 = N222 & N307 ;
  buffer buf_n2340( .i (n2339), .o (n2340) );
  buffer buf_n2035( .i (n2034), .o (n2035) );
  buffer buf_n2036( .i (n2035), .o (n2036) );
  buffer buf_n2037( .i (n2036), .o (n2037) );
  assign n2342 = ~N256 & n2037 ;
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n2031( .i (n2030), .o (n2031) );
  buffer buf_n2032( .i (n2031), .o (n2032) );
  assign n2343 = N256 & N273 ;
  buffer buf_n2344( .i (n2343), .o (n2344) );
  assign n2345 = n2032 | n2344 ;
  assign n2346 = ~N222 & n2031 ;
  assign n2347 = n2344 & n2346 ;
  assign n2348 = n2345 & ~n2347 ;
  buffer buf_n2349( .i (n2348), .o (n2349) );
  assign n2354 = ~n2342 & n2349 ;
  buffer buf_n2355( .i (n2354), .o (n2355) );
  assign n2357 = ~n2340 & n2355 ;
  buffer buf_n2358( .i (n2357), .o (n2358) );
  buffer buf_n2341( .i (n2340), .o (n2341) );
  buffer buf_n2356( .i (n2355), .o (n2356) );
  assign n2359 = n2341 & ~n2356 ;
  assign n2360 = n2358 | n2359 ;
  buffer buf_n2361( .i (n2360), .o (n2361) );
  assign n2363 = n2337 | n2361 ;
  buffer buf_n2364( .i (n2363), .o (n2364) );
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2362( .i (n2361), .o (n2362) );
  assign n2369 = n2338 & n2362 ;
  assign n2370 = n2364 & ~n2369 ;
  buffer buf_n2371( .i (n2370), .o (n2371) );
  assign n2373 = ~n2334 & n2371 ;
  buffer buf_n2374( .i (n2373), .o (n2374) );
  buffer buf_n2335( .i (n2334), .o (n2335) );
  buffer buf_n2372( .i (n2371), .o (n2372) );
  assign n2375 = n2335 & ~n2372 ;
  assign n2376 = n2374 | n2375 ;
  buffer buf_n2377( .i (n2376), .o (n2377) );
  assign n2379 = n2331 | n2377 ;
  buffer buf_n2380( .i (n2379), .o (n2380) );
  buffer buf_n2332( .i (n2331), .o (n2332) );
  buffer buf_n2378( .i (n2377), .o (n2378) );
  assign n2385 = n2332 & n2378 ;
  assign n2386 = n2380 & ~n2385 ;
  buffer buf_n2387( .i (n2386), .o (n2387) );
  assign n2389 = ~n2328 & n2387 ;
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2329( .i (n2328), .o (n2329) );
  buffer buf_n2388( .i (n2387), .o (n2388) );
  assign n2391 = n2329 & ~n2388 ;
  assign n2392 = n2390 | n2391 ;
  buffer buf_n2393( .i (n2392), .o (n2393) );
  assign n2395 = n2325 | n2393 ;
  buffer buf_n2396( .i (n2395), .o (n2396) );
  buffer buf_n2326( .i (n2325), .o (n2326) );
  buffer buf_n2394( .i (n2393), .o (n2394) );
  assign n2401 = n2326 & n2394 ;
  assign n2402 = n2396 & ~n2401 ;
  buffer buf_n2403( .i (n2402), .o (n2403) );
  assign n2405 = ~n2322 & n2403 ;
  buffer buf_n2406( .i (n2405), .o (n2406) );
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2404( .i (n2403), .o (n2404) );
  assign n2407 = n2323 & ~n2404 ;
  assign n2408 = n2406 | n2407 ;
  buffer buf_n2409( .i (n2408), .o (n2409) );
  assign n2411 = n2319 | n2409 ;
  buffer buf_n2412( .i (n2411), .o (n2412) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  assign n2417 = n2320 & n2410 ;
  assign n2418 = n2412 & ~n2417 ;
  buffer buf_n2419( .i (n2418), .o (n2419) );
  assign n2421 = ~n2316 & n2419 ;
  buffer buf_n2422( .i (n2421), .o (n2422) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  buffer buf_n2420( .i (n2419), .o (n2420) );
  assign n2423 = n2317 & ~n2420 ;
  assign n2424 = n2422 | n2423 ;
  buffer buf_n2425( .i (n2424), .o (n2425) );
  assign n2427 = n2313 | n2425 ;
  buffer buf_n2428( .i (n2427), .o (n2428) );
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2426( .i (n2425), .o (n2426) );
  assign n2433 = n2314 & n2426 ;
  assign n2434 = n2428 & ~n2433 ;
  buffer buf_n2435( .i (n2434), .o (n2435) );
  assign n2437 = ~n2310 & n2435 ;
  buffer buf_n2438( .i (n2437), .o (n2438) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2436( .i (n2435), .o (n2436) );
  assign n2439 = n2311 & ~n2436 ;
  assign n2440 = n2438 | n2439 ;
  buffer buf_n2441( .i (n2440), .o (n2441) );
  assign n2443 = n2307 | n2441 ;
  buffer buf_n2444( .i (n2443), .o (n2444) );
  buffer buf_n2308( .i (n2307), .o (n2308) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  assign n2449 = n2308 & n2442 ;
  assign n2450 = n2444 & ~n2449 ;
  buffer buf_n2451( .i (n2450), .o (n2451) );
  assign n2453 = ~n2304 & n2451 ;
  buffer buf_n2454( .i (n2453), .o (n2454) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2452( .i (n2451), .o (n2452) );
  assign n2455 = n2305 & ~n2452 ;
  assign n2456 = n2454 | n2455 ;
  buffer buf_n2457( .i (n2456), .o (n2457) );
  assign n2459 = n2301 | n2457 ;
  buffer buf_n2460( .i (n2459), .o (n2460) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2458( .i (n2457), .o (n2458) );
  assign n2465 = n2302 & n2458 ;
  assign n2466 = n2460 & ~n2465 ;
  buffer buf_n2467( .i (n2466), .o (n2467) );
  assign n2469 = ~n2298 & n2467 ;
  buffer buf_n2470( .i (n2469), .o (n2470) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2468( .i (n2467), .o (n2468) );
  assign n2471 = n2299 & ~n2468 ;
  assign n2472 = n2470 | n2471 ;
  buffer buf_n2473( .i (n2472), .o (n2473) );
  assign n2475 = n2295 | n2473 ;
  buffer buf_n2476( .i (n2475), .o (n2476) );
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n2474( .i (n2473), .o (n2474) );
  assign n2481 = n2296 & n2474 ;
  assign n2482 = n2476 & ~n2481 ;
  buffer buf_n2483( .i (n2482), .o (n2483) );
  assign n2485 = ~n2292 & n2483 ;
  buffer buf_n2486( .i (n2485), .o (n2486) );
  buffer buf_n2293( .i (n2292), .o (n2293) );
  buffer buf_n2484( .i (n2483), .o (n2484) );
  assign n2487 = n2293 & ~n2484 ;
  assign n2488 = n2486 | n2487 ;
  buffer buf_n2489( .i (n2488), .o (n2489) );
  assign n2491 = n2289 | n2489 ;
  buffer buf_n2492( .i (n2491), .o (n2492) );
  buffer buf_n2290( .i (n2289), .o (n2290) );
  buffer buf_n2490( .i (n2489), .o (n2490) );
  assign n2497 = n2290 & n2490 ;
  assign n2498 = n2492 & ~n2497 ;
  buffer buf_n2499( .i (n2498), .o (n2499) );
  assign n2501 = ~n2286 & n2499 ;
  buffer buf_n2502( .i (n2501), .o (n2502) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2500( .i (n2499), .o (n2500) );
  assign n2503 = n2287 & ~n2500 ;
  assign n2504 = n2502 | n2503 ;
  buffer buf_n2505( .i (n2504), .o (n2505) );
  assign n2507 = n2283 | n2505 ;
  buffer buf_n2508( .i (n2507), .o (n2508) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2506( .i (n2505), .o (n2506) );
  assign n2513 = n2284 & n2506 ;
  assign n2514 = n2508 & ~n2513 ;
  buffer buf_n2515( .i (n2514), .o (n2515) );
  assign n2517 = ~n2280 & n2515 ;
  buffer buf_n2518( .i (n2517), .o (n2518) );
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2516( .i (n2515), .o (n2516) );
  assign n2519 = n2281 & ~n2516 ;
  assign n2520 = n2518 | n2519 ;
  buffer buf_n2521( .i (n2520), .o (n2521) );
  assign n2523 = n2277 | n2521 ;
  buffer buf_n2524( .i (n2523), .o (n2524) );
  buffer buf_n2278( .i (n2277), .o (n2278) );
  buffer buf_n2522( .i (n2521), .o (n2522) );
  assign n2529 = n2278 & n2522 ;
  assign n2530 = n2524 & ~n2529 ;
  buffer buf_n2531( .i (n2530), .o (n2531) );
  assign n2533 = ~n2274 & n2531 ;
  buffer buf_n2534( .i (n2533), .o (n2534) );
  buffer buf_n2275( .i (n2274), .o (n2275) );
  buffer buf_n2532( .i (n2531), .o (n2532) );
  assign n2535 = n2275 & ~n2532 ;
  assign n2536 = n2534 | n2535 ;
  buffer buf_n2537( .i (n2536), .o (n2537) );
  assign n2539 = n2271 | n2537 ;
  buffer buf_n2540( .i (n2539), .o (n2540) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2538( .i (n2537), .o (n2538) );
  assign n2545 = n2272 & n2538 ;
  assign n2546 = n2540 & ~n2545 ;
  buffer buf_n2547( .i (n2546), .o (n2547) );
  assign n2551 = ~n2266 & n2547 ;
  buffer buf_n2552( .i (n2551), .o (n2552) );
  buffer buf_n2553( .i (n2552), .o (n2553) );
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  buffer buf_n2269( .i (n2268), .o (n2269) );
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  assign n2555 = n2269 & ~n2550 ;
  assign n2556 = n2554 | n2555 ;
  buffer buf_n2557( .i (n2556), .o (n2557) );
  assign n2559 = n2263 | n2557 ;
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  buffer buf_n2558( .i (n2557), .o (n2558) );
  assign n2565 = n2264 & n2558 ;
  assign n2566 = n2560 & ~n2565 ;
  buffer buf_n2567( .i (n2566), .o (n2567) );
  assign n2569 = ~n2260 & n2567 ;
  buffer buf_n2570( .i (n2569), .o (n2570) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2568( .i (n2567), .o (n2568) );
  assign n2571 = n2261 & ~n2568 ;
  assign n2572 = n2570 | n2571 ;
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  buffer buf_n2563( .i (n2562), .o (n2563) );
  buffer buf_n2564( .i (n2563), .o (n2564) );
  assign n2573 = n2564 & ~n2570 ;
  buffer buf_n2574( .i (n2573), .o (n2574) );
  assign n2576 = N18 & N528 ;
  buffer buf_n2577( .i (n2576), .o (n2577) );
  buffer buf_n2541( .i (n2540), .o (n2541) );
  buffer buf_n2542( .i (n2541), .o (n2542) );
  buffer buf_n2543( .i (n2542), .o (n2543) );
  buffer buf_n2544( .i (n2543), .o (n2544) );
  assign n2581 = n2544 & ~n2552 ;
  buffer buf_n2582( .i (n2581), .o (n2582) );
  assign n2584 = N35 & N511 ;
  buffer buf_n2585( .i (n2584), .o (n2585) );
  buffer buf_n2525( .i (n2524), .o (n2525) );
  buffer buf_n2526( .i (n2525), .o (n2526) );
  buffer buf_n2527( .i (n2526), .o (n2527) );
  buffer buf_n2528( .i (n2527), .o (n2528) );
  assign n2587 = n2528 & ~n2534 ;
  buffer buf_n2588( .i (n2587), .o (n2588) );
  assign n2590 = N494 & N52 ;
  buffer buf_n2591( .i (n2590), .o (n2591) );
  buffer buf_n2509( .i (n2508), .o (n2509) );
  buffer buf_n2510( .i (n2509), .o (n2510) );
  buffer buf_n2511( .i (n2510), .o (n2511) );
  buffer buf_n2512( .i (n2511), .o (n2512) );
  assign n2593 = n2512 & ~n2518 ;
  buffer buf_n2594( .i (n2593), .o (n2594) );
  assign n2596 = N477 & N69 ;
  buffer buf_n2597( .i (n2596), .o (n2597) );
  buffer buf_n2493( .i (n2492), .o (n2493) );
  buffer buf_n2494( .i (n2493), .o (n2494) );
  buffer buf_n2495( .i (n2494), .o (n2495) );
  buffer buf_n2496( .i (n2495), .o (n2496) );
  assign n2599 = n2496 & ~n2502 ;
  buffer buf_n2600( .i (n2599), .o (n2600) );
  assign n2602 = N460 & N86 ;
  buffer buf_n2603( .i (n2602), .o (n2603) );
  buffer buf_n2477( .i (n2476), .o (n2477) );
  buffer buf_n2478( .i (n2477), .o (n2478) );
  buffer buf_n2479( .i (n2478), .o (n2479) );
  buffer buf_n2480( .i (n2479), .o (n2480) );
  assign n2605 = n2480 & ~n2486 ;
  buffer buf_n2606( .i (n2605), .o (n2606) );
  assign n2608 = N103 & N443 ;
  buffer buf_n2609( .i (n2608), .o (n2609) );
  buffer buf_n2461( .i (n2460), .o (n2461) );
  buffer buf_n2462( .i (n2461), .o (n2462) );
  buffer buf_n2463( .i (n2462), .o (n2463) );
  buffer buf_n2464( .i (n2463), .o (n2464) );
  assign n2611 = n2464 & ~n2470 ;
  buffer buf_n2612( .i (n2611), .o (n2612) );
  assign n2614 = N120 & N426 ;
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2445( .i (n2444), .o (n2445) );
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n2448( .i (n2447), .o (n2448) );
  assign n2617 = n2448 & ~n2454 ;
  buffer buf_n2618( .i (n2617), .o (n2618) );
  assign n2620 = N137 & N409 ;
  buffer buf_n2621( .i (n2620), .o (n2621) );
  buffer buf_n2429( .i (n2428), .o (n2429) );
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  buffer buf_n2432( .i (n2431), .o (n2432) );
  assign n2623 = n2432 & ~n2438 ;
  buffer buf_n2624( .i (n2623), .o (n2624) );
  assign n2626 = N154 & N392 ;
  buffer buf_n2627( .i (n2626), .o (n2627) );
  buffer buf_n2413( .i (n2412), .o (n2413) );
  buffer buf_n2414( .i (n2413), .o (n2414) );
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n2416( .i (n2415), .o (n2416) );
  assign n2629 = n2416 & ~n2422 ;
  buffer buf_n2630( .i (n2629), .o (n2630) );
  assign n2632 = N171 & N375 ;
  buffer buf_n2633( .i (n2632), .o (n2633) );
  buffer buf_n2397( .i (n2396), .o (n2397) );
  buffer buf_n2398( .i (n2397), .o (n2398) );
  buffer buf_n2399( .i (n2398), .o (n2399) );
  buffer buf_n2400( .i (n2399), .o (n2400) );
  assign n2635 = n2400 & ~n2406 ;
  buffer buf_n2636( .i (n2635), .o (n2636) );
  assign n2638 = N188 & N358 ;
  buffer buf_n2639( .i (n2638), .o (n2639) );
  buffer buf_n2381( .i (n2380), .o (n2381) );
  buffer buf_n2382( .i (n2381), .o (n2382) );
  buffer buf_n2383( .i (n2382), .o (n2383) );
  buffer buf_n2384( .i (n2383), .o (n2384) );
  assign n2641 = n2384 & ~n2390 ;
  buffer buf_n2642( .i (n2641), .o (n2642) );
  assign n2644 = N205 & N341 ;
  buffer buf_n2645( .i (n2644), .o (n2645) );
  buffer buf_n2365( .i (n2364), .o (n2365) );
  buffer buf_n2366( .i (n2365), .o (n2366) );
  buffer buf_n2367( .i (n2366), .o (n2367) );
  buffer buf_n2368( .i (n2367), .o (n2368) );
  assign n2647 = n2368 & ~n2374 ;
  buffer buf_n2648( .i (n2647), .o (n2648) );
  assign n2650 = N222 & N324 ;
  buffer buf_n2651( .i (n2650), .o (n2651) );
  buffer buf_n2350( .i (n2349), .o (n2350) );
  buffer buf_n2351( .i (n2350), .o (n2351) );
  buffer buf_n2352( .i (n2351), .o (n2352) );
  buffer buf_n2353( .i (n2352), .o (n2353) );
  assign n2653 = n2353 & ~n2358 ;
  buffer buf_n2654( .i (n2653), .o (n2654) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  assign n2656 = N256 & N290 ;
  buffer buf_n2657( .i (n2656), .o (n2657) );
  assign n2662 = ~n2044 & n2657 ;
  buffer buf_n2663( .i (n2662), .o (n2663) );
  assign n2665 = N239 & N307 ;
  buffer buf_n2666( .i (n2665), .o (n2666) );
  assign n2668 = n2663 & ~n2666 ;
  buffer buf_n2669( .i (n2668), .o (n2669) );
  buffer buf_n2664( .i (n2663), .o (n2664) );
  buffer buf_n2667( .i (n2666), .o (n2667) );
  assign n2670 = ~n2664 & n2667 ;
  assign n2671 = n2669 | n2670 ;
  buffer buf_n2672( .i (n2671), .o (n2672) );
  assign n2674 = n2654 | n2672 ;
  buffer buf_n2675( .i (n2674), .o (n2675) );
  buffer buf_n2655( .i (n2654), .o (n2655) );
  buffer buf_n2673( .i (n2672), .o (n2673) );
  assign n2680 = n2655 & n2673 ;
  assign n2681 = n2675 & ~n2680 ;
  buffer buf_n2682( .i (n2681), .o (n2682) );
  assign n2684 = ~n2651 & n2682 ;
  buffer buf_n2685( .i (n2684), .o (n2685) );
  buffer buf_n2652( .i (n2651), .o (n2652) );
  buffer buf_n2683( .i (n2682), .o (n2683) );
  assign n2686 = n2652 & ~n2683 ;
  assign n2687 = n2685 | n2686 ;
  buffer buf_n2688( .i (n2687), .o (n2688) );
  assign n2690 = n2648 | n2688 ;
  buffer buf_n2691( .i (n2690), .o (n2691) );
  buffer buf_n2649( .i (n2648), .o (n2649) );
  buffer buf_n2689( .i (n2688), .o (n2689) );
  assign n2696 = n2649 & n2689 ;
  assign n2697 = n2691 & ~n2696 ;
  buffer buf_n2698( .i (n2697), .o (n2698) );
  assign n2700 = ~n2645 & n2698 ;
  buffer buf_n2701( .i (n2700), .o (n2701) );
  buffer buf_n2646( .i (n2645), .o (n2646) );
  buffer buf_n2699( .i (n2698), .o (n2699) );
  assign n2702 = n2646 & ~n2699 ;
  assign n2703 = n2701 | n2702 ;
  buffer buf_n2704( .i (n2703), .o (n2704) );
  assign n2706 = n2642 | n2704 ;
  buffer buf_n2707( .i (n2706), .o (n2707) );
  buffer buf_n2643( .i (n2642), .o (n2643) );
  buffer buf_n2705( .i (n2704), .o (n2705) );
  assign n2712 = n2643 & n2705 ;
  assign n2713 = n2707 & ~n2712 ;
  buffer buf_n2714( .i (n2713), .o (n2714) );
  assign n2716 = ~n2639 & n2714 ;
  buffer buf_n2717( .i (n2716), .o (n2717) );
  buffer buf_n2640( .i (n2639), .o (n2640) );
  buffer buf_n2715( .i (n2714), .o (n2715) );
  assign n2718 = n2640 & ~n2715 ;
  assign n2719 = n2717 | n2718 ;
  buffer buf_n2720( .i (n2719), .o (n2720) );
  assign n2722 = n2636 | n2720 ;
  buffer buf_n2723( .i (n2722), .o (n2723) );
  buffer buf_n2637( .i (n2636), .o (n2637) );
  buffer buf_n2721( .i (n2720), .o (n2721) );
  assign n2728 = n2637 & n2721 ;
  assign n2729 = n2723 & ~n2728 ;
  buffer buf_n2730( .i (n2729), .o (n2730) );
  assign n2732 = ~n2633 & n2730 ;
  buffer buf_n2733( .i (n2732), .o (n2733) );
  buffer buf_n2634( .i (n2633), .o (n2634) );
  buffer buf_n2731( .i (n2730), .o (n2731) );
  assign n2734 = n2634 & ~n2731 ;
  assign n2735 = n2733 | n2734 ;
  buffer buf_n2736( .i (n2735), .o (n2736) );
  assign n2738 = n2630 | n2736 ;
  buffer buf_n2739( .i (n2738), .o (n2739) );
  buffer buf_n2631( .i (n2630), .o (n2631) );
  buffer buf_n2737( .i (n2736), .o (n2737) );
  assign n2744 = n2631 & n2737 ;
  assign n2745 = n2739 & ~n2744 ;
  buffer buf_n2746( .i (n2745), .o (n2746) );
  assign n2748 = ~n2627 & n2746 ;
  buffer buf_n2749( .i (n2748), .o (n2749) );
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2747( .i (n2746), .o (n2747) );
  assign n2750 = n2628 & ~n2747 ;
  assign n2751 = n2749 | n2750 ;
  buffer buf_n2752( .i (n2751), .o (n2752) );
  assign n2754 = n2624 | n2752 ;
  buffer buf_n2755( .i (n2754), .o (n2755) );
  buffer buf_n2625( .i (n2624), .o (n2625) );
  buffer buf_n2753( .i (n2752), .o (n2753) );
  assign n2760 = n2625 & n2753 ;
  assign n2761 = n2755 & ~n2760 ;
  buffer buf_n2762( .i (n2761), .o (n2762) );
  assign n2764 = ~n2621 & n2762 ;
  buffer buf_n2765( .i (n2764), .o (n2765) );
  buffer buf_n2622( .i (n2621), .o (n2622) );
  buffer buf_n2763( .i (n2762), .o (n2763) );
  assign n2766 = n2622 & ~n2763 ;
  assign n2767 = n2765 | n2766 ;
  buffer buf_n2768( .i (n2767), .o (n2768) );
  assign n2770 = n2618 | n2768 ;
  buffer buf_n2771( .i (n2770), .o (n2771) );
  buffer buf_n2619( .i (n2618), .o (n2619) );
  buffer buf_n2769( .i (n2768), .o (n2769) );
  assign n2776 = n2619 & n2769 ;
  assign n2777 = n2771 & ~n2776 ;
  buffer buf_n2778( .i (n2777), .o (n2778) );
  assign n2780 = ~n2615 & n2778 ;
  buffer buf_n2781( .i (n2780), .o (n2781) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  buffer buf_n2779( .i (n2778), .o (n2779) );
  assign n2782 = n2616 & ~n2779 ;
  assign n2783 = n2781 | n2782 ;
  buffer buf_n2784( .i (n2783), .o (n2784) );
  assign n2786 = n2612 | n2784 ;
  buffer buf_n2787( .i (n2786), .o (n2787) );
  buffer buf_n2613( .i (n2612), .o (n2613) );
  buffer buf_n2785( .i (n2784), .o (n2785) );
  assign n2792 = n2613 & n2785 ;
  assign n2793 = n2787 & ~n2792 ;
  buffer buf_n2794( .i (n2793), .o (n2794) );
  assign n2796 = ~n2609 & n2794 ;
  buffer buf_n2797( .i (n2796), .o (n2797) );
  buffer buf_n2610( .i (n2609), .o (n2610) );
  buffer buf_n2795( .i (n2794), .o (n2795) );
  assign n2798 = n2610 & ~n2795 ;
  assign n2799 = n2797 | n2798 ;
  buffer buf_n2800( .i (n2799), .o (n2800) );
  assign n2802 = n2606 | n2800 ;
  buffer buf_n2803( .i (n2802), .o (n2803) );
  buffer buf_n2607( .i (n2606), .o (n2607) );
  buffer buf_n2801( .i (n2800), .o (n2801) );
  assign n2808 = n2607 & n2801 ;
  assign n2809 = n2803 & ~n2808 ;
  buffer buf_n2810( .i (n2809), .o (n2810) );
  assign n2812 = ~n2603 & n2810 ;
  buffer buf_n2813( .i (n2812), .o (n2813) );
  buffer buf_n2604( .i (n2603), .o (n2604) );
  buffer buf_n2811( .i (n2810), .o (n2811) );
  assign n2814 = n2604 & ~n2811 ;
  assign n2815 = n2813 | n2814 ;
  buffer buf_n2816( .i (n2815), .o (n2816) );
  assign n2818 = n2600 | n2816 ;
  buffer buf_n2819( .i (n2818), .o (n2819) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  buffer buf_n2817( .i (n2816), .o (n2817) );
  assign n2824 = n2601 & n2817 ;
  assign n2825 = n2819 & ~n2824 ;
  buffer buf_n2826( .i (n2825), .o (n2826) );
  assign n2828 = ~n2597 & n2826 ;
  buffer buf_n2829( .i (n2828), .o (n2829) );
  buffer buf_n2598( .i (n2597), .o (n2598) );
  buffer buf_n2827( .i (n2826), .o (n2827) );
  assign n2830 = n2598 & ~n2827 ;
  assign n2831 = n2829 | n2830 ;
  buffer buf_n2832( .i (n2831), .o (n2832) );
  assign n2834 = n2594 | n2832 ;
  buffer buf_n2835( .i (n2834), .o (n2835) );
  buffer buf_n2595( .i (n2594), .o (n2595) );
  buffer buf_n2833( .i (n2832), .o (n2833) );
  assign n2840 = n2595 & n2833 ;
  assign n2841 = n2835 & ~n2840 ;
  buffer buf_n2842( .i (n2841), .o (n2842) );
  assign n2844 = ~n2591 & n2842 ;
  buffer buf_n2845( .i (n2844), .o (n2845) );
  buffer buf_n2592( .i (n2591), .o (n2592) );
  buffer buf_n2843( .i (n2842), .o (n2843) );
  assign n2846 = n2592 & ~n2843 ;
  assign n2847 = n2845 | n2846 ;
  buffer buf_n2848( .i (n2847), .o (n2848) );
  assign n2850 = n2588 | n2848 ;
  buffer buf_n2851( .i (n2850), .o (n2851) );
  buffer buf_n2589( .i (n2588), .o (n2589) );
  buffer buf_n2849( .i (n2848), .o (n2849) );
  assign n2856 = n2589 & n2849 ;
  assign n2857 = n2851 & ~n2856 ;
  buffer buf_n2858( .i (n2857), .o (n2858) );
  assign n2860 = ~n2585 & n2858 ;
  buffer buf_n2861( .i (n2860), .o (n2861) );
  buffer buf_n2586( .i (n2585), .o (n2586) );
  buffer buf_n2859( .i (n2858), .o (n2859) );
  assign n2862 = n2586 & ~n2859 ;
  assign n2863 = n2861 | n2862 ;
  buffer buf_n2864( .i (n2863), .o (n2864) );
  assign n2866 = n2582 | n2864 ;
  buffer buf_n2867( .i (n2866), .o (n2867) );
  buffer buf_n2583( .i (n2582), .o (n2583) );
  buffer buf_n2865( .i (n2864), .o (n2865) );
  assign n2872 = n2583 & n2865 ;
  assign n2873 = n2867 & ~n2872 ;
  buffer buf_n2874( .i (n2873), .o (n2874) );
  assign n2878 = ~n2577 & n2874 ;
  buffer buf_n2879( .i (n2878), .o (n2879) );
  buffer buf_n2880( .i (n2879), .o (n2880) );
  buffer buf_n2881( .i (n2880), .o (n2881) );
  buffer buf_n2578( .i (n2577), .o (n2578) );
  buffer buf_n2579( .i (n2578), .o (n2579) );
  buffer buf_n2580( .i (n2579), .o (n2580) );
  buffer buf_n2875( .i (n2874), .o (n2875) );
  buffer buf_n2876( .i (n2875), .o (n2876) );
  buffer buf_n2877( .i (n2876), .o (n2877) );
  assign n2882 = n2580 & ~n2877 ;
  assign n2883 = n2881 | n2882 ;
  buffer buf_n2884( .i (n2883), .o (n2884) );
  assign n2886 = n2574 & n2884 ;
  buffer buf_n2887( .i (n2886), .o (n2887) );
  buffer buf_n2575( .i (n2574), .o (n2575) );
  buffer buf_n2885( .i (n2884), .o (n2885) );
  assign n2889 = n2575 | n2885 ;
  assign n2890 = ~n2887 & n2889 ;
  buffer buf_n2868( .i (n2867), .o (n2868) );
  buffer buf_n2869( .i (n2868), .o (n2869) );
  buffer buf_n2870( .i (n2869), .o (n2870) );
  buffer buf_n2871( .i (n2870), .o (n2871) );
  assign n2891 = n2871 & ~n2879 ;
  buffer buf_n2892( .i (n2891), .o (n2892) );
  assign n2894 = N35 & N528 ;
  buffer buf_n2895( .i (n2894), .o (n2895) );
  buffer buf_n2852( .i (n2851), .o (n2852) );
  buffer buf_n2853( .i (n2852), .o (n2853) );
  buffer buf_n2854( .i (n2853), .o (n2854) );
  buffer buf_n2855( .i (n2854), .o (n2855) );
  assign n2897 = n2855 & ~n2861 ;
  buffer buf_n2898( .i (n2897), .o (n2898) );
  assign n2900 = N511 & N52 ;
  buffer buf_n2901( .i (n2900), .o (n2901) );
  buffer buf_n2836( .i (n2835), .o (n2836) );
  buffer buf_n2837( .i (n2836), .o (n2837) );
  buffer buf_n2838( .i (n2837), .o (n2838) );
  buffer buf_n2839( .i (n2838), .o (n2839) );
  assign n2903 = n2839 & ~n2845 ;
  buffer buf_n2904( .i (n2903), .o (n2904) );
  assign n2906 = N494 & N69 ;
  buffer buf_n2907( .i (n2906), .o (n2907) );
  buffer buf_n2820( .i (n2819), .o (n2820) );
  buffer buf_n2821( .i (n2820), .o (n2821) );
  buffer buf_n2822( .i (n2821), .o (n2822) );
  buffer buf_n2823( .i (n2822), .o (n2823) );
  assign n2909 = n2823 & ~n2829 ;
  buffer buf_n2910( .i (n2909), .o (n2910) );
  assign n2912 = N477 & N86 ;
  buffer buf_n2913( .i (n2912), .o (n2913) );
  buffer buf_n2804( .i (n2803), .o (n2804) );
  buffer buf_n2805( .i (n2804), .o (n2805) );
  buffer buf_n2806( .i (n2805), .o (n2806) );
  buffer buf_n2807( .i (n2806), .o (n2807) );
  assign n2915 = n2807 & ~n2813 ;
  buffer buf_n2916( .i (n2915), .o (n2916) );
  assign n2918 = N103 & N460 ;
  buffer buf_n2919( .i (n2918), .o (n2919) );
  buffer buf_n2788( .i (n2787), .o (n2788) );
  buffer buf_n2789( .i (n2788), .o (n2789) );
  buffer buf_n2790( .i (n2789), .o (n2790) );
  buffer buf_n2791( .i (n2790), .o (n2791) );
  assign n2921 = n2791 & ~n2797 ;
  buffer buf_n2922( .i (n2921), .o (n2922) );
  assign n2924 = N120 & N443 ;
  buffer buf_n2925( .i (n2924), .o (n2925) );
  buffer buf_n2772( .i (n2771), .o (n2772) );
  buffer buf_n2773( .i (n2772), .o (n2773) );
  buffer buf_n2774( .i (n2773), .o (n2774) );
  buffer buf_n2775( .i (n2774), .o (n2775) );
  assign n2927 = n2775 & ~n2781 ;
  buffer buf_n2928( .i (n2927), .o (n2928) );
  assign n2930 = N137 & N426 ;
  buffer buf_n2931( .i (n2930), .o (n2931) );
  buffer buf_n2756( .i (n2755), .o (n2756) );
  buffer buf_n2757( .i (n2756), .o (n2757) );
  buffer buf_n2758( .i (n2757), .o (n2758) );
  buffer buf_n2759( .i (n2758), .o (n2759) );
  assign n2933 = n2759 & ~n2765 ;
  buffer buf_n2934( .i (n2933), .o (n2934) );
  assign n2936 = N154 & N409 ;
  buffer buf_n2937( .i (n2936), .o (n2937) );
  buffer buf_n2740( .i (n2739), .o (n2740) );
  buffer buf_n2741( .i (n2740), .o (n2741) );
  buffer buf_n2742( .i (n2741), .o (n2742) );
  buffer buf_n2743( .i (n2742), .o (n2743) );
  assign n2939 = n2743 & ~n2749 ;
  buffer buf_n2940( .i (n2939), .o (n2940) );
  assign n2942 = N171 & N392 ;
  buffer buf_n2943( .i (n2942), .o (n2943) );
  buffer buf_n2724( .i (n2723), .o (n2724) );
  buffer buf_n2725( .i (n2724), .o (n2725) );
  buffer buf_n2726( .i (n2725), .o (n2726) );
  buffer buf_n2727( .i (n2726), .o (n2727) );
  assign n2945 = n2727 & ~n2733 ;
  buffer buf_n2946( .i (n2945), .o (n2946) );
  assign n2948 = N188 & N375 ;
  buffer buf_n2949( .i (n2948), .o (n2949) );
  buffer buf_n2708( .i (n2707), .o (n2708) );
  buffer buf_n2709( .i (n2708), .o (n2709) );
  buffer buf_n2710( .i (n2709), .o (n2710) );
  buffer buf_n2711( .i (n2710), .o (n2711) );
  assign n2951 = n2711 & ~n2717 ;
  buffer buf_n2952( .i (n2951), .o (n2952) );
  assign n2954 = N205 & N358 ;
  buffer buf_n2955( .i (n2954), .o (n2955) );
  buffer buf_n2692( .i (n2691), .o (n2692) );
  buffer buf_n2693( .i (n2692), .o (n2693) );
  buffer buf_n2694( .i (n2693), .o (n2694) );
  buffer buf_n2695( .i (n2694), .o (n2695) );
  assign n2957 = n2695 & ~n2701 ;
  buffer buf_n2958( .i (n2957), .o (n2958) );
  assign n2960 = N222 & N341 ;
  buffer buf_n2961( .i (n2960), .o (n2961) );
  buffer buf_n2676( .i (n2675), .o (n2676) );
  buffer buf_n2677( .i (n2676), .o (n2677) );
  buffer buf_n2678( .i (n2677), .o (n2678) );
  buffer buf_n2679( .i (n2678), .o (n2679) );
  assign n2963 = n2679 & ~n2685 ;
  buffer buf_n2964( .i (n2963), .o (n2964) );
  assign n2966 = N239 & N324 ;
  buffer buf_n2967( .i (n2966), .o (n2967) );
  assign n2969 = N256 & N307 ;
  buffer buf_n2970( .i (n2969), .o (n2970) );
  buffer buf_n2658( .i (n2657), .o (n2658) );
  buffer buf_n2659( .i (n2658), .o (n2659) );
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2660), .o (n2661) );
  assign n2972 = n2661 & ~n2669 ;
  buffer buf_n2973( .i (n2972), .o (n2973) );
  assign n2975 = n2970 | n2973 ;
  buffer buf_n2976( .i (n2975), .o (n2976) );
  buffer buf_n2971( .i (n2970), .o (n2971) );
  buffer buf_n2974( .i (n2973), .o (n2974) );
  assign n2985 = n2971 & n2974 ;
  assign n2986 = n2976 & ~n2985 ;
  buffer buf_n2987( .i (n2986), .o (n2987) );
  assign n2989 = ~n2967 & n2987 ;
  buffer buf_n2990( .i (n2989), .o (n2990) );
  buffer buf_n2968( .i (n2967), .o (n2968) );
  buffer buf_n2988( .i (n2987), .o (n2988) );
  assign n2995 = n2968 & ~n2988 ;
  assign n2996 = n2990 | n2995 ;
  buffer buf_n2997( .i (n2996), .o (n2997) );
  assign n2999 = n2964 | n2997 ;
  buffer buf_n3000( .i (n2999), .o (n3000) );
  buffer buf_n2965( .i (n2964), .o (n2965) );
  buffer buf_n2998( .i (n2997), .o (n2998) );
  assign n3009 = n2965 & n2998 ;
  assign n3010 = n3000 & ~n3009 ;
  buffer buf_n3011( .i (n3010), .o (n3011) );
  assign n3013 = ~n2961 & n3011 ;
  buffer buf_n3014( .i (n3013), .o (n3014) );
  buffer buf_n2962( .i (n2961), .o (n2962) );
  buffer buf_n3012( .i (n3011), .o (n3012) );
  assign n3019 = n2962 & ~n3012 ;
  assign n3020 = n3014 | n3019 ;
  buffer buf_n3021( .i (n3020), .o (n3021) );
  assign n3023 = n2958 | n3021 ;
  buffer buf_n3024( .i (n3023), .o (n3024) );
  buffer buf_n2959( .i (n2958), .o (n2959) );
  buffer buf_n3022( .i (n3021), .o (n3022) );
  assign n3033 = n2959 & n3022 ;
  assign n3034 = n3024 & ~n3033 ;
  buffer buf_n3035( .i (n3034), .o (n3035) );
  assign n3037 = ~n2955 & n3035 ;
  buffer buf_n3038( .i (n3037), .o (n3038) );
  buffer buf_n2956( .i (n2955), .o (n2956) );
  buffer buf_n3036( .i (n3035), .o (n3036) );
  assign n3043 = n2956 & ~n3036 ;
  assign n3044 = n3038 | n3043 ;
  buffer buf_n3045( .i (n3044), .o (n3045) );
  assign n3047 = n2952 | n3045 ;
  buffer buf_n3048( .i (n3047), .o (n3048) );
  buffer buf_n2953( .i (n2952), .o (n2953) );
  buffer buf_n3046( .i (n3045), .o (n3046) );
  assign n3057 = n2953 & n3046 ;
  assign n3058 = n3048 & ~n3057 ;
  buffer buf_n3059( .i (n3058), .o (n3059) );
  assign n3061 = ~n2949 & n3059 ;
  buffer buf_n3062( .i (n3061), .o (n3062) );
  buffer buf_n2950( .i (n2949), .o (n2950) );
  buffer buf_n3060( .i (n3059), .o (n3060) );
  assign n3067 = n2950 & ~n3060 ;
  assign n3068 = n3062 | n3067 ;
  buffer buf_n3069( .i (n3068), .o (n3069) );
  assign n3071 = n2946 | n3069 ;
  buffer buf_n3072( .i (n3071), .o (n3072) );
  buffer buf_n2947( .i (n2946), .o (n2947) );
  buffer buf_n3070( .i (n3069), .o (n3070) );
  assign n3081 = n2947 & n3070 ;
  assign n3082 = n3072 & ~n3081 ;
  buffer buf_n3083( .i (n3082), .o (n3083) );
  assign n3085 = ~n2943 & n3083 ;
  buffer buf_n3086( .i (n3085), .o (n3086) );
  buffer buf_n2944( .i (n2943), .o (n2944) );
  buffer buf_n3084( .i (n3083), .o (n3084) );
  assign n3091 = n2944 & ~n3084 ;
  assign n3092 = n3086 | n3091 ;
  buffer buf_n3093( .i (n3092), .o (n3093) );
  assign n3095 = n2940 | n3093 ;
  buffer buf_n3096( .i (n3095), .o (n3096) );
  buffer buf_n2941( .i (n2940), .o (n2941) );
  buffer buf_n3094( .i (n3093), .o (n3094) );
  assign n3105 = n2941 & n3094 ;
  assign n3106 = n3096 & ~n3105 ;
  buffer buf_n3107( .i (n3106), .o (n3107) );
  assign n3109 = ~n2937 & n3107 ;
  buffer buf_n3110( .i (n3109), .o (n3110) );
  buffer buf_n2938( .i (n2937), .o (n2938) );
  buffer buf_n3108( .i (n3107), .o (n3108) );
  assign n3115 = n2938 & ~n3108 ;
  assign n3116 = n3110 | n3115 ;
  buffer buf_n3117( .i (n3116), .o (n3117) );
  assign n3119 = n2934 | n3117 ;
  buffer buf_n3120( .i (n3119), .o (n3120) );
  buffer buf_n2935( .i (n2934), .o (n2935) );
  buffer buf_n3118( .i (n3117), .o (n3118) );
  assign n3129 = n2935 & n3118 ;
  assign n3130 = n3120 & ~n3129 ;
  buffer buf_n3131( .i (n3130), .o (n3131) );
  assign n3133 = ~n2931 & n3131 ;
  buffer buf_n3134( .i (n3133), .o (n3134) );
  buffer buf_n2932( .i (n2931), .o (n2932) );
  buffer buf_n3132( .i (n3131), .o (n3132) );
  assign n3139 = n2932 & ~n3132 ;
  assign n3140 = n3134 | n3139 ;
  buffer buf_n3141( .i (n3140), .o (n3141) );
  assign n3143 = n2928 | n3141 ;
  buffer buf_n3144( .i (n3143), .o (n3144) );
  buffer buf_n2929( .i (n2928), .o (n2929) );
  buffer buf_n3142( .i (n3141), .o (n3142) );
  assign n3153 = n2929 & n3142 ;
  assign n3154 = n3144 & ~n3153 ;
  buffer buf_n3155( .i (n3154), .o (n3155) );
  assign n3157 = ~n2925 & n3155 ;
  buffer buf_n3158( .i (n3157), .o (n3158) );
  buffer buf_n2926( .i (n2925), .o (n2926) );
  buffer buf_n3156( .i (n3155), .o (n3156) );
  assign n3163 = n2926 & ~n3156 ;
  assign n3164 = n3158 | n3163 ;
  buffer buf_n3165( .i (n3164), .o (n3165) );
  assign n3167 = n2922 | n3165 ;
  buffer buf_n3168( .i (n3167), .o (n3168) );
  buffer buf_n2923( .i (n2922), .o (n2923) );
  buffer buf_n3166( .i (n3165), .o (n3166) );
  assign n3177 = n2923 & n3166 ;
  assign n3178 = n3168 & ~n3177 ;
  buffer buf_n3179( .i (n3178), .o (n3179) );
  assign n3181 = ~n2919 & n3179 ;
  buffer buf_n3182( .i (n3181), .o (n3182) );
  buffer buf_n2920( .i (n2919), .o (n2920) );
  buffer buf_n3180( .i (n3179), .o (n3180) );
  assign n3187 = n2920 & ~n3180 ;
  assign n3188 = n3182 | n3187 ;
  buffer buf_n3189( .i (n3188), .o (n3189) );
  assign n3191 = n2916 | n3189 ;
  buffer buf_n3192( .i (n3191), .o (n3192) );
  buffer buf_n2917( .i (n2916), .o (n2917) );
  buffer buf_n3190( .i (n3189), .o (n3190) );
  assign n3201 = n2917 & n3190 ;
  assign n3202 = n3192 & ~n3201 ;
  buffer buf_n3203( .i (n3202), .o (n3203) );
  assign n3205 = ~n2913 & n3203 ;
  buffer buf_n3206( .i (n3205), .o (n3206) );
  buffer buf_n2914( .i (n2913), .o (n2914) );
  buffer buf_n3204( .i (n3203), .o (n3204) );
  assign n3211 = n2914 & ~n3204 ;
  assign n3212 = n3206 | n3211 ;
  buffer buf_n3213( .i (n3212), .o (n3213) );
  assign n3215 = n2910 | n3213 ;
  buffer buf_n3216( .i (n3215), .o (n3216) );
  buffer buf_n2911( .i (n2910), .o (n2911) );
  buffer buf_n3214( .i (n3213), .o (n3214) );
  assign n3225 = n2911 & n3214 ;
  assign n3226 = n3216 & ~n3225 ;
  buffer buf_n3227( .i (n3226), .o (n3227) );
  assign n3229 = ~n2907 & n3227 ;
  buffer buf_n3230( .i (n3229), .o (n3230) );
  buffer buf_n2908( .i (n2907), .o (n2908) );
  buffer buf_n3228( .i (n3227), .o (n3228) );
  assign n3235 = n2908 & ~n3228 ;
  assign n3236 = n3230 | n3235 ;
  buffer buf_n3237( .i (n3236), .o (n3237) );
  assign n3239 = n2904 | n3237 ;
  buffer buf_n3240( .i (n3239), .o (n3240) );
  buffer buf_n2905( .i (n2904), .o (n2905) );
  buffer buf_n3238( .i (n3237), .o (n3238) );
  assign n3249 = n2905 & n3238 ;
  assign n3250 = n3240 & ~n3249 ;
  buffer buf_n3251( .i (n3250), .o (n3251) );
  assign n3253 = ~n2901 & n3251 ;
  buffer buf_n3254( .i (n3253), .o (n3254) );
  buffer buf_n2902( .i (n2901), .o (n2902) );
  buffer buf_n3252( .i (n3251), .o (n3252) );
  assign n3259 = n2902 & ~n3252 ;
  assign n3260 = n3254 | n3259 ;
  buffer buf_n3261( .i (n3260), .o (n3261) );
  assign n3263 = n2898 | n3261 ;
  buffer buf_n3264( .i (n3263), .o (n3264) );
  buffer buf_n2899( .i (n2898), .o (n2899) );
  buffer buf_n3262( .i (n3261), .o (n3262) );
  assign n3273 = n2899 & n3262 ;
  assign n3274 = n3264 & ~n3273 ;
  buffer buf_n3275( .i (n3274), .o (n3275) );
  assign n3277 = ~n2895 & n3275 ;
  buffer buf_n3278( .i (n3277), .o (n3278) );
  buffer buf_n2896( .i (n2895), .o (n2896) );
  buffer buf_n3276( .i (n3275), .o (n3276) );
  assign n3283 = n2896 & ~n3276 ;
  assign n3284 = n3278 | n3283 ;
  buffer buf_n3285( .i (n3284), .o (n3285) );
  assign n3287 = n2892 | n3285 ;
  buffer buf_n3288( .i (n3287), .o (n3288) );
  buffer buf_n2893( .i (n2892), .o (n2893) );
  buffer buf_n3286( .i (n3285), .o (n3286) );
  assign n3293 = n2893 & n3286 ;
  assign n3294 = n3288 & ~n3293 ;
  buffer buf_n3295( .i (n3294), .o (n3295) );
  assign n3297 = ~n2887 & n3295 ;
  buffer buf_n3298( .i (n3297), .o (n3298) );
  buffer buf_n2888( .i (n2887), .o (n2888) );
  buffer buf_n3296( .i (n3295), .o (n3296) );
  assign n3299 = n2888 & ~n3296 ;
  assign n3300 = n3298 | n3299 ;
  buffer buf_n3289( .i (n3288), .o (n3289) );
  buffer buf_n3290( .i (n3289), .o (n3290) );
  buffer buf_n3291( .i (n3290), .o (n3291) );
  buffer buf_n3292( .i (n3291), .o (n3292) );
  assign n3301 = n3292 & ~n3298 ;
  buffer buf_n3302( .i (n3301), .o (n3302) );
  buffer buf_n3265( .i (n3264), .o (n3265) );
  buffer buf_n3266( .i (n3265), .o (n3266) );
  buffer buf_n3267( .i (n3266), .o (n3267) );
  buffer buf_n3268( .i (n3267), .o (n3268) );
  buffer buf_n3269( .i (n3268), .o (n3269) );
  buffer buf_n3270( .i (n3269), .o (n3270) );
  buffer buf_n3271( .i (n3270), .o (n3271) );
  buffer buf_n3272( .i (n3271), .o (n3272) );
  buffer buf_n3279( .i (n3278), .o (n3279) );
  buffer buf_n3280( .i (n3279), .o (n3280) );
  buffer buf_n3281( .i (n3280), .o (n3281) );
  buffer buf_n3282( .i (n3281), .o (n3282) );
  assign n3304 = n3272 & ~n3282 ;
  buffer buf_n3305( .i (n3304), .o (n3305) );
  assign n3307 = N52 & N528 ;
  buffer buf_n3308( .i (n3307), .o (n3308) );
  buffer buf_n3241( .i (n3240), .o (n3241) );
  buffer buf_n3242( .i (n3241), .o (n3242) );
  buffer buf_n3243( .i (n3242), .o (n3243) );
  buffer buf_n3244( .i (n3243), .o (n3244) );
  buffer buf_n3245( .i (n3244), .o (n3245) );
  buffer buf_n3246( .i (n3245), .o (n3246) );
  buffer buf_n3247( .i (n3246), .o (n3247) );
  buffer buf_n3248( .i (n3247), .o (n3248) );
  buffer buf_n3255( .i (n3254), .o (n3255) );
  buffer buf_n3256( .i (n3255), .o (n3256) );
  buffer buf_n3257( .i (n3256), .o (n3257) );
  buffer buf_n3258( .i (n3257), .o (n3258) );
  assign n3310 = n3248 & ~n3258 ;
  buffer buf_n3311( .i (n3310), .o (n3311) );
  assign n3313 = N511 & N69 ;
  buffer buf_n3314( .i (n3313), .o (n3314) );
  buffer buf_n3217( .i (n3216), .o (n3217) );
  buffer buf_n3218( .i (n3217), .o (n3218) );
  buffer buf_n3219( .i (n3218), .o (n3219) );
  buffer buf_n3220( .i (n3219), .o (n3220) );
  buffer buf_n3221( .i (n3220), .o (n3221) );
  buffer buf_n3222( .i (n3221), .o (n3222) );
  buffer buf_n3223( .i (n3222), .o (n3223) );
  buffer buf_n3224( .i (n3223), .o (n3224) );
  buffer buf_n3231( .i (n3230), .o (n3231) );
  buffer buf_n3232( .i (n3231), .o (n3232) );
  buffer buf_n3233( .i (n3232), .o (n3233) );
  buffer buf_n3234( .i (n3233), .o (n3234) );
  assign n3316 = n3224 & ~n3234 ;
  buffer buf_n3317( .i (n3316), .o (n3317) );
  assign n3319 = N494 & N86 ;
  buffer buf_n3320( .i (n3319), .o (n3320) );
  buffer buf_n3193( .i (n3192), .o (n3193) );
  buffer buf_n3194( .i (n3193), .o (n3194) );
  buffer buf_n3195( .i (n3194), .o (n3195) );
  buffer buf_n3196( .i (n3195), .o (n3196) );
  buffer buf_n3197( .i (n3196), .o (n3197) );
  buffer buf_n3198( .i (n3197), .o (n3198) );
  buffer buf_n3199( .i (n3198), .o (n3199) );
  buffer buf_n3200( .i (n3199), .o (n3200) );
  buffer buf_n3207( .i (n3206), .o (n3207) );
  buffer buf_n3208( .i (n3207), .o (n3208) );
  buffer buf_n3209( .i (n3208), .o (n3209) );
  buffer buf_n3210( .i (n3209), .o (n3210) );
  assign n3322 = n3200 & ~n3210 ;
  buffer buf_n3323( .i (n3322), .o (n3323) );
  assign n3325 = N103 & N477 ;
  buffer buf_n3326( .i (n3325), .o (n3326) );
  buffer buf_n3169( .i (n3168), .o (n3169) );
  buffer buf_n3170( .i (n3169), .o (n3170) );
  buffer buf_n3171( .i (n3170), .o (n3171) );
  buffer buf_n3172( .i (n3171), .o (n3172) );
  buffer buf_n3173( .i (n3172), .o (n3173) );
  buffer buf_n3174( .i (n3173), .o (n3174) );
  buffer buf_n3175( .i (n3174), .o (n3175) );
  buffer buf_n3176( .i (n3175), .o (n3176) );
  buffer buf_n3183( .i (n3182), .o (n3183) );
  buffer buf_n3184( .i (n3183), .o (n3184) );
  buffer buf_n3185( .i (n3184), .o (n3185) );
  buffer buf_n3186( .i (n3185), .o (n3186) );
  assign n3328 = n3176 & ~n3186 ;
  buffer buf_n3329( .i (n3328), .o (n3329) );
  assign n3331 = N120 & N460 ;
  buffer buf_n3332( .i (n3331), .o (n3332) );
  buffer buf_n3145( .i (n3144), .o (n3145) );
  buffer buf_n3146( .i (n3145), .o (n3146) );
  buffer buf_n3147( .i (n3146), .o (n3147) );
  buffer buf_n3148( .i (n3147), .o (n3148) );
  buffer buf_n3149( .i (n3148), .o (n3149) );
  buffer buf_n3150( .i (n3149), .o (n3150) );
  buffer buf_n3151( .i (n3150), .o (n3151) );
  buffer buf_n3152( .i (n3151), .o (n3152) );
  buffer buf_n3159( .i (n3158), .o (n3159) );
  buffer buf_n3160( .i (n3159), .o (n3160) );
  buffer buf_n3161( .i (n3160), .o (n3161) );
  buffer buf_n3162( .i (n3161), .o (n3162) );
  assign n3334 = n3152 & ~n3162 ;
  buffer buf_n3335( .i (n3334), .o (n3335) );
  assign n3337 = N137 & N443 ;
  buffer buf_n3338( .i (n3337), .o (n3338) );
  buffer buf_n3121( .i (n3120), .o (n3121) );
  buffer buf_n3122( .i (n3121), .o (n3122) );
  buffer buf_n3123( .i (n3122), .o (n3123) );
  buffer buf_n3124( .i (n3123), .o (n3124) );
  buffer buf_n3125( .i (n3124), .o (n3125) );
  buffer buf_n3126( .i (n3125), .o (n3126) );
  buffer buf_n3127( .i (n3126), .o (n3127) );
  buffer buf_n3128( .i (n3127), .o (n3128) );
  buffer buf_n3135( .i (n3134), .o (n3135) );
  buffer buf_n3136( .i (n3135), .o (n3136) );
  buffer buf_n3137( .i (n3136), .o (n3137) );
  buffer buf_n3138( .i (n3137), .o (n3138) );
  assign n3340 = n3128 & ~n3138 ;
  buffer buf_n3341( .i (n3340), .o (n3341) );
  assign n3343 = N154 & N426 ;
  buffer buf_n3344( .i (n3343), .o (n3344) );
  buffer buf_n3097( .i (n3096), .o (n3097) );
  buffer buf_n3098( .i (n3097), .o (n3098) );
  buffer buf_n3099( .i (n3098), .o (n3099) );
  buffer buf_n3100( .i (n3099), .o (n3100) );
  buffer buf_n3101( .i (n3100), .o (n3101) );
  buffer buf_n3102( .i (n3101), .o (n3102) );
  buffer buf_n3103( .i (n3102), .o (n3103) );
  buffer buf_n3104( .i (n3103), .o (n3104) );
  buffer buf_n3111( .i (n3110), .o (n3111) );
  buffer buf_n3112( .i (n3111), .o (n3112) );
  buffer buf_n3113( .i (n3112), .o (n3113) );
  buffer buf_n3114( .i (n3113), .o (n3114) );
  assign n3346 = n3104 & ~n3114 ;
  buffer buf_n3347( .i (n3346), .o (n3347) );
  assign n3349 = N171 & N409 ;
  buffer buf_n3350( .i (n3349), .o (n3350) );
  buffer buf_n3073( .i (n3072), .o (n3073) );
  buffer buf_n3074( .i (n3073), .o (n3074) );
  buffer buf_n3075( .i (n3074), .o (n3075) );
  buffer buf_n3076( .i (n3075), .o (n3076) );
  buffer buf_n3077( .i (n3076), .o (n3077) );
  buffer buf_n3078( .i (n3077), .o (n3078) );
  buffer buf_n3079( .i (n3078), .o (n3079) );
  buffer buf_n3080( .i (n3079), .o (n3080) );
  buffer buf_n3087( .i (n3086), .o (n3087) );
  buffer buf_n3088( .i (n3087), .o (n3088) );
  buffer buf_n3089( .i (n3088), .o (n3089) );
  buffer buf_n3090( .i (n3089), .o (n3090) );
  assign n3352 = n3080 & ~n3090 ;
  buffer buf_n3353( .i (n3352), .o (n3353) );
  assign n3355 = N188 & N392 ;
  buffer buf_n3356( .i (n3355), .o (n3356) );
  buffer buf_n3049( .i (n3048), .o (n3049) );
  buffer buf_n3050( .i (n3049), .o (n3050) );
  buffer buf_n3051( .i (n3050), .o (n3051) );
  buffer buf_n3052( .i (n3051), .o (n3052) );
  buffer buf_n3053( .i (n3052), .o (n3053) );
  buffer buf_n3054( .i (n3053), .o (n3054) );
  buffer buf_n3055( .i (n3054), .o (n3055) );
  buffer buf_n3056( .i (n3055), .o (n3056) );
  buffer buf_n3063( .i (n3062), .o (n3063) );
  buffer buf_n3064( .i (n3063), .o (n3064) );
  buffer buf_n3065( .i (n3064), .o (n3065) );
  buffer buf_n3066( .i (n3065), .o (n3066) );
  assign n3358 = n3056 & ~n3066 ;
  buffer buf_n3359( .i (n3358), .o (n3359) );
  assign n3361 = N205 & N375 ;
  buffer buf_n3362( .i (n3361), .o (n3362) );
  buffer buf_n3025( .i (n3024), .o (n3025) );
  buffer buf_n3026( .i (n3025), .o (n3026) );
  buffer buf_n3027( .i (n3026), .o (n3027) );
  buffer buf_n3028( .i (n3027), .o (n3028) );
  buffer buf_n3029( .i (n3028), .o (n3029) );
  buffer buf_n3030( .i (n3029), .o (n3030) );
  buffer buf_n3031( .i (n3030), .o (n3031) );
  buffer buf_n3032( .i (n3031), .o (n3032) );
  buffer buf_n3039( .i (n3038), .o (n3039) );
  buffer buf_n3040( .i (n3039), .o (n3040) );
  buffer buf_n3041( .i (n3040), .o (n3041) );
  buffer buf_n3042( .i (n3041), .o (n3042) );
  assign n3364 = n3032 & ~n3042 ;
  buffer buf_n3365( .i (n3364), .o (n3365) );
  assign n3367 = N222 & N358 ;
  buffer buf_n3368( .i (n3367), .o (n3368) );
  buffer buf_n3001( .i (n3000), .o (n3001) );
  buffer buf_n3002( .i (n3001), .o (n3002) );
  buffer buf_n3003( .i (n3002), .o (n3003) );
  buffer buf_n3004( .i (n3003), .o (n3004) );
  buffer buf_n3005( .i (n3004), .o (n3005) );
  buffer buf_n3006( .i (n3005), .o (n3006) );
  buffer buf_n3007( .i (n3006), .o (n3007) );
  buffer buf_n3008( .i (n3007), .o (n3008) );
  buffer buf_n3015( .i (n3014), .o (n3015) );
  buffer buf_n3016( .i (n3015), .o (n3016) );
  buffer buf_n3017( .i (n3016), .o (n3017) );
  buffer buf_n3018( .i (n3017), .o (n3018) );
  assign n3370 = n3008 & ~n3018 ;
  buffer buf_n3371( .i (n3370), .o (n3371) );
  assign n3373 = N239 & N341 ;
  buffer buf_n3374( .i (n3373), .o (n3374) );
  assign n3376 = N256 & N324 ;
  buffer buf_n3377( .i (n3376), .o (n3377) );
  buffer buf_n2977( .i (n2976), .o (n2977) );
  buffer buf_n2978( .i (n2977), .o (n2978) );
  buffer buf_n2979( .i (n2978), .o (n2979) );
  buffer buf_n2980( .i (n2979), .o (n2980) );
  buffer buf_n2981( .i (n2980), .o (n2981) );
  buffer buf_n2982( .i (n2981), .o (n2982) );
  buffer buf_n2983( .i (n2982), .o (n2983) );
  buffer buf_n2984( .i (n2983), .o (n2984) );
  buffer buf_n2991( .i (n2990), .o (n2991) );
  buffer buf_n2992( .i (n2991), .o (n2992) );
  buffer buf_n2993( .i (n2992), .o (n2993) );
  buffer buf_n2994( .i (n2993), .o (n2994) );
  assign n3379 = n2984 & ~n2994 ;
  buffer buf_n3380( .i (n3379), .o (n3380) );
  assign n3382 = n3377 | n3380 ;
  buffer buf_n3383( .i (n3382), .o (n3383) );
  buffer buf_n3378( .i (n3377), .o (n3378) );
  buffer buf_n3381( .i (n3380), .o (n3381) );
  assign n3392 = n3378 & n3381 ;
  assign n3393 = n3383 & ~n3392 ;
  buffer buf_n3394( .i (n3393), .o (n3394) );
  assign n3396 = ~n3374 & n3394 ;
  buffer buf_n3397( .i (n3396), .o (n3397) );
  buffer buf_n3375( .i (n3374), .o (n3375) );
  buffer buf_n3395( .i (n3394), .o (n3395) );
  assign n3402 = n3375 & ~n3395 ;
  assign n3403 = n3397 | n3402 ;
  buffer buf_n3404( .i (n3403), .o (n3404) );
  assign n3406 = n3371 | n3404 ;
  buffer buf_n3407( .i (n3406), .o (n3407) );
  buffer buf_n3372( .i (n3371), .o (n3372) );
  buffer buf_n3405( .i (n3404), .o (n3405) );
  assign n3416 = n3372 & n3405 ;
  assign n3417 = n3407 & ~n3416 ;
  buffer buf_n3418( .i (n3417), .o (n3418) );
  assign n3420 = ~n3368 & n3418 ;
  buffer buf_n3421( .i (n3420), .o (n3421) );
  buffer buf_n3369( .i (n3368), .o (n3369) );
  buffer buf_n3419( .i (n3418), .o (n3419) );
  assign n3426 = n3369 & ~n3419 ;
  assign n3427 = n3421 | n3426 ;
  buffer buf_n3428( .i (n3427), .o (n3428) );
  assign n3430 = n3365 | n3428 ;
  buffer buf_n3431( .i (n3430), .o (n3431) );
  buffer buf_n3366( .i (n3365), .o (n3366) );
  buffer buf_n3429( .i (n3428), .o (n3429) );
  assign n3440 = n3366 & n3429 ;
  assign n3441 = n3431 & ~n3440 ;
  buffer buf_n3442( .i (n3441), .o (n3442) );
  assign n3444 = ~n3362 & n3442 ;
  buffer buf_n3445( .i (n3444), .o (n3445) );
  buffer buf_n3363( .i (n3362), .o (n3363) );
  buffer buf_n3443( .i (n3442), .o (n3443) );
  assign n3450 = n3363 & ~n3443 ;
  assign n3451 = n3445 | n3450 ;
  buffer buf_n3452( .i (n3451), .o (n3452) );
  assign n3454 = n3359 | n3452 ;
  buffer buf_n3455( .i (n3454), .o (n3455) );
  buffer buf_n3360( .i (n3359), .o (n3360) );
  buffer buf_n3453( .i (n3452), .o (n3453) );
  assign n3464 = n3360 & n3453 ;
  assign n3465 = n3455 & ~n3464 ;
  buffer buf_n3466( .i (n3465), .o (n3466) );
  assign n3468 = ~n3356 & n3466 ;
  buffer buf_n3469( .i (n3468), .o (n3469) );
  buffer buf_n3357( .i (n3356), .o (n3357) );
  buffer buf_n3467( .i (n3466), .o (n3467) );
  assign n3474 = n3357 & ~n3467 ;
  assign n3475 = n3469 | n3474 ;
  buffer buf_n3476( .i (n3475), .o (n3476) );
  assign n3478 = n3353 | n3476 ;
  buffer buf_n3479( .i (n3478), .o (n3479) );
  buffer buf_n3354( .i (n3353), .o (n3354) );
  buffer buf_n3477( .i (n3476), .o (n3477) );
  assign n3488 = n3354 & n3477 ;
  assign n3489 = n3479 & ~n3488 ;
  buffer buf_n3490( .i (n3489), .o (n3490) );
  assign n3492 = ~n3350 & n3490 ;
  buffer buf_n3493( .i (n3492), .o (n3493) );
  buffer buf_n3351( .i (n3350), .o (n3351) );
  buffer buf_n3491( .i (n3490), .o (n3491) );
  assign n3498 = n3351 & ~n3491 ;
  assign n3499 = n3493 | n3498 ;
  buffer buf_n3500( .i (n3499), .o (n3500) );
  assign n3502 = n3347 | n3500 ;
  buffer buf_n3503( .i (n3502), .o (n3503) );
  buffer buf_n3348( .i (n3347), .o (n3348) );
  buffer buf_n3501( .i (n3500), .o (n3501) );
  assign n3512 = n3348 & n3501 ;
  assign n3513 = n3503 & ~n3512 ;
  buffer buf_n3514( .i (n3513), .o (n3514) );
  assign n3516 = ~n3344 & n3514 ;
  buffer buf_n3517( .i (n3516), .o (n3517) );
  buffer buf_n3345( .i (n3344), .o (n3345) );
  buffer buf_n3515( .i (n3514), .o (n3515) );
  assign n3522 = n3345 & ~n3515 ;
  assign n3523 = n3517 | n3522 ;
  buffer buf_n3524( .i (n3523), .o (n3524) );
  assign n3526 = n3341 | n3524 ;
  buffer buf_n3527( .i (n3526), .o (n3527) );
  buffer buf_n3342( .i (n3341), .o (n3342) );
  buffer buf_n3525( .i (n3524), .o (n3525) );
  assign n3536 = n3342 & n3525 ;
  assign n3537 = n3527 & ~n3536 ;
  buffer buf_n3538( .i (n3537), .o (n3538) );
  assign n3540 = ~n3338 & n3538 ;
  buffer buf_n3541( .i (n3540), .o (n3541) );
  buffer buf_n3339( .i (n3338), .o (n3339) );
  buffer buf_n3539( .i (n3538), .o (n3539) );
  assign n3546 = n3339 & ~n3539 ;
  assign n3547 = n3541 | n3546 ;
  buffer buf_n3548( .i (n3547), .o (n3548) );
  assign n3550 = n3335 | n3548 ;
  buffer buf_n3551( .i (n3550), .o (n3551) );
  buffer buf_n3336( .i (n3335), .o (n3336) );
  buffer buf_n3549( .i (n3548), .o (n3549) );
  assign n3560 = n3336 & n3549 ;
  assign n3561 = n3551 & ~n3560 ;
  buffer buf_n3562( .i (n3561), .o (n3562) );
  assign n3564 = ~n3332 & n3562 ;
  buffer buf_n3565( .i (n3564), .o (n3565) );
  buffer buf_n3333( .i (n3332), .o (n3333) );
  buffer buf_n3563( .i (n3562), .o (n3563) );
  assign n3570 = n3333 & ~n3563 ;
  assign n3571 = n3565 | n3570 ;
  buffer buf_n3572( .i (n3571), .o (n3572) );
  assign n3574 = n3329 | n3572 ;
  buffer buf_n3575( .i (n3574), .o (n3575) );
  buffer buf_n3330( .i (n3329), .o (n3330) );
  buffer buf_n3573( .i (n3572), .o (n3573) );
  assign n3584 = n3330 & n3573 ;
  assign n3585 = n3575 & ~n3584 ;
  buffer buf_n3586( .i (n3585), .o (n3586) );
  assign n3588 = ~n3326 & n3586 ;
  buffer buf_n3589( .i (n3588), .o (n3589) );
  buffer buf_n3327( .i (n3326), .o (n3327) );
  buffer buf_n3587( .i (n3586), .o (n3587) );
  assign n3594 = n3327 & ~n3587 ;
  assign n3595 = n3589 | n3594 ;
  buffer buf_n3596( .i (n3595), .o (n3596) );
  assign n3598 = n3323 | n3596 ;
  buffer buf_n3599( .i (n3598), .o (n3599) );
  buffer buf_n3324( .i (n3323), .o (n3324) );
  buffer buf_n3597( .i (n3596), .o (n3597) );
  assign n3608 = n3324 & n3597 ;
  assign n3609 = n3599 & ~n3608 ;
  buffer buf_n3610( .i (n3609), .o (n3610) );
  assign n3612 = ~n3320 & n3610 ;
  buffer buf_n3613( .i (n3612), .o (n3613) );
  buffer buf_n3321( .i (n3320), .o (n3321) );
  buffer buf_n3611( .i (n3610), .o (n3611) );
  assign n3618 = n3321 & ~n3611 ;
  assign n3619 = n3613 | n3618 ;
  buffer buf_n3620( .i (n3619), .o (n3620) );
  assign n3622 = n3317 | n3620 ;
  buffer buf_n3623( .i (n3622), .o (n3623) );
  buffer buf_n3318( .i (n3317), .o (n3318) );
  buffer buf_n3621( .i (n3620), .o (n3621) );
  assign n3632 = n3318 & n3621 ;
  assign n3633 = n3623 & ~n3632 ;
  buffer buf_n3634( .i (n3633), .o (n3634) );
  assign n3636 = ~n3314 & n3634 ;
  buffer buf_n3637( .i (n3636), .o (n3637) );
  buffer buf_n3315( .i (n3314), .o (n3315) );
  buffer buf_n3635( .i (n3634), .o (n3635) );
  assign n3642 = n3315 & ~n3635 ;
  assign n3643 = n3637 | n3642 ;
  buffer buf_n3644( .i (n3643), .o (n3644) );
  assign n3646 = n3311 | n3644 ;
  buffer buf_n3647( .i (n3646), .o (n3647) );
  buffer buf_n3312( .i (n3311), .o (n3312) );
  buffer buf_n3645( .i (n3644), .o (n3645) );
  assign n3656 = n3312 & n3645 ;
  assign n3657 = n3647 & ~n3656 ;
  buffer buf_n3658( .i (n3657), .o (n3658) );
  assign n3660 = ~n3308 & n3658 ;
  buffer buf_n3661( .i (n3660), .o (n3661) );
  buffer buf_n3309( .i (n3308), .o (n3309) );
  buffer buf_n3659( .i (n3658), .o (n3659) );
  assign n3666 = n3309 & ~n3659 ;
  assign n3667 = n3661 | n3666 ;
  buffer buf_n3668( .i (n3667), .o (n3668) );
  assign n3670 = n3305 | n3668 ;
  buffer buf_n3671( .i (n3670), .o (n3671) );
  buffer buf_n3306( .i (n3305), .o (n3306) );
  buffer buf_n3669( .i (n3668), .o (n3669) );
  assign n3676 = n3306 & n3669 ;
  assign n3677 = n3671 & ~n3676 ;
  buffer buf_n3678( .i (n3677), .o (n3678) );
  assign n3680 = ~n3302 & n3678 ;
  buffer buf_n3681( .i (n3680), .o (n3681) );
  buffer buf_n3303( .i (n3302), .o (n3303) );
  buffer buf_n3679( .i (n3678), .o (n3679) );
  assign n3682 = n3303 & ~n3679 ;
  assign n3683 = n3681 | n3682 ;
  buffer buf_n3672( .i (n3671), .o (n3672) );
  buffer buf_n3673( .i (n3672), .o (n3673) );
  buffer buf_n3674( .i (n3673), .o (n3674) );
  buffer buf_n3675( .i (n3674), .o (n3675) );
  assign n3684 = n3675 & ~n3681 ;
  buffer buf_n3685( .i (n3684), .o (n3685) );
  buffer buf_n3648( .i (n3647), .o (n3648) );
  buffer buf_n3649( .i (n3648), .o (n3649) );
  buffer buf_n3650( .i (n3649), .o (n3650) );
  buffer buf_n3651( .i (n3650), .o (n3651) );
  buffer buf_n3652( .i (n3651), .o (n3652) );
  buffer buf_n3653( .i (n3652), .o (n3653) );
  buffer buf_n3654( .i (n3653), .o (n3654) );
  buffer buf_n3655( .i (n3654), .o (n3655) );
  buffer buf_n3662( .i (n3661), .o (n3662) );
  buffer buf_n3663( .i (n3662), .o (n3663) );
  buffer buf_n3664( .i (n3663), .o (n3664) );
  buffer buf_n3665( .i (n3664), .o (n3665) );
  assign n3687 = n3655 & ~n3665 ;
  buffer buf_n3688( .i (n3687), .o (n3688) );
  assign n3690 = N528 & N69 ;
  buffer buf_n3691( .i (n3690), .o (n3691) );
  buffer buf_n3624( .i (n3623), .o (n3624) );
  buffer buf_n3625( .i (n3624), .o (n3625) );
  buffer buf_n3626( .i (n3625), .o (n3626) );
  buffer buf_n3627( .i (n3626), .o (n3627) );
  buffer buf_n3628( .i (n3627), .o (n3628) );
  buffer buf_n3629( .i (n3628), .o (n3629) );
  buffer buf_n3630( .i (n3629), .o (n3630) );
  buffer buf_n3631( .i (n3630), .o (n3631) );
  buffer buf_n3638( .i (n3637), .o (n3638) );
  buffer buf_n3639( .i (n3638), .o (n3639) );
  buffer buf_n3640( .i (n3639), .o (n3640) );
  buffer buf_n3641( .i (n3640), .o (n3641) );
  assign n3693 = n3631 & ~n3641 ;
  buffer buf_n3694( .i (n3693), .o (n3694) );
  assign n3696 = N511 & N86 ;
  buffer buf_n3697( .i (n3696), .o (n3697) );
  buffer buf_n3600( .i (n3599), .o (n3600) );
  buffer buf_n3601( .i (n3600), .o (n3601) );
  buffer buf_n3602( .i (n3601), .o (n3602) );
  buffer buf_n3603( .i (n3602), .o (n3603) );
  buffer buf_n3604( .i (n3603), .o (n3604) );
  buffer buf_n3605( .i (n3604), .o (n3605) );
  buffer buf_n3606( .i (n3605), .o (n3606) );
  buffer buf_n3607( .i (n3606), .o (n3607) );
  buffer buf_n3614( .i (n3613), .o (n3614) );
  buffer buf_n3615( .i (n3614), .o (n3615) );
  buffer buf_n3616( .i (n3615), .o (n3616) );
  buffer buf_n3617( .i (n3616), .o (n3617) );
  assign n3699 = n3607 & ~n3617 ;
  buffer buf_n3700( .i (n3699), .o (n3700) );
  assign n3702 = N103 & N494 ;
  buffer buf_n3703( .i (n3702), .o (n3703) );
  buffer buf_n3576( .i (n3575), .o (n3576) );
  buffer buf_n3577( .i (n3576), .o (n3577) );
  buffer buf_n3578( .i (n3577), .o (n3578) );
  buffer buf_n3579( .i (n3578), .o (n3579) );
  buffer buf_n3580( .i (n3579), .o (n3580) );
  buffer buf_n3581( .i (n3580), .o (n3581) );
  buffer buf_n3582( .i (n3581), .o (n3582) );
  buffer buf_n3583( .i (n3582), .o (n3583) );
  buffer buf_n3590( .i (n3589), .o (n3590) );
  buffer buf_n3591( .i (n3590), .o (n3591) );
  buffer buf_n3592( .i (n3591), .o (n3592) );
  buffer buf_n3593( .i (n3592), .o (n3593) );
  assign n3705 = n3583 & ~n3593 ;
  buffer buf_n3706( .i (n3705), .o (n3706) );
  assign n3708 = N120 & N477 ;
  buffer buf_n3709( .i (n3708), .o (n3709) );
  buffer buf_n3552( .i (n3551), .o (n3552) );
  buffer buf_n3553( .i (n3552), .o (n3553) );
  buffer buf_n3554( .i (n3553), .o (n3554) );
  buffer buf_n3555( .i (n3554), .o (n3555) );
  buffer buf_n3556( .i (n3555), .o (n3556) );
  buffer buf_n3557( .i (n3556), .o (n3557) );
  buffer buf_n3558( .i (n3557), .o (n3558) );
  buffer buf_n3559( .i (n3558), .o (n3559) );
  buffer buf_n3566( .i (n3565), .o (n3566) );
  buffer buf_n3567( .i (n3566), .o (n3567) );
  buffer buf_n3568( .i (n3567), .o (n3568) );
  buffer buf_n3569( .i (n3568), .o (n3569) );
  assign n3711 = n3559 & ~n3569 ;
  buffer buf_n3712( .i (n3711), .o (n3712) );
  assign n3714 = N137 & N460 ;
  buffer buf_n3715( .i (n3714), .o (n3715) );
  buffer buf_n3528( .i (n3527), .o (n3528) );
  buffer buf_n3529( .i (n3528), .o (n3529) );
  buffer buf_n3530( .i (n3529), .o (n3530) );
  buffer buf_n3531( .i (n3530), .o (n3531) );
  buffer buf_n3532( .i (n3531), .o (n3532) );
  buffer buf_n3533( .i (n3532), .o (n3533) );
  buffer buf_n3534( .i (n3533), .o (n3534) );
  buffer buf_n3535( .i (n3534), .o (n3535) );
  buffer buf_n3542( .i (n3541), .o (n3542) );
  buffer buf_n3543( .i (n3542), .o (n3543) );
  buffer buf_n3544( .i (n3543), .o (n3544) );
  buffer buf_n3545( .i (n3544), .o (n3545) );
  assign n3717 = n3535 & ~n3545 ;
  buffer buf_n3718( .i (n3717), .o (n3718) );
  assign n3720 = N154 & N443 ;
  buffer buf_n3721( .i (n3720), .o (n3721) );
  buffer buf_n3504( .i (n3503), .o (n3504) );
  buffer buf_n3505( .i (n3504), .o (n3505) );
  buffer buf_n3506( .i (n3505), .o (n3506) );
  buffer buf_n3507( .i (n3506), .o (n3507) );
  buffer buf_n3508( .i (n3507), .o (n3508) );
  buffer buf_n3509( .i (n3508), .o (n3509) );
  buffer buf_n3510( .i (n3509), .o (n3510) );
  buffer buf_n3511( .i (n3510), .o (n3511) );
  buffer buf_n3518( .i (n3517), .o (n3518) );
  buffer buf_n3519( .i (n3518), .o (n3519) );
  buffer buf_n3520( .i (n3519), .o (n3520) );
  buffer buf_n3521( .i (n3520), .o (n3521) );
  assign n3723 = n3511 & ~n3521 ;
  buffer buf_n3724( .i (n3723), .o (n3724) );
  assign n3726 = N171 & N426 ;
  buffer buf_n3727( .i (n3726), .o (n3727) );
  buffer buf_n3480( .i (n3479), .o (n3480) );
  buffer buf_n3481( .i (n3480), .o (n3481) );
  buffer buf_n3482( .i (n3481), .o (n3482) );
  buffer buf_n3483( .i (n3482), .o (n3483) );
  buffer buf_n3484( .i (n3483), .o (n3484) );
  buffer buf_n3485( .i (n3484), .o (n3485) );
  buffer buf_n3486( .i (n3485), .o (n3486) );
  buffer buf_n3487( .i (n3486), .o (n3487) );
  buffer buf_n3494( .i (n3493), .o (n3494) );
  buffer buf_n3495( .i (n3494), .o (n3495) );
  buffer buf_n3496( .i (n3495), .o (n3496) );
  buffer buf_n3497( .i (n3496), .o (n3497) );
  assign n3729 = n3487 & ~n3497 ;
  buffer buf_n3730( .i (n3729), .o (n3730) );
  assign n3732 = N188 & N409 ;
  buffer buf_n3733( .i (n3732), .o (n3733) );
  buffer buf_n3456( .i (n3455), .o (n3456) );
  buffer buf_n3457( .i (n3456), .o (n3457) );
  buffer buf_n3458( .i (n3457), .o (n3458) );
  buffer buf_n3459( .i (n3458), .o (n3459) );
  buffer buf_n3460( .i (n3459), .o (n3460) );
  buffer buf_n3461( .i (n3460), .o (n3461) );
  buffer buf_n3462( .i (n3461), .o (n3462) );
  buffer buf_n3463( .i (n3462), .o (n3463) );
  buffer buf_n3470( .i (n3469), .o (n3470) );
  buffer buf_n3471( .i (n3470), .o (n3471) );
  buffer buf_n3472( .i (n3471), .o (n3472) );
  buffer buf_n3473( .i (n3472), .o (n3473) );
  assign n3735 = n3463 & ~n3473 ;
  buffer buf_n3736( .i (n3735), .o (n3736) );
  assign n3738 = N205 & N392 ;
  buffer buf_n3739( .i (n3738), .o (n3739) );
  buffer buf_n3432( .i (n3431), .o (n3432) );
  buffer buf_n3433( .i (n3432), .o (n3433) );
  buffer buf_n3434( .i (n3433), .o (n3434) );
  buffer buf_n3435( .i (n3434), .o (n3435) );
  buffer buf_n3436( .i (n3435), .o (n3436) );
  buffer buf_n3437( .i (n3436), .o (n3437) );
  buffer buf_n3438( .i (n3437), .o (n3438) );
  buffer buf_n3439( .i (n3438), .o (n3439) );
  buffer buf_n3446( .i (n3445), .o (n3446) );
  buffer buf_n3447( .i (n3446), .o (n3447) );
  buffer buf_n3448( .i (n3447), .o (n3448) );
  buffer buf_n3449( .i (n3448), .o (n3449) );
  assign n3741 = n3439 & ~n3449 ;
  buffer buf_n3742( .i (n3741), .o (n3742) );
  assign n3744 = N222 & N375 ;
  buffer buf_n3745( .i (n3744), .o (n3745) );
  buffer buf_n3408( .i (n3407), .o (n3408) );
  buffer buf_n3409( .i (n3408), .o (n3409) );
  buffer buf_n3410( .i (n3409), .o (n3410) );
  buffer buf_n3411( .i (n3410), .o (n3411) );
  buffer buf_n3412( .i (n3411), .o (n3412) );
  buffer buf_n3413( .i (n3412), .o (n3413) );
  buffer buf_n3414( .i (n3413), .o (n3414) );
  buffer buf_n3415( .i (n3414), .o (n3415) );
  buffer buf_n3422( .i (n3421), .o (n3422) );
  buffer buf_n3423( .i (n3422), .o (n3423) );
  buffer buf_n3424( .i (n3423), .o (n3424) );
  buffer buf_n3425( .i (n3424), .o (n3425) );
  assign n3747 = n3415 & ~n3425 ;
  buffer buf_n3748( .i (n3747), .o (n3748) );
  assign n3750 = N239 & N358 ;
  buffer buf_n3751( .i (n3750), .o (n3751) );
  assign n3753 = N256 & N341 ;
  buffer buf_n3754( .i (n3753), .o (n3754) );
  buffer buf_n3384( .i (n3383), .o (n3384) );
  buffer buf_n3385( .i (n3384), .o (n3385) );
  buffer buf_n3386( .i (n3385), .o (n3386) );
  buffer buf_n3387( .i (n3386), .o (n3387) );
  buffer buf_n3388( .i (n3387), .o (n3388) );
  buffer buf_n3389( .i (n3388), .o (n3389) );
  buffer buf_n3390( .i (n3389), .o (n3390) );
  buffer buf_n3391( .i (n3390), .o (n3391) );
  buffer buf_n3398( .i (n3397), .o (n3398) );
  buffer buf_n3399( .i (n3398), .o (n3399) );
  buffer buf_n3400( .i (n3399), .o (n3400) );
  buffer buf_n3401( .i (n3400), .o (n3401) );
  assign n3756 = n3391 & ~n3401 ;
  buffer buf_n3757( .i (n3756), .o (n3757) );
  assign n3759 = n3754 | n3757 ;
  buffer buf_n3760( .i (n3759), .o (n3760) );
  buffer buf_n3755( .i (n3754), .o (n3755) );
  buffer buf_n3758( .i (n3757), .o (n3758) );
  assign n3769 = n3755 & n3758 ;
  assign n3770 = n3760 & ~n3769 ;
  buffer buf_n3771( .i (n3770), .o (n3771) );
  assign n3773 = ~n3751 & n3771 ;
  buffer buf_n3774( .i (n3773), .o (n3774) );
  buffer buf_n3752( .i (n3751), .o (n3752) );
  buffer buf_n3772( .i (n3771), .o (n3772) );
  assign n3779 = n3752 & ~n3772 ;
  assign n3780 = n3774 | n3779 ;
  buffer buf_n3781( .i (n3780), .o (n3781) );
  assign n3783 = n3748 | n3781 ;
  buffer buf_n3784( .i (n3783), .o (n3784) );
  buffer buf_n3749( .i (n3748), .o (n3749) );
  buffer buf_n3782( .i (n3781), .o (n3782) );
  assign n3793 = n3749 & n3782 ;
  assign n3794 = n3784 & ~n3793 ;
  buffer buf_n3795( .i (n3794), .o (n3795) );
  assign n3797 = ~n3745 & n3795 ;
  buffer buf_n3798( .i (n3797), .o (n3798) );
  buffer buf_n3746( .i (n3745), .o (n3746) );
  buffer buf_n3796( .i (n3795), .o (n3796) );
  assign n3803 = n3746 & ~n3796 ;
  assign n3804 = n3798 | n3803 ;
  buffer buf_n3805( .i (n3804), .o (n3805) );
  assign n3807 = n3742 | n3805 ;
  buffer buf_n3808( .i (n3807), .o (n3808) );
  buffer buf_n3743( .i (n3742), .o (n3743) );
  buffer buf_n3806( .i (n3805), .o (n3806) );
  assign n3817 = n3743 & n3806 ;
  assign n3818 = n3808 & ~n3817 ;
  buffer buf_n3819( .i (n3818), .o (n3819) );
  assign n3821 = ~n3739 & n3819 ;
  buffer buf_n3822( .i (n3821), .o (n3822) );
  buffer buf_n3740( .i (n3739), .o (n3740) );
  buffer buf_n3820( .i (n3819), .o (n3820) );
  assign n3827 = n3740 & ~n3820 ;
  assign n3828 = n3822 | n3827 ;
  buffer buf_n3829( .i (n3828), .o (n3829) );
  assign n3831 = n3736 | n3829 ;
  buffer buf_n3832( .i (n3831), .o (n3832) );
  buffer buf_n3737( .i (n3736), .o (n3737) );
  buffer buf_n3830( .i (n3829), .o (n3830) );
  assign n3841 = n3737 & n3830 ;
  assign n3842 = n3832 & ~n3841 ;
  buffer buf_n3843( .i (n3842), .o (n3843) );
  assign n3845 = ~n3733 & n3843 ;
  buffer buf_n3846( .i (n3845), .o (n3846) );
  buffer buf_n3734( .i (n3733), .o (n3734) );
  buffer buf_n3844( .i (n3843), .o (n3844) );
  assign n3851 = n3734 & ~n3844 ;
  assign n3852 = n3846 | n3851 ;
  buffer buf_n3853( .i (n3852), .o (n3853) );
  assign n3855 = n3730 | n3853 ;
  buffer buf_n3856( .i (n3855), .o (n3856) );
  buffer buf_n3731( .i (n3730), .o (n3731) );
  buffer buf_n3854( .i (n3853), .o (n3854) );
  assign n3865 = n3731 & n3854 ;
  assign n3866 = n3856 & ~n3865 ;
  buffer buf_n3867( .i (n3866), .o (n3867) );
  assign n3869 = ~n3727 & n3867 ;
  buffer buf_n3870( .i (n3869), .o (n3870) );
  buffer buf_n3728( .i (n3727), .o (n3728) );
  buffer buf_n3868( .i (n3867), .o (n3868) );
  assign n3875 = n3728 & ~n3868 ;
  assign n3876 = n3870 | n3875 ;
  buffer buf_n3877( .i (n3876), .o (n3877) );
  assign n3879 = n3724 | n3877 ;
  buffer buf_n3880( .i (n3879), .o (n3880) );
  buffer buf_n3725( .i (n3724), .o (n3725) );
  buffer buf_n3878( .i (n3877), .o (n3878) );
  assign n3889 = n3725 & n3878 ;
  assign n3890 = n3880 & ~n3889 ;
  buffer buf_n3891( .i (n3890), .o (n3891) );
  assign n3893 = ~n3721 & n3891 ;
  buffer buf_n3894( .i (n3893), .o (n3894) );
  buffer buf_n3722( .i (n3721), .o (n3722) );
  buffer buf_n3892( .i (n3891), .o (n3892) );
  assign n3899 = n3722 & ~n3892 ;
  assign n3900 = n3894 | n3899 ;
  buffer buf_n3901( .i (n3900), .o (n3901) );
  assign n3903 = n3718 | n3901 ;
  buffer buf_n3904( .i (n3903), .o (n3904) );
  buffer buf_n3719( .i (n3718), .o (n3719) );
  buffer buf_n3902( .i (n3901), .o (n3902) );
  assign n3913 = n3719 & n3902 ;
  assign n3914 = n3904 & ~n3913 ;
  buffer buf_n3915( .i (n3914), .o (n3915) );
  assign n3917 = ~n3715 & n3915 ;
  buffer buf_n3918( .i (n3917), .o (n3918) );
  buffer buf_n3716( .i (n3715), .o (n3716) );
  buffer buf_n3916( .i (n3915), .o (n3916) );
  assign n3923 = n3716 & ~n3916 ;
  assign n3924 = n3918 | n3923 ;
  buffer buf_n3925( .i (n3924), .o (n3925) );
  assign n3927 = n3712 | n3925 ;
  buffer buf_n3928( .i (n3927), .o (n3928) );
  buffer buf_n3713( .i (n3712), .o (n3713) );
  buffer buf_n3926( .i (n3925), .o (n3926) );
  assign n3937 = n3713 & n3926 ;
  assign n3938 = n3928 & ~n3937 ;
  buffer buf_n3939( .i (n3938), .o (n3939) );
  assign n3941 = ~n3709 & n3939 ;
  buffer buf_n3942( .i (n3941), .o (n3942) );
  buffer buf_n3710( .i (n3709), .o (n3710) );
  buffer buf_n3940( .i (n3939), .o (n3940) );
  assign n3947 = n3710 & ~n3940 ;
  assign n3948 = n3942 | n3947 ;
  buffer buf_n3949( .i (n3948), .o (n3949) );
  assign n3951 = n3706 | n3949 ;
  buffer buf_n3952( .i (n3951), .o (n3952) );
  buffer buf_n3707( .i (n3706), .o (n3707) );
  buffer buf_n3950( .i (n3949), .o (n3950) );
  assign n3961 = n3707 & n3950 ;
  assign n3962 = n3952 & ~n3961 ;
  buffer buf_n3963( .i (n3962), .o (n3963) );
  assign n3965 = ~n3703 & n3963 ;
  buffer buf_n3966( .i (n3965), .o (n3966) );
  buffer buf_n3704( .i (n3703), .o (n3704) );
  buffer buf_n3964( .i (n3963), .o (n3964) );
  assign n3971 = n3704 & ~n3964 ;
  assign n3972 = n3966 | n3971 ;
  buffer buf_n3973( .i (n3972), .o (n3973) );
  assign n3975 = n3700 | n3973 ;
  buffer buf_n3976( .i (n3975), .o (n3976) );
  buffer buf_n3701( .i (n3700), .o (n3701) );
  buffer buf_n3974( .i (n3973), .o (n3974) );
  assign n3985 = n3701 & n3974 ;
  assign n3986 = n3976 & ~n3985 ;
  buffer buf_n3987( .i (n3986), .o (n3987) );
  assign n3989 = ~n3697 & n3987 ;
  buffer buf_n3990( .i (n3989), .o (n3990) );
  buffer buf_n3698( .i (n3697), .o (n3698) );
  buffer buf_n3988( .i (n3987), .o (n3988) );
  assign n3995 = n3698 & ~n3988 ;
  assign n3996 = n3990 | n3995 ;
  buffer buf_n3997( .i (n3996), .o (n3997) );
  assign n3999 = n3694 | n3997 ;
  buffer buf_n4000( .i (n3999), .o (n4000) );
  buffer buf_n3695( .i (n3694), .o (n3695) );
  buffer buf_n3998( .i (n3997), .o (n3998) );
  assign n4009 = n3695 & n3998 ;
  assign n4010 = n4000 & ~n4009 ;
  buffer buf_n4011( .i (n4010), .o (n4011) );
  assign n4013 = ~n3691 & n4011 ;
  buffer buf_n4014( .i (n4013), .o (n4014) );
  buffer buf_n3692( .i (n3691), .o (n3692) );
  buffer buf_n4012( .i (n4011), .o (n4012) );
  assign n4019 = n3692 & ~n4012 ;
  assign n4020 = n4014 | n4019 ;
  buffer buf_n4021( .i (n4020), .o (n4021) );
  assign n4023 = n3688 | n4021 ;
  buffer buf_n4024( .i (n4023), .o (n4024) );
  buffer buf_n3689( .i (n3688), .o (n3689) );
  buffer buf_n4022( .i (n4021), .o (n4022) );
  assign n4029 = n3689 & n4022 ;
  assign n4030 = n4024 & ~n4029 ;
  buffer buf_n4031( .i (n4030), .o (n4031) );
  assign n4033 = ~n3685 & n4031 ;
  buffer buf_n4034( .i (n4033), .o (n4034) );
  buffer buf_n3686( .i (n3685), .o (n3686) );
  buffer buf_n4032( .i (n4031), .o (n4032) );
  assign n4035 = n3686 & ~n4032 ;
  assign n4036 = n4034 | n4035 ;
  buffer buf_n4025( .i (n4024), .o (n4025) );
  buffer buf_n4026( .i (n4025), .o (n4026) );
  buffer buf_n4027( .i (n4026), .o (n4027) );
  buffer buf_n4028( .i (n4027), .o (n4028) );
  assign n4037 = n4028 & ~n4034 ;
  buffer buf_n4038( .i (n4037), .o (n4038) );
  buffer buf_n4001( .i (n4000), .o (n4001) );
  buffer buf_n4002( .i (n4001), .o (n4002) );
  buffer buf_n4003( .i (n4002), .o (n4003) );
  buffer buf_n4004( .i (n4003), .o (n4004) );
  buffer buf_n4005( .i (n4004), .o (n4005) );
  buffer buf_n4006( .i (n4005), .o (n4006) );
  buffer buf_n4007( .i (n4006), .o (n4007) );
  buffer buf_n4008( .i (n4007), .o (n4008) );
  buffer buf_n4015( .i (n4014), .o (n4015) );
  buffer buf_n4016( .i (n4015), .o (n4016) );
  buffer buf_n4017( .i (n4016), .o (n4017) );
  buffer buf_n4018( .i (n4017), .o (n4018) );
  assign n4040 = n4008 & ~n4018 ;
  buffer buf_n4041( .i (n4040), .o (n4041) );
  assign n4043 = N528 & N86 ;
  buffer buf_n4044( .i (n4043), .o (n4044) );
  buffer buf_n3977( .i (n3976), .o (n3977) );
  buffer buf_n3978( .i (n3977), .o (n3978) );
  buffer buf_n3979( .i (n3978), .o (n3979) );
  buffer buf_n3980( .i (n3979), .o (n3980) );
  buffer buf_n3981( .i (n3980), .o (n3981) );
  buffer buf_n3982( .i (n3981), .o (n3982) );
  buffer buf_n3983( .i (n3982), .o (n3983) );
  buffer buf_n3984( .i (n3983), .o (n3984) );
  buffer buf_n3991( .i (n3990), .o (n3991) );
  buffer buf_n3992( .i (n3991), .o (n3992) );
  buffer buf_n3993( .i (n3992), .o (n3993) );
  buffer buf_n3994( .i (n3993), .o (n3994) );
  assign n4046 = n3984 & ~n3994 ;
  buffer buf_n4047( .i (n4046), .o (n4047) );
  assign n4049 = N103 & N511 ;
  buffer buf_n4050( .i (n4049), .o (n4050) );
  buffer buf_n3953( .i (n3952), .o (n3953) );
  buffer buf_n3954( .i (n3953), .o (n3954) );
  buffer buf_n3955( .i (n3954), .o (n3955) );
  buffer buf_n3956( .i (n3955), .o (n3956) );
  buffer buf_n3957( .i (n3956), .o (n3957) );
  buffer buf_n3958( .i (n3957), .o (n3958) );
  buffer buf_n3959( .i (n3958), .o (n3959) );
  buffer buf_n3960( .i (n3959), .o (n3960) );
  buffer buf_n3967( .i (n3966), .o (n3967) );
  buffer buf_n3968( .i (n3967), .o (n3968) );
  buffer buf_n3969( .i (n3968), .o (n3969) );
  buffer buf_n3970( .i (n3969), .o (n3970) );
  assign n4052 = n3960 & ~n3970 ;
  buffer buf_n4053( .i (n4052), .o (n4053) );
  assign n4055 = N120 & N494 ;
  buffer buf_n4056( .i (n4055), .o (n4056) );
  buffer buf_n3929( .i (n3928), .o (n3929) );
  buffer buf_n3930( .i (n3929), .o (n3930) );
  buffer buf_n3931( .i (n3930), .o (n3931) );
  buffer buf_n3932( .i (n3931), .o (n3932) );
  buffer buf_n3933( .i (n3932), .o (n3933) );
  buffer buf_n3934( .i (n3933), .o (n3934) );
  buffer buf_n3935( .i (n3934), .o (n3935) );
  buffer buf_n3936( .i (n3935), .o (n3936) );
  buffer buf_n3943( .i (n3942), .o (n3943) );
  buffer buf_n3944( .i (n3943), .o (n3944) );
  buffer buf_n3945( .i (n3944), .o (n3945) );
  buffer buf_n3946( .i (n3945), .o (n3946) );
  assign n4058 = n3936 & ~n3946 ;
  buffer buf_n4059( .i (n4058), .o (n4059) );
  assign n4061 = N137 & N477 ;
  buffer buf_n4062( .i (n4061), .o (n4062) );
  buffer buf_n3905( .i (n3904), .o (n3905) );
  buffer buf_n3906( .i (n3905), .o (n3906) );
  buffer buf_n3907( .i (n3906), .o (n3907) );
  buffer buf_n3908( .i (n3907), .o (n3908) );
  buffer buf_n3909( .i (n3908), .o (n3909) );
  buffer buf_n3910( .i (n3909), .o (n3910) );
  buffer buf_n3911( .i (n3910), .o (n3911) );
  buffer buf_n3912( .i (n3911), .o (n3912) );
  buffer buf_n3919( .i (n3918), .o (n3919) );
  buffer buf_n3920( .i (n3919), .o (n3920) );
  buffer buf_n3921( .i (n3920), .o (n3921) );
  buffer buf_n3922( .i (n3921), .o (n3922) );
  assign n4064 = n3912 & ~n3922 ;
  buffer buf_n4065( .i (n4064), .o (n4065) );
  assign n4067 = N154 & N460 ;
  buffer buf_n4068( .i (n4067), .o (n4068) );
  buffer buf_n3881( .i (n3880), .o (n3881) );
  buffer buf_n3882( .i (n3881), .o (n3882) );
  buffer buf_n3883( .i (n3882), .o (n3883) );
  buffer buf_n3884( .i (n3883), .o (n3884) );
  buffer buf_n3885( .i (n3884), .o (n3885) );
  buffer buf_n3886( .i (n3885), .o (n3886) );
  buffer buf_n3887( .i (n3886), .o (n3887) );
  buffer buf_n3888( .i (n3887), .o (n3888) );
  buffer buf_n3895( .i (n3894), .o (n3895) );
  buffer buf_n3896( .i (n3895), .o (n3896) );
  buffer buf_n3897( .i (n3896), .o (n3897) );
  buffer buf_n3898( .i (n3897), .o (n3898) );
  assign n4070 = n3888 & ~n3898 ;
  buffer buf_n4071( .i (n4070), .o (n4071) );
  assign n4073 = N171 & N443 ;
  buffer buf_n4074( .i (n4073), .o (n4074) );
  buffer buf_n3857( .i (n3856), .o (n3857) );
  buffer buf_n3858( .i (n3857), .o (n3858) );
  buffer buf_n3859( .i (n3858), .o (n3859) );
  buffer buf_n3860( .i (n3859), .o (n3860) );
  buffer buf_n3861( .i (n3860), .o (n3861) );
  buffer buf_n3862( .i (n3861), .o (n3862) );
  buffer buf_n3863( .i (n3862), .o (n3863) );
  buffer buf_n3864( .i (n3863), .o (n3864) );
  buffer buf_n3871( .i (n3870), .o (n3871) );
  buffer buf_n3872( .i (n3871), .o (n3872) );
  buffer buf_n3873( .i (n3872), .o (n3873) );
  buffer buf_n3874( .i (n3873), .o (n3874) );
  assign n4076 = n3864 & ~n3874 ;
  buffer buf_n4077( .i (n4076), .o (n4077) );
  assign n4079 = N188 & N426 ;
  buffer buf_n4080( .i (n4079), .o (n4080) );
  buffer buf_n3833( .i (n3832), .o (n3833) );
  buffer buf_n3834( .i (n3833), .o (n3834) );
  buffer buf_n3835( .i (n3834), .o (n3835) );
  buffer buf_n3836( .i (n3835), .o (n3836) );
  buffer buf_n3837( .i (n3836), .o (n3837) );
  buffer buf_n3838( .i (n3837), .o (n3838) );
  buffer buf_n3839( .i (n3838), .o (n3839) );
  buffer buf_n3840( .i (n3839), .o (n3840) );
  buffer buf_n3847( .i (n3846), .o (n3847) );
  buffer buf_n3848( .i (n3847), .o (n3848) );
  buffer buf_n3849( .i (n3848), .o (n3849) );
  buffer buf_n3850( .i (n3849), .o (n3850) );
  assign n4082 = n3840 & ~n3850 ;
  buffer buf_n4083( .i (n4082), .o (n4083) );
  assign n4085 = N205 & N409 ;
  buffer buf_n4086( .i (n4085), .o (n4086) );
  buffer buf_n3809( .i (n3808), .o (n3809) );
  buffer buf_n3810( .i (n3809), .o (n3810) );
  buffer buf_n3811( .i (n3810), .o (n3811) );
  buffer buf_n3812( .i (n3811), .o (n3812) );
  buffer buf_n3813( .i (n3812), .o (n3813) );
  buffer buf_n3814( .i (n3813), .o (n3814) );
  buffer buf_n3815( .i (n3814), .o (n3815) );
  buffer buf_n3816( .i (n3815), .o (n3816) );
  buffer buf_n3823( .i (n3822), .o (n3823) );
  buffer buf_n3824( .i (n3823), .o (n3824) );
  buffer buf_n3825( .i (n3824), .o (n3825) );
  buffer buf_n3826( .i (n3825), .o (n3826) );
  assign n4088 = n3816 & ~n3826 ;
  buffer buf_n4089( .i (n4088), .o (n4089) );
  assign n4091 = N222 & N392 ;
  buffer buf_n4092( .i (n4091), .o (n4092) );
  buffer buf_n3785( .i (n3784), .o (n3785) );
  buffer buf_n3786( .i (n3785), .o (n3786) );
  buffer buf_n3787( .i (n3786), .o (n3787) );
  buffer buf_n3788( .i (n3787), .o (n3788) );
  buffer buf_n3789( .i (n3788), .o (n3789) );
  buffer buf_n3790( .i (n3789), .o (n3790) );
  buffer buf_n3791( .i (n3790), .o (n3791) );
  buffer buf_n3792( .i (n3791), .o (n3792) );
  buffer buf_n3799( .i (n3798), .o (n3799) );
  buffer buf_n3800( .i (n3799), .o (n3800) );
  buffer buf_n3801( .i (n3800), .o (n3801) );
  buffer buf_n3802( .i (n3801), .o (n3802) );
  assign n4094 = n3792 & ~n3802 ;
  buffer buf_n4095( .i (n4094), .o (n4095) );
  assign n4097 = N239 & N375 ;
  buffer buf_n4098( .i (n4097), .o (n4098) );
  assign n4100 = N256 & N358 ;
  buffer buf_n4101( .i (n4100), .o (n4101) );
  buffer buf_n3761( .i (n3760), .o (n3761) );
  buffer buf_n3762( .i (n3761), .o (n3762) );
  buffer buf_n3763( .i (n3762), .o (n3763) );
  buffer buf_n3764( .i (n3763), .o (n3764) );
  buffer buf_n3765( .i (n3764), .o (n3765) );
  buffer buf_n3766( .i (n3765), .o (n3766) );
  buffer buf_n3767( .i (n3766), .o (n3767) );
  buffer buf_n3768( .i (n3767), .o (n3768) );
  buffer buf_n3775( .i (n3774), .o (n3775) );
  buffer buf_n3776( .i (n3775), .o (n3776) );
  buffer buf_n3777( .i (n3776), .o (n3777) );
  buffer buf_n3778( .i (n3777), .o (n3778) );
  assign n4103 = n3768 & ~n3778 ;
  buffer buf_n4104( .i (n4103), .o (n4104) );
  assign n4106 = n4101 | n4104 ;
  buffer buf_n4107( .i (n4106), .o (n4107) );
  buffer buf_n4102( .i (n4101), .o (n4102) );
  buffer buf_n4105( .i (n4104), .o (n4105) );
  assign n4116 = n4102 & n4105 ;
  assign n4117 = n4107 & ~n4116 ;
  buffer buf_n4118( .i (n4117), .o (n4118) );
  assign n4120 = ~n4098 & n4118 ;
  buffer buf_n4121( .i (n4120), .o (n4121) );
  buffer buf_n4099( .i (n4098), .o (n4099) );
  buffer buf_n4119( .i (n4118), .o (n4119) );
  assign n4126 = n4099 & ~n4119 ;
  assign n4127 = n4121 | n4126 ;
  buffer buf_n4128( .i (n4127), .o (n4128) );
  assign n4130 = n4095 | n4128 ;
  buffer buf_n4131( .i (n4130), .o (n4131) );
  buffer buf_n4096( .i (n4095), .o (n4096) );
  buffer buf_n4129( .i (n4128), .o (n4129) );
  assign n4140 = n4096 & n4129 ;
  assign n4141 = n4131 & ~n4140 ;
  buffer buf_n4142( .i (n4141), .o (n4142) );
  assign n4144 = ~n4092 & n4142 ;
  buffer buf_n4145( .i (n4144), .o (n4145) );
  buffer buf_n4093( .i (n4092), .o (n4093) );
  buffer buf_n4143( .i (n4142), .o (n4143) );
  assign n4150 = n4093 & ~n4143 ;
  assign n4151 = n4145 | n4150 ;
  buffer buf_n4152( .i (n4151), .o (n4152) );
  assign n4154 = n4089 | n4152 ;
  buffer buf_n4155( .i (n4154), .o (n4155) );
  buffer buf_n4090( .i (n4089), .o (n4090) );
  buffer buf_n4153( .i (n4152), .o (n4153) );
  assign n4164 = n4090 & n4153 ;
  assign n4165 = n4155 & ~n4164 ;
  buffer buf_n4166( .i (n4165), .o (n4166) );
  assign n4168 = ~n4086 & n4166 ;
  buffer buf_n4169( .i (n4168), .o (n4169) );
  buffer buf_n4087( .i (n4086), .o (n4087) );
  buffer buf_n4167( .i (n4166), .o (n4167) );
  assign n4174 = n4087 & ~n4167 ;
  assign n4175 = n4169 | n4174 ;
  buffer buf_n4176( .i (n4175), .o (n4176) );
  assign n4178 = n4083 | n4176 ;
  buffer buf_n4179( .i (n4178), .o (n4179) );
  buffer buf_n4084( .i (n4083), .o (n4084) );
  buffer buf_n4177( .i (n4176), .o (n4177) );
  assign n4188 = n4084 & n4177 ;
  assign n4189 = n4179 & ~n4188 ;
  buffer buf_n4190( .i (n4189), .o (n4190) );
  assign n4192 = ~n4080 & n4190 ;
  buffer buf_n4193( .i (n4192), .o (n4193) );
  buffer buf_n4081( .i (n4080), .o (n4081) );
  buffer buf_n4191( .i (n4190), .o (n4191) );
  assign n4198 = n4081 & ~n4191 ;
  assign n4199 = n4193 | n4198 ;
  buffer buf_n4200( .i (n4199), .o (n4200) );
  assign n4202 = n4077 | n4200 ;
  buffer buf_n4203( .i (n4202), .o (n4203) );
  buffer buf_n4078( .i (n4077), .o (n4078) );
  buffer buf_n4201( .i (n4200), .o (n4201) );
  assign n4212 = n4078 & n4201 ;
  assign n4213 = n4203 & ~n4212 ;
  buffer buf_n4214( .i (n4213), .o (n4214) );
  assign n4216 = ~n4074 & n4214 ;
  buffer buf_n4217( .i (n4216), .o (n4217) );
  buffer buf_n4075( .i (n4074), .o (n4075) );
  buffer buf_n4215( .i (n4214), .o (n4215) );
  assign n4222 = n4075 & ~n4215 ;
  assign n4223 = n4217 | n4222 ;
  buffer buf_n4224( .i (n4223), .o (n4224) );
  assign n4226 = n4071 | n4224 ;
  buffer buf_n4227( .i (n4226), .o (n4227) );
  buffer buf_n4072( .i (n4071), .o (n4072) );
  buffer buf_n4225( .i (n4224), .o (n4225) );
  assign n4236 = n4072 & n4225 ;
  assign n4237 = n4227 & ~n4236 ;
  buffer buf_n4238( .i (n4237), .o (n4238) );
  assign n4240 = ~n4068 & n4238 ;
  buffer buf_n4241( .i (n4240), .o (n4241) );
  buffer buf_n4069( .i (n4068), .o (n4069) );
  buffer buf_n4239( .i (n4238), .o (n4239) );
  assign n4246 = n4069 & ~n4239 ;
  assign n4247 = n4241 | n4246 ;
  buffer buf_n4248( .i (n4247), .o (n4248) );
  assign n4250 = n4065 | n4248 ;
  buffer buf_n4251( .i (n4250), .o (n4251) );
  buffer buf_n4066( .i (n4065), .o (n4066) );
  buffer buf_n4249( .i (n4248), .o (n4249) );
  assign n4260 = n4066 & n4249 ;
  assign n4261 = n4251 & ~n4260 ;
  buffer buf_n4262( .i (n4261), .o (n4262) );
  assign n4264 = ~n4062 & n4262 ;
  buffer buf_n4265( .i (n4264), .o (n4265) );
  buffer buf_n4063( .i (n4062), .o (n4063) );
  buffer buf_n4263( .i (n4262), .o (n4263) );
  assign n4270 = n4063 & ~n4263 ;
  assign n4271 = n4265 | n4270 ;
  buffer buf_n4272( .i (n4271), .o (n4272) );
  assign n4274 = n4059 | n4272 ;
  buffer buf_n4275( .i (n4274), .o (n4275) );
  buffer buf_n4060( .i (n4059), .o (n4060) );
  buffer buf_n4273( .i (n4272), .o (n4273) );
  assign n4284 = n4060 & n4273 ;
  assign n4285 = n4275 & ~n4284 ;
  buffer buf_n4286( .i (n4285), .o (n4286) );
  assign n4288 = ~n4056 & n4286 ;
  buffer buf_n4289( .i (n4288), .o (n4289) );
  buffer buf_n4057( .i (n4056), .o (n4057) );
  buffer buf_n4287( .i (n4286), .o (n4287) );
  assign n4294 = n4057 & ~n4287 ;
  assign n4295 = n4289 | n4294 ;
  buffer buf_n4296( .i (n4295), .o (n4296) );
  assign n4298 = n4053 | n4296 ;
  buffer buf_n4299( .i (n4298), .o (n4299) );
  buffer buf_n4054( .i (n4053), .o (n4054) );
  buffer buf_n4297( .i (n4296), .o (n4297) );
  assign n4308 = n4054 & n4297 ;
  assign n4309 = n4299 & ~n4308 ;
  buffer buf_n4310( .i (n4309), .o (n4310) );
  assign n4312 = ~n4050 & n4310 ;
  buffer buf_n4313( .i (n4312), .o (n4313) );
  buffer buf_n4051( .i (n4050), .o (n4051) );
  buffer buf_n4311( .i (n4310), .o (n4311) );
  assign n4318 = n4051 & ~n4311 ;
  assign n4319 = n4313 | n4318 ;
  buffer buf_n4320( .i (n4319), .o (n4320) );
  assign n4322 = n4047 | n4320 ;
  buffer buf_n4323( .i (n4322), .o (n4323) );
  buffer buf_n4048( .i (n4047), .o (n4048) );
  buffer buf_n4321( .i (n4320), .o (n4321) );
  assign n4332 = n4048 & n4321 ;
  assign n4333 = n4323 & ~n4332 ;
  buffer buf_n4334( .i (n4333), .o (n4334) );
  assign n4336 = ~n4044 & n4334 ;
  buffer buf_n4337( .i (n4336), .o (n4337) );
  buffer buf_n4045( .i (n4044), .o (n4045) );
  buffer buf_n4335( .i (n4334), .o (n4335) );
  assign n4342 = n4045 & ~n4335 ;
  assign n4343 = n4337 | n4342 ;
  buffer buf_n4344( .i (n4343), .o (n4344) );
  assign n4346 = n4041 | n4344 ;
  buffer buf_n4347( .i (n4346), .o (n4347) );
  buffer buf_n4042( .i (n4041), .o (n4042) );
  buffer buf_n4345( .i (n4344), .o (n4345) );
  assign n4352 = n4042 & n4345 ;
  assign n4353 = n4347 & ~n4352 ;
  buffer buf_n4354( .i (n4353), .o (n4354) );
  assign n4356 = ~n4038 & n4354 ;
  buffer buf_n4357( .i (n4356), .o (n4357) );
  buffer buf_n4039( .i (n4038), .o (n4039) );
  buffer buf_n4355( .i (n4354), .o (n4355) );
  assign n4358 = n4039 & ~n4355 ;
  assign n4359 = n4357 | n4358 ;
  buffer buf_n4348( .i (n4347), .o (n4348) );
  buffer buf_n4349( .i (n4348), .o (n4349) );
  buffer buf_n4350( .i (n4349), .o (n4350) );
  buffer buf_n4351( .i (n4350), .o (n4351) );
  assign n4360 = n4351 & ~n4357 ;
  buffer buf_n4361( .i (n4360), .o (n4361) );
  buffer buf_n4324( .i (n4323), .o (n4324) );
  buffer buf_n4325( .i (n4324), .o (n4325) );
  buffer buf_n4326( .i (n4325), .o (n4326) );
  buffer buf_n4327( .i (n4326), .o (n4327) );
  buffer buf_n4328( .i (n4327), .o (n4328) );
  buffer buf_n4329( .i (n4328), .o (n4329) );
  buffer buf_n4330( .i (n4329), .o (n4330) );
  buffer buf_n4331( .i (n4330), .o (n4331) );
  buffer buf_n4338( .i (n4337), .o (n4338) );
  buffer buf_n4339( .i (n4338), .o (n4339) );
  buffer buf_n4340( .i (n4339), .o (n4340) );
  buffer buf_n4341( .i (n4340), .o (n4341) );
  assign n4363 = n4331 & ~n4341 ;
  buffer buf_n4364( .i (n4363), .o (n4364) );
  assign n4366 = N103 & N528 ;
  buffer buf_n4367( .i (n4366), .o (n4367) );
  buffer buf_n4300( .i (n4299), .o (n4300) );
  buffer buf_n4301( .i (n4300), .o (n4301) );
  buffer buf_n4302( .i (n4301), .o (n4302) );
  buffer buf_n4303( .i (n4302), .o (n4303) );
  buffer buf_n4304( .i (n4303), .o (n4304) );
  buffer buf_n4305( .i (n4304), .o (n4305) );
  buffer buf_n4306( .i (n4305), .o (n4306) );
  buffer buf_n4307( .i (n4306), .o (n4307) );
  buffer buf_n4314( .i (n4313), .o (n4314) );
  buffer buf_n4315( .i (n4314), .o (n4315) );
  buffer buf_n4316( .i (n4315), .o (n4316) );
  buffer buf_n4317( .i (n4316), .o (n4317) );
  assign n4369 = n4307 & ~n4317 ;
  buffer buf_n4370( .i (n4369), .o (n4370) );
  assign n4372 = N120 & N511 ;
  buffer buf_n4373( .i (n4372), .o (n4373) );
  buffer buf_n4276( .i (n4275), .o (n4276) );
  buffer buf_n4277( .i (n4276), .o (n4277) );
  buffer buf_n4278( .i (n4277), .o (n4278) );
  buffer buf_n4279( .i (n4278), .o (n4279) );
  buffer buf_n4280( .i (n4279), .o (n4280) );
  buffer buf_n4281( .i (n4280), .o (n4281) );
  buffer buf_n4282( .i (n4281), .o (n4282) );
  buffer buf_n4283( .i (n4282), .o (n4283) );
  buffer buf_n4290( .i (n4289), .o (n4290) );
  buffer buf_n4291( .i (n4290), .o (n4291) );
  buffer buf_n4292( .i (n4291), .o (n4292) );
  buffer buf_n4293( .i (n4292), .o (n4293) );
  assign n4375 = n4283 & ~n4293 ;
  buffer buf_n4376( .i (n4375), .o (n4376) );
  assign n4378 = N137 & N494 ;
  buffer buf_n4379( .i (n4378), .o (n4379) );
  buffer buf_n4252( .i (n4251), .o (n4252) );
  buffer buf_n4253( .i (n4252), .o (n4253) );
  buffer buf_n4254( .i (n4253), .o (n4254) );
  buffer buf_n4255( .i (n4254), .o (n4255) );
  buffer buf_n4256( .i (n4255), .o (n4256) );
  buffer buf_n4257( .i (n4256), .o (n4257) );
  buffer buf_n4258( .i (n4257), .o (n4258) );
  buffer buf_n4259( .i (n4258), .o (n4259) );
  buffer buf_n4266( .i (n4265), .o (n4266) );
  buffer buf_n4267( .i (n4266), .o (n4267) );
  buffer buf_n4268( .i (n4267), .o (n4268) );
  buffer buf_n4269( .i (n4268), .o (n4269) );
  assign n4381 = n4259 & ~n4269 ;
  buffer buf_n4382( .i (n4381), .o (n4382) );
  assign n4384 = N154 & N477 ;
  buffer buf_n4385( .i (n4384), .o (n4385) );
  buffer buf_n4228( .i (n4227), .o (n4228) );
  buffer buf_n4229( .i (n4228), .o (n4229) );
  buffer buf_n4230( .i (n4229), .o (n4230) );
  buffer buf_n4231( .i (n4230), .o (n4231) );
  buffer buf_n4232( .i (n4231), .o (n4232) );
  buffer buf_n4233( .i (n4232), .o (n4233) );
  buffer buf_n4234( .i (n4233), .o (n4234) );
  buffer buf_n4235( .i (n4234), .o (n4235) );
  buffer buf_n4242( .i (n4241), .o (n4242) );
  buffer buf_n4243( .i (n4242), .o (n4243) );
  buffer buf_n4244( .i (n4243), .o (n4244) );
  buffer buf_n4245( .i (n4244), .o (n4245) );
  assign n4387 = n4235 & ~n4245 ;
  buffer buf_n4388( .i (n4387), .o (n4388) );
  assign n4390 = N171 & N460 ;
  buffer buf_n4391( .i (n4390), .o (n4391) );
  buffer buf_n4204( .i (n4203), .o (n4204) );
  buffer buf_n4205( .i (n4204), .o (n4205) );
  buffer buf_n4206( .i (n4205), .o (n4206) );
  buffer buf_n4207( .i (n4206), .o (n4207) );
  buffer buf_n4208( .i (n4207), .o (n4208) );
  buffer buf_n4209( .i (n4208), .o (n4209) );
  buffer buf_n4210( .i (n4209), .o (n4210) );
  buffer buf_n4211( .i (n4210), .o (n4211) );
  buffer buf_n4218( .i (n4217), .o (n4218) );
  buffer buf_n4219( .i (n4218), .o (n4219) );
  buffer buf_n4220( .i (n4219), .o (n4220) );
  buffer buf_n4221( .i (n4220), .o (n4221) );
  assign n4393 = n4211 & ~n4221 ;
  buffer buf_n4394( .i (n4393), .o (n4394) );
  assign n4396 = N188 & N443 ;
  buffer buf_n4397( .i (n4396), .o (n4397) );
  buffer buf_n4180( .i (n4179), .o (n4180) );
  buffer buf_n4181( .i (n4180), .o (n4181) );
  buffer buf_n4182( .i (n4181), .o (n4182) );
  buffer buf_n4183( .i (n4182), .o (n4183) );
  buffer buf_n4184( .i (n4183), .o (n4184) );
  buffer buf_n4185( .i (n4184), .o (n4185) );
  buffer buf_n4186( .i (n4185), .o (n4186) );
  buffer buf_n4187( .i (n4186), .o (n4187) );
  buffer buf_n4194( .i (n4193), .o (n4194) );
  buffer buf_n4195( .i (n4194), .o (n4195) );
  buffer buf_n4196( .i (n4195), .o (n4196) );
  buffer buf_n4197( .i (n4196), .o (n4197) );
  assign n4399 = n4187 & ~n4197 ;
  buffer buf_n4400( .i (n4399), .o (n4400) );
  assign n4402 = N205 & N426 ;
  buffer buf_n4403( .i (n4402), .o (n4403) );
  buffer buf_n4156( .i (n4155), .o (n4156) );
  buffer buf_n4157( .i (n4156), .o (n4157) );
  buffer buf_n4158( .i (n4157), .o (n4158) );
  buffer buf_n4159( .i (n4158), .o (n4159) );
  buffer buf_n4160( .i (n4159), .o (n4160) );
  buffer buf_n4161( .i (n4160), .o (n4161) );
  buffer buf_n4162( .i (n4161), .o (n4162) );
  buffer buf_n4163( .i (n4162), .o (n4163) );
  buffer buf_n4170( .i (n4169), .o (n4170) );
  buffer buf_n4171( .i (n4170), .o (n4171) );
  buffer buf_n4172( .i (n4171), .o (n4172) );
  buffer buf_n4173( .i (n4172), .o (n4173) );
  assign n4405 = n4163 & ~n4173 ;
  buffer buf_n4406( .i (n4405), .o (n4406) );
  assign n4408 = N222 & N409 ;
  buffer buf_n4409( .i (n4408), .o (n4409) );
  buffer buf_n4132( .i (n4131), .o (n4132) );
  buffer buf_n4133( .i (n4132), .o (n4133) );
  buffer buf_n4134( .i (n4133), .o (n4134) );
  buffer buf_n4135( .i (n4134), .o (n4135) );
  buffer buf_n4136( .i (n4135), .o (n4136) );
  buffer buf_n4137( .i (n4136), .o (n4137) );
  buffer buf_n4138( .i (n4137), .o (n4138) );
  buffer buf_n4139( .i (n4138), .o (n4139) );
  buffer buf_n4146( .i (n4145), .o (n4146) );
  buffer buf_n4147( .i (n4146), .o (n4147) );
  buffer buf_n4148( .i (n4147), .o (n4148) );
  buffer buf_n4149( .i (n4148), .o (n4149) );
  assign n4411 = n4139 & ~n4149 ;
  buffer buf_n4412( .i (n4411), .o (n4412) );
  assign n4414 = N239 & N392 ;
  buffer buf_n4415( .i (n4414), .o (n4415) );
  assign n4417 = N256 & N375 ;
  buffer buf_n4418( .i (n4417), .o (n4418) );
  buffer buf_n4108( .i (n4107), .o (n4108) );
  buffer buf_n4109( .i (n4108), .o (n4109) );
  buffer buf_n4110( .i (n4109), .o (n4110) );
  buffer buf_n4111( .i (n4110), .o (n4111) );
  buffer buf_n4112( .i (n4111), .o (n4112) );
  buffer buf_n4113( .i (n4112), .o (n4113) );
  buffer buf_n4114( .i (n4113), .o (n4114) );
  buffer buf_n4115( .i (n4114), .o (n4115) );
  buffer buf_n4122( .i (n4121), .o (n4122) );
  buffer buf_n4123( .i (n4122), .o (n4123) );
  buffer buf_n4124( .i (n4123), .o (n4124) );
  buffer buf_n4125( .i (n4124), .o (n4125) );
  assign n4420 = n4115 & ~n4125 ;
  buffer buf_n4421( .i (n4420), .o (n4421) );
  assign n4423 = n4418 | n4421 ;
  buffer buf_n4424( .i (n4423), .o (n4424) );
  buffer buf_n4419( .i (n4418), .o (n4419) );
  buffer buf_n4422( .i (n4421), .o (n4422) );
  assign n4433 = n4419 & n4422 ;
  assign n4434 = n4424 & ~n4433 ;
  buffer buf_n4435( .i (n4434), .o (n4435) );
  assign n4437 = ~n4415 & n4435 ;
  buffer buf_n4438( .i (n4437), .o (n4438) );
  buffer buf_n4416( .i (n4415), .o (n4416) );
  buffer buf_n4436( .i (n4435), .o (n4436) );
  assign n4443 = n4416 & ~n4436 ;
  assign n4444 = n4438 | n4443 ;
  buffer buf_n4445( .i (n4444), .o (n4445) );
  assign n4447 = n4412 | n4445 ;
  buffer buf_n4448( .i (n4447), .o (n4448) );
  buffer buf_n4413( .i (n4412), .o (n4413) );
  buffer buf_n4446( .i (n4445), .o (n4446) );
  assign n4457 = n4413 & n4446 ;
  assign n4458 = n4448 & ~n4457 ;
  buffer buf_n4459( .i (n4458), .o (n4459) );
  assign n4461 = ~n4409 & n4459 ;
  buffer buf_n4462( .i (n4461), .o (n4462) );
  buffer buf_n4410( .i (n4409), .o (n4410) );
  buffer buf_n4460( .i (n4459), .o (n4460) );
  assign n4467 = n4410 & ~n4460 ;
  assign n4468 = n4462 | n4467 ;
  buffer buf_n4469( .i (n4468), .o (n4469) );
  assign n4471 = n4406 | n4469 ;
  buffer buf_n4472( .i (n4471), .o (n4472) );
  buffer buf_n4407( .i (n4406), .o (n4407) );
  buffer buf_n4470( .i (n4469), .o (n4470) );
  assign n4481 = n4407 & n4470 ;
  assign n4482 = n4472 & ~n4481 ;
  buffer buf_n4483( .i (n4482), .o (n4483) );
  assign n4485 = ~n4403 & n4483 ;
  buffer buf_n4486( .i (n4485), .o (n4486) );
  buffer buf_n4404( .i (n4403), .o (n4404) );
  buffer buf_n4484( .i (n4483), .o (n4484) );
  assign n4491 = n4404 & ~n4484 ;
  assign n4492 = n4486 | n4491 ;
  buffer buf_n4493( .i (n4492), .o (n4493) );
  assign n4495 = n4400 | n4493 ;
  buffer buf_n4496( .i (n4495), .o (n4496) );
  buffer buf_n4401( .i (n4400), .o (n4401) );
  buffer buf_n4494( .i (n4493), .o (n4494) );
  assign n4505 = n4401 & n4494 ;
  assign n4506 = n4496 & ~n4505 ;
  buffer buf_n4507( .i (n4506), .o (n4507) );
  assign n4509 = ~n4397 & n4507 ;
  buffer buf_n4510( .i (n4509), .o (n4510) );
  buffer buf_n4398( .i (n4397), .o (n4398) );
  buffer buf_n4508( .i (n4507), .o (n4508) );
  assign n4515 = n4398 & ~n4508 ;
  assign n4516 = n4510 | n4515 ;
  buffer buf_n4517( .i (n4516), .o (n4517) );
  assign n4519 = n4394 | n4517 ;
  buffer buf_n4520( .i (n4519), .o (n4520) );
  buffer buf_n4395( .i (n4394), .o (n4395) );
  buffer buf_n4518( .i (n4517), .o (n4518) );
  assign n4529 = n4395 & n4518 ;
  assign n4530 = n4520 & ~n4529 ;
  buffer buf_n4531( .i (n4530), .o (n4531) );
  assign n4533 = ~n4391 & n4531 ;
  buffer buf_n4534( .i (n4533), .o (n4534) );
  buffer buf_n4392( .i (n4391), .o (n4392) );
  buffer buf_n4532( .i (n4531), .o (n4532) );
  assign n4539 = n4392 & ~n4532 ;
  assign n4540 = n4534 | n4539 ;
  buffer buf_n4541( .i (n4540), .o (n4541) );
  assign n4543 = n4388 | n4541 ;
  buffer buf_n4544( .i (n4543), .o (n4544) );
  buffer buf_n4389( .i (n4388), .o (n4389) );
  buffer buf_n4542( .i (n4541), .o (n4542) );
  assign n4553 = n4389 & n4542 ;
  assign n4554 = n4544 & ~n4553 ;
  buffer buf_n4555( .i (n4554), .o (n4555) );
  assign n4557 = ~n4385 & n4555 ;
  buffer buf_n4558( .i (n4557), .o (n4558) );
  buffer buf_n4386( .i (n4385), .o (n4386) );
  buffer buf_n4556( .i (n4555), .o (n4556) );
  assign n4563 = n4386 & ~n4556 ;
  assign n4564 = n4558 | n4563 ;
  buffer buf_n4565( .i (n4564), .o (n4565) );
  assign n4567 = n4382 | n4565 ;
  buffer buf_n4568( .i (n4567), .o (n4568) );
  buffer buf_n4383( .i (n4382), .o (n4383) );
  buffer buf_n4566( .i (n4565), .o (n4566) );
  assign n4577 = n4383 & n4566 ;
  assign n4578 = n4568 & ~n4577 ;
  buffer buf_n4579( .i (n4578), .o (n4579) );
  assign n4581 = ~n4379 & n4579 ;
  buffer buf_n4582( .i (n4581), .o (n4582) );
  buffer buf_n4380( .i (n4379), .o (n4380) );
  buffer buf_n4580( .i (n4579), .o (n4580) );
  assign n4587 = n4380 & ~n4580 ;
  assign n4588 = n4582 | n4587 ;
  buffer buf_n4589( .i (n4588), .o (n4589) );
  assign n4591 = n4376 | n4589 ;
  buffer buf_n4592( .i (n4591), .o (n4592) );
  buffer buf_n4377( .i (n4376), .o (n4377) );
  buffer buf_n4590( .i (n4589), .o (n4590) );
  assign n4601 = n4377 & n4590 ;
  assign n4602 = n4592 & ~n4601 ;
  buffer buf_n4603( .i (n4602), .o (n4603) );
  assign n4605 = ~n4373 & n4603 ;
  buffer buf_n4606( .i (n4605), .o (n4606) );
  buffer buf_n4374( .i (n4373), .o (n4374) );
  buffer buf_n4604( .i (n4603), .o (n4604) );
  assign n4611 = n4374 & ~n4604 ;
  assign n4612 = n4606 | n4611 ;
  buffer buf_n4613( .i (n4612), .o (n4613) );
  assign n4615 = n4370 | n4613 ;
  buffer buf_n4616( .i (n4615), .o (n4616) );
  buffer buf_n4371( .i (n4370), .o (n4371) );
  buffer buf_n4614( .i (n4613), .o (n4614) );
  assign n4625 = n4371 & n4614 ;
  assign n4626 = n4616 & ~n4625 ;
  buffer buf_n4627( .i (n4626), .o (n4627) );
  assign n4629 = ~n4367 & n4627 ;
  buffer buf_n4630( .i (n4629), .o (n4630) );
  buffer buf_n4368( .i (n4367), .o (n4368) );
  buffer buf_n4628( .i (n4627), .o (n4628) );
  assign n4635 = n4368 & ~n4628 ;
  assign n4636 = n4630 | n4635 ;
  buffer buf_n4637( .i (n4636), .o (n4637) );
  assign n4639 = n4364 | n4637 ;
  buffer buf_n4640( .i (n4639), .o (n4640) );
  buffer buf_n4365( .i (n4364), .o (n4365) );
  buffer buf_n4638( .i (n4637), .o (n4638) );
  assign n4645 = n4365 & n4638 ;
  assign n4646 = n4640 & ~n4645 ;
  buffer buf_n4647( .i (n4646), .o (n4647) );
  assign n4649 = ~n4361 & n4647 ;
  buffer buf_n4650( .i (n4649), .o (n4650) );
  buffer buf_n4362( .i (n4361), .o (n4362) );
  buffer buf_n4648( .i (n4647), .o (n4648) );
  assign n4651 = n4362 & ~n4648 ;
  assign n4652 = n4650 | n4651 ;
  buffer buf_n4641( .i (n4640), .o (n4641) );
  buffer buf_n4642( .i (n4641), .o (n4642) );
  buffer buf_n4643( .i (n4642), .o (n4643) );
  buffer buf_n4644( .i (n4643), .o (n4644) );
  assign n4653 = n4644 & ~n4650 ;
  buffer buf_n4654( .i (n4653), .o (n4654) );
  buffer buf_n4617( .i (n4616), .o (n4617) );
  buffer buf_n4618( .i (n4617), .o (n4618) );
  buffer buf_n4619( .i (n4618), .o (n4619) );
  buffer buf_n4620( .i (n4619), .o (n4620) );
  buffer buf_n4621( .i (n4620), .o (n4621) );
  buffer buf_n4622( .i (n4621), .o (n4622) );
  buffer buf_n4623( .i (n4622), .o (n4623) );
  buffer buf_n4624( .i (n4623), .o (n4624) );
  buffer buf_n4631( .i (n4630), .o (n4631) );
  buffer buf_n4632( .i (n4631), .o (n4632) );
  buffer buf_n4633( .i (n4632), .o (n4633) );
  buffer buf_n4634( .i (n4633), .o (n4634) );
  assign n4656 = n4624 & ~n4634 ;
  buffer buf_n4657( .i (n4656), .o (n4657) );
  assign n4659 = N120 & N528 ;
  buffer buf_n4660( .i (n4659), .o (n4660) );
  buffer buf_n4593( .i (n4592), .o (n4593) );
  buffer buf_n4594( .i (n4593), .o (n4594) );
  buffer buf_n4595( .i (n4594), .o (n4595) );
  buffer buf_n4596( .i (n4595), .o (n4596) );
  buffer buf_n4597( .i (n4596), .o (n4597) );
  buffer buf_n4598( .i (n4597), .o (n4598) );
  buffer buf_n4599( .i (n4598), .o (n4599) );
  buffer buf_n4600( .i (n4599), .o (n4600) );
  buffer buf_n4607( .i (n4606), .o (n4607) );
  buffer buf_n4608( .i (n4607), .o (n4608) );
  buffer buf_n4609( .i (n4608), .o (n4609) );
  buffer buf_n4610( .i (n4609), .o (n4610) );
  assign n4662 = n4600 & ~n4610 ;
  buffer buf_n4663( .i (n4662), .o (n4663) );
  assign n4665 = N137 & N511 ;
  buffer buf_n4666( .i (n4665), .o (n4666) );
  buffer buf_n4569( .i (n4568), .o (n4569) );
  buffer buf_n4570( .i (n4569), .o (n4570) );
  buffer buf_n4571( .i (n4570), .o (n4571) );
  buffer buf_n4572( .i (n4571), .o (n4572) );
  buffer buf_n4573( .i (n4572), .o (n4573) );
  buffer buf_n4574( .i (n4573), .o (n4574) );
  buffer buf_n4575( .i (n4574), .o (n4575) );
  buffer buf_n4576( .i (n4575), .o (n4576) );
  buffer buf_n4583( .i (n4582), .o (n4583) );
  buffer buf_n4584( .i (n4583), .o (n4584) );
  buffer buf_n4585( .i (n4584), .o (n4585) );
  buffer buf_n4586( .i (n4585), .o (n4586) );
  assign n4668 = n4576 & ~n4586 ;
  buffer buf_n4669( .i (n4668), .o (n4669) );
  assign n4671 = N154 & N494 ;
  buffer buf_n4672( .i (n4671), .o (n4672) );
  buffer buf_n4545( .i (n4544), .o (n4545) );
  buffer buf_n4546( .i (n4545), .o (n4546) );
  buffer buf_n4547( .i (n4546), .o (n4547) );
  buffer buf_n4548( .i (n4547), .o (n4548) );
  buffer buf_n4549( .i (n4548), .o (n4549) );
  buffer buf_n4550( .i (n4549), .o (n4550) );
  buffer buf_n4551( .i (n4550), .o (n4551) );
  buffer buf_n4552( .i (n4551), .o (n4552) );
  buffer buf_n4559( .i (n4558), .o (n4559) );
  buffer buf_n4560( .i (n4559), .o (n4560) );
  buffer buf_n4561( .i (n4560), .o (n4561) );
  buffer buf_n4562( .i (n4561), .o (n4562) );
  assign n4674 = n4552 & ~n4562 ;
  buffer buf_n4675( .i (n4674), .o (n4675) );
  assign n4677 = N171 & N477 ;
  buffer buf_n4678( .i (n4677), .o (n4678) );
  buffer buf_n4521( .i (n4520), .o (n4521) );
  buffer buf_n4522( .i (n4521), .o (n4522) );
  buffer buf_n4523( .i (n4522), .o (n4523) );
  buffer buf_n4524( .i (n4523), .o (n4524) );
  buffer buf_n4525( .i (n4524), .o (n4525) );
  buffer buf_n4526( .i (n4525), .o (n4526) );
  buffer buf_n4527( .i (n4526), .o (n4527) );
  buffer buf_n4528( .i (n4527), .o (n4528) );
  buffer buf_n4535( .i (n4534), .o (n4535) );
  buffer buf_n4536( .i (n4535), .o (n4536) );
  buffer buf_n4537( .i (n4536), .o (n4537) );
  buffer buf_n4538( .i (n4537), .o (n4538) );
  assign n4680 = n4528 & ~n4538 ;
  buffer buf_n4681( .i (n4680), .o (n4681) );
  assign n4683 = N188 & N460 ;
  buffer buf_n4684( .i (n4683), .o (n4684) );
  buffer buf_n4497( .i (n4496), .o (n4497) );
  buffer buf_n4498( .i (n4497), .o (n4498) );
  buffer buf_n4499( .i (n4498), .o (n4499) );
  buffer buf_n4500( .i (n4499), .o (n4500) );
  buffer buf_n4501( .i (n4500), .o (n4501) );
  buffer buf_n4502( .i (n4501), .o (n4502) );
  buffer buf_n4503( .i (n4502), .o (n4503) );
  buffer buf_n4504( .i (n4503), .o (n4504) );
  buffer buf_n4511( .i (n4510), .o (n4511) );
  buffer buf_n4512( .i (n4511), .o (n4512) );
  buffer buf_n4513( .i (n4512), .o (n4513) );
  buffer buf_n4514( .i (n4513), .o (n4514) );
  assign n4686 = n4504 & ~n4514 ;
  buffer buf_n4687( .i (n4686), .o (n4687) );
  assign n4689 = N205 & N443 ;
  buffer buf_n4690( .i (n4689), .o (n4690) );
  buffer buf_n4473( .i (n4472), .o (n4473) );
  buffer buf_n4474( .i (n4473), .o (n4474) );
  buffer buf_n4475( .i (n4474), .o (n4475) );
  buffer buf_n4476( .i (n4475), .o (n4476) );
  buffer buf_n4477( .i (n4476), .o (n4477) );
  buffer buf_n4478( .i (n4477), .o (n4478) );
  buffer buf_n4479( .i (n4478), .o (n4479) );
  buffer buf_n4480( .i (n4479), .o (n4480) );
  buffer buf_n4487( .i (n4486), .o (n4487) );
  buffer buf_n4488( .i (n4487), .o (n4488) );
  buffer buf_n4489( .i (n4488), .o (n4489) );
  buffer buf_n4490( .i (n4489), .o (n4490) );
  assign n4692 = n4480 & ~n4490 ;
  buffer buf_n4693( .i (n4692), .o (n4693) );
  assign n4695 = N222 & N426 ;
  buffer buf_n4696( .i (n4695), .o (n4696) );
  buffer buf_n4449( .i (n4448), .o (n4449) );
  buffer buf_n4450( .i (n4449), .o (n4450) );
  buffer buf_n4451( .i (n4450), .o (n4451) );
  buffer buf_n4452( .i (n4451), .o (n4452) );
  buffer buf_n4453( .i (n4452), .o (n4453) );
  buffer buf_n4454( .i (n4453), .o (n4454) );
  buffer buf_n4455( .i (n4454), .o (n4455) );
  buffer buf_n4456( .i (n4455), .o (n4456) );
  buffer buf_n4463( .i (n4462), .o (n4463) );
  buffer buf_n4464( .i (n4463), .o (n4464) );
  buffer buf_n4465( .i (n4464), .o (n4465) );
  buffer buf_n4466( .i (n4465), .o (n4466) );
  assign n4698 = n4456 & ~n4466 ;
  buffer buf_n4699( .i (n4698), .o (n4699) );
  assign n4701 = N239 & N409 ;
  buffer buf_n4702( .i (n4701), .o (n4702) );
  assign n4704 = N256 & N392 ;
  buffer buf_n4705( .i (n4704), .o (n4705) );
  buffer buf_n4425( .i (n4424), .o (n4425) );
  buffer buf_n4426( .i (n4425), .o (n4426) );
  buffer buf_n4427( .i (n4426), .o (n4427) );
  buffer buf_n4428( .i (n4427), .o (n4428) );
  buffer buf_n4429( .i (n4428), .o (n4429) );
  buffer buf_n4430( .i (n4429), .o (n4430) );
  buffer buf_n4431( .i (n4430), .o (n4431) );
  buffer buf_n4432( .i (n4431), .o (n4432) );
  buffer buf_n4439( .i (n4438), .o (n4439) );
  buffer buf_n4440( .i (n4439), .o (n4440) );
  buffer buf_n4441( .i (n4440), .o (n4441) );
  buffer buf_n4442( .i (n4441), .o (n4442) );
  assign n4707 = n4432 & ~n4442 ;
  buffer buf_n4708( .i (n4707), .o (n4708) );
  assign n4710 = n4705 | n4708 ;
  buffer buf_n4711( .i (n4710), .o (n4711) );
  buffer buf_n4706( .i (n4705), .o (n4706) );
  buffer buf_n4709( .i (n4708), .o (n4709) );
  assign n4720 = n4706 & n4709 ;
  assign n4721 = n4711 & ~n4720 ;
  buffer buf_n4722( .i (n4721), .o (n4722) );
  assign n4724 = ~n4702 & n4722 ;
  buffer buf_n4725( .i (n4724), .o (n4725) );
  buffer buf_n4703( .i (n4702), .o (n4703) );
  buffer buf_n4723( .i (n4722), .o (n4723) );
  assign n4730 = n4703 & ~n4723 ;
  assign n4731 = n4725 | n4730 ;
  buffer buf_n4732( .i (n4731), .o (n4732) );
  assign n4734 = n4699 | n4732 ;
  buffer buf_n4735( .i (n4734), .o (n4735) );
  buffer buf_n4700( .i (n4699), .o (n4700) );
  buffer buf_n4733( .i (n4732), .o (n4733) );
  assign n4744 = n4700 & n4733 ;
  assign n4745 = n4735 & ~n4744 ;
  buffer buf_n4746( .i (n4745), .o (n4746) );
  assign n4748 = ~n4696 & n4746 ;
  buffer buf_n4749( .i (n4748), .o (n4749) );
  buffer buf_n4697( .i (n4696), .o (n4697) );
  buffer buf_n4747( .i (n4746), .o (n4747) );
  assign n4754 = n4697 & ~n4747 ;
  assign n4755 = n4749 | n4754 ;
  buffer buf_n4756( .i (n4755), .o (n4756) );
  assign n4758 = n4693 | n4756 ;
  buffer buf_n4759( .i (n4758), .o (n4759) );
  buffer buf_n4694( .i (n4693), .o (n4694) );
  buffer buf_n4757( .i (n4756), .o (n4757) );
  assign n4768 = n4694 & n4757 ;
  assign n4769 = n4759 & ~n4768 ;
  buffer buf_n4770( .i (n4769), .o (n4770) );
  assign n4772 = ~n4690 & n4770 ;
  buffer buf_n4773( .i (n4772), .o (n4773) );
  buffer buf_n4691( .i (n4690), .o (n4691) );
  buffer buf_n4771( .i (n4770), .o (n4771) );
  assign n4778 = n4691 & ~n4771 ;
  assign n4779 = n4773 | n4778 ;
  buffer buf_n4780( .i (n4779), .o (n4780) );
  assign n4782 = n4687 | n4780 ;
  buffer buf_n4783( .i (n4782), .o (n4783) );
  buffer buf_n4688( .i (n4687), .o (n4688) );
  buffer buf_n4781( .i (n4780), .o (n4781) );
  assign n4792 = n4688 & n4781 ;
  assign n4793 = n4783 & ~n4792 ;
  buffer buf_n4794( .i (n4793), .o (n4794) );
  assign n4796 = ~n4684 & n4794 ;
  buffer buf_n4797( .i (n4796), .o (n4797) );
  buffer buf_n4685( .i (n4684), .o (n4685) );
  buffer buf_n4795( .i (n4794), .o (n4795) );
  assign n4802 = n4685 & ~n4795 ;
  assign n4803 = n4797 | n4802 ;
  buffer buf_n4804( .i (n4803), .o (n4804) );
  assign n4806 = n4681 | n4804 ;
  buffer buf_n4807( .i (n4806), .o (n4807) );
  buffer buf_n4682( .i (n4681), .o (n4682) );
  buffer buf_n4805( .i (n4804), .o (n4805) );
  assign n4816 = n4682 & n4805 ;
  assign n4817 = n4807 & ~n4816 ;
  buffer buf_n4818( .i (n4817), .o (n4818) );
  assign n4820 = ~n4678 & n4818 ;
  buffer buf_n4821( .i (n4820), .o (n4821) );
  buffer buf_n4679( .i (n4678), .o (n4679) );
  buffer buf_n4819( .i (n4818), .o (n4819) );
  assign n4826 = n4679 & ~n4819 ;
  assign n4827 = n4821 | n4826 ;
  buffer buf_n4828( .i (n4827), .o (n4828) );
  assign n4830 = n4675 | n4828 ;
  buffer buf_n4831( .i (n4830), .o (n4831) );
  buffer buf_n4676( .i (n4675), .o (n4676) );
  buffer buf_n4829( .i (n4828), .o (n4829) );
  assign n4840 = n4676 & n4829 ;
  assign n4841 = n4831 & ~n4840 ;
  buffer buf_n4842( .i (n4841), .o (n4842) );
  assign n4844 = ~n4672 & n4842 ;
  buffer buf_n4845( .i (n4844), .o (n4845) );
  buffer buf_n4673( .i (n4672), .o (n4673) );
  buffer buf_n4843( .i (n4842), .o (n4843) );
  assign n4850 = n4673 & ~n4843 ;
  assign n4851 = n4845 | n4850 ;
  buffer buf_n4852( .i (n4851), .o (n4852) );
  assign n4854 = n4669 | n4852 ;
  buffer buf_n4855( .i (n4854), .o (n4855) );
  buffer buf_n4670( .i (n4669), .o (n4670) );
  buffer buf_n4853( .i (n4852), .o (n4853) );
  assign n4864 = n4670 & n4853 ;
  assign n4865 = n4855 & ~n4864 ;
  buffer buf_n4866( .i (n4865), .o (n4866) );
  assign n4868 = ~n4666 & n4866 ;
  buffer buf_n4869( .i (n4868), .o (n4869) );
  buffer buf_n4667( .i (n4666), .o (n4667) );
  buffer buf_n4867( .i (n4866), .o (n4867) );
  assign n4874 = n4667 & ~n4867 ;
  assign n4875 = n4869 | n4874 ;
  buffer buf_n4876( .i (n4875), .o (n4876) );
  assign n4878 = n4663 | n4876 ;
  buffer buf_n4879( .i (n4878), .o (n4879) );
  buffer buf_n4664( .i (n4663), .o (n4664) );
  buffer buf_n4877( .i (n4876), .o (n4877) );
  assign n4888 = n4664 & n4877 ;
  assign n4889 = n4879 & ~n4888 ;
  buffer buf_n4890( .i (n4889), .o (n4890) );
  assign n4892 = ~n4660 & n4890 ;
  buffer buf_n4893( .i (n4892), .o (n4893) );
  buffer buf_n4661( .i (n4660), .o (n4661) );
  buffer buf_n4891( .i (n4890), .o (n4891) );
  assign n4898 = n4661 & ~n4891 ;
  assign n4899 = n4893 | n4898 ;
  buffer buf_n4900( .i (n4899), .o (n4900) );
  assign n4902 = n4657 | n4900 ;
  buffer buf_n4903( .i (n4902), .o (n4903) );
  buffer buf_n4658( .i (n4657), .o (n4658) );
  buffer buf_n4901( .i (n4900), .o (n4901) );
  assign n4908 = n4658 & n4901 ;
  assign n4909 = n4903 & ~n4908 ;
  buffer buf_n4910( .i (n4909), .o (n4910) );
  assign n4912 = ~n4654 & n4910 ;
  buffer buf_n4913( .i (n4912), .o (n4913) );
  buffer buf_n4655( .i (n4654), .o (n4655) );
  buffer buf_n4911( .i (n4910), .o (n4911) );
  assign n4914 = n4655 & ~n4911 ;
  assign n4915 = n4913 | n4914 ;
  buffer buf_n4904( .i (n4903), .o (n4904) );
  buffer buf_n4905( .i (n4904), .o (n4905) );
  buffer buf_n4906( .i (n4905), .o (n4906) );
  buffer buf_n4907( .i (n4906), .o (n4907) );
  assign n4916 = n4907 & ~n4913 ;
  buffer buf_n4917( .i (n4916), .o (n4917) );
  buffer buf_n4880( .i (n4879), .o (n4880) );
  buffer buf_n4881( .i (n4880), .o (n4881) );
  buffer buf_n4882( .i (n4881), .o (n4882) );
  buffer buf_n4883( .i (n4882), .o (n4883) );
  buffer buf_n4884( .i (n4883), .o (n4884) );
  buffer buf_n4885( .i (n4884), .o (n4885) );
  buffer buf_n4886( .i (n4885), .o (n4886) );
  buffer buf_n4887( .i (n4886), .o (n4887) );
  buffer buf_n4894( .i (n4893), .o (n4894) );
  buffer buf_n4895( .i (n4894), .o (n4895) );
  buffer buf_n4896( .i (n4895), .o (n4896) );
  buffer buf_n4897( .i (n4896), .o (n4897) );
  assign n4919 = n4887 & ~n4897 ;
  buffer buf_n4920( .i (n4919), .o (n4920) );
  assign n4922 = N137 & N528 ;
  buffer buf_n4923( .i (n4922), .o (n4923) );
  buffer buf_n4856( .i (n4855), .o (n4856) );
  buffer buf_n4857( .i (n4856), .o (n4857) );
  buffer buf_n4858( .i (n4857), .o (n4858) );
  buffer buf_n4859( .i (n4858), .o (n4859) );
  buffer buf_n4860( .i (n4859), .o (n4860) );
  buffer buf_n4861( .i (n4860), .o (n4861) );
  buffer buf_n4862( .i (n4861), .o (n4862) );
  buffer buf_n4863( .i (n4862), .o (n4863) );
  buffer buf_n4870( .i (n4869), .o (n4870) );
  buffer buf_n4871( .i (n4870), .o (n4871) );
  buffer buf_n4872( .i (n4871), .o (n4872) );
  buffer buf_n4873( .i (n4872), .o (n4873) );
  assign n4925 = n4863 & ~n4873 ;
  buffer buf_n4926( .i (n4925), .o (n4926) );
  assign n4928 = N154 & N511 ;
  buffer buf_n4929( .i (n4928), .o (n4929) );
  buffer buf_n4832( .i (n4831), .o (n4832) );
  buffer buf_n4833( .i (n4832), .o (n4833) );
  buffer buf_n4834( .i (n4833), .o (n4834) );
  buffer buf_n4835( .i (n4834), .o (n4835) );
  buffer buf_n4836( .i (n4835), .o (n4836) );
  buffer buf_n4837( .i (n4836), .o (n4837) );
  buffer buf_n4838( .i (n4837), .o (n4838) );
  buffer buf_n4839( .i (n4838), .o (n4839) );
  buffer buf_n4846( .i (n4845), .o (n4846) );
  buffer buf_n4847( .i (n4846), .o (n4847) );
  buffer buf_n4848( .i (n4847), .o (n4848) );
  buffer buf_n4849( .i (n4848), .o (n4849) );
  assign n4931 = n4839 & ~n4849 ;
  buffer buf_n4932( .i (n4931), .o (n4932) );
  assign n4934 = N171 & N494 ;
  buffer buf_n4935( .i (n4934), .o (n4935) );
  buffer buf_n4808( .i (n4807), .o (n4808) );
  buffer buf_n4809( .i (n4808), .o (n4809) );
  buffer buf_n4810( .i (n4809), .o (n4810) );
  buffer buf_n4811( .i (n4810), .o (n4811) );
  buffer buf_n4812( .i (n4811), .o (n4812) );
  buffer buf_n4813( .i (n4812), .o (n4813) );
  buffer buf_n4814( .i (n4813), .o (n4814) );
  buffer buf_n4815( .i (n4814), .o (n4815) );
  buffer buf_n4822( .i (n4821), .o (n4822) );
  buffer buf_n4823( .i (n4822), .o (n4823) );
  buffer buf_n4824( .i (n4823), .o (n4824) );
  buffer buf_n4825( .i (n4824), .o (n4825) );
  assign n4937 = n4815 & ~n4825 ;
  buffer buf_n4938( .i (n4937), .o (n4938) );
  assign n4940 = N188 & N477 ;
  buffer buf_n4941( .i (n4940), .o (n4941) );
  buffer buf_n4784( .i (n4783), .o (n4784) );
  buffer buf_n4785( .i (n4784), .o (n4785) );
  buffer buf_n4786( .i (n4785), .o (n4786) );
  buffer buf_n4787( .i (n4786), .o (n4787) );
  buffer buf_n4788( .i (n4787), .o (n4788) );
  buffer buf_n4789( .i (n4788), .o (n4789) );
  buffer buf_n4790( .i (n4789), .o (n4790) );
  buffer buf_n4791( .i (n4790), .o (n4791) );
  buffer buf_n4798( .i (n4797), .o (n4798) );
  buffer buf_n4799( .i (n4798), .o (n4799) );
  buffer buf_n4800( .i (n4799), .o (n4800) );
  buffer buf_n4801( .i (n4800), .o (n4801) );
  assign n4943 = n4791 & ~n4801 ;
  buffer buf_n4944( .i (n4943), .o (n4944) );
  assign n4946 = N205 & N460 ;
  buffer buf_n4947( .i (n4946), .o (n4947) );
  buffer buf_n4760( .i (n4759), .o (n4760) );
  buffer buf_n4761( .i (n4760), .o (n4761) );
  buffer buf_n4762( .i (n4761), .o (n4762) );
  buffer buf_n4763( .i (n4762), .o (n4763) );
  buffer buf_n4764( .i (n4763), .o (n4764) );
  buffer buf_n4765( .i (n4764), .o (n4765) );
  buffer buf_n4766( .i (n4765), .o (n4766) );
  buffer buf_n4767( .i (n4766), .o (n4767) );
  buffer buf_n4774( .i (n4773), .o (n4774) );
  buffer buf_n4775( .i (n4774), .o (n4775) );
  buffer buf_n4776( .i (n4775), .o (n4776) );
  buffer buf_n4777( .i (n4776), .o (n4777) );
  assign n4949 = n4767 & ~n4777 ;
  buffer buf_n4950( .i (n4949), .o (n4950) );
  assign n4952 = N222 & N443 ;
  buffer buf_n4953( .i (n4952), .o (n4953) );
  buffer buf_n4736( .i (n4735), .o (n4736) );
  buffer buf_n4737( .i (n4736), .o (n4737) );
  buffer buf_n4738( .i (n4737), .o (n4738) );
  buffer buf_n4739( .i (n4738), .o (n4739) );
  buffer buf_n4740( .i (n4739), .o (n4740) );
  buffer buf_n4741( .i (n4740), .o (n4741) );
  buffer buf_n4742( .i (n4741), .o (n4742) );
  buffer buf_n4743( .i (n4742), .o (n4743) );
  buffer buf_n4750( .i (n4749), .o (n4750) );
  buffer buf_n4751( .i (n4750), .o (n4751) );
  buffer buf_n4752( .i (n4751), .o (n4752) );
  buffer buf_n4753( .i (n4752), .o (n4753) );
  assign n4955 = n4743 & ~n4753 ;
  buffer buf_n4956( .i (n4955), .o (n4956) );
  assign n4958 = N239 & N426 ;
  buffer buf_n4959( .i (n4958), .o (n4959) );
  assign n4961 = N256 & N409 ;
  buffer buf_n4962( .i (n4961), .o (n4962) );
  buffer buf_n4712( .i (n4711), .o (n4712) );
  buffer buf_n4713( .i (n4712), .o (n4713) );
  buffer buf_n4714( .i (n4713), .o (n4714) );
  buffer buf_n4715( .i (n4714), .o (n4715) );
  buffer buf_n4716( .i (n4715), .o (n4716) );
  buffer buf_n4717( .i (n4716), .o (n4717) );
  buffer buf_n4718( .i (n4717), .o (n4718) );
  buffer buf_n4719( .i (n4718), .o (n4719) );
  buffer buf_n4726( .i (n4725), .o (n4726) );
  buffer buf_n4727( .i (n4726), .o (n4727) );
  buffer buf_n4728( .i (n4727), .o (n4728) );
  buffer buf_n4729( .i (n4728), .o (n4729) );
  assign n4964 = n4719 & ~n4729 ;
  buffer buf_n4965( .i (n4964), .o (n4965) );
  assign n4967 = n4962 | n4965 ;
  buffer buf_n4968( .i (n4967), .o (n4968) );
  buffer buf_n4963( .i (n4962), .o (n4963) );
  buffer buf_n4966( .i (n4965), .o (n4966) );
  assign n4977 = n4963 & n4966 ;
  assign n4978 = n4968 & ~n4977 ;
  buffer buf_n4979( .i (n4978), .o (n4979) );
  assign n4981 = ~n4959 & n4979 ;
  buffer buf_n4982( .i (n4981), .o (n4982) );
  buffer buf_n4960( .i (n4959), .o (n4960) );
  buffer buf_n4980( .i (n4979), .o (n4980) );
  assign n4987 = n4960 & ~n4980 ;
  assign n4988 = n4982 | n4987 ;
  buffer buf_n4989( .i (n4988), .o (n4989) );
  assign n4991 = n4956 | n4989 ;
  buffer buf_n4992( .i (n4991), .o (n4992) );
  buffer buf_n4957( .i (n4956), .o (n4957) );
  buffer buf_n4990( .i (n4989), .o (n4990) );
  assign n5001 = n4957 & n4990 ;
  assign n5002 = n4992 & ~n5001 ;
  buffer buf_n5003( .i (n5002), .o (n5003) );
  assign n5005 = ~n4953 & n5003 ;
  buffer buf_n5006( .i (n5005), .o (n5006) );
  buffer buf_n4954( .i (n4953), .o (n4954) );
  buffer buf_n5004( .i (n5003), .o (n5004) );
  assign n5011 = n4954 & ~n5004 ;
  assign n5012 = n5006 | n5011 ;
  buffer buf_n5013( .i (n5012), .o (n5013) );
  assign n5015 = n4950 | n5013 ;
  buffer buf_n5016( .i (n5015), .o (n5016) );
  buffer buf_n4951( .i (n4950), .o (n4951) );
  buffer buf_n5014( .i (n5013), .o (n5014) );
  assign n5025 = n4951 & n5014 ;
  assign n5026 = n5016 & ~n5025 ;
  buffer buf_n5027( .i (n5026), .o (n5027) );
  assign n5029 = ~n4947 & n5027 ;
  buffer buf_n5030( .i (n5029), .o (n5030) );
  buffer buf_n4948( .i (n4947), .o (n4948) );
  buffer buf_n5028( .i (n5027), .o (n5028) );
  assign n5035 = n4948 & ~n5028 ;
  assign n5036 = n5030 | n5035 ;
  buffer buf_n5037( .i (n5036), .o (n5037) );
  assign n5039 = n4944 | n5037 ;
  buffer buf_n5040( .i (n5039), .o (n5040) );
  buffer buf_n4945( .i (n4944), .o (n4945) );
  buffer buf_n5038( .i (n5037), .o (n5038) );
  assign n5049 = n4945 & n5038 ;
  assign n5050 = n5040 & ~n5049 ;
  buffer buf_n5051( .i (n5050), .o (n5051) );
  assign n5053 = ~n4941 & n5051 ;
  buffer buf_n5054( .i (n5053), .o (n5054) );
  buffer buf_n4942( .i (n4941), .o (n4942) );
  buffer buf_n5052( .i (n5051), .o (n5052) );
  assign n5059 = n4942 & ~n5052 ;
  assign n5060 = n5054 | n5059 ;
  buffer buf_n5061( .i (n5060), .o (n5061) );
  assign n5063 = n4938 | n5061 ;
  buffer buf_n5064( .i (n5063), .o (n5064) );
  buffer buf_n4939( .i (n4938), .o (n4939) );
  buffer buf_n5062( .i (n5061), .o (n5062) );
  assign n5073 = n4939 & n5062 ;
  assign n5074 = n5064 & ~n5073 ;
  buffer buf_n5075( .i (n5074), .o (n5075) );
  assign n5077 = ~n4935 & n5075 ;
  buffer buf_n5078( .i (n5077), .o (n5078) );
  buffer buf_n4936( .i (n4935), .o (n4936) );
  buffer buf_n5076( .i (n5075), .o (n5076) );
  assign n5083 = n4936 & ~n5076 ;
  assign n5084 = n5078 | n5083 ;
  buffer buf_n5085( .i (n5084), .o (n5085) );
  assign n5087 = n4932 | n5085 ;
  buffer buf_n5088( .i (n5087), .o (n5088) );
  buffer buf_n4933( .i (n4932), .o (n4933) );
  buffer buf_n5086( .i (n5085), .o (n5086) );
  assign n5097 = n4933 & n5086 ;
  assign n5098 = n5088 & ~n5097 ;
  buffer buf_n5099( .i (n5098), .o (n5099) );
  assign n5101 = ~n4929 & n5099 ;
  buffer buf_n5102( .i (n5101), .o (n5102) );
  buffer buf_n4930( .i (n4929), .o (n4930) );
  buffer buf_n5100( .i (n5099), .o (n5100) );
  assign n5107 = n4930 & ~n5100 ;
  assign n5108 = n5102 | n5107 ;
  buffer buf_n5109( .i (n5108), .o (n5109) );
  assign n5111 = n4926 | n5109 ;
  buffer buf_n5112( .i (n5111), .o (n5112) );
  buffer buf_n4927( .i (n4926), .o (n4927) );
  buffer buf_n5110( .i (n5109), .o (n5110) );
  assign n5121 = n4927 & n5110 ;
  assign n5122 = n5112 & ~n5121 ;
  buffer buf_n5123( .i (n5122), .o (n5123) );
  assign n5125 = ~n4923 & n5123 ;
  buffer buf_n5126( .i (n5125), .o (n5126) );
  buffer buf_n4924( .i (n4923), .o (n4924) );
  buffer buf_n5124( .i (n5123), .o (n5124) );
  assign n5131 = n4924 & ~n5124 ;
  assign n5132 = n5126 | n5131 ;
  buffer buf_n5133( .i (n5132), .o (n5133) );
  assign n5135 = n4920 | n5133 ;
  buffer buf_n5136( .i (n5135), .o (n5136) );
  buffer buf_n4921( .i (n4920), .o (n4921) );
  buffer buf_n5134( .i (n5133), .o (n5134) );
  assign n5141 = n4921 & n5134 ;
  assign n5142 = n5136 & ~n5141 ;
  buffer buf_n5143( .i (n5142), .o (n5143) );
  assign n5145 = ~n4917 & n5143 ;
  buffer buf_n5146( .i (n5145), .o (n5146) );
  buffer buf_n4918( .i (n4917), .o (n4918) );
  buffer buf_n5144( .i (n5143), .o (n5144) );
  assign n5147 = n4918 & ~n5144 ;
  assign n5148 = n5146 | n5147 ;
  buffer buf_n5137( .i (n5136), .o (n5137) );
  buffer buf_n5138( .i (n5137), .o (n5138) );
  buffer buf_n5139( .i (n5138), .o (n5139) );
  buffer buf_n5140( .i (n5139), .o (n5140) );
  assign n5149 = n5140 & ~n5146 ;
  buffer buf_n5150( .i (n5149), .o (n5150) );
  buffer buf_n5113( .i (n5112), .o (n5113) );
  buffer buf_n5114( .i (n5113), .o (n5114) );
  buffer buf_n5115( .i (n5114), .o (n5115) );
  buffer buf_n5116( .i (n5115), .o (n5116) );
  buffer buf_n5117( .i (n5116), .o (n5117) );
  buffer buf_n5118( .i (n5117), .o (n5118) );
  buffer buf_n5119( .i (n5118), .o (n5119) );
  buffer buf_n5120( .i (n5119), .o (n5120) );
  buffer buf_n5127( .i (n5126), .o (n5127) );
  buffer buf_n5128( .i (n5127), .o (n5128) );
  buffer buf_n5129( .i (n5128), .o (n5129) );
  buffer buf_n5130( .i (n5129), .o (n5130) );
  assign n5152 = n5120 & ~n5130 ;
  buffer buf_n5153( .i (n5152), .o (n5153) );
  assign n5155 = N154 & N528 ;
  buffer buf_n5156( .i (n5155), .o (n5156) );
  buffer buf_n5089( .i (n5088), .o (n5089) );
  buffer buf_n5090( .i (n5089), .o (n5090) );
  buffer buf_n5091( .i (n5090), .o (n5091) );
  buffer buf_n5092( .i (n5091), .o (n5092) );
  buffer buf_n5093( .i (n5092), .o (n5093) );
  buffer buf_n5094( .i (n5093), .o (n5094) );
  buffer buf_n5095( .i (n5094), .o (n5095) );
  buffer buf_n5096( .i (n5095), .o (n5096) );
  buffer buf_n5103( .i (n5102), .o (n5103) );
  buffer buf_n5104( .i (n5103), .o (n5104) );
  buffer buf_n5105( .i (n5104), .o (n5105) );
  buffer buf_n5106( .i (n5105), .o (n5106) );
  assign n5158 = n5096 & ~n5106 ;
  buffer buf_n5159( .i (n5158), .o (n5159) );
  assign n5161 = N171 & N511 ;
  buffer buf_n5162( .i (n5161), .o (n5162) );
  buffer buf_n5065( .i (n5064), .o (n5065) );
  buffer buf_n5066( .i (n5065), .o (n5066) );
  buffer buf_n5067( .i (n5066), .o (n5067) );
  buffer buf_n5068( .i (n5067), .o (n5068) );
  buffer buf_n5069( .i (n5068), .o (n5069) );
  buffer buf_n5070( .i (n5069), .o (n5070) );
  buffer buf_n5071( .i (n5070), .o (n5071) );
  buffer buf_n5072( .i (n5071), .o (n5072) );
  buffer buf_n5079( .i (n5078), .o (n5079) );
  buffer buf_n5080( .i (n5079), .o (n5080) );
  buffer buf_n5081( .i (n5080), .o (n5081) );
  buffer buf_n5082( .i (n5081), .o (n5082) );
  assign n5164 = n5072 & ~n5082 ;
  buffer buf_n5165( .i (n5164), .o (n5165) );
  assign n5167 = N188 & N494 ;
  buffer buf_n5168( .i (n5167), .o (n5168) );
  buffer buf_n5041( .i (n5040), .o (n5041) );
  buffer buf_n5042( .i (n5041), .o (n5042) );
  buffer buf_n5043( .i (n5042), .o (n5043) );
  buffer buf_n5044( .i (n5043), .o (n5044) );
  buffer buf_n5045( .i (n5044), .o (n5045) );
  buffer buf_n5046( .i (n5045), .o (n5046) );
  buffer buf_n5047( .i (n5046), .o (n5047) );
  buffer buf_n5048( .i (n5047), .o (n5048) );
  buffer buf_n5055( .i (n5054), .o (n5055) );
  buffer buf_n5056( .i (n5055), .o (n5056) );
  buffer buf_n5057( .i (n5056), .o (n5057) );
  buffer buf_n5058( .i (n5057), .o (n5058) );
  assign n5170 = n5048 & ~n5058 ;
  buffer buf_n5171( .i (n5170), .o (n5171) );
  assign n5173 = N205 & N477 ;
  buffer buf_n5174( .i (n5173), .o (n5174) );
  buffer buf_n5017( .i (n5016), .o (n5017) );
  buffer buf_n5018( .i (n5017), .o (n5018) );
  buffer buf_n5019( .i (n5018), .o (n5019) );
  buffer buf_n5020( .i (n5019), .o (n5020) );
  buffer buf_n5021( .i (n5020), .o (n5021) );
  buffer buf_n5022( .i (n5021), .o (n5022) );
  buffer buf_n5023( .i (n5022), .o (n5023) );
  buffer buf_n5024( .i (n5023), .o (n5024) );
  buffer buf_n5031( .i (n5030), .o (n5031) );
  buffer buf_n5032( .i (n5031), .o (n5032) );
  buffer buf_n5033( .i (n5032), .o (n5033) );
  buffer buf_n5034( .i (n5033), .o (n5034) );
  assign n5176 = n5024 & ~n5034 ;
  buffer buf_n5177( .i (n5176), .o (n5177) );
  assign n5179 = N222 & N460 ;
  buffer buf_n5180( .i (n5179), .o (n5180) );
  buffer buf_n4993( .i (n4992), .o (n4993) );
  buffer buf_n4994( .i (n4993), .o (n4994) );
  buffer buf_n4995( .i (n4994), .o (n4995) );
  buffer buf_n4996( .i (n4995), .o (n4996) );
  buffer buf_n4997( .i (n4996), .o (n4997) );
  buffer buf_n4998( .i (n4997), .o (n4998) );
  buffer buf_n4999( .i (n4998), .o (n4999) );
  buffer buf_n5000( .i (n4999), .o (n5000) );
  buffer buf_n5007( .i (n5006), .o (n5007) );
  buffer buf_n5008( .i (n5007), .o (n5008) );
  buffer buf_n5009( .i (n5008), .o (n5009) );
  buffer buf_n5010( .i (n5009), .o (n5010) );
  assign n5182 = n5000 & ~n5010 ;
  buffer buf_n5183( .i (n5182), .o (n5183) );
  assign n5185 = N239 & N443 ;
  buffer buf_n5186( .i (n5185), .o (n5186) );
  assign n5188 = N256 & N426 ;
  buffer buf_n5189( .i (n5188), .o (n5189) );
  buffer buf_n4969( .i (n4968), .o (n4969) );
  buffer buf_n4970( .i (n4969), .o (n4970) );
  buffer buf_n4971( .i (n4970), .o (n4971) );
  buffer buf_n4972( .i (n4971), .o (n4972) );
  buffer buf_n4973( .i (n4972), .o (n4973) );
  buffer buf_n4974( .i (n4973), .o (n4974) );
  buffer buf_n4975( .i (n4974), .o (n4975) );
  buffer buf_n4976( .i (n4975), .o (n4976) );
  buffer buf_n4983( .i (n4982), .o (n4983) );
  buffer buf_n4984( .i (n4983), .o (n4984) );
  buffer buf_n4985( .i (n4984), .o (n4985) );
  buffer buf_n4986( .i (n4985), .o (n4986) );
  assign n5191 = n4976 & ~n4986 ;
  buffer buf_n5192( .i (n5191), .o (n5192) );
  assign n5194 = n5189 | n5192 ;
  buffer buf_n5195( .i (n5194), .o (n5195) );
  buffer buf_n5190( .i (n5189), .o (n5190) );
  buffer buf_n5193( .i (n5192), .o (n5193) );
  assign n5204 = n5190 & n5193 ;
  assign n5205 = n5195 & ~n5204 ;
  buffer buf_n5206( .i (n5205), .o (n5206) );
  assign n5208 = ~n5186 & n5206 ;
  buffer buf_n5209( .i (n5208), .o (n5209) );
  buffer buf_n5187( .i (n5186), .o (n5187) );
  buffer buf_n5207( .i (n5206), .o (n5207) );
  assign n5214 = n5187 & ~n5207 ;
  assign n5215 = n5209 | n5214 ;
  buffer buf_n5216( .i (n5215), .o (n5216) );
  assign n5218 = n5183 | n5216 ;
  buffer buf_n5219( .i (n5218), .o (n5219) );
  buffer buf_n5184( .i (n5183), .o (n5184) );
  buffer buf_n5217( .i (n5216), .o (n5217) );
  assign n5228 = n5184 & n5217 ;
  assign n5229 = n5219 & ~n5228 ;
  buffer buf_n5230( .i (n5229), .o (n5230) );
  assign n5232 = ~n5180 & n5230 ;
  buffer buf_n5233( .i (n5232), .o (n5233) );
  buffer buf_n5181( .i (n5180), .o (n5181) );
  buffer buf_n5231( .i (n5230), .o (n5231) );
  assign n5238 = n5181 & ~n5231 ;
  assign n5239 = n5233 | n5238 ;
  buffer buf_n5240( .i (n5239), .o (n5240) );
  assign n5242 = n5177 | n5240 ;
  buffer buf_n5243( .i (n5242), .o (n5243) );
  buffer buf_n5178( .i (n5177), .o (n5178) );
  buffer buf_n5241( .i (n5240), .o (n5241) );
  assign n5252 = n5178 & n5241 ;
  assign n5253 = n5243 & ~n5252 ;
  buffer buf_n5254( .i (n5253), .o (n5254) );
  assign n5256 = ~n5174 & n5254 ;
  buffer buf_n5257( .i (n5256), .o (n5257) );
  buffer buf_n5175( .i (n5174), .o (n5175) );
  buffer buf_n5255( .i (n5254), .o (n5255) );
  assign n5262 = n5175 & ~n5255 ;
  assign n5263 = n5257 | n5262 ;
  buffer buf_n5264( .i (n5263), .o (n5264) );
  assign n5266 = n5171 | n5264 ;
  buffer buf_n5267( .i (n5266), .o (n5267) );
  buffer buf_n5172( .i (n5171), .o (n5172) );
  buffer buf_n5265( .i (n5264), .o (n5265) );
  assign n5276 = n5172 & n5265 ;
  assign n5277 = n5267 & ~n5276 ;
  buffer buf_n5278( .i (n5277), .o (n5278) );
  assign n5280 = ~n5168 & n5278 ;
  buffer buf_n5281( .i (n5280), .o (n5281) );
  buffer buf_n5169( .i (n5168), .o (n5169) );
  buffer buf_n5279( .i (n5278), .o (n5279) );
  assign n5286 = n5169 & ~n5279 ;
  assign n5287 = n5281 | n5286 ;
  buffer buf_n5288( .i (n5287), .o (n5288) );
  assign n5290 = n5165 | n5288 ;
  buffer buf_n5291( .i (n5290), .o (n5291) );
  buffer buf_n5166( .i (n5165), .o (n5166) );
  buffer buf_n5289( .i (n5288), .o (n5289) );
  assign n5300 = n5166 & n5289 ;
  assign n5301 = n5291 & ~n5300 ;
  buffer buf_n5302( .i (n5301), .o (n5302) );
  assign n5304 = ~n5162 & n5302 ;
  buffer buf_n5305( .i (n5304), .o (n5305) );
  buffer buf_n5163( .i (n5162), .o (n5163) );
  buffer buf_n5303( .i (n5302), .o (n5303) );
  assign n5310 = n5163 & ~n5303 ;
  assign n5311 = n5305 | n5310 ;
  buffer buf_n5312( .i (n5311), .o (n5312) );
  assign n5314 = n5159 | n5312 ;
  buffer buf_n5315( .i (n5314), .o (n5315) );
  buffer buf_n5160( .i (n5159), .o (n5160) );
  buffer buf_n5313( .i (n5312), .o (n5313) );
  assign n5324 = n5160 & n5313 ;
  assign n5325 = n5315 & ~n5324 ;
  buffer buf_n5326( .i (n5325), .o (n5326) );
  assign n5328 = ~n5156 & n5326 ;
  buffer buf_n5329( .i (n5328), .o (n5329) );
  buffer buf_n5157( .i (n5156), .o (n5157) );
  buffer buf_n5327( .i (n5326), .o (n5327) );
  assign n5334 = n5157 & ~n5327 ;
  assign n5335 = n5329 | n5334 ;
  buffer buf_n5336( .i (n5335), .o (n5336) );
  assign n5338 = n5153 | n5336 ;
  buffer buf_n5339( .i (n5338), .o (n5339) );
  buffer buf_n5154( .i (n5153), .o (n5154) );
  buffer buf_n5337( .i (n5336), .o (n5337) );
  assign n5344 = n5154 & n5337 ;
  assign n5345 = n5339 & ~n5344 ;
  buffer buf_n5346( .i (n5345), .o (n5346) );
  assign n5348 = ~n5150 & n5346 ;
  buffer buf_n5349( .i (n5348), .o (n5349) );
  buffer buf_n5151( .i (n5150), .o (n5151) );
  buffer buf_n5347( .i (n5346), .o (n5347) );
  assign n5350 = n5151 & ~n5347 ;
  assign n5351 = n5349 | n5350 ;
  buffer buf_n5340( .i (n5339), .o (n5340) );
  buffer buf_n5341( .i (n5340), .o (n5341) );
  buffer buf_n5342( .i (n5341), .o (n5342) );
  buffer buf_n5343( .i (n5342), .o (n5343) );
  assign n5352 = n5343 & ~n5349 ;
  buffer buf_n5353( .i (n5352), .o (n5353) );
  buffer buf_n5316( .i (n5315), .o (n5316) );
  buffer buf_n5317( .i (n5316), .o (n5317) );
  buffer buf_n5318( .i (n5317), .o (n5318) );
  buffer buf_n5319( .i (n5318), .o (n5319) );
  buffer buf_n5320( .i (n5319), .o (n5320) );
  buffer buf_n5321( .i (n5320), .o (n5321) );
  buffer buf_n5322( .i (n5321), .o (n5322) );
  buffer buf_n5323( .i (n5322), .o (n5323) );
  buffer buf_n5330( .i (n5329), .o (n5330) );
  buffer buf_n5331( .i (n5330), .o (n5331) );
  buffer buf_n5332( .i (n5331), .o (n5332) );
  buffer buf_n5333( .i (n5332), .o (n5333) );
  assign n5355 = n5323 & ~n5333 ;
  buffer buf_n5356( .i (n5355), .o (n5356) );
  assign n5358 = N171 & N528 ;
  buffer buf_n5359( .i (n5358), .o (n5359) );
  buffer buf_n5292( .i (n5291), .o (n5292) );
  buffer buf_n5293( .i (n5292), .o (n5293) );
  buffer buf_n5294( .i (n5293), .o (n5294) );
  buffer buf_n5295( .i (n5294), .o (n5295) );
  buffer buf_n5296( .i (n5295), .o (n5296) );
  buffer buf_n5297( .i (n5296), .o (n5297) );
  buffer buf_n5298( .i (n5297), .o (n5298) );
  buffer buf_n5299( .i (n5298), .o (n5299) );
  buffer buf_n5306( .i (n5305), .o (n5306) );
  buffer buf_n5307( .i (n5306), .o (n5307) );
  buffer buf_n5308( .i (n5307), .o (n5308) );
  buffer buf_n5309( .i (n5308), .o (n5309) );
  assign n5361 = n5299 & ~n5309 ;
  buffer buf_n5362( .i (n5361), .o (n5362) );
  assign n5364 = N188 & N511 ;
  buffer buf_n5365( .i (n5364), .o (n5365) );
  buffer buf_n5268( .i (n5267), .o (n5268) );
  buffer buf_n5269( .i (n5268), .o (n5269) );
  buffer buf_n5270( .i (n5269), .o (n5270) );
  buffer buf_n5271( .i (n5270), .o (n5271) );
  buffer buf_n5272( .i (n5271), .o (n5272) );
  buffer buf_n5273( .i (n5272), .o (n5273) );
  buffer buf_n5274( .i (n5273), .o (n5274) );
  buffer buf_n5275( .i (n5274), .o (n5275) );
  buffer buf_n5282( .i (n5281), .o (n5282) );
  buffer buf_n5283( .i (n5282), .o (n5283) );
  buffer buf_n5284( .i (n5283), .o (n5284) );
  buffer buf_n5285( .i (n5284), .o (n5285) );
  assign n5367 = n5275 & ~n5285 ;
  buffer buf_n5368( .i (n5367), .o (n5368) );
  assign n5370 = N205 & N494 ;
  buffer buf_n5371( .i (n5370), .o (n5371) );
  buffer buf_n5244( .i (n5243), .o (n5244) );
  buffer buf_n5245( .i (n5244), .o (n5245) );
  buffer buf_n5246( .i (n5245), .o (n5246) );
  buffer buf_n5247( .i (n5246), .o (n5247) );
  buffer buf_n5248( .i (n5247), .o (n5248) );
  buffer buf_n5249( .i (n5248), .o (n5249) );
  buffer buf_n5250( .i (n5249), .o (n5250) );
  buffer buf_n5251( .i (n5250), .o (n5251) );
  buffer buf_n5258( .i (n5257), .o (n5258) );
  buffer buf_n5259( .i (n5258), .o (n5259) );
  buffer buf_n5260( .i (n5259), .o (n5260) );
  buffer buf_n5261( .i (n5260), .o (n5261) );
  assign n5373 = n5251 & ~n5261 ;
  buffer buf_n5374( .i (n5373), .o (n5374) );
  assign n5376 = N222 & N477 ;
  buffer buf_n5377( .i (n5376), .o (n5377) );
  buffer buf_n5220( .i (n5219), .o (n5220) );
  buffer buf_n5221( .i (n5220), .o (n5221) );
  buffer buf_n5222( .i (n5221), .o (n5222) );
  buffer buf_n5223( .i (n5222), .o (n5223) );
  buffer buf_n5224( .i (n5223), .o (n5224) );
  buffer buf_n5225( .i (n5224), .o (n5225) );
  buffer buf_n5226( .i (n5225), .o (n5226) );
  buffer buf_n5227( .i (n5226), .o (n5227) );
  buffer buf_n5234( .i (n5233), .o (n5234) );
  buffer buf_n5235( .i (n5234), .o (n5235) );
  buffer buf_n5236( .i (n5235), .o (n5236) );
  buffer buf_n5237( .i (n5236), .o (n5237) );
  assign n5379 = n5227 & ~n5237 ;
  buffer buf_n5380( .i (n5379), .o (n5380) );
  assign n5382 = N239 & N460 ;
  buffer buf_n5383( .i (n5382), .o (n5383) );
  assign n5385 = N256 & N443 ;
  buffer buf_n5386( .i (n5385), .o (n5386) );
  buffer buf_n5196( .i (n5195), .o (n5196) );
  buffer buf_n5197( .i (n5196), .o (n5197) );
  buffer buf_n5198( .i (n5197), .o (n5198) );
  buffer buf_n5199( .i (n5198), .o (n5199) );
  buffer buf_n5200( .i (n5199), .o (n5200) );
  buffer buf_n5201( .i (n5200), .o (n5201) );
  buffer buf_n5202( .i (n5201), .o (n5202) );
  buffer buf_n5203( .i (n5202), .o (n5203) );
  buffer buf_n5210( .i (n5209), .o (n5210) );
  buffer buf_n5211( .i (n5210), .o (n5211) );
  buffer buf_n5212( .i (n5211), .o (n5212) );
  buffer buf_n5213( .i (n5212), .o (n5213) );
  assign n5388 = n5203 & ~n5213 ;
  buffer buf_n5389( .i (n5388), .o (n5389) );
  assign n5391 = n5386 | n5389 ;
  buffer buf_n5392( .i (n5391), .o (n5392) );
  buffer buf_n5387( .i (n5386), .o (n5387) );
  buffer buf_n5390( .i (n5389), .o (n5390) );
  assign n5401 = n5387 & n5390 ;
  assign n5402 = n5392 & ~n5401 ;
  buffer buf_n5403( .i (n5402), .o (n5403) );
  assign n5405 = ~n5383 & n5403 ;
  buffer buf_n5406( .i (n5405), .o (n5406) );
  buffer buf_n5384( .i (n5383), .o (n5384) );
  buffer buf_n5404( .i (n5403), .o (n5404) );
  assign n5411 = n5384 & ~n5404 ;
  assign n5412 = n5406 | n5411 ;
  buffer buf_n5413( .i (n5412), .o (n5413) );
  assign n5415 = n5380 | n5413 ;
  buffer buf_n5416( .i (n5415), .o (n5416) );
  buffer buf_n5381( .i (n5380), .o (n5381) );
  buffer buf_n5414( .i (n5413), .o (n5414) );
  assign n5425 = n5381 & n5414 ;
  assign n5426 = n5416 & ~n5425 ;
  buffer buf_n5427( .i (n5426), .o (n5427) );
  assign n5429 = ~n5377 & n5427 ;
  buffer buf_n5430( .i (n5429), .o (n5430) );
  buffer buf_n5378( .i (n5377), .o (n5378) );
  buffer buf_n5428( .i (n5427), .o (n5428) );
  assign n5435 = n5378 & ~n5428 ;
  assign n5436 = n5430 | n5435 ;
  buffer buf_n5437( .i (n5436), .o (n5437) );
  assign n5439 = n5374 | n5437 ;
  buffer buf_n5440( .i (n5439), .o (n5440) );
  buffer buf_n5375( .i (n5374), .o (n5375) );
  buffer buf_n5438( .i (n5437), .o (n5438) );
  assign n5449 = n5375 & n5438 ;
  assign n5450 = n5440 & ~n5449 ;
  buffer buf_n5451( .i (n5450), .o (n5451) );
  assign n5453 = ~n5371 & n5451 ;
  buffer buf_n5454( .i (n5453), .o (n5454) );
  buffer buf_n5372( .i (n5371), .o (n5372) );
  buffer buf_n5452( .i (n5451), .o (n5452) );
  assign n5459 = n5372 & ~n5452 ;
  assign n5460 = n5454 | n5459 ;
  buffer buf_n5461( .i (n5460), .o (n5461) );
  assign n5463 = n5368 | n5461 ;
  buffer buf_n5464( .i (n5463), .o (n5464) );
  buffer buf_n5369( .i (n5368), .o (n5369) );
  buffer buf_n5462( .i (n5461), .o (n5462) );
  assign n5473 = n5369 & n5462 ;
  assign n5474 = n5464 & ~n5473 ;
  buffer buf_n5475( .i (n5474), .o (n5475) );
  assign n5477 = ~n5365 & n5475 ;
  buffer buf_n5478( .i (n5477), .o (n5478) );
  buffer buf_n5366( .i (n5365), .o (n5366) );
  buffer buf_n5476( .i (n5475), .o (n5476) );
  assign n5483 = n5366 & ~n5476 ;
  assign n5484 = n5478 | n5483 ;
  buffer buf_n5485( .i (n5484), .o (n5485) );
  assign n5487 = n5362 | n5485 ;
  buffer buf_n5488( .i (n5487), .o (n5488) );
  buffer buf_n5363( .i (n5362), .o (n5363) );
  buffer buf_n5486( .i (n5485), .o (n5486) );
  assign n5497 = n5363 & n5486 ;
  assign n5498 = n5488 & ~n5497 ;
  buffer buf_n5499( .i (n5498), .o (n5499) );
  assign n5501 = ~n5359 & n5499 ;
  buffer buf_n5502( .i (n5501), .o (n5502) );
  buffer buf_n5360( .i (n5359), .o (n5360) );
  buffer buf_n5500( .i (n5499), .o (n5500) );
  assign n5507 = n5360 & ~n5500 ;
  assign n5508 = n5502 | n5507 ;
  buffer buf_n5509( .i (n5508), .o (n5509) );
  assign n5511 = n5356 | n5509 ;
  buffer buf_n5512( .i (n5511), .o (n5512) );
  buffer buf_n5357( .i (n5356), .o (n5357) );
  buffer buf_n5510( .i (n5509), .o (n5510) );
  assign n5517 = n5357 & n5510 ;
  assign n5518 = n5512 & ~n5517 ;
  buffer buf_n5519( .i (n5518), .o (n5519) );
  assign n5521 = ~n5353 & n5519 ;
  buffer buf_n5522( .i (n5521), .o (n5522) );
  buffer buf_n5354( .i (n5353), .o (n5354) );
  buffer buf_n5520( .i (n5519), .o (n5520) );
  assign n5523 = n5354 & ~n5520 ;
  assign n5524 = n5522 | n5523 ;
  buffer buf_n5513( .i (n5512), .o (n5513) );
  buffer buf_n5514( .i (n5513), .o (n5514) );
  buffer buf_n5515( .i (n5514), .o (n5515) );
  buffer buf_n5516( .i (n5515), .o (n5516) );
  assign n5525 = n5516 & ~n5522 ;
  buffer buf_n5526( .i (n5525), .o (n5526) );
  buffer buf_n5489( .i (n5488), .o (n5489) );
  buffer buf_n5490( .i (n5489), .o (n5490) );
  buffer buf_n5491( .i (n5490), .o (n5491) );
  buffer buf_n5492( .i (n5491), .o (n5492) );
  buffer buf_n5493( .i (n5492), .o (n5493) );
  buffer buf_n5494( .i (n5493), .o (n5494) );
  buffer buf_n5495( .i (n5494), .o (n5495) );
  buffer buf_n5496( .i (n5495), .o (n5496) );
  buffer buf_n5503( .i (n5502), .o (n5503) );
  buffer buf_n5504( .i (n5503), .o (n5504) );
  buffer buf_n5505( .i (n5504), .o (n5505) );
  buffer buf_n5506( .i (n5505), .o (n5506) );
  assign n5528 = n5496 & ~n5506 ;
  buffer buf_n5529( .i (n5528), .o (n5529) );
  assign n5531 = N188 & N528 ;
  buffer buf_n5532( .i (n5531), .o (n5532) );
  buffer buf_n5465( .i (n5464), .o (n5465) );
  buffer buf_n5466( .i (n5465), .o (n5466) );
  buffer buf_n5467( .i (n5466), .o (n5467) );
  buffer buf_n5468( .i (n5467), .o (n5468) );
  buffer buf_n5469( .i (n5468), .o (n5469) );
  buffer buf_n5470( .i (n5469), .o (n5470) );
  buffer buf_n5471( .i (n5470), .o (n5471) );
  buffer buf_n5472( .i (n5471), .o (n5472) );
  buffer buf_n5479( .i (n5478), .o (n5479) );
  buffer buf_n5480( .i (n5479), .o (n5480) );
  buffer buf_n5481( .i (n5480), .o (n5481) );
  buffer buf_n5482( .i (n5481), .o (n5482) );
  assign n5534 = n5472 & ~n5482 ;
  buffer buf_n5535( .i (n5534), .o (n5535) );
  assign n5537 = N205 & N511 ;
  buffer buf_n5538( .i (n5537), .o (n5538) );
  buffer buf_n5441( .i (n5440), .o (n5441) );
  buffer buf_n5442( .i (n5441), .o (n5442) );
  buffer buf_n5443( .i (n5442), .o (n5443) );
  buffer buf_n5444( .i (n5443), .o (n5444) );
  buffer buf_n5445( .i (n5444), .o (n5445) );
  buffer buf_n5446( .i (n5445), .o (n5446) );
  buffer buf_n5447( .i (n5446), .o (n5447) );
  buffer buf_n5448( .i (n5447), .o (n5448) );
  buffer buf_n5455( .i (n5454), .o (n5455) );
  buffer buf_n5456( .i (n5455), .o (n5456) );
  buffer buf_n5457( .i (n5456), .o (n5457) );
  buffer buf_n5458( .i (n5457), .o (n5458) );
  assign n5540 = n5448 & ~n5458 ;
  buffer buf_n5541( .i (n5540), .o (n5541) );
  assign n5543 = N222 & N494 ;
  buffer buf_n5544( .i (n5543), .o (n5544) );
  buffer buf_n5417( .i (n5416), .o (n5417) );
  buffer buf_n5418( .i (n5417), .o (n5418) );
  buffer buf_n5419( .i (n5418), .o (n5419) );
  buffer buf_n5420( .i (n5419), .o (n5420) );
  buffer buf_n5421( .i (n5420), .o (n5421) );
  buffer buf_n5422( .i (n5421), .o (n5422) );
  buffer buf_n5423( .i (n5422), .o (n5423) );
  buffer buf_n5424( .i (n5423), .o (n5424) );
  buffer buf_n5431( .i (n5430), .o (n5431) );
  buffer buf_n5432( .i (n5431), .o (n5432) );
  buffer buf_n5433( .i (n5432), .o (n5433) );
  buffer buf_n5434( .i (n5433), .o (n5434) );
  assign n5546 = n5424 & ~n5434 ;
  buffer buf_n5547( .i (n5546), .o (n5547) );
  assign n5549 = N239 & N477 ;
  buffer buf_n5550( .i (n5549), .o (n5550) );
  assign n5552 = N256 & N460 ;
  buffer buf_n5553( .i (n5552), .o (n5553) );
  buffer buf_n5393( .i (n5392), .o (n5393) );
  buffer buf_n5394( .i (n5393), .o (n5394) );
  buffer buf_n5395( .i (n5394), .o (n5395) );
  buffer buf_n5396( .i (n5395), .o (n5396) );
  buffer buf_n5397( .i (n5396), .o (n5397) );
  buffer buf_n5398( .i (n5397), .o (n5398) );
  buffer buf_n5399( .i (n5398), .o (n5399) );
  buffer buf_n5400( .i (n5399), .o (n5400) );
  buffer buf_n5407( .i (n5406), .o (n5407) );
  buffer buf_n5408( .i (n5407), .o (n5408) );
  buffer buf_n5409( .i (n5408), .o (n5409) );
  buffer buf_n5410( .i (n5409), .o (n5410) );
  assign n5555 = n5400 & ~n5410 ;
  buffer buf_n5556( .i (n5555), .o (n5556) );
  assign n5558 = n5553 | n5556 ;
  buffer buf_n5559( .i (n5558), .o (n5559) );
  buffer buf_n5554( .i (n5553), .o (n5554) );
  buffer buf_n5557( .i (n5556), .o (n5557) );
  assign n5568 = n5554 & n5557 ;
  assign n5569 = n5559 & ~n5568 ;
  buffer buf_n5570( .i (n5569), .o (n5570) );
  assign n5572 = ~n5550 & n5570 ;
  buffer buf_n5573( .i (n5572), .o (n5573) );
  buffer buf_n5551( .i (n5550), .o (n5551) );
  buffer buf_n5571( .i (n5570), .o (n5571) );
  assign n5578 = n5551 & ~n5571 ;
  assign n5579 = n5573 | n5578 ;
  buffer buf_n5580( .i (n5579), .o (n5580) );
  assign n5582 = n5547 | n5580 ;
  buffer buf_n5583( .i (n5582), .o (n5583) );
  buffer buf_n5548( .i (n5547), .o (n5548) );
  buffer buf_n5581( .i (n5580), .o (n5581) );
  assign n5592 = n5548 & n5581 ;
  assign n5593 = n5583 & ~n5592 ;
  buffer buf_n5594( .i (n5593), .o (n5594) );
  assign n5596 = ~n5544 & n5594 ;
  buffer buf_n5597( .i (n5596), .o (n5597) );
  buffer buf_n5545( .i (n5544), .o (n5545) );
  buffer buf_n5595( .i (n5594), .o (n5595) );
  assign n5602 = n5545 & ~n5595 ;
  assign n5603 = n5597 | n5602 ;
  buffer buf_n5604( .i (n5603), .o (n5604) );
  assign n5606 = n5541 | n5604 ;
  buffer buf_n5607( .i (n5606), .o (n5607) );
  buffer buf_n5542( .i (n5541), .o (n5542) );
  buffer buf_n5605( .i (n5604), .o (n5605) );
  assign n5616 = n5542 & n5605 ;
  assign n5617 = n5607 & ~n5616 ;
  buffer buf_n5618( .i (n5617), .o (n5618) );
  assign n5620 = ~n5538 & n5618 ;
  buffer buf_n5621( .i (n5620), .o (n5621) );
  buffer buf_n5539( .i (n5538), .o (n5539) );
  buffer buf_n5619( .i (n5618), .o (n5619) );
  assign n5626 = n5539 & ~n5619 ;
  assign n5627 = n5621 | n5626 ;
  buffer buf_n5628( .i (n5627), .o (n5628) );
  assign n5630 = n5535 | n5628 ;
  buffer buf_n5631( .i (n5630), .o (n5631) );
  buffer buf_n5536( .i (n5535), .o (n5536) );
  buffer buf_n5629( .i (n5628), .o (n5629) );
  assign n5640 = n5536 & n5629 ;
  assign n5641 = n5631 & ~n5640 ;
  buffer buf_n5642( .i (n5641), .o (n5642) );
  assign n5644 = ~n5532 & n5642 ;
  buffer buf_n5645( .i (n5644), .o (n5645) );
  buffer buf_n5533( .i (n5532), .o (n5533) );
  buffer buf_n5643( .i (n5642), .o (n5643) );
  assign n5650 = n5533 & ~n5643 ;
  assign n5651 = n5645 | n5650 ;
  buffer buf_n5652( .i (n5651), .o (n5652) );
  assign n5654 = n5529 | n5652 ;
  buffer buf_n5655( .i (n5654), .o (n5655) );
  buffer buf_n5530( .i (n5529), .o (n5530) );
  buffer buf_n5653( .i (n5652), .o (n5653) );
  assign n5660 = n5530 & n5653 ;
  assign n5661 = n5655 & ~n5660 ;
  buffer buf_n5662( .i (n5661), .o (n5662) );
  assign n5664 = ~n5526 & n5662 ;
  buffer buf_n5665( .i (n5664), .o (n5665) );
  buffer buf_n5527( .i (n5526), .o (n5527) );
  buffer buf_n5663( .i (n5662), .o (n5663) );
  assign n5666 = n5527 & ~n5663 ;
  assign n5667 = n5665 | n5666 ;
  buffer buf_n5656( .i (n5655), .o (n5656) );
  buffer buf_n5657( .i (n5656), .o (n5657) );
  buffer buf_n5658( .i (n5657), .o (n5658) );
  buffer buf_n5659( .i (n5658), .o (n5659) );
  assign n5668 = n5659 & ~n5665 ;
  buffer buf_n5669( .i (n5668), .o (n5669) );
  buffer buf_n5632( .i (n5631), .o (n5632) );
  buffer buf_n5633( .i (n5632), .o (n5633) );
  buffer buf_n5634( .i (n5633), .o (n5634) );
  buffer buf_n5635( .i (n5634), .o (n5635) );
  buffer buf_n5636( .i (n5635), .o (n5636) );
  buffer buf_n5637( .i (n5636), .o (n5637) );
  buffer buf_n5638( .i (n5637), .o (n5638) );
  buffer buf_n5639( .i (n5638), .o (n5639) );
  buffer buf_n5646( .i (n5645), .o (n5646) );
  buffer buf_n5647( .i (n5646), .o (n5647) );
  buffer buf_n5648( .i (n5647), .o (n5648) );
  buffer buf_n5649( .i (n5648), .o (n5649) );
  assign n5671 = n5639 & ~n5649 ;
  buffer buf_n5672( .i (n5671), .o (n5672) );
  assign n5674 = N205 & N528 ;
  buffer buf_n5675( .i (n5674), .o (n5675) );
  buffer buf_n5608( .i (n5607), .o (n5608) );
  buffer buf_n5609( .i (n5608), .o (n5609) );
  buffer buf_n5610( .i (n5609), .o (n5610) );
  buffer buf_n5611( .i (n5610), .o (n5611) );
  buffer buf_n5612( .i (n5611), .o (n5612) );
  buffer buf_n5613( .i (n5612), .o (n5613) );
  buffer buf_n5614( .i (n5613), .o (n5614) );
  buffer buf_n5615( .i (n5614), .o (n5615) );
  buffer buf_n5622( .i (n5621), .o (n5622) );
  buffer buf_n5623( .i (n5622), .o (n5623) );
  buffer buf_n5624( .i (n5623), .o (n5624) );
  buffer buf_n5625( .i (n5624), .o (n5625) );
  assign n5677 = n5615 & ~n5625 ;
  buffer buf_n5678( .i (n5677), .o (n5678) );
  assign n5680 = N222 & N511 ;
  buffer buf_n5681( .i (n5680), .o (n5681) );
  buffer buf_n5584( .i (n5583), .o (n5584) );
  buffer buf_n5585( .i (n5584), .o (n5585) );
  buffer buf_n5586( .i (n5585), .o (n5586) );
  buffer buf_n5587( .i (n5586), .o (n5587) );
  buffer buf_n5588( .i (n5587), .o (n5588) );
  buffer buf_n5589( .i (n5588), .o (n5589) );
  buffer buf_n5590( .i (n5589), .o (n5590) );
  buffer buf_n5591( .i (n5590), .o (n5591) );
  buffer buf_n5598( .i (n5597), .o (n5598) );
  buffer buf_n5599( .i (n5598), .o (n5599) );
  buffer buf_n5600( .i (n5599), .o (n5600) );
  buffer buf_n5601( .i (n5600), .o (n5601) );
  assign n5683 = n5591 & ~n5601 ;
  buffer buf_n5684( .i (n5683), .o (n5684) );
  assign n5686 = N239 & N494 ;
  buffer buf_n5687( .i (n5686), .o (n5687) );
  assign n5689 = N256 & N477 ;
  buffer buf_n5690( .i (n5689), .o (n5690) );
  buffer buf_n5560( .i (n5559), .o (n5560) );
  buffer buf_n5561( .i (n5560), .o (n5561) );
  buffer buf_n5562( .i (n5561), .o (n5562) );
  buffer buf_n5563( .i (n5562), .o (n5563) );
  buffer buf_n5564( .i (n5563), .o (n5564) );
  buffer buf_n5565( .i (n5564), .o (n5565) );
  buffer buf_n5566( .i (n5565), .o (n5566) );
  buffer buf_n5567( .i (n5566), .o (n5567) );
  buffer buf_n5574( .i (n5573), .o (n5574) );
  buffer buf_n5575( .i (n5574), .o (n5575) );
  buffer buf_n5576( .i (n5575), .o (n5576) );
  buffer buf_n5577( .i (n5576), .o (n5577) );
  assign n5692 = n5567 & ~n5577 ;
  buffer buf_n5693( .i (n5692), .o (n5693) );
  assign n5695 = n5690 | n5693 ;
  buffer buf_n5696( .i (n5695), .o (n5696) );
  buffer buf_n5691( .i (n5690), .o (n5691) );
  buffer buf_n5694( .i (n5693), .o (n5694) );
  assign n5705 = n5691 & n5694 ;
  assign n5706 = n5696 & ~n5705 ;
  buffer buf_n5707( .i (n5706), .o (n5707) );
  assign n5709 = ~n5687 & n5707 ;
  buffer buf_n5710( .i (n5709), .o (n5710) );
  buffer buf_n5688( .i (n5687), .o (n5688) );
  buffer buf_n5708( .i (n5707), .o (n5708) );
  assign n5715 = n5688 & ~n5708 ;
  assign n5716 = n5710 | n5715 ;
  buffer buf_n5717( .i (n5716), .o (n5717) );
  assign n5719 = n5684 | n5717 ;
  buffer buf_n5720( .i (n5719), .o (n5720) );
  buffer buf_n5685( .i (n5684), .o (n5685) );
  buffer buf_n5718( .i (n5717), .o (n5718) );
  assign n5729 = n5685 & n5718 ;
  assign n5730 = n5720 & ~n5729 ;
  buffer buf_n5731( .i (n5730), .o (n5731) );
  assign n5733 = ~n5681 & n5731 ;
  buffer buf_n5734( .i (n5733), .o (n5734) );
  buffer buf_n5682( .i (n5681), .o (n5682) );
  buffer buf_n5732( .i (n5731), .o (n5732) );
  assign n5739 = n5682 & ~n5732 ;
  assign n5740 = n5734 | n5739 ;
  buffer buf_n5741( .i (n5740), .o (n5741) );
  assign n5743 = n5678 | n5741 ;
  buffer buf_n5744( .i (n5743), .o (n5744) );
  buffer buf_n5679( .i (n5678), .o (n5679) );
  buffer buf_n5742( .i (n5741), .o (n5742) );
  assign n5753 = n5679 & n5742 ;
  assign n5754 = n5744 & ~n5753 ;
  buffer buf_n5755( .i (n5754), .o (n5755) );
  assign n5757 = ~n5675 & n5755 ;
  buffer buf_n5758( .i (n5757), .o (n5758) );
  buffer buf_n5676( .i (n5675), .o (n5676) );
  buffer buf_n5756( .i (n5755), .o (n5756) );
  assign n5763 = n5676 & ~n5756 ;
  assign n5764 = n5758 | n5763 ;
  buffer buf_n5765( .i (n5764), .o (n5765) );
  assign n5767 = n5672 | n5765 ;
  buffer buf_n5768( .i (n5767), .o (n5768) );
  buffer buf_n5673( .i (n5672), .o (n5673) );
  buffer buf_n5766( .i (n5765), .o (n5766) );
  assign n5773 = n5673 & n5766 ;
  assign n5774 = n5768 & ~n5773 ;
  buffer buf_n5775( .i (n5774), .o (n5775) );
  assign n5777 = ~n5669 & n5775 ;
  buffer buf_n5778( .i (n5777), .o (n5778) );
  buffer buf_n5670( .i (n5669), .o (n5670) );
  buffer buf_n5776( .i (n5775), .o (n5776) );
  assign n5779 = n5670 & ~n5776 ;
  assign n5780 = n5778 | n5779 ;
  buffer buf_n5769( .i (n5768), .o (n5769) );
  buffer buf_n5770( .i (n5769), .o (n5770) );
  buffer buf_n5771( .i (n5770), .o (n5771) );
  buffer buf_n5772( .i (n5771), .o (n5772) );
  assign n5781 = n5772 & ~n5778 ;
  buffer buf_n5782( .i (n5781), .o (n5782) );
  buffer buf_n5745( .i (n5744), .o (n5745) );
  buffer buf_n5746( .i (n5745), .o (n5746) );
  buffer buf_n5747( .i (n5746), .o (n5747) );
  buffer buf_n5748( .i (n5747), .o (n5748) );
  buffer buf_n5749( .i (n5748), .o (n5749) );
  buffer buf_n5750( .i (n5749), .o (n5750) );
  buffer buf_n5751( .i (n5750), .o (n5751) );
  buffer buf_n5752( .i (n5751), .o (n5752) );
  buffer buf_n5759( .i (n5758), .o (n5759) );
  buffer buf_n5760( .i (n5759), .o (n5760) );
  buffer buf_n5761( .i (n5760), .o (n5761) );
  buffer buf_n5762( .i (n5761), .o (n5762) );
  assign n5784 = n5752 & ~n5762 ;
  buffer buf_n5785( .i (n5784), .o (n5785) );
  assign n5787 = N222 & N528 ;
  buffer buf_n5788( .i (n5787), .o (n5788) );
  buffer buf_n5721( .i (n5720), .o (n5721) );
  buffer buf_n5722( .i (n5721), .o (n5722) );
  buffer buf_n5723( .i (n5722), .o (n5723) );
  buffer buf_n5724( .i (n5723), .o (n5724) );
  buffer buf_n5725( .i (n5724), .o (n5725) );
  buffer buf_n5726( .i (n5725), .o (n5726) );
  buffer buf_n5727( .i (n5726), .o (n5727) );
  buffer buf_n5728( .i (n5727), .o (n5728) );
  buffer buf_n5735( .i (n5734), .o (n5735) );
  buffer buf_n5736( .i (n5735), .o (n5736) );
  buffer buf_n5737( .i (n5736), .o (n5737) );
  buffer buf_n5738( .i (n5737), .o (n5738) );
  assign n5790 = n5728 & ~n5738 ;
  buffer buf_n5791( .i (n5790), .o (n5791) );
  assign n5793 = N239 & N511 ;
  buffer buf_n5794( .i (n5793), .o (n5794) );
  assign n5796 = N256 & N494 ;
  buffer buf_n5797( .i (n5796), .o (n5797) );
  buffer buf_n5697( .i (n5696), .o (n5697) );
  buffer buf_n5698( .i (n5697), .o (n5698) );
  buffer buf_n5699( .i (n5698), .o (n5699) );
  buffer buf_n5700( .i (n5699), .o (n5700) );
  buffer buf_n5701( .i (n5700), .o (n5701) );
  buffer buf_n5702( .i (n5701), .o (n5702) );
  buffer buf_n5703( .i (n5702), .o (n5703) );
  buffer buf_n5704( .i (n5703), .o (n5704) );
  buffer buf_n5711( .i (n5710), .o (n5711) );
  buffer buf_n5712( .i (n5711), .o (n5712) );
  buffer buf_n5713( .i (n5712), .o (n5713) );
  buffer buf_n5714( .i (n5713), .o (n5714) );
  assign n5799 = n5704 & ~n5714 ;
  buffer buf_n5800( .i (n5799), .o (n5800) );
  assign n5802 = n5797 | n5800 ;
  buffer buf_n5803( .i (n5802), .o (n5803) );
  buffer buf_n5798( .i (n5797), .o (n5798) );
  buffer buf_n5801( .i (n5800), .o (n5801) );
  assign n5812 = n5798 & n5801 ;
  assign n5813 = n5803 & ~n5812 ;
  buffer buf_n5814( .i (n5813), .o (n5814) );
  assign n5816 = ~n5794 & n5814 ;
  buffer buf_n5817( .i (n5816), .o (n5817) );
  buffer buf_n5795( .i (n5794), .o (n5795) );
  buffer buf_n5815( .i (n5814), .o (n5815) );
  assign n5822 = n5795 & ~n5815 ;
  assign n5823 = n5817 | n5822 ;
  buffer buf_n5824( .i (n5823), .o (n5824) );
  assign n5826 = n5791 | n5824 ;
  buffer buf_n5827( .i (n5826), .o (n5827) );
  buffer buf_n5792( .i (n5791), .o (n5792) );
  buffer buf_n5825( .i (n5824), .o (n5825) );
  assign n5836 = n5792 & n5825 ;
  assign n5837 = n5827 & ~n5836 ;
  buffer buf_n5838( .i (n5837), .o (n5838) );
  assign n5840 = ~n5788 & n5838 ;
  buffer buf_n5841( .i (n5840), .o (n5841) );
  buffer buf_n5789( .i (n5788), .o (n5789) );
  buffer buf_n5839( .i (n5838), .o (n5839) );
  assign n5846 = n5789 & ~n5839 ;
  assign n5847 = n5841 | n5846 ;
  buffer buf_n5848( .i (n5847), .o (n5848) );
  assign n5850 = n5785 | n5848 ;
  buffer buf_n5851( .i (n5850), .o (n5851) );
  buffer buf_n5786( .i (n5785), .o (n5786) );
  buffer buf_n5849( .i (n5848), .o (n5849) );
  assign n5856 = n5786 & n5849 ;
  assign n5857 = n5851 & ~n5856 ;
  buffer buf_n5858( .i (n5857), .o (n5858) );
  assign n5860 = ~n5782 & n5858 ;
  buffer buf_n5861( .i (n5860), .o (n5861) );
  buffer buf_n5783( .i (n5782), .o (n5783) );
  buffer buf_n5859( .i (n5858), .o (n5859) );
  assign n5862 = n5783 & ~n5859 ;
  assign n5863 = n5861 | n5862 ;
  buffer buf_n5852( .i (n5851), .o (n5852) );
  buffer buf_n5853( .i (n5852), .o (n5853) );
  buffer buf_n5854( .i (n5853), .o (n5854) );
  buffer buf_n5855( .i (n5854), .o (n5855) );
  assign n5864 = n5855 & ~n5861 ;
  buffer buf_n5865( .i (n5864), .o (n5865) );
  buffer buf_n5828( .i (n5827), .o (n5828) );
  buffer buf_n5829( .i (n5828), .o (n5829) );
  buffer buf_n5830( .i (n5829), .o (n5830) );
  buffer buf_n5831( .i (n5830), .o (n5831) );
  buffer buf_n5832( .i (n5831), .o (n5832) );
  buffer buf_n5833( .i (n5832), .o (n5833) );
  buffer buf_n5834( .i (n5833), .o (n5834) );
  buffer buf_n5835( .i (n5834), .o (n5835) );
  buffer buf_n5842( .i (n5841), .o (n5842) );
  buffer buf_n5843( .i (n5842), .o (n5843) );
  buffer buf_n5844( .i (n5843), .o (n5844) );
  buffer buf_n5845( .i (n5844), .o (n5845) );
  assign n5867 = n5835 & ~n5845 ;
  buffer buf_n5868( .i (n5867), .o (n5868) );
  assign n5870 = N239 & N528 ;
  buffer buf_n5871( .i (n5870), .o (n5871) );
  assign n5873 = N256 & N511 ;
  buffer buf_n5874( .i (n5873), .o (n5874) );
  buffer buf_n5804( .i (n5803), .o (n5804) );
  buffer buf_n5805( .i (n5804), .o (n5805) );
  buffer buf_n5806( .i (n5805), .o (n5806) );
  buffer buf_n5807( .i (n5806), .o (n5807) );
  buffer buf_n5808( .i (n5807), .o (n5808) );
  buffer buf_n5809( .i (n5808), .o (n5809) );
  buffer buf_n5810( .i (n5809), .o (n5810) );
  buffer buf_n5811( .i (n5810), .o (n5811) );
  buffer buf_n5818( .i (n5817), .o (n5818) );
  buffer buf_n5819( .i (n5818), .o (n5819) );
  buffer buf_n5820( .i (n5819), .o (n5820) );
  buffer buf_n5821( .i (n5820), .o (n5821) );
  assign n5876 = n5811 & ~n5821 ;
  buffer buf_n5877( .i (n5876), .o (n5877) );
  assign n5879 = n5874 | n5877 ;
  buffer buf_n5880( .i (n5879), .o (n5880) );
  buffer buf_n5875( .i (n5874), .o (n5875) );
  buffer buf_n5878( .i (n5877), .o (n5878) );
  assign n5889 = n5875 & n5878 ;
  assign n5890 = n5880 & ~n5889 ;
  buffer buf_n5891( .i (n5890), .o (n5891) );
  assign n5893 = ~n5871 & n5891 ;
  buffer buf_n5894( .i (n5893), .o (n5894) );
  buffer buf_n5872( .i (n5871), .o (n5872) );
  buffer buf_n5892( .i (n5891), .o (n5892) );
  assign n5899 = n5872 & ~n5892 ;
  assign n5900 = n5894 | n5899 ;
  buffer buf_n5901( .i (n5900), .o (n5901) );
  assign n5903 = n5868 | n5901 ;
  buffer buf_n5904( .i (n5903), .o (n5904) );
  buffer buf_n5869( .i (n5868), .o (n5869) );
  buffer buf_n5902( .i (n5901), .o (n5902) );
  assign n5909 = n5869 & n5902 ;
  assign n5910 = n5904 & ~n5909 ;
  buffer buf_n5911( .i (n5910), .o (n5911) );
  assign n5913 = ~n5865 & n5911 ;
  buffer buf_n5914( .i (n5913), .o (n5914) );
  buffer buf_n5866( .i (n5865), .o (n5866) );
  buffer buf_n5912( .i (n5911), .o (n5912) );
  assign n5915 = n5866 & ~n5912 ;
  assign n5916 = n5914 | n5915 ;
  assign n5917 = N256 & N528 ;
  buffer buf_n5918( .i (n5917), .o (n5918) );
  buffer buf_n5881( .i (n5880), .o (n5881) );
  buffer buf_n5882( .i (n5881), .o (n5882) );
  buffer buf_n5883( .i (n5882), .o (n5883) );
  buffer buf_n5884( .i (n5883), .o (n5884) );
  buffer buf_n5885( .i (n5884), .o (n5885) );
  buffer buf_n5886( .i (n5885), .o (n5886) );
  buffer buf_n5887( .i (n5886), .o (n5887) );
  buffer buf_n5888( .i (n5887), .o (n5888) );
  buffer buf_n5895( .i (n5894), .o (n5895) );
  buffer buf_n5896( .i (n5895), .o (n5896) );
  buffer buf_n5897( .i (n5896), .o (n5897) );
  buffer buf_n5898( .i (n5897), .o (n5898) );
  assign n5920 = n5888 & ~n5898 ;
  buffer buf_n5921( .i (n5920), .o (n5921) );
  assign n5923 = n5918 | n5921 ;
  buffer buf_n5924( .i (n5923), .o (n5924) );
  buffer buf_n5925( .i (n5924), .o (n5925) );
  buffer buf_n5926( .i (n5925), .o (n5926) );
  buffer buf_n5927( .i (n5926), .o (n5927) );
  buffer buf_n5928( .i (n5927), .o (n5928) );
  buffer buf_n5905( .i (n5904), .o (n5905) );
  buffer buf_n5906( .i (n5905), .o (n5906) );
  buffer buf_n5907( .i (n5906), .o (n5907) );
  buffer buf_n5908( .i (n5907), .o (n5908) );
  assign n5929 = n5908 & ~n5914 ;
  buffer buf_n5930( .i (n5929), .o (n5930) );
  buffer buf_n5919( .i (n5918), .o (n5919) );
  buffer buf_n5922( .i (n5921), .o (n5922) );
  assign n5932 = n5919 & n5922 ;
  assign n5933 = n5924 & ~n5932 ;
  buffer buf_n5934( .i (n5933), .o (n5934) );
  assign n5936 = ~n5930 & n5934 ;
  buffer buf_n5937( .i (n5936), .o (n5937) );
  assign n5938 = n5928 & ~n5937 ;
  buffer buf_n5931( .i (n5930), .o (n5931) );
  buffer buf_n5935( .i (n5934), .o (n5935) );
  assign n5939 = n5931 & ~n5935 ;
  assign n5940 = n5937 | n5939 ;
  assign N1581 = n48 ;
  assign N1901 = n80 ;
  assign N2223 = n140 ;
  assign N2548 = n222 ;
  assign N2877 = n326 ;
  assign N3211 = n452 ;
  assign N3552 = n600 ;
  assign N3895 = n770 ;
  assign N4241 = n962 ;
  assign N4591 = n1176 ;
  assign N4946 = n1412 ;
  assign N5308 = n1670 ;
  assign N545 = n37 ;
  assign N5672 = n1950 ;
  assign N5971 = n2258 ;
  assign N6123 = n2572 ;
  assign N6150 = n2890 ;
  assign N6160 = n3300 ;
  assign N6170 = n3683 ;
  assign N6180 = n4036 ;
  assign N6190 = n4359 ;
  assign N6200 = n4652 ;
  assign N6210 = n4915 ;
  assign N6220 = n5148 ;
  assign N6230 = n5351 ;
  assign N6240 = n5524 ;
  assign N6250 = n5667 ;
  assign N6260 = n5780 ;
  assign N6270 = n5863 ;
  assign N6280 = n5916 ;
  assign N6287 = n5938 ;
  assign N6288 = n5940 ;
endmodule
