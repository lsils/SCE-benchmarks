module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 ;
  wire n2 , n4 , n6 , n8 , n10 , n12 , n13 , n15 , n17 , n19 , n21 , n23 , n24 , n26 , n27 , n29 , n31 , n32 , n34 , n36 , n38 , n39 , n41 , n43 , n45 , n47 , n49 , n51 , n52 , n54 , n56 , n57 , n59 , n61 , n63 , n65 , n67 , n68 , n70 , n72 , n73 , n75 , n77 , n79 , n80 , n82 , n83 , n85 , n87 , n89 , n91 , n93 , n94 , n96 , n97 , n99 , n100 , n102 , n104 , n105 , n107 , n109 , n110 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 ;
  buffer buf_n96( .i (x41), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n41( .i (x17), .o (n41) );
  buffer buf_n54( .i (x23), .o (n54) );
  assign n113 = n41 & n54 ;
  assign n114 = n97 & n113 ;
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n38( .i (x16), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n34( .i (x14), .o (n34) );
  buffer buf_n75( .i (x32), .o (n75) );
  assign n116 = n34 | n75 ;
  assign n117 = n39 | n116 ;
  buffer buf_n118( .i (n117), .o (n118) );
  assign n119 = n115 & n118 ;
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  assign n122 = n41 | n54 ;
  assign n123 = n97 | n122 ;
  buffer buf_n124( .i (n123), .o (n124) );
  assign n125 = n34 & n75 ;
  assign n126 = n39 & n125 ;
  buffer buf_n127( .i (n126), .o (n127) );
  assign n128 = n124 & n127 ;
  buffer buf_n129( .i (n128), .o (n129) );
  assign n130 = ( n41 & n54 ) | ( n41 & n96 ) | ( n54 & n96 ) ;
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  assign n133 = ( n34 & n38 ) | ( n34 & n75 ) | ( n38 & n75 ) ;
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  assign n136 = n132 & n135 ;
  buffer buf_n137( .i (n136), .o (n137) );
  assign n138 = n129 & n137 ;
  assign n139 = n121 & n138 ;
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n12( .i (x5), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n70( .i (x30), .o (n70) );
  buffer buf_n85( .i (x36), .o (n85) );
  assign n141 = n70 & n85 ;
  assign n142 = n13 & n141 ;
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n99( .i (x42), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n43( .i (x18), .o (n43) );
  buffer buf_n89( .i (x38), .o (n89) );
  assign n144 = n43 | n89 ;
  assign n145 = n100 | n144 ;
  buffer buf_n146( .i (n145), .o (n146) );
  assign n147 = n143 | n146 ;
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  assign n150 = ( n12 & n70 ) | ( n12 & n85 ) | ( n70 & n85 ) ;
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  assign n153 = ( n43 & n89 ) | ( n43 & n99 ) | ( n89 & n99 ) ;
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  assign n156 = n152 | n155 ;
  buffer buf_n157( .i (n156), .o (n157) );
  assign n158 = n70 | n85 ;
  assign n159 = n13 | n158 ;
  buffer buf_n160( .i (n159), .o (n160) );
  assign n161 = n43 & n89 ;
  assign n162 = n100 & n161 ;
  buffer buf_n163( .i (n162), .o (n163) );
  assign n164 = n160 | n163 ;
  buffer buf_n165( .i (n164), .o (n165) );
  assign n166 = n157 | n165 ;
  assign n167 = n149 | n166 ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = n140 & n168 ;
  buffer buf_n170( .i (n169), .o (n170) );
  assign n171 = n115 | n118 ;
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  assign n174 = n124 | n127 ;
  buffer buf_n175( .i (n174), .o (n175) );
  assign n176 = n132 | n135 ;
  buffer buf_n177( .i (n176), .o (n177) );
  assign n178 = n175 & n177 ;
  assign n179 = n173 & n178 ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = n143 & n146 ;
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  assign n184 = n152 & n155 ;
  buffer buf_n185( .i (n184), .o (n185) );
  assign n186 = n160 & n163 ;
  buffer buf_n187( .i (n186), .o (n187) );
  assign n188 = n185 | n187 ;
  assign n189 = n183 | n188 ;
  buffer buf_n190( .i (n189), .o (n190) );
  assign n191 = n180 & n190 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = n170 & n192 ;
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  assign n196 = ( n120 & n129 ) | ( n120 & n137 ) | ( n129 & n137 ) ;
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  assign n199 = ( n148 & n157 ) | ( n148 & n165 ) | ( n157 & n165 ) ;
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  assign n202 = n198 & n201 ;
  buffer buf_n203( .i (n202), .o (n203) );
  assign n204 = ( n172 & n175 ) | ( n172 & n177 ) | ( n175 & n177 ) ;
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  assign n207 = ( n182 & n185 ) | ( n182 & n187 ) | ( n185 & n187 ) ;
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  assign n210 = n206 & n209 ;
  buffer buf_n211( .i (n210), .o (n211) );
  assign n212 = n203 & n211 ;
  buffer buf_n213( .i (n212), .o (n213) );
  assign n214 = n129 | n137 ;
  assign n215 = n121 | n214 ;
  buffer buf_n216( .i (n215), .o (n216) );
  assign n217 = n157 & n165 ;
  assign n218 = n149 & n217 ;
  buffer buf_n219( .i (n218), .o (n219) );
  assign n220 = n216 & n219 ;
  buffer buf_n221( .i (n220), .o (n221) );
  assign n222 = n175 | n177 ;
  assign n223 = n173 | n222 ;
  buffer buf_n224( .i (n223), .o (n224) );
  assign n225 = n185 & n187 ;
  assign n226 = n183 & n225 ;
  buffer buf_n227( .i (n226), .o (n227) );
  assign n228 = n224 & n227 ;
  buffer buf_n229( .i (n228), .o (n229) );
  assign n230 = n221 & n229 ;
  buffer buf_n231( .i (n230), .o (n231) );
  assign n232 = n213 & n231 ;
  assign n233 = n195 & n232 ;
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n109( .i (x46), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n17( .i (x7), .o (n17) );
  buffer buf_n61( .i (x26), .o (n61) );
  assign n235 = n17 & n61 ;
  assign n236 = n110 & n235 ;
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n79( .i (x34), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n6( .i (x2), .o (n6) );
  buffer buf_n65( .i (x28), .o (n65) );
  assign n238 = n6 | n65 ;
  assign n239 = n80 | n238 ;
  buffer buf_n240( .i (n239), .o (n240) );
  assign n241 = n237 & n240 ;
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  assign n244 = n17 | n61 ;
  assign n245 = n110 | n244 ;
  buffer buf_n246( .i (n245), .o (n246) );
  assign n247 = n6 & n65 ;
  assign n248 = n80 & n247 ;
  buffer buf_n249( .i (n248), .o (n249) );
  assign n250 = n246 & n249 ;
  buffer buf_n251( .i (n250), .o (n251) );
  assign n252 = ( n17 & n61 ) | ( n17 & n109 ) | ( n61 & n109 ) ;
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  assign n255 = ( n6 & n65 ) | ( n6 & n79 ) | ( n65 & n79 ) ;
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  assign n258 = n254 & n257 ;
  buffer buf_n259( .i (n258), .o (n259) );
  assign n260 = n251 | n259 ;
  assign n261 = n243 | n260 ;
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n8( .i (x3), .o (n8) );
  buffer buf_n56( .i (x24), .o (n56) );
  assign n263 = ( n2 & n8 ) | ( n2 & n56 ) | ( n8 & n56 ) ;
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n19( .i (x8), .o (n19) );
  buffer buf_n51( .i (x22), .o (n51) );
  buffer buf_n87( .i (x37), .o (n87) );
  assign n266 = ( n19 & n51 ) | ( n19 & n87 ) | ( n51 & n87 ) ;
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  assign n269 = n265 | n268 ;
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n57( .i (n56), .o (n57) );
  assign n271 = n2 & n8 ;
  assign n272 = n57 & n271 ;
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n52( .i (n51), .o (n52) );
  assign n274 = n19 | n87 ;
  assign n275 = n52 | n274 ;
  buffer buf_n276( .i (n275), .o (n276) );
  assign n277 = n273 | n276 ;
  buffer buf_n278( .i (n277), .o (n278) );
  assign n279 = n270 & n278 ;
  assign n280 = n19 & n87 ;
  assign n281 = n52 & n280 ;
  buffer buf_n282( .i (n281), .o (n282) );
  assign n283 = n2 | n8 ;
  assign n284 = n57 | n283 ;
  buffer buf_n285( .i (n284), .o (n285) );
  assign n286 = n282 | n285 ;
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  assign n289 = n279 & n288 ;
  buffer buf_n290( .i (n289), .o (n290) );
  assign n291 = n262 | n290 ;
  buffer buf_n292( .i (n291), .o (n292) );
  assign n293 = n237 | n240 ;
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = n246 | n249 ;
  buffer buf_n297( .i (n296), .o (n297) );
  assign n298 = n254 | n257 ;
  buffer buf_n299( .i (n298), .o (n299) );
  assign n300 = n297 | n299 ;
  assign n301 = n295 | n300 ;
  buffer buf_n302( .i (n301), .o (n302) );
  assign n303 = n265 & n268 ;
  buffer buf_n304( .i (n303), .o (n304) );
  assign n305 = n273 & n276 ;
  buffer buf_n306( .i (n305), .o (n306) );
  assign n307 = n304 & n306 ;
  assign n308 = n282 & n285 ;
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  assign n311 = n307 & n310 ;
  buffer buf_n312( .i (n311), .o (n312) );
  assign n313 = n302 | n312 ;
  buffer buf_n314( .i (n313), .o (n314) );
  assign n315 = n292 | n314 ;
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  assign n318 = n251 & n259 ;
  assign n319 = n243 & n318 ;
  buffer buf_n320( .i (n319), .o (n320) );
  assign n321 = n270 | n278 ;
  assign n322 = n288 | n321 ;
  buffer buf_n323( .i (n322), .o (n323) );
  assign n324 = n320 | n323 ;
  buffer buf_n325( .i (n324), .o (n325) );
  assign n326 = n297 & n299 ;
  assign n327 = n295 & n326 ;
  buffer buf_n328( .i (n327), .o (n328) );
  assign n329 = n304 | n306 ;
  assign n330 = n310 | n329 ;
  buffer buf_n331( .i (n330), .o (n331) );
  assign n332 = n328 | n331 ;
  buffer buf_n333( .i (n332), .o (n333) );
  assign n334 = n325 | n333 ;
  buffer buf_n335( .i (n334), .o (n335) );
  assign n336 = ( n242 & n251 ) | ( n242 & n259 ) | ( n251 & n259 ) ;
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  assign n339 = ( n270 & n278 ) | ( n270 & n287 ) | ( n278 & n287 ) ;
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  assign n342 = n338 | n341 ;
  buffer buf_n343( .i (n342), .o (n343) );
  assign n344 = ( n294 & n297 ) | ( n294 & n299 ) | ( n297 & n299 ) ;
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  assign n347 = ( n304 & n306 ) | ( n304 & n309 ) | ( n306 & n309 ) ;
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  assign n350 = n346 | n349 ;
  buffer buf_n351( .i (n350), .o (n351) );
  assign n352 = n343 | n351 ;
  buffer buf_n353( .i (n352), .o (n353) );
  assign n354 = n335 | n353 ;
  assign n355 = n317 | n354 ;
  buffer buf_n356( .i (n355), .o (n356) );
  assign n357 = n234 & n356 ;
  buffer buf_n358( .i (n357), .o (n358) );
  assign n359 = n140 | n168 ;
  buffer buf_n360( .i (n359), .o (n360) );
  assign n361 = n180 | n190 ;
  buffer buf_n362( .i (n361), .o (n362) );
  assign n363 = n360 & n362 ;
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  assign n366 = n216 | n219 ;
  buffer buf_n367( .i (n366), .o (n367) );
  assign n368 = n224 | n227 ;
  buffer buf_n369( .i (n368), .o (n369) );
  assign n370 = n367 & n369 ;
  buffer buf_n371( .i (n370), .o (n371) );
  assign n372 = n198 | n201 ;
  buffer buf_n373( .i (n372), .o (n373) );
  assign n374 = n206 | n209 ;
  buffer buf_n375( .i (n374), .o (n375) );
  assign n376 = n373 & n375 ;
  buffer buf_n377( .i (n376), .o (n377) );
  assign n378 = n371 & n377 ;
  assign n379 = n365 & n378 ;
  buffer buf_n380( .i (n379), .o (n380) );
  assign n381 = n262 & n290 ;
  buffer buf_n382( .i (n381), .o (n382) );
  assign n383 = n302 & n312 ;
  buffer buf_n384( .i (n383), .o (n384) );
  assign n385 = n382 | n384 ;
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  assign n388 = n320 & n323 ;
  buffer buf_n389( .i (n388), .o (n389) );
  assign n390 = n328 & n331 ;
  buffer buf_n391( .i (n390), .o (n391) );
  assign n392 = n389 | n391 ;
  buffer buf_n393( .i (n392), .o (n393) );
  assign n394 = n338 & n341 ;
  buffer buf_n395( .i (n394), .o (n395) );
  assign n396 = n346 & n349 ;
  buffer buf_n397( .i (n396), .o (n397) );
  assign n398 = n395 | n397 ;
  buffer buf_n399( .i (n398), .o (n399) );
  assign n400 = n393 | n399 ;
  assign n401 = n387 | n400 ;
  buffer buf_n402( .i (n401), .o (n402) );
  assign n403 = n380 & n402 ;
  buffer buf_n404( .i (n403), .o (n404) );
  assign n405 = n358 & n404 ;
  buffer buf_n406( .i (n405), .o (n406) );
  assign n407 = n170 | n192 ;
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  assign n410 = n203 | n211 ;
  buffer buf_n411( .i (n410), .o (n411) );
  assign n412 = n221 | n229 ;
  buffer buf_n413( .i (n412), .o (n413) );
  assign n414 = n411 & n413 ;
  assign n415 = n409 & n414 ;
  buffer buf_n416( .i (n415), .o (n416) );
  assign n417 = n292 & n314 ;
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  assign n420 = n325 & n333 ;
  buffer buf_n421( .i (n420), .o (n421) );
  assign n422 = n343 & n351 ;
  buffer buf_n423( .i (n422), .o (n423) );
  assign n424 = n421 | n423 ;
  assign n425 = n419 | n424 ;
  buffer buf_n426( .i (n425), .o (n426) );
  assign n427 = n416 & n426 ;
  buffer buf_n428( .i (n427), .o (n428) );
  assign n429 = n360 | n362 ;
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  assign n432 = n367 | n369 ;
  buffer buf_n433( .i (n432), .o (n433) );
  assign n434 = n373 | n375 ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n436 = n433 & n435 ;
  assign n437 = n431 & n436 ;
  buffer buf_n438( .i (n437), .o (n438) );
  assign n439 = n382 & n384 ;
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  assign n442 = n389 & n391 ;
  buffer buf_n443( .i (n442), .o (n443) );
  assign n444 = n395 & n397 ;
  buffer buf_n445( .i (n444), .o (n445) );
  assign n446 = n443 | n445 ;
  assign n447 = n441 | n446 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = n438 & n448 ;
  buffer buf_n450( .i (n449), .o (n450) );
  assign n451 = n428 & n450 ;
  buffer buf_n452( .i (n451), .o (n452) );
  assign n453 = n406 & n452 ;
  buffer buf_n454( .i (n453), .o (n454) );
  assign n455 = ( n194 & n213 ) | ( n194 & n231 ) | ( n213 & n231 ) ;
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  assign n458 = ( n316 & n335 ) | ( n316 & n353 ) | ( n335 & n353 ) ;
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  assign n461 = n457 & n460 ;
  buffer buf_n462( .i (n461), .o (n462) );
  assign n463 = ( n364 & n371 ) | ( n364 & n377 ) | ( n371 & n377 ) ;
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  assign n466 = ( n386 & n393 ) | ( n386 & n399 ) | ( n393 & n399 ) ;
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  assign n469 = n465 & n468 ;
  buffer buf_n470( .i (n469), .o (n470) );
  assign n471 = n462 & n470 ;
  buffer buf_n472( .i (n471), .o (n472) );
  assign n473 = ( n408 & n411 ) | ( n408 & n413 ) | ( n411 & n413 ) ;
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  assign n476 = ( n418 & n421 ) | ( n418 & n423 ) | ( n421 & n423 ) ;
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  assign n479 = n475 & n478 ;
  buffer buf_n480( .i (n479), .o (n480) );
  assign n481 = ( n430 & n433 ) | ( n430 & n435 ) | ( n433 & n435 ) ;
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  assign n484 = ( n440 & n443 ) | ( n440 & n445 ) | ( n443 & n445 ) ;
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  assign n487 = n483 & n486 ;
  buffer buf_n488( .i (n487), .o (n488) );
  assign n489 = n480 & n488 ;
  buffer buf_n490( .i (n489), .o (n490) );
  assign n491 = n472 & n490 ;
  buffer buf_n492( .i (n491), .o (n492) );
  assign n493 = n454 & n492 ;
  assign n494 = n213 | n231 ;
  assign n495 = n195 | n494 ;
  buffer buf_n496( .i (n495), .o (n496) );
  assign n497 = n335 & n353 ;
  assign n498 = n317 & n497 ;
  buffer buf_n499( .i (n498), .o (n499) );
  assign n500 = n496 & n499 ;
  buffer buf_n501( .i (n500), .o (n501) );
  assign n502 = n371 | n377 ;
  assign n503 = n365 | n502 ;
  buffer buf_n504( .i (n503), .o (n504) );
  assign n505 = n393 & n399 ;
  assign n506 = n387 & n505 ;
  buffer buf_n507( .i (n506), .o (n507) );
  assign n508 = n504 & n507 ;
  buffer buf_n509( .i (n508), .o (n509) );
  assign n510 = n501 & n509 ;
  buffer buf_n511( .i (n510), .o (n511) );
  assign n512 = n411 | n413 ;
  assign n513 = n409 | n512 ;
  buffer buf_n514( .i (n513), .o (n514) );
  assign n515 = n421 & n423 ;
  assign n516 = n419 & n515 ;
  buffer buf_n517( .i (n516), .o (n517) );
  assign n518 = n514 & n517 ;
  buffer buf_n519( .i (n518), .o (n519) );
  assign n520 = n433 | n435 ;
  assign n521 = n431 | n520 ;
  buffer buf_n522( .i (n521), .o (n522) );
  assign n523 = n443 & n445 ;
  assign n524 = n441 & n523 ;
  buffer buf_n525( .i (n524), .o (n525) );
  assign n526 = n522 & n525 ;
  buffer buf_n527( .i (n526), .o (n527) );
  assign n528 = n519 & n527 ;
  buffer buf_n529( .i (n528), .o (n529) );
  assign n530 = n511 & n529 ;
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  assign n533 = n493 & n532 ;
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n31( .i (x13), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n21( .i (x9), .o (n21) );
  buffer buf_n91( .i (x39), .o (n91) );
  assign n535 = n21 & n91 ;
  assign n536 = n32 & n535 ;
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n26( .i (x11), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n15( .i (x6), .o (n15) );
  buffer buf_n47( .i (x20), .o (n47) );
  assign n538 = n15 | n47 ;
  assign n539 = n27 | n538 ;
  buffer buf_n540( .i (n539), .o (n540) );
  assign n541 = n537 & n540 ;
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  assign n544 = n21 | n91 ;
  assign n545 = n32 | n544 ;
  buffer buf_n546( .i (n545), .o (n546) );
  assign n547 = n15 & n47 ;
  assign n548 = n27 & n547 ;
  buffer buf_n549( .i (n548), .o (n549) );
  assign n550 = n546 & n549 ;
  buffer buf_n551( .i (n550), .o (n551) );
  assign n552 = ( n21 & n31 ) | ( n21 & n91 ) | ( n31 & n91 ) ;
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  assign n555 = ( n15 & n26 ) | ( n15 & n47 ) | ( n26 & n47 ) ;
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  assign n558 = n554 & n557 ;
  buffer buf_n559( .i (n558), .o (n559) );
  assign n560 = n551 & n559 ;
  assign n561 = n543 & n560 ;
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n82( .i (x35), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n4( .i (x1), .o (n4) );
  buffer buf_n36( .i (x15), .o (n36) );
  assign n563 = n4 & n36 ;
  assign n564 = n83 & n563 ;
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n23( .i (x10), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n102( .i (x43), .o (n102) );
  buffer buf_n107( .i (x45), .o (n107) );
  assign n566 = n102 | n107 ;
  assign n567 = n24 | n566 ;
  buffer buf_n568( .i (n567), .o (n568) );
  assign n569 = n565 | n568 ;
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  assign n572 = n4 | n36 ;
  assign n573 = n83 | n572 ;
  buffer buf_n574( .i (n573), .o (n574) );
  assign n575 = n102 & n107 ;
  assign n576 = n24 & n575 ;
  buffer buf_n577( .i (n576), .o (n577) );
  assign n578 = n574 | n577 ;
  buffer buf_n579( .i (n578), .o (n579) );
  assign n580 = ( n4 & n36 ) | ( n4 & n82 ) | ( n36 & n82 ) ;
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  assign n583 = ( n23 & n102 ) | ( n23 & n107 ) | ( n102 & n107 ) ;
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  assign n586 = n582 | n585 ;
  buffer buf_n587( .i (n586), .o (n587) );
  assign n588 = n579 | n587 ;
  assign n589 = n571 | n588 ;
  buffer buf_n590( .i (n589), .o (n590) );
  assign n591 = n562 & n590 ;
  buffer buf_n592( .i (n591), .o (n592) );
  assign n593 = n537 | n540 ;
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  assign n596 = n546 | n549 ;
  buffer buf_n597( .i (n596), .o (n597) );
  assign n598 = n554 | n557 ;
  buffer buf_n599( .i (n598), .o (n599) );
  assign n600 = n597 & n599 ;
  assign n601 = n595 & n600 ;
  buffer buf_n602( .i (n601), .o (n602) );
  assign n603 = n565 & n568 ;
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  assign n606 = n574 & n577 ;
  buffer buf_n607( .i (n606), .o (n607) );
  assign n608 = n582 & n585 ;
  buffer buf_n609( .i (n608), .o (n609) );
  assign n610 = n607 | n609 ;
  assign n611 = n605 | n610 ;
  buffer buf_n612( .i (n611), .o (n612) );
  assign n613 = n602 & n612 ;
  buffer buf_n614( .i (n613), .o (n614) );
  assign n615 = n592 & n614 ;
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  assign n618 = n551 | n559 ;
  assign n619 = n543 | n618 ;
  buffer buf_n620( .i (n619), .o (n620) );
  assign n621 = n579 & n587 ;
  assign n622 = n571 & n621 ;
  buffer buf_n623( .i (n622), .o (n623) );
  assign n624 = n620 & n623 ;
  buffer buf_n625( .i (n624), .o (n625) );
  assign n626 = n597 | n599 ;
  assign n627 = n595 | n626 ;
  buffer buf_n628( .i (n627), .o (n628) );
  assign n629 = n607 & n609 ;
  assign n630 = n605 & n629 ;
  buffer buf_n631( .i (n630), .o (n631) );
  assign n632 = n628 & n631 ;
  buffer buf_n633( .i (n632), .o (n633) );
  assign n634 = n625 & n633 ;
  buffer buf_n635( .i (n634), .o (n635) );
  assign n636 = ( n542 & n551 ) | ( n542 & n559 ) | ( n551 & n559 ) ;
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  assign n639 = ( n570 & n579 ) | ( n570 & n587 ) | ( n579 & n587 ) ;
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  assign n642 = n638 & n641 ;
  buffer buf_n643( .i (n642), .o (n643) );
  assign n644 = ( n594 & n597 ) | ( n594 & n599 ) | ( n597 & n599 ) ;
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  assign n647 = ( n604 & n607 ) | ( n604 & n609 ) | ( n607 & n609 ) ;
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  assign n650 = n646 & n649 ;
  buffer buf_n651( .i (n650), .o (n651) );
  assign n652 = n643 & n651 ;
  buffer buf_n653( .i (n652), .o (n653) );
  assign n654 = n635 & n653 ;
  assign n655 = n617 & n654 ;
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n72( .i (x31), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n77( .i (x33), .o (n77) );
  buffer buf_n112( .i (x47), .o (n112) );
  assign n657 = n77 & n112 ;
  assign n658 = n73 & n657 ;
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n67( .i (x29), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n10( .i (x4), .o (n10) );
  buffer buf_n45( .i (x19), .o (n45) );
  assign n660 = n10 | n45 ;
  assign n661 = n68 | n660 ;
  buffer buf_n662( .i (n661), .o (n662) );
  assign n663 = n659 | n662 ;
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  assign n666 = n77 | n112 ;
  assign n667 = n73 | n666 ;
  buffer buf_n668( .i (n667), .o (n668) );
  assign n669 = n10 & n45 ;
  assign n670 = n68 & n669 ;
  buffer buf_n671( .i (n670), .o (n671) );
  assign n672 = n668 | n671 ;
  buffer buf_n673( .i (n672), .o (n673) );
  assign n674 = ( n72 & n77 ) | ( n72 & n112 ) | ( n77 & n112 ) ;
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  assign n677 = ( n10 & n45 ) | ( n10 & n67 ) | ( n45 & n67 ) ;
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  assign n680 = n676 | n679 ;
  buffer buf_n681( .i (n680), .o (n681) );
  assign n682 = n673 & n681 ;
  assign n683 = n665 & n682 ;
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n104( .i (x44), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n29( .i (x12), .o (n29) );
  buffer buf_n63( .i (x27), .o (n63) );
  assign n685 = n29 & n63 ;
  assign n686 = n105 & n685 ;
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n93( .i (x40), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n49( .i (x21), .o (n49) );
  buffer buf_n59( .i (x25), .o (n59) );
  assign n688 = n49 | n59 ;
  assign n689 = n94 | n688 ;
  buffer buf_n690( .i (n689), .o (n690) );
  assign n691 = n687 & n690 ;
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  assign n694 = n29 | n63 ;
  assign n695 = n105 | n694 ;
  buffer buf_n696( .i (n695), .o (n696) );
  assign n697 = n49 & n59 ;
  assign n698 = n94 & n697 ;
  buffer buf_n699( .i (n698), .o (n699) );
  assign n700 = n696 & n699 ;
  buffer buf_n701( .i (n700), .o (n701) );
  assign n702 = ( n29 & n63 ) | ( n29 & n104 ) | ( n63 & n104 ) ;
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  assign n705 = ( n49 & n59 ) | ( n49 & n93 ) | ( n59 & n93 ) ;
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  assign n708 = n704 & n707 ;
  buffer buf_n709( .i (n708), .o (n709) );
  assign n710 = n701 | n709 ;
  assign n711 = n693 | n710 ;
  buffer buf_n712( .i (n711), .o (n712) );
  assign n713 = n684 | n712 ;
  buffer buf_n714( .i (n713), .o (n714) );
  assign n715 = n659 & n662 ;
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  assign n718 = n668 & n671 ;
  buffer buf_n719( .i (n718), .o (n719) );
  assign n720 = n676 & n679 ;
  buffer buf_n721( .i (n720), .o (n721) );
  assign n722 = n719 & n721 ;
  assign n723 = n717 & n722 ;
  buffer buf_n724( .i (n723), .o (n724) );
  assign n725 = n696 | n699 ;
  buffer buf_n726( .i (n725), .o (n726) );
  assign n727 = n704 | n707 ;
  buffer buf_n728( .i (n727), .o (n728) );
  assign n729 = n726 | n728 ;
  assign n730 = n687 | n690 ;
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  assign n733 = n729 | n732 ;
  buffer buf_n734( .i (n733), .o (n734) );
  assign n735 = n724 | n734 ;
  buffer buf_n736( .i (n735), .o (n736) );
  assign n737 = n714 | n736 ;
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  assign n740 = n673 | n681 ;
  assign n741 = n665 | n740 ;
  buffer buf_n742( .i (n741), .o (n742) );
  assign n743 = n701 & n709 ;
  assign n744 = n693 & n743 ;
  buffer buf_n745( .i (n744), .o (n745) );
  assign n746 = n742 | n745 ;
  buffer buf_n747( .i (n746), .o (n747) );
  assign n748 = n719 | n721 ;
  assign n749 = n717 | n748 ;
  buffer buf_n750( .i (n749), .o (n750) );
  assign n751 = n726 & n728 ;
  assign n752 = n732 & n751 ;
  buffer buf_n753( .i (n752), .o (n753) );
  assign n754 = n750 | n753 ;
  buffer buf_n755( .i (n754), .o (n755) );
  assign n756 = n747 | n755 ;
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = ( n664 & n673 ) | ( n664 & n681 ) | ( n673 & n681 ) ;
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  assign n761 = ( n692 & n701 ) | ( n692 & n709 ) | ( n701 & n709 ) ;
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  assign n764 = n760 | n763 ;
  buffer buf_n765( .i (n764), .o (n765) );
  assign n766 = ( n716 & n719 ) | ( n716 & n721 ) | ( n719 & n721 ) ;
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  assign n769 = ( n726 & n728 ) | ( n726 & n731 ) | ( n728 & n731 ) ;
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  assign n772 = n768 | n771 ;
  buffer buf_n773( .i (n772), .o (n773) );
  assign n774 = n765 | n773 ;
  buffer buf_n775( .i (n774), .o (n775) );
  assign n776 = n757 | n775 ;
  assign n777 = n739 | n776 ;
  buffer buf_n778( .i (n777), .o (n778) );
  assign n779 = n656 | n778 ;
  buffer buf_n780( .i (n779), .o (n780) );
  assign n781 = n562 | n590 ;
  buffer buf_n782( .i (n781), .o (n782) );
  assign n783 = n602 | n612 ;
  buffer buf_n784( .i (n783), .o (n784) );
  assign n785 = n782 & n784 ;
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  assign n788 = n638 | n641 ;
  buffer buf_n789( .i (n788), .o (n789) );
  assign n790 = n646 | n649 ;
  buffer buf_n791( .i (n790), .o (n791) );
  assign n792 = n789 & n791 ;
  buffer buf_n793( .i (n792), .o (n793) );
  assign n794 = n620 | n623 ;
  buffer buf_n795( .i (n794), .o (n795) );
  assign n796 = n628 | n631 ;
  buffer buf_n797( .i (n796), .o (n797) );
  assign n798 = n795 & n797 ;
  buffer buf_n799( .i (n798), .o (n799) );
  assign n800 = n793 & n799 ;
  assign n801 = n787 & n800 ;
  buffer buf_n802( .i (n801), .o (n802) );
  assign n803 = n684 & n712 ;
  buffer buf_n804( .i (n803), .o (n804) );
  assign n805 = n724 & n734 ;
  buffer buf_n806( .i (n805), .o (n806) );
  assign n807 = n804 | n806 ;
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  assign n810 = n742 & n745 ;
  buffer buf_n811( .i (n810), .o (n811) );
  assign n812 = n750 & n753 ;
  buffer buf_n813( .i (n812), .o (n813) );
  assign n814 = n811 | n813 ;
  buffer buf_n815( .i (n814), .o (n815) );
  assign n816 = n760 & n763 ;
  buffer buf_n817( .i (n816), .o (n817) );
  assign n818 = n768 & n771 ;
  buffer buf_n819( .i (n818), .o (n819) );
  assign n820 = n817 | n819 ;
  buffer buf_n821( .i (n820), .o (n821) );
  assign n822 = n815 | n821 ;
  assign n823 = n809 | n822 ;
  buffer buf_n824( .i (n823), .o (n824) );
  assign n825 = n802 | n824 ;
  buffer buf_n826( .i (n825), .o (n826) );
  assign n827 = n780 | n826 ;
  buffer buf_n828( .i (n827), .o (n828) );
  assign n829 = n625 | n633 ;
  buffer buf_n830( .i (n829), .o (n830) );
  assign n831 = n643 | n651 ;
  buffer buf_n832( .i (n831), .o (n832) );
  assign n833 = n830 & n832 ;
  assign n834 = n592 | n614 ;
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  assign n837 = n833 & n836 ;
  buffer buf_n838( .i (n837), .o (n838) );
  assign n839 = n714 & n736 ;
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  assign n842 = n747 & n755 ;
  buffer buf_n843( .i (n842), .o (n843) );
  assign n844 = n765 & n773 ;
  buffer buf_n845( .i (n844), .o (n845) );
  assign n846 = n843 | n845 ;
  assign n847 = n841 | n846 ;
  buffer buf_n848( .i (n847), .o (n848) );
  assign n849 = n838 | n848 ;
  buffer buf_n850( .i (n849), .o (n850) );
  assign n851 = n782 | n784 ;
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  assign n854 = n789 | n791 ;
  buffer buf_n855( .i (n854), .o (n855) );
  assign n856 = n795 | n797 ;
  buffer buf_n857( .i (n856), .o (n857) );
  assign n858 = n855 & n857 ;
  assign n859 = n853 & n858 ;
  buffer buf_n860( .i (n859), .o (n860) );
  assign n861 = n804 & n806 ;
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  assign n864 = n811 & n813 ;
  buffer buf_n865( .i (n864), .o (n865) );
  assign n866 = n817 & n819 ;
  buffer buf_n867( .i (n866), .o (n867) );
  assign n868 = n865 | n867 ;
  assign n869 = n863 | n868 ;
  buffer buf_n870( .i (n869), .o (n870) );
  assign n871 = n860 | n870 ;
  buffer buf_n872( .i (n871), .o (n872) );
  assign n873 = n850 | n872 ;
  buffer buf_n874( .i (n873), .o (n874) );
  assign n875 = n828 | n874 ;
  buffer buf_n876( .i (n875), .o (n876) );
  assign n877 = ( n616 & n635 ) | ( n616 & n653 ) | ( n635 & n653 ) ;
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  assign n880 = ( n738 & n757 ) | ( n738 & n775 ) | ( n757 & n775 ) ;
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  assign n883 = n879 | n882 ;
  buffer buf_n884( .i (n883), .o (n884) );
  assign n885 = ( n786 & n793 ) | ( n786 & n799 ) | ( n793 & n799 ) ;
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  assign n888 = ( n808 & n815 ) | ( n808 & n821 ) | ( n815 & n821 ) ;
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  assign n891 = n887 | n890 ;
  buffer buf_n892( .i (n891), .o (n892) );
  assign n893 = n884 | n892 ;
  buffer buf_n894( .i (n893), .o (n894) );
  assign n895 = ( n830 & n832 ) | ( n830 & n835 ) | ( n832 & n835 ) ;
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  assign n898 = ( n840 & n843 ) | ( n840 & n845 ) | ( n843 & n845 ) ;
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  assign n901 = n897 | n900 ;
  buffer buf_n902( .i (n901), .o (n902) );
  assign n903 = ( n852 & n855 ) | ( n852 & n857 ) | ( n855 & n857 ) ;
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  assign n906 = ( n862 & n865 ) | ( n862 & n867 ) | ( n865 & n867 ) ;
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  assign n909 = n905 | n908 ;
  buffer buf_n910( .i (n909), .o (n910) );
  assign n911 = n902 | n910 ;
  buffer buf_n912( .i (n911), .o (n912) );
  assign n913 = n894 | n912 ;
  buffer buf_n914( .i (n913), .o (n914) );
  assign n915 = n876 | n914 ;
  assign n916 = n635 | n653 ;
  assign n917 = n617 | n916 ;
  buffer buf_n918( .i (n917), .o (n918) );
  assign n919 = n757 & n775 ;
  assign n920 = n739 & n919 ;
  buffer buf_n921( .i (n920), .o (n921) );
  assign n922 = n918 | n921 ;
  buffer buf_n923( .i (n922), .o (n923) );
  assign n924 = n793 | n799 ;
  assign n925 = n787 | n924 ;
  buffer buf_n926( .i (n925), .o (n926) );
  assign n927 = n815 & n821 ;
  assign n928 = n809 & n927 ;
  buffer buf_n929( .i (n928), .o (n929) );
  assign n930 = n926 | n929 ;
  buffer buf_n931( .i (n930), .o (n931) );
  assign n932 = n923 | n931 ;
  buffer buf_n933( .i (n932), .o (n933) );
  assign n934 = n830 | n832 ;
  assign n935 = n836 | n934 ;
  buffer buf_n936( .i (n935), .o (n936) );
  assign n937 = n843 & n845 ;
  assign n938 = n841 & n937 ;
  buffer buf_n939( .i (n938), .o (n939) );
  assign n940 = n936 | n939 ;
  buffer buf_n941( .i (n940), .o (n941) );
  assign n942 = n855 | n857 ;
  assign n943 = n853 | n942 ;
  buffer buf_n944( .i (n943), .o (n944) );
  assign n945 = n865 & n867 ;
  assign n946 = n863 & n945 ;
  buffer buf_n947( .i (n946), .o (n947) );
  assign n948 = n944 | n947 ;
  buffer buf_n949( .i (n948), .o (n949) );
  assign n950 = n941 | n949 ;
  buffer buf_n951( .i (n950), .o (n951) );
  assign n952 = n933 | n951 ;
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  assign n955 = n915 | n954 ;
  buffer buf_n956( .i (n955), .o (n956) );
  assign n957 = n534 | n956 ;
  buffer buf_n958( .i (n957), .o (n958) );
  assign n959 = n234 | n356 ;
  buffer buf_n960( .i (n959), .o (n960) );
  assign n961 = n380 | n402 ;
  buffer buf_n962( .i (n961), .o (n962) );
  assign n963 = n960 & n962 ;
  buffer buf_n964( .i (n963), .o (n964) );
  assign n965 = n416 | n426 ;
  buffer buf_n966( .i (n965), .o (n966) );
  assign n967 = n438 | n448 ;
  buffer buf_n968( .i (n967), .o (n968) );
  assign n969 = n966 & n968 ;
  buffer buf_n970( .i (n969), .o (n970) );
  assign n971 = n964 & n970 ;
  buffer buf_n972( .i (n971), .o (n972) );
  assign n973 = n457 | n460 ;
  buffer buf_n974( .i (n973), .o (n974) );
  assign n975 = n465 | n468 ;
  buffer buf_n976( .i (n975), .o (n976) );
  assign n977 = n974 & n976 ;
  buffer buf_n978( .i (n977), .o (n978) );
  assign n979 = n475 | n478 ;
  buffer buf_n980( .i (n979), .o (n980) );
  assign n981 = n483 | n486 ;
  buffer buf_n982( .i (n981), .o (n982) );
  assign n983 = n980 & n982 ;
  buffer buf_n984( .i (n983), .o (n984) );
  assign n985 = n978 & n984 ;
  buffer buf_n986( .i (n985), .o (n986) );
  assign n987 = n972 & n986 ;
  assign n988 = n496 | n499 ;
  buffer buf_n989( .i (n988), .o (n989) );
  assign n990 = n504 | n507 ;
  buffer buf_n991( .i (n990), .o (n991) );
  assign n992 = n989 & n991 ;
  buffer buf_n993( .i (n992), .o (n993) );
  assign n994 = n514 | n517 ;
  buffer buf_n995( .i (n994), .o (n995) );
  assign n996 = n522 | n525 ;
  buffer buf_n997( .i (n996), .o (n997) );
  assign n998 = n995 & n997 ;
  buffer buf_n999( .i (n998), .o (n999) );
  assign n1000 = n993 & n999 ;
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  assign n1003 = n987 & n1002 ;
  buffer buf_n1004( .i (n1003), .o (n1004) );
  assign n1005 = n656 & n778 ;
  buffer buf_n1006( .i (n1005), .o (n1006) );
  assign n1007 = n802 & n824 ;
  buffer buf_n1008( .i (n1007), .o (n1008) );
  assign n1009 = n1006 | n1008 ;
  buffer buf_n1010( .i (n1009), .o (n1010) );
  assign n1011 = n838 & n848 ;
  buffer buf_n1012( .i (n1011), .o (n1012) );
  assign n1013 = n860 & n870 ;
  buffer buf_n1014( .i (n1013), .o (n1014) );
  assign n1015 = n1012 | n1014 ;
  buffer buf_n1016( .i (n1015), .o (n1016) );
  assign n1017 = n1010 | n1016 ;
  buffer buf_n1018( .i (n1017), .o (n1018) );
  assign n1019 = n879 & n882 ;
  buffer buf_n1020( .i (n1019), .o (n1020) );
  assign n1021 = n887 & n890 ;
  buffer buf_n1022( .i (n1021), .o (n1022) );
  assign n1023 = n1020 | n1022 ;
  buffer buf_n1024( .i (n1023), .o (n1024) );
  assign n1025 = n897 & n900 ;
  buffer buf_n1026( .i (n1025), .o (n1026) );
  assign n1027 = n905 & n908 ;
  buffer buf_n1028( .i (n1027), .o (n1028) );
  assign n1029 = n1026 | n1028 ;
  buffer buf_n1030( .i (n1029), .o (n1030) );
  assign n1031 = n1024 | n1030 ;
  buffer buf_n1032( .i (n1031), .o (n1032) );
  assign n1033 = n1018 | n1032 ;
  assign n1034 = n918 & n921 ;
  buffer buf_n1035( .i (n1034), .o (n1035) );
  assign n1036 = n926 & n929 ;
  buffer buf_n1037( .i (n1036), .o (n1037) );
  assign n1038 = n1035 | n1037 ;
  buffer buf_n1039( .i (n1038), .o (n1039) );
  assign n1040 = n936 & n939 ;
  buffer buf_n1041( .i (n1040), .o (n1041) );
  assign n1042 = n944 & n947 ;
  buffer buf_n1043( .i (n1042), .o (n1043) );
  assign n1044 = n1041 | n1043 ;
  buffer buf_n1045( .i (n1044), .o (n1045) );
  assign n1046 = n1039 | n1045 ;
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  assign n1049 = n1033 | n1048 ;
  buffer buf_n1050( .i (n1049), .o (n1050) );
  assign n1051 = n1004 | n1050 ;
  buffer buf_n1052( .i (n1051), .o (n1052) );
  assign n1053 = n958 | n1052 ;
  buffer buf_n1054( .i (n1053), .o (n1054) );
  assign n1055 = n358 | n404 ;
  buffer buf_n1056( .i (n1055), .o (n1056) );
  assign n1057 = n428 | n450 ;
  buffer buf_n1058( .i (n1057), .o (n1058) );
  assign n1059 = n1056 & n1058 ;
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1061 = n462 | n470 ;
  buffer buf_n1062( .i (n1061), .o (n1062) );
  assign n1063 = n480 | n488 ;
  buffer buf_n1064( .i (n1063), .o (n1064) );
  assign n1065 = n1062 & n1064 ;
  buffer buf_n1066( .i (n1065), .o (n1066) );
  assign n1067 = n1060 & n1066 ;
  assign n1068 = n501 | n509 ;
  buffer buf_n1069( .i (n1068), .o (n1069) );
  assign n1070 = n519 | n527 ;
  buffer buf_n1071( .i (n1070), .o (n1071) );
  assign n1072 = n1069 & n1071 ;
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  assign n1075 = n1067 & n1074 ;
  buffer buf_n1076( .i (n1075), .o (n1076) );
  assign n1077 = n780 & n826 ;
  buffer buf_n1078( .i (n1077), .o (n1078) );
  assign n1079 = n850 & n872 ;
  buffer buf_n1080( .i (n1079), .o (n1080) );
  assign n1081 = n1078 | n1080 ;
  buffer buf_n1082( .i (n1081), .o (n1082) );
  assign n1083 = n884 & n892 ;
  buffer buf_n1084( .i (n1083), .o (n1084) );
  assign n1085 = n902 & n910 ;
  buffer buf_n1086( .i (n1085), .o (n1086) );
  assign n1087 = n1084 | n1086 ;
  buffer buf_n1088( .i (n1087), .o (n1088) );
  assign n1089 = n1082 | n1088 ;
  assign n1090 = n923 & n931 ;
  buffer buf_n1091( .i (n1090), .o (n1091) );
  assign n1092 = n941 & n949 ;
  buffer buf_n1093( .i (n1092), .o (n1093) );
  assign n1094 = n1091 | n1093 ;
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  assign n1097 = n1089 | n1096 ;
  buffer buf_n1098( .i (n1097), .o (n1098) );
  assign n1099 = n1076 | n1098 ;
  buffer buf_n1100( .i (n1099), .o (n1100) );
  assign n1101 = n960 | n962 ;
  buffer buf_n1102( .i (n1101), .o (n1102) );
  assign n1103 = n966 | n968 ;
  buffer buf_n1104( .i (n1103), .o (n1104) );
  assign n1105 = n1102 & n1104 ;
  buffer buf_n1106( .i (n1105), .o (n1106) );
  assign n1107 = n974 | n976 ;
  buffer buf_n1108( .i (n1107), .o (n1108) );
  assign n1109 = n980 | n982 ;
  buffer buf_n1110( .i (n1109), .o (n1110) );
  assign n1111 = n1108 & n1110 ;
  buffer buf_n1112( .i (n1111), .o (n1112) );
  assign n1113 = n1106 & n1112 ;
  assign n1114 = n989 | n991 ;
  buffer buf_n1115( .i (n1114), .o (n1115) );
  assign n1116 = n995 | n997 ;
  buffer buf_n1117( .i (n1116), .o (n1117) );
  assign n1118 = n1115 & n1117 ;
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  assign n1121 = n1113 & n1120 ;
  buffer buf_n1122( .i (n1121), .o (n1122) );
  assign n1123 = n1006 & n1008 ;
  buffer buf_n1124( .i (n1123), .o (n1124) );
  assign n1125 = n1012 & n1014 ;
  buffer buf_n1126( .i (n1125), .o (n1126) );
  assign n1127 = n1124 | n1126 ;
  buffer buf_n1128( .i (n1127), .o (n1128) );
  assign n1129 = n1020 & n1022 ;
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n1131 = n1026 & n1028 ;
  buffer buf_n1132( .i (n1131), .o (n1132) );
  assign n1133 = n1130 | n1132 ;
  buffer buf_n1134( .i (n1133), .o (n1134) );
  assign n1135 = n1128 | n1134 ;
  assign n1136 = n1035 & n1037 ;
  buffer buf_n1137( .i (n1136), .o (n1137) );
  assign n1138 = n1041 & n1043 ;
  buffer buf_n1139( .i (n1138), .o (n1139) );
  assign n1140 = n1137 | n1139 ;
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  assign n1143 = n1135 | n1142 ;
  buffer buf_n1144( .i (n1143), .o (n1144) );
  assign n1145 = n1122 | n1144 ;
  buffer buf_n1146( .i (n1145), .o (n1146) );
  assign n1147 = n1100 | n1146 ;
  buffer buf_n1148( .i (n1147), .o (n1148) );
  assign n1149 = n1054 | n1148 ;
  buffer buf_n1150( .i (n1149), .o (n1150) );
  assign n1151 = n406 | n452 ;
  buffer buf_n1152( .i (n1151), .o (n1152) );
  assign n1153 = n472 | n490 ;
  buffer buf_n1154( .i (n1153), .o (n1154) );
  assign n1155 = n1152 & n1154 ;
  assign n1156 = n511 | n529 ;
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  assign n1159 = n1155 & n1158 ;
  buffer buf_n1160( .i (n1159), .o (n1160) );
  assign n1161 = n828 & n874 ;
  buffer buf_n1162( .i (n1161), .o (n1162) );
  assign n1163 = n894 & n912 ;
  buffer buf_n1164( .i (n1163), .o (n1164) );
  assign n1165 = n1162 | n1164 ;
  assign n1166 = n933 & n951 ;
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  assign n1169 = n1165 | n1168 ;
  buffer buf_n1170( .i (n1169), .o (n1170) );
  assign n1171 = n1160 | n1170 ;
  buffer buf_n1172( .i (n1171), .o (n1172) );
  assign n1173 = n964 | n970 ;
  buffer buf_n1174( .i (n1173), .o (n1174) );
  assign n1175 = n978 | n984 ;
  buffer buf_n1176( .i (n1175), .o (n1176) );
  assign n1177 = n1174 & n1176 ;
  assign n1178 = n993 | n999 ;
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  assign n1181 = n1177 & n1180 ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  assign n1183 = n1010 & n1016 ;
  buffer buf_n1184( .i (n1183), .o (n1184) );
  assign n1185 = n1024 & n1030 ;
  buffer buf_n1186( .i (n1185), .o (n1186) );
  assign n1187 = n1184 | n1186 ;
  assign n1188 = n1039 & n1045 ;
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  assign n1191 = n1187 | n1190 ;
  buffer buf_n1192( .i (n1191), .o (n1192) );
  assign n1193 = n1182 | n1192 ;
  buffer buf_n1194( .i (n1193), .o (n1194) );
  assign n1195 = n1172 | n1194 ;
  buffer buf_n1196( .i (n1195), .o (n1196) );
  assign n1197 = n1056 | n1058 ;
  buffer buf_n1198( .i (n1197), .o (n1198) );
  assign n1199 = n1062 | n1064 ;
  buffer buf_n1200( .i (n1199), .o (n1200) );
  assign n1201 = n1198 & n1200 ;
  assign n1202 = n1069 | n1071 ;
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  assign n1205 = n1201 & n1204 ;
  buffer buf_n1206( .i (n1205), .o (n1206) );
  assign n1207 = n1078 & n1080 ;
  buffer buf_n1208( .i (n1207), .o (n1208) );
  assign n1209 = n1084 & n1086 ;
  buffer buf_n1210( .i (n1209), .o (n1210) );
  assign n1211 = n1208 | n1210 ;
  assign n1212 = n1091 & n1093 ;
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  assign n1215 = n1211 | n1214 ;
  buffer buf_n1216( .i (n1215), .o (n1216) );
  assign n1217 = n1206 | n1216 ;
  buffer buf_n1218( .i (n1217), .o (n1218) );
  assign n1219 = n1102 | n1104 ;
  buffer buf_n1220( .i (n1219), .o (n1220) );
  assign n1221 = n1108 | n1110 ;
  buffer buf_n1222( .i (n1221), .o (n1222) );
  assign n1223 = n1220 & n1222 ;
  assign n1224 = n1115 | n1117 ;
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  assign n1227 = n1223 & n1226 ;
  buffer buf_n1228( .i (n1227), .o (n1228) );
  assign n1229 = n1124 & n1126 ;
  buffer buf_n1230( .i (n1229), .o (n1230) );
  assign n1231 = n1130 & n1132 ;
  buffer buf_n1232( .i (n1231), .o (n1232) );
  assign n1233 = n1230 | n1232 ;
  assign n1234 = n1137 & n1139 ;
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  assign n1237 = n1233 | n1236 ;
  buffer buf_n1238( .i (n1237), .o (n1238) );
  assign n1239 = n1228 | n1238 ;
  buffer buf_n1240( .i (n1239), .o (n1240) );
  assign n1241 = n1218 | n1240 ;
  buffer buf_n1242( .i (n1241), .o (n1242) );
  assign n1243 = n1196 | n1242 ;
  buffer buf_n1244( .i (n1243), .o (n1244) );
  assign n1245 = n1150 | n1244 ;
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n1247( .i (n1246), .o (n1247) );
  assign n1248 = ( n454 & n492 ) | ( n454 & n531 ) | ( n492 & n531 ) ;
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  assign n1251 = ( n876 & n914 ) | ( n876 & n953 ) | ( n914 & n953 ) ;
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  assign n1254 = n1250 | n1253 ;
  buffer buf_n1255( .i (n1254), .o (n1255) );
  assign n1256 = ( n972 & n986 ) | ( n972 & n1001 ) | ( n986 & n1001 ) ;
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  assign n1259 = ( n1018 & n1032 ) | ( n1018 & n1047 ) | ( n1032 & n1047 ) ;
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  assign n1262 = n1258 | n1261 ;
  buffer buf_n1263( .i (n1262), .o (n1263) );
  assign n1264 = n1255 | n1263 ;
  buffer buf_n1265( .i (n1264), .o (n1265) );
  assign n1266 = ( n1060 & n1066 ) | ( n1060 & n1073 ) | ( n1066 & n1073 ) ;
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  assign n1269 = ( n1082 & n1088 ) | ( n1082 & n1095 ) | ( n1088 & n1095 ) ;
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  assign n1272 = n1268 | n1271 ;
  buffer buf_n1273( .i (n1272), .o (n1273) );
  assign n1274 = ( n1106 & n1112 ) | ( n1106 & n1119 ) | ( n1112 & n1119 ) ;
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  assign n1277 = ( n1128 & n1134 ) | ( n1128 & n1141 ) | ( n1134 & n1141 ) ;
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  assign n1280 = n1276 | n1279 ;
  buffer buf_n1281( .i (n1280), .o (n1281) );
  assign n1282 = n1273 | n1281 ;
  buffer buf_n1283( .i (n1282), .o (n1283) );
  assign n1284 = n1265 | n1283 ;
  buffer buf_n1285( .i (n1284), .o (n1285) );
  assign n1286 = ( n1152 & n1154 ) | ( n1152 & n1157 ) | ( n1154 & n1157 ) ;
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  assign n1289 = ( n1162 & n1164 ) | ( n1162 & n1167 ) | ( n1164 & n1167 ) ;
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  assign n1292 = n1288 | n1291 ;
  buffer buf_n1293( .i (n1292), .o (n1293) );
  assign n1294 = ( n1174 & n1176 ) | ( n1174 & n1179 ) | ( n1176 & n1179 ) ;
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  assign n1297 = ( n1184 & n1186 ) | ( n1184 & n1189 ) | ( n1186 & n1189 ) ;
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  assign n1300 = n1296 | n1299 ;
  buffer buf_n1301( .i (n1300), .o (n1301) );
  assign n1302 = n1293 | n1301 ;
  buffer buf_n1303( .i (n1302), .o (n1303) );
  assign n1304 = ( n1198 & n1200 ) | ( n1198 & n1203 ) | ( n1200 & n1203 ) ;
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  assign n1307 = ( n1208 & n1210 ) | ( n1208 & n1213 ) | ( n1210 & n1213 ) ;
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  assign n1310 = n1306 | n1309 ;
  buffer buf_n1311( .i (n1310), .o (n1311) );
  assign n1312 = ( n1220 & n1222 ) | ( n1220 & n1225 ) | ( n1222 & n1225 ) ;
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  assign n1315 = ( n1230 & n1232 ) | ( n1230 & n1235 ) | ( n1232 & n1235 ) ;
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  assign n1318 = n1314 | n1317 ;
  buffer buf_n1319( .i (n1318), .o (n1319) );
  assign n1320 = n1311 | n1319 ;
  buffer buf_n1321( .i (n1320), .o (n1321) );
  assign n1322 = n1303 | n1321 ;
  buffer buf_n1323( .i (n1322), .o (n1323) );
  assign n1324 = n1285 | n1323 ;
  buffer buf_n1325( .i (n1324), .o (n1325) );
  assign n1326 = n454 | n492 ;
  assign n1327 = n532 | n1326 ;
  buffer buf_n1328( .i (n1327), .o (n1328) );
  assign n1329 = n876 & n914 ;
  assign n1330 = n954 & n1329 ;
  buffer buf_n1331( .i (n1330), .o (n1331) );
  assign n1332 = n1328 | n1331 ;
  buffer buf_n1333( .i (n1332), .o (n1333) );
  assign n1334 = n972 | n986 ;
  assign n1335 = n1002 | n1334 ;
  buffer buf_n1336( .i (n1335), .o (n1336) );
  assign n1337 = n1018 & n1032 ;
  assign n1338 = n1048 & n1337 ;
  buffer buf_n1339( .i (n1338), .o (n1339) );
  assign n1340 = n1336 | n1339 ;
  buffer buf_n1341( .i (n1340), .o (n1341) );
  assign n1342 = n1333 | n1341 ;
  buffer buf_n1343( .i (n1342), .o (n1343) );
  assign n1344 = n1060 | n1066 ;
  assign n1345 = n1074 | n1344 ;
  buffer buf_n1346( .i (n1345), .o (n1346) );
  assign n1347 = n1082 & n1088 ;
  assign n1348 = n1096 & n1347 ;
  buffer buf_n1349( .i (n1348), .o (n1349) );
  assign n1350 = n1346 | n1349 ;
  buffer buf_n1351( .i (n1350), .o (n1351) );
  assign n1352 = n1106 | n1112 ;
  assign n1353 = n1120 | n1352 ;
  buffer buf_n1354( .i (n1353), .o (n1354) );
  assign n1355 = n1128 & n1134 ;
  assign n1356 = n1142 & n1355 ;
  buffer buf_n1357( .i (n1356), .o (n1357) );
  assign n1358 = n1354 | n1357 ;
  buffer buf_n1359( .i (n1358), .o (n1359) );
  assign n1360 = n1351 | n1359 ;
  buffer buf_n1361( .i (n1360), .o (n1361) );
  assign n1362 = n1343 | n1361 ;
  buffer buf_n1363( .i (n1362), .o (n1363) );
  assign n1364 = n1152 | n1154 ;
  assign n1365 = n1158 | n1364 ;
  buffer buf_n1366( .i (n1365), .o (n1366) );
  assign n1367 = n1162 & n1164 ;
  assign n1368 = n1168 & n1367 ;
  buffer buf_n1369( .i (n1368), .o (n1369) );
  assign n1370 = n1366 | n1369 ;
  buffer buf_n1371( .i (n1370), .o (n1371) );
  assign n1372 = n1174 | n1176 ;
  assign n1373 = n1180 | n1372 ;
  buffer buf_n1374( .i (n1373), .o (n1374) );
  assign n1375 = n1184 & n1186 ;
  assign n1376 = n1190 & n1375 ;
  buffer buf_n1377( .i (n1376), .o (n1377) );
  assign n1378 = n1374 | n1377 ;
  buffer buf_n1379( .i (n1378), .o (n1379) );
  assign n1380 = n1371 | n1379 ;
  buffer buf_n1381( .i (n1380), .o (n1381) );
  assign n1382 = n1198 | n1200 ;
  assign n1383 = n1204 | n1382 ;
  buffer buf_n1384( .i (n1383), .o (n1384) );
  assign n1385 = n1208 & n1210 ;
  assign n1386 = n1214 & n1385 ;
  buffer buf_n1387( .i (n1386), .o (n1387) );
  assign n1388 = n1384 | n1387 ;
  buffer buf_n1389( .i (n1388), .o (n1389) );
  assign n1390 = n1220 | n1222 ;
  assign n1391 = n1226 | n1390 ;
  buffer buf_n1392( .i (n1391), .o (n1392) );
  assign n1393 = n1230 & n1232 ;
  assign n1394 = n1236 & n1393 ;
  buffer buf_n1395( .i (n1394), .o (n1395) );
  assign n1396 = n1392 | n1395 ;
  buffer buf_n1397( .i (n1396), .o (n1397) );
  assign n1398 = n1389 | n1397 ;
  buffer buf_n1399( .i (n1398), .o (n1399) );
  assign n1400 = n1381 | n1399 ;
  buffer buf_n1401( .i (n1400), .o (n1401) );
  assign n1402 = n1363 | n1401 ;
  buffer buf_n1403( .i (n1402), .o (n1403) );
  assign n1404 = n1325 | n1403 ;
  assign n1405 = n1247 | n1404 ;
  assign n1406 = n1150 & n1244 ;
  buffer buf_n1407( .i (n1406), .o (n1407) );
  assign n1409 = n1285 & n1323 ;
  buffer buf_n1410( .i (n1409), .o (n1410) );
  assign n1411 = n1363 & n1401 ;
  buffer buf_n1412( .i (n1411), .o (n1412) );
  assign n1413 = ( n1407 & n1410 ) | ( n1407 & n1412 ) | ( n1410 & n1412 ) ;
  buffer buf_n1414( .i (n1413), .o (n1414) );
  assign n1415 = n1054 & n1148 ;
  buffer buf_n1416( .i (n1415), .o (n1416) );
  assign n1417 = n1196 & n1242 ;
  buffer buf_n1418( .i (n1417), .o (n1418) );
  assign n1419 = n1416 | n1418 ;
  buffer buf_n1420( .i (n1419), .o (n1420) );
  assign n1422 = n1265 & n1283 ;
  buffer buf_n1423( .i (n1422), .o (n1423) );
  assign n1424 = n1303 & n1321 ;
  buffer buf_n1425( .i (n1424), .o (n1425) );
  assign n1426 = n1423 | n1425 ;
  buffer buf_n1427( .i (n1426), .o (n1427) );
  assign n1428 = n1343 & n1361 ;
  buffer buf_n1429( .i (n1428), .o (n1429) );
  assign n1430 = n1381 & n1399 ;
  buffer buf_n1431( .i (n1430), .o (n1431) );
  assign n1432 = n1429 | n1431 ;
  buffer buf_n1433( .i (n1432), .o (n1433) );
  assign n1434 = ( n1420 & n1427 ) | ( n1420 & n1433 ) | ( n1427 & n1433 ) ;
  buffer buf_n1435( .i (n1434), .o (n1435) );
  assign n1436 = n534 & n956 ;
  buffer buf_n1437( .i (n1436), .o (n1437) );
  assign n1438 = n1004 & n1050 ;
  buffer buf_n1439( .i (n1438), .o (n1439) );
  assign n1440 = n1437 & n1439 ;
  buffer buf_n1441( .i (n1440), .o (n1441) );
  assign n1442 = n1076 & n1098 ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  assign n1444 = n1122 & n1144 ;
  buffer buf_n1445( .i (n1444), .o (n1445) );
  assign n1446 = n1443 & n1445 ;
  buffer buf_n1447( .i (n1446), .o (n1447) );
  assign n1448 = n1441 | n1447 ;
  buffer buf_n1449( .i (n1448), .o (n1449) );
  assign n1450 = n1160 & n1170 ;
  buffer buf_n1451( .i (n1450), .o (n1451) );
  assign n1452 = n1182 & n1192 ;
  buffer buf_n1453( .i (n1452), .o (n1453) );
  assign n1454 = n1451 & n1453 ;
  buffer buf_n1455( .i (n1454), .o (n1455) );
  assign n1456 = n1206 & n1216 ;
  buffer buf_n1457( .i (n1456), .o (n1457) );
  assign n1458 = n1228 & n1238 ;
  buffer buf_n1459( .i (n1458), .o (n1459) );
  assign n1460 = n1457 & n1459 ;
  buffer buf_n1461( .i (n1460), .o (n1461) );
  assign n1462 = n1455 | n1461 ;
  buffer buf_n1463( .i (n1462), .o (n1463) );
  assign n1464 = n1449 | n1463 ;
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  assign n1467 = n1250 & n1253 ;
  buffer buf_n1468( .i (n1467), .o (n1468) );
  assign n1469 = n1258 & n1261 ;
  buffer buf_n1470( .i (n1469), .o (n1470) );
  assign n1471 = n1468 & n1470 ;
  buffer buf_n1472( .i (n1471), .o (n1472) );
  assign n1473 = n1268 & n1271 ;
  buffer buf_n1474( .i (n1473), .o (n1474) );
  assign n1475 = n1276 & n1279 ;
  buffer buf_n1476( .i (n1475), .o (n1476) );
  assign n1477 = n1474 & n1476 ;
  buffer buf_n1478( .i (n1477), .o (n1478) );
  assign n1479 = n1472 | n1478 ;
  buffer buf_n1480( .i (n1479), .o (n1480) );
  assign n1481 = n1288 & n1291 ;
  buffer buf_n1482( .i (n1481), .o (n1482) );
  assign n1483 = n1296 & n1299 ;
  buffer buf_n1484( .i (n1483), .o (n1484) );
  assign n1485 = n1482 & n1484 ;
  buffer buf_n1486( .i (n1485), .o (n1486) );
  assign n1487 = n1306 & n1309 ;
  buffer buf_n1488( .i (n1487), .o (n1488) );
  assign n1489 = n1314 & n1317 ;
  buffer buf_n1490( .i (n1489), .o (n1490) );
  assign n1491 = n1488 & n1490 ;
  buffer buf_n1492( .i (n1491), .o (n1492) );
  assign n1493 = n1486 | n1492 ;
  buffer buf_n1494( .i (n1493), .o (n1494) );
  assign n1495 = n1480 | n1494 ;
  buffer buf_n1496( .i (n1495), .o (n1496) );
  assign n1497 = n1328 & n1331 ;
  buffer buf_n1498( .i (n1497), .o (n1498) );
  assign n1499 = n1336 & n1339 ;
  buffer buf_n1500( .i (n1499), .o (n1500) );
  assign n1501 = n1498 & n1500 ;
  buffer buf_n1502( .i (n1501), .o (n1502) );
  assign n1503 = n1346 & n1349 ;
  buffer buf_n1504( .i (n1503), .o (n1504) );
  assign n1505 = n1354 & n1357 ;
  buffer buf_n1506( .i (n1505), .o (n1506) );
  assign n1507 = n1504 & n1506 ;
  buffer buf_n1508( .i (n1507), .o (n1508) );
  assign n1509 = n1502 | n1508 ;
  buffer buf_n1510( .i (n1509), .o (n1510) );
  assign n1511 = n1366 & n1369 ;
  buffer buf_n1512( .i (n1511), .o (n1512) );
  assign n1513 = n1374 & n1377 ;
  buffer buf_n1514( .i (n1513), .o (n1514) );
  assign n1515 = n1512 & n1514 ;
  buffer buf_n1516( .i (n1515), .o (n1516) );
  assign n1517 = n1384 & n1387 ;
  buffer buf_n1518( .i (n1517), .o (n1518) );
  assign n1519 = n1392 & n1395 ;
  buffer buf_n1520( .i (n1519), .o (n1520) );
  assign n1521 = n1518 & n1520 ;
  buffer buf_n1522( .i (n1521), .o (n1522) );
  assign n1523 = n1516 | n1522 ;
  buffer buf_n1524( .i (n1523), .o (n1524) );
  assign n1525 = n1510 | n1524 ;
  buffer buf_n1526( .i (n1525), .o (n1526) );
  assign n1527 = n1496 | n1526 ;
  assign n1528 = n1466 | n1527 ;
  assign n1529 = n1449 & n1463 ;
  buffer buf_n1530( .i (n1529), .o (n1530) );
  assign n1532 = n1480 & n1494 ;
  buffer buf_n1533( .i (n1532), .o (n1533) );
  assign n1534 = n1510 & n1524 ;
  buffer buf_n1535( .i (n1534), .o (n1535) );
  assign n1536 = ( n1530 & n1533 ) | ( n1530 & n1535 ) | ( n1533 & n1535 ) ;
  buffer buf_n1537( .i (n1536), .o (n1537) );
  assign n1538 = n1441 & n1447 ;
  buffer buf_n1539( .i (n1538), .o (n1539) );
  assign n1540 = n1455 & n1461 ;
  buffer buf_n1541( .i (n1540), .o (n1541) );
  assign n1542 = n1539 | n1541 ;
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  assign n1545 = n1472 & n1478 ;
  buffer buf_n1546( .i (n1545), .o (n1546) );
  assign n1547 = n1486 & n1492 ;
  buffer buf_n1548( .i (n1547), .o (n1548) );
  assign n1549 = n1546 | n1548 ;
  buffer buf_n1550( .i (n1549), .o (n1550) );
  assign n1551 = n1502 & n1508 ;
  buffer buf_n1552( .i (n1551), .o (n1552) );
  assign n1553 = n1516 & n1522 ;
  buffer buf_n1554( .i (n1553), .o (n1554) );
  assign n1555 = n1552 | n1554 ;
  buffer buf_n1556( .i (n1555), .o (n1556) );
  assign n1557 = n1550 | n1556 ;
  assign n1558 = n1544 | n1557 ;
  assign n1559 = n958 & n1052 ;
  buffer buf_n1560( .i (n1559), .o (n1560) );
  assign n1561 = n1100 & n1146 ;
  buffer buf_n1562( .i (n1561), .o (n1562) );
  assign n1563 = n1560 | n1562 ;
  buffer buf_n1564( .i (n1563), .o (n1564) );
  assign n1565 = n1172 & n1194 ;
  buffer buf_n1566( .i (n1565), .o (n1566) );
  assign n1567 = n1218 & n1240 ;
  buffer buf_n1568( .i (n1567), .o (n1568) );
  assign n1569 = n1566 | n1568 ;
  buffer buf_n1570( .i (n1569), .o (n1570) );
  assign n1571 = n1564 & n1570 ;
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  assign n1574 = n1255 & n1263 ;
  buffer buf_n1575( .i (n1574), .o (n1575) );
  assign n1576 = n1273 & n1281 ;
  buffer buf_n1577( .i (n1576), .o (n1577) );
  assign n1578 = n1575 | n1577 ;
  buffer buf_n1579( .i (n1578), .o (n1579) );
  assign n1580 = n1293 & n1301 ;
  buffer buf_n1581( .i (n1580), .o (n1581) );
  assign n1582 = n1311 & n1319 ;
  buffer buf_n1583( .i (n1582), .o (n1583) );
  assign n1584 = n1581 | n1583 ;
  buffer buf_n1585( .i (n1584), .o (n1585) );
  assign n1586 = n1579 & n1585 ;
  buffer buf_n1587( .i (n1586), .o (n1587) );
  assign n1588 = n1333 & n1341 ;
  buffer buf_n1589( .i (n1588), .o (n1589) );
  assign n1590 = n1351 & n1359 ;
  buffer buf_n1591( .i (n1590), .o (n1591) );
  assign n1592 = n1589 | n1591 ;
  buffer buf_n1593( .i (n1592), .o (n1593) );
  assign n1594 = n1371 & n1379 ;
  buffer buf_n1595( .i (n1594), .o (n1595) );
  assign n1596 = n1389 & n1397 ;
  buffer buf_n1597( .i (n1596), .o (n1597) );
  assign n1598 = n1595 | n1597 ;
  buffer buf_n1599( .i (n1598), .o (n1599) );
  assign n1600 = n1593 & n1599 ;
  buffer buf_n1601( .i (n1600), .o (n1601) );
  assign n1602 = n1587 | n1601 ;
  assign n1603 = n1573 | n1602 ;
  assign n1604 = n1437 | n1439 ;
  buffer buf_n1605( .i (n1604), .o (n1605) );
  assign n1606 = n1443 | n1445 ;
  buffer buf_n1607( .i (n1606), .o (n1607) );
  assign n1608 = n1605 & n1607 ;
  buffer buf_n1609( .i (n1608), .o (n1609) );
  assign n1610 = n1451 | n1453 ;
  buffer buf_n1611( .i (n1610), .o (n1611) );
  assign n1612 = n1457 | n1459 ;
  buffer buf_n1613( .i (n1612), .o (n1613) );
  assign n1614 = n1611 & n1613 ;
  buffer buf_n1615( .i (n1614), .o (n1615) );
  assign n1616 = n1609 | n1615 ;
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  assign n1619 = n1468 | n1470 ;
  buffer buf_n1620( .i (n1619), .o (n1620) );
  assign n1621 = n1474 | n1476 ;
  buffer buf_n1622( .i (n1621), .o (n1622) );
  assign n1623 = n1620 & n1622 ;
  buffer buf_n1624( .i (n1623), .o (n1624) );
  assign n1625 = n1482 | n1484 ;
  buffer buf_n1626( .i (n1625), .o (n1626) );
  assign n1627 = n1488 | n1490 ;
  buffer buf_n1628( .i (n1627), .o (n1628) );
  assign n1629 = n1626 & n1628 ;
  buffer buf_n1630( .i (n1629), .o (n1630) );
  assign n1631 = n1624 | n1630 ;
  buffer buf_n1632( .i (n1631), .o (n1632) );
  assign n1633 = n1498 | n1500 ;
  buffer buf_n1634( .i (n1633), .o (n1634) );
  assign n1635 = n1504 | n1506 ;
  buffer buf_n1636( .i (n1635), .o (n1636) );
  assign n1637 = n1634 & n1636 ;
  buffer buf_n1638( .i (n1637), .o (n1638) );
  assign n1639 = n1512 | n1514 ;
  buffer buf_n1640( .i (n1639), .o (n1640) );
  assign n1641 = n1518 | n1520 ;
  buffer buf_n1642( .i (n1641), .o (n1642) );
  assign n1643 = n1640 & n1642 ;
  buffer buf_n1644( .i (n1643), .o (n1644) );
  assign n1645 = n1638 | n1644 ;
  buffer buf_n1646( .i (n1645), .o (n1646) );
  assign n1647 = n1632 | n1646 ;
  assign n1648 = n1618 | n1647 ;
  assign n1649 = n1560 & n1562 ;
  buffer buf_n1650( .i (n1649), .o (n1650) );
  assign n1651 = n1566 & n1568 ;
  buffer buf_n1652( .i (n1651), .o (n1652) );
  assign n1653 = n1650 | n1652 ;
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  assign n1656 = n1575 & n1577 ;
  buffer buf_n1657( .i (n1656), .o (n1657) );
  assign n1658 = n1581 & n1583 ;
  buffer buf_n1659( .i (n1658), .o (n1659) );
  assign n1660 = n1657 | n1659 ;
  buffer buf_n1661( .i (n1660), .o (n1661) );
  assign n1662 = n1589 & n1591 ;
  buffer buf_n1663( .i (n1662), .o (n1663) );
  assign n1664 = n1595 & n1597 ;
  buffer buf_n1665( .i (n1664), .o (n1665) );
  assign n1666 = n1663 | n1665 ;
  buffer buf_n1667( .i (n1666), .o (n1667) );
  assign n1668 = n1661 | n1667 ;
  assign n1669 = n1655 | n1668 ;
  assign n1670 = n1650 & n1652 ;
  buffer buf_n1671( .i (n1670), .o (n1671) );
  assign n1673 = n1657 & n1659 ;
  buffer buf_n1674( .i (n1673), .o (n1674) );
  assign n1675 = n1663 & n1665 ;
  buffer buf_n1676( .i (n1675), .o (n1676) );
  assign n1677 = ( n1671 & n1674 ) | ( n1671 & n1676 ) | ( n1674 & n1676 ) ;
  buffer buf_n1678( .i (n1677), .o (n1678) );
  assign n1679 = n1609 & n1615 ;
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  assign n1682 = n1624 & n1630 ;
  buffer buf_n1683( .i (n1682), .o (n1683) );
  assign n1684 = n1638 & n1644 ;
  buffer buf_n1685( .i (n1684), .o (n1685) );
  assign n1686 = n1683 & n1685 ;
  assign n1687 = n1681 & n1686 ;
  assign n1688 = ( n1617 & n1632 ) | ( n1617 & n1646 ) | ( n1632 & n1646 ) ;
  buffer buf_n1689( .i (n1688), .o (n1689) );
  assign n1690 = n1539 & n1541 ;
  buffer buf_n1691( .i (n1690), .o (n1691) );
  assign n1693 = n1546 & n1548 ;
  buffer buf_n1694( .i (n1693), .o (n1694) );
  assign n1695 = n1552 & n1554 ;
  buffer buf_n1696( .i (n1695), .o (n1696) );
  assign n1697 = ( n1691 & n1694 ) | ( n1691 & n1696 ) | ( n1694 & n1696 ) ;
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  assign n1699 = n1410 & n1412 ;
  assign n1700 = n1408 & n1699 ;
  buffer buf_n1692( .i (n1691), .o (n1692) );
  assign n1701 = n1694 & n1696 ;
  assign n1702 = n1692 & n1701 ;
  assign n1703 = ( n1654 & n1661 ) | ( n1654 & n1667 ) | ( n1661 & n1667 ) ;
  buffer buf_n1704( .i (n1703), .o (n1704) );
  assign n1705 = n1496 & n1526 ;
  assign n1706 = n1466 & n1705 ;
  assign n1707 = n1416 & n1418 ;
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  assign n1710 = n1423 & n1425 ;
  buffer buf_n1711( .i (n1710), .o (n1711) );
  assign n1712 = n1429 & n1431 ;
  buffer buf_n1713( .i (n1712), .o (n1713) );
  assign n1714 = n1711 & n1713 ;
  assign n1715 = n1709 & n1714 ;
  assign n1716 = n1694 | n1696 ;
  assign n1717 = n1692 | n1716 ;
  assign n1718 = n1605 | n1607 ;
  buffer buf_n1719( .i (n1718), .o (n1719) );
  assign n1720 = n1611 | n1613 ;
  buffer buf_n1721( .i (n1720), .o (n1721) );
  assign n1722 = n1719 & n1721 ;
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  assign n1725 = n1620 | n1622 ;
  buffer buf_n1726( .i (n1725), .o (n1726) );
  assign n1727 = n1626 | n1628 ;
  buffer buf_n1728( .i (n1727), .o (n1728) );
  assign n1729 = n1726 & n1728 ;
  buffer buf_n1730( .i (n1729), .o (n1730) );
  assign n1731 = n1634 | n1636 ;
  buffer buf_n1732( .i (n1731), .o (n1732) );
  assign n1733 = n1640 | n1642 ;
  buffer buf_n1734( .i (n1733), .o (n1734) );
  assign n1735 = n1732 & n1734 ;
  buffer buf_n1736( .i (n1735), .o (n1736) );
  assign n1737 = n1730 | n1736 ;
  assign n1738 = n1724 | n1737 ;
  buffer buf_n1421( .i (n1420), .o (n1421) );
  assign n1739 = n1427 | n1433 ;
  assign n1740 = n1421 | n1739 ;
  assign n1741 = n1564 | n1570 ;
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  assign n1744 = n1579 | n1585 ;
  buffer buf_n1745( .i (n1744), .o (n1745) );
  assign n1746 = n1593 | n1599 ;
  buffer buf_n1747( .i (n1746), .o (n1747) );
  assign n1748 = n1745 & n1747 ;
  assign n1749 = n1743 & n1748 ;
  assign n1750 = ( n1572 & n1587 ) | ( n1572 & n1601 ) | ( n1587 & n1601 ) ;
  buffer buf_n1751( .i (n1750), .o (n1751) );
  assign n1752 = ( n1742 & n1745 ) | ( n1742 & n1747 ) | ( n1745 & n1747 ) ;
  buffer buf_n1753( .i (n1752), .o (n1753) );
  assign n1754 = ( n1680 & n1683 ) | ( n1680 & n1685 ) | ( n1683 & n1685 ) ;
  buffer buf_n1755( .i (n1754), .o (n1755) );
  assign n1756 = n1719 | n1721 ;
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  assign n1759 = n1726 | n1728 ;
  buffer buf_n1760( .i (n1759), .o (n1760) );
  assign n1761 = n1732 | n1734 ;
  buffer buf_n1762( .i (n1761), .o (n1762) );
  assign n1763 = n1760 & n1762 ;
  assign n1764 = n1758 & n1763 ;
  assign n1765 = n1745 | n1747 ;
  assign n1766 = n1743 | n1765 ;
  assign n1767 = n1427 & n1433 ;
  assign n1768 = n1421 & n1767 ;
  assign n1769 = n1661 & n1667 ;
  assign n1770 = n1655 & n1769 ;
  assign n1771 = ( n1246 & n1325 ) | ( n1246 & n1403 ) | ( n1325 & n1403 ) ;
  buffer buf_n1772( .i (n1771), .o (n1772) );
  assign n1773 = ( n1543 & n1550 ) | ( n1543 & n1556 ) | ( n1550 & n1556 ) ;
  buffer buf_n1774( .i (n1773), .o (n1774) );
  assign n1775 = n1683 | n1685 ;
  assign n1776 = n1681 | n1775 ;
  assign n1777 = ( n1708 & n1711 ) | ( n1708 & n1713 ) | ( n1711 & n1713 ) ;
  buffer buf_n1778( .i (n1777), .o (n1778) );
  assign n1779 = ( n1757 & n1760 ) | ( n1757 & n1762 ) | ( n1760 & n1762 ) ;
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  assign n1781 = n1533 & n1535 ;
  assign n1782 = n1531 & n1781 ;
  assign n1783 = n1711 | n1713 ;
  assign n1784 = n1709 | n1783 ;
  assign n1785 = n1730 & n1736 ;
  assign n1786 = n1724 & n1785 ;
  assign n1787 = n1632 & n1646 ;
  assign n1788 = n1618 & n1787 ;
  assign n1789 = n1587 & n1601 ;
  assign n1790 = n1573 & n1789 ;
  assign n1791 = n1533 | n1535 ;
  assign n1792 = n1531 | n1791 ;
  buffer buf_n1672( .i (n1671), .o (n1672) );
  assign n1793 = n1674 | n1676 ;
  assign n1794 = n1672 | n1793 ;
  assign n1795 = n1674 & n1676 ;
  assign n1796 = n1672 & n1795 ;
  assign n1797 = ( n1723 & n1730 ) | ( n1723 & n1736 ) | ( n1730 & n1736 ) ;
  buffer buf_n1798( .i (n1797), .o (n1798) );
  assign n1799 = n1760 | n1762 ;
  assign n1800 = n1758 | n1799 ;
  assign n1801 = ( n1465 & n1496 ) | ( n1465 & n1526 ) | ( n1496 & n1526 ) ;
  buffer buf_n1802( .i (n1801), .o (n1802) );
  assign n1803 = n1550 & n1556 ;
  assign n1804 = n1544 & n1803 ;
  assign n1805 = n1325 & n1403 ;
  assign n1806 = n1247 & n1805 ;
  assign n1807 = n1410 | n1412 ;
  assign n1808 = n1408 | n1807 ;
  assign y0 = n1405 ;
  assign y1 = n1414 ;
  assign y2 = n1435 ;
  assign y3 = n1528 ;
  assign y4 = n1537 ;
  assign y5 = n1558 ;
  assign y6 = n1603 ;
  assign y7 = n1648 ;
  assign y8 = n1669 ;
  assign y9 = n1678 ;
  assign y10 = n1687 ;
  assign y11 = n1689 ;
  assign y12 = n1698 ;
  assign y13 = n1700 ;
  assign y14 = n1702 ;
  assign y15 = n1704 ;
  assign y16 = n1706 ;
  assign y17 = n1715 ;
  assign y18 = n1717 ;
  assign y19 = n1738 ;
  assign y20 = n1740 ;
  assign y21 = n1749 ;
  assign y22 = n1751 ;
  assign y23 = n1753 ;
  assign y24 = n1755 ;
  assign y25 = n1764 ;
  assign y26 = n1766 ;
  assign y27 = n1768 ;
  assign y28 = n1770 ;
  assign y29 = n1772 ;
  assign y30 = n1774 ;
  assign y31 = n1776 ;
  assign y32 = n1778 ;
  assign y33 = n1780 ;
  assign y34 = n1782 ;
  assign y35 = n1784 ;
  assign y36 = n1786 ;
  assign y37 = n1788 ;
  assign y38 = n1790 ;
  assign y39 = n1792 ;
  assign y40 = n1794 ;
  assign y41 = n1796 ;
  assign y42 = n1798 ;
  assign y43 = n1800 ;
  assign y44 = n1802 ;
  assign y45 = n1804 ;
  assign y46 = n1806 ;
  assign y47 = n1808 ;
endmodule
