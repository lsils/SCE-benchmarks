module top( in_6_ , in_15_ , in_13_ , in_14_ , in_2_ , in_10_ , in_24_ , in_8_ , in_22_ , in_20_ , in_7_ , in_25_ , in_5_ , in_4_ , in_23_ , in_27_ , in_1_ , in_0_ , in_16_ , in_30_ , in_26_ , in_12_ , in_11_ , in_17_ , in_19_ , in_18_ , in_21_ , in_31_ , in_29_ , in_28_ , in_9_ , in_3_ , out_2_ , out_1_ , out_3_ , out_0_ , out_5_ , out_4_ );
  input in_6_ , in_15_ , in_13_ , in_14_ , in_2_ , in_10_ , in_24_ , in_8_ , in_22_ , in_20_ , in_7_ , in_25_ , in_5_ , in_4_ , in_23_ , in_27_ , in_1_ , in_0_ , in_16_ , in_30_ , in_26_ , in_12_ , in_11_ , in_17_ , in_19_ , in_18_ , in_21_ , in_31_ , in_29_ , in_28_ , in_9_ , in_3_ ;
  output out_2_ , out_1_ , out_3_ , out_0_ , out_5_ , out_4_ ;
  wire n33 , n41 , n45 , n47 , n49 , n55 , n57 , n59 , n63 , n65 , n67 , n73 , n75 , n77 , n81 , n87 , n89 , n91 , n101 , n103 , n105 , n107 , n109 , n111 , n113 , n121 , n125 , n127 , n129 , n135 , n137 , n139 , n143 , n145 , n147 , n153 , n155 , n157 , n161 , n167 , n169 , n171 , n181 , n183 , n185 , n187 , n189 , n191 , n193 , n194 , n195 , n197 , n199 , n201 , n203 , n205 , n210 , n211 , n212 , n215 , n217 , n224 , n230 , n232 , n234 , n240 , n242 , n244 , n245 , n246 , n248 , n253 , n254 , n255 , n256 , n258 , n261 , n262 , n263 , n265 , n266 , n267 ;
  assign n33 = in_29_ | in_28_ ;
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  assign n41 = in_20_ | in_21_ ;
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  assign n45 = in_16_ | in_17_ ;
  buffer buf_n46( .i (n45), .o (n46) );
  assign n47 = in_19_ & in_18_ ;
  buffer buf_n48( .i (n47), .o (n48) );
  assign n49 = ( n42 & n46 ) | ( n42 & n48 ) | ( n46 & n48 ) ;
  buffer buf_n50( .i (n49), .o (n50) );
  assign n55 = ( ~n42 & n46 ) | ( ~n42 & n48 ) | ( n46 & n48 ) ;
  buffer buf_n56( .i (n55), .o (n56) );
  assign n57 = ( n44 & ~n50 ) | ( n44 & n56 ) | ( ~n50 & n56 ) ;
  buffer buf_n58( .i (n57), .o (n58) );
  assign n59 = in_27_ & in_26_ ;
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  assign n63 = in_22_ & in_23_ ;
  buffer buf_n64( .i (n63), .o (n64) );
  assign n65 = in_24_ | in_25_ ;
  buffer buf_n66( .i (n65), .o (n66) );
  assign n67 = ( n60 & n64 ) | ( n60 & n66 ) | ( n64 & n66 ) ;
  buffer buf_n68( .i (n67), .o (n68) );
  assign n73 = ( ~n60 & n64 ) | ( ~n60 & n66 ) | ( n64 & n66 ) ;
  buffer buf_n74( .i (n73), .o (n74) );
  assign n75 = ( n62 & ~n68 ) | ( n62 & n74 ) | ( ~n68 & n74 ) ;
  buffer buf_n76( .i (n75), .o (n76) );
  assign n77 = ( n38 & n58 ) | ( n38 & n76 ) | ( n58 & n76 ) ;
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  assign n81 = ( n54 & n72 ) | ( n54 & n78 ) | ( n72 & n78 ) ;
  buffer buf_n82( .i (n81), .o (n82) );
  assign n87 = ( n54 & n72 ) | ( n54 & ~n78 ) | ( n72 & ~n78 ) ;
  buffer buf_n88( .i (n87), .o (n88) );
  assign n89 = ( n80 & ~n82 ) | ( n80 & n88 ) | ( ~n82 & n88 ) ;
  buffer buf_n90( .i (n89), .o (n90) );
  assign n91 = in_30_ & in_31_ ;
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  assign n101 = ( ~n38 & n58 ) | ( ~n38 & n76 ) | ( n58 & n76 ) ;
  buffer buf_n102( .i (n101), .o (n102) );
  assign n103 = ( n40 & ~n78 ) | ( n40 & n102 ) | ( ~n78 & n102 ) ;
  buffer buf_n104( .i (n103), .o (n104) );
  assign n105 = n100 & n104 ;
  buffer buf_n106( .i (n105), .o (n106) );
  assign n107 = n90 & n106 ;
  buffer buf_n108( .i (n107), .o (n108) );
  assign n109 = n90 | n106 ;
  buffer buf_n110( .i (n109), .o (n110) );
  assign n111 = ~n108 & n110 ;
  buffer buf_n112( .i (n111), .o (n112) );
  assign n113 = in_13_ | in_12_ ;
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  assign n121 = in_5_ | in_4_ ;
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  assign n125 = in_1_ | in_0_ ;
  buffer buf_n126( .i (n125), .o (n126) );
  assign n127 = in_2_ & in_3_ ;
  buffer buf_n128( .i (n127), .o (n128) );
  assign n129 = ( n122 & n126 ) | ( n122 & n128 ) | ( n126 & n128 ) ;
  buffer buf_n130( .i (n129), .o (n130) );
  assign n135 = ( ~n122 & n126 ) | ( ~n122 & n128 ) | ( n126 & n128 ) ;
  buffer buf_n136( .i (n135), .o (n136) );
  assign n137 = ( n124 & ~n130 ) | ( n124 & n136 ) | ( ~n130 & n136 ) ;
  buffer buf_n138( .i (n137), .o (n138) );
  assign n139 = in_10_ & in_11_ ;
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  assign n143 = in_6_ & in_7_ ;
  buffer buf_n144( .i (n143), .o (n144) );
  assign n145 = in_8_ | in_9_ ;
  buffer buf_n146( .i (n145), .o (n146) );
  assign n147 = ( n140 & n144 ) | ( n140 & n146 ) | ( n144 & n146 ) ;
  buffer buf_n148( .i (n147), .o (n148) );
  assign n153 = ( ~n140 & n144 ) | ( ~n140 & n146 ) | ( n144 & n146 ) ;
  buffer buf_n154( .i (n153), .o (n154) );
  assign n155 = ( n142 & ~n148 ) | ( n142 & n154 ) | ( ~n148 & n154 ) ;
  buffer buf_n156( .i (n155), .o (n156) );
  assign n157 = ( n118 & n138 ) | ( n118 & n156 ) | ( n138 & n156 ) ;
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  assign n161 = ( n134 & n152 ) | ( n134 & n158 ) | ( n152 & n158 ) ;
  buffer buf_n162( .i (n161), .o (n162) );
  assign n167 = ( n134 & n152 ) | ( n134 & ~n158 ) | ( n152 & ~n158 ) ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = ( n160 & ~n162 ) | ( n160 & n168 ) | ( ~n162 & n168 ) ;
  buffer buf_n170( .i (n169), .o (n170) );
  assign n171 = in_15_ & in_14_ ;
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  assign n181 = ( ~n118 & n138 ) | ( ~n118 & n156 ) | ( n138 & n156 ) ;
  buffer buf_n182( .i (n181), .o (n182) );
  assign n183 = ( n120 & ~n158 ) | ( n120 & n182 ) | ( ~n158 & n182 ) ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n185 = n180 & n184 ;
  buffer buf_n186( .i (n185), .o (n186) );
  assign n187 = n170 & n186 ;
  buffer buf_n188( .i (n187), .o (n188) );
  assign n189 = n170 | n186 ;
  buffer buf_n190( .i (n189), .o (n190) );
  assign n191 = ~n188 & n190 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = n112 & n192 ;
  assign n194 = n112 | n192 ;
  assign n195 = ~n193 & n194 ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n197 = n100 | n104 ;
  buffer buf_n198( .i (n197), .o (n198) );
  assign n199 = ~n106 & n198 ;
  buffer buf_n200( .i (n199), .o (n200) );
  assign n201 = n180 | n184 ;
  buffer buf_n202( .i (n201), .o (n202) );
  assign n203 = ~n186 & n202 ;
  buffer buf_n204( .i (n203), .o (n204) );
  assign n205 = n200 & n204 ;
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  assign n210 = n196 & n209 ;
  assign n211 = n196 | n209 ;
  assign n212 = ~n210 & n211 ;
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n215 = n200 | n204 ;
  buffer buf_n216( .i (n215), .o (n216) );
  assign n217 = ~n206 & n216 ;
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  assign n224 = n86 & n108 ;
  buffer buf_n225( .i (n224), .o (n225) );
  assign n230 = n86 | n108 ;
  buffer buf_n231( .i (n230), .o (n231) );
  assign n232 = ~n225 & n231 ;
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  assign n234 = n166 & n188 ;
  buffer buf_n235( .i (n234), .o (n235) );
  assign n240 = n166 | n188 ;
  buffer buf_n241( .i (n240), .o (n241) );
  assign n242 = ~n235 & n241 ;
  buffer buf_n243( .i (n242), .o (n243) );
  assign n244 = n233 & n243 ;
  assign n245 = n233 | n243 ;
  assign n246 = ~n244 & n245 ;
  buffer buf_n247( .i (n246), .o (n247) );
  assign n248 = ( n112 & n192 ) | ( n112 & n206 ) | ( n192 & n206 ) ;
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  assign n253 = n247 & n252 ;
  assign n254 = n247 | n252 ;
  assign n255 = ~n253 & n254 ;
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  assign n256 = ( n233 & n243 ) | ( n233 & n249 ) | ( n243 & n249 ) ;
  buffer buf_n257( .i (n256), .o (n257) );
  assign n258 = ( n229 & n239 ) | ( n229 & n257 ) | ( n239 & n257 ) ;
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  assign n261 = n226 | n236 ;
  assign n262 = n226 & n236 ;
  assign n263 = n261 & ~n262 ;
  buffer buf_n264( .i (n263), .o (n264) );
  assign n265 = n257 & n264 ;
  assign n266 = n257 | n264 ;
  assign n267 = ~n265 & n266 ;
  buffer buf_n268( .i (n267), .o (n268) );
  assign out_2_ = n214 ;
  assign out_1_ = n223 ;
  assign out_3_ = n255 ;
  assign out_0_ = 1'b0 ;
  assign out_5_ = n260 ;
  assign out_4_ = n268 ;
endmodule
