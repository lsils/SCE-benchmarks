module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( N1 , N102 , N105 , N108 , N11 , N112 , N115 , N14 , N17 , N21 , N24 , N27 , N30 , N34 , N37 , N4 , N40 , N43 , N47 , N50 , N53 , N56 , N60 , N63 , N66 , N69 , N73 , N76 , N79 , N8 , N82 , N86 , N89 , N92 , N95 , N99 , N223 , N329 , N370 , N421 , N430 , N431 , N432 );
  input N1 , N102 , N105 , N108 , N11 , N112 , N115 , N14 , N17 , N21 , N24 , N27 , N30 , N34 , N37 , N4 , N40 , N43 , N47 , N50 , N53 , N56 , N60 , N63 , N66 , N69 , N73 , N76 , N79 , N8 , N82 , N86 , N89 , N92 , N95 , N99 ;
  output N223 , N329 , N370 , N421 , N430 , N431 , N432 ;
  wire n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 ;
  assign n37 = ~N24 & N30 ;
  buffer buf_n38( .i (n37), .o (n38) );
  assign n44 = ~N102 & N108 ;
  assign n45 = n38 | n44 ;
  assign n46 = ~N1 & N4 ;
  assign n47 = ~N89 & N95 ;
  assign n48 = ~N76 & N82 ;
  assign n49 = n47 | n48 ;
  assign n50 = n46 | n49 ;
  assign n51 = ~N63 & N69 ;
  buffer buf_n52( .i (n51), .o (n52) );
  assign n59 = ~N37 & N43 ;
  assign n60 = n52 | n59 ;
  assign n61 = ~N50 & N56 ;
  assign n62 = ~N11 & N17 ;
  assign n63 = n61 | n62 ;
  assign n64 = n60 | n63 ;
  assign n65 = n50 | n64 ;
  assign n66 = n45 | n65 ;
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  assign n97 = N102 & n68 ;
  assign n98 = N108 & ~n97 ;
  buffer buf_n99( .i (n98), .o (n99) );
  assign n107 = ~N112 & n99 ;
  assign n108 = N76 & n68 ;
  assign n109 = N82 & ~n108 ;
  buffer buf_n110( .i (n109), .o (n110) );
  assign n119 = ~N86 & n110 ;
  assign n120 = n107 | n119 ;
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  assign n121 = N30 & ~n68 ;
  assign n122 = n43 | n121 ;
  buffer buf_n123( .i (n122), .o (n123) );
  assign n133 = ~N34 & n123 ;
  buffer buf_n134( .i (n67), .o (n134) );
  assign n135 = N11 & n134 ;
  assign n136 = N17 & ~n135 ;
  buffer buf_n137( .i (n136), .o (n137) );
  assign n146 = ~N21 & n137 ;
  assign n147 = n133 | n146 ;
  assign n148 = n120 | n147 ;
  assign n149 = N1 & n134 ;
  assign n150 = N4 & ~n149 ;
  buffer buf_n151( .i (n150), .o (n151) );
  assign n160 = ~N8 & n151 ;
  assign n161 = N89 & n134 ;
  assign n162 = N95 & ~n161 ;
  buffer buf_n163( .i (n162), .o (n163) );
  assign n172 = ~N99 & n163 ;
  assign n173 = n160 | n172 ;
  assign n174 = N50 & n134 ;
  assign n175 = N56 & ~n174 ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n183 = ~N60 & n176 ;
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  assign n184 = N69 & ~n67 ;
  assign n185 = n58 | n184 ;
  buffer buf_n186( .i (n185), .o (n186) );
  assign n195 = ~N73 & n186 ;
  assign n196 = N37 & n67 ;
  assign n197 = N43 & ~n196 ;
  buffer buf_n198( .i (n197), .o (n198) );
  assign n207 = ~N47 & n198 ;
  assign n208 = n195 | n207 ;
  assign n209 = n183 | n208 ;
  assign n210 = n173 | n209 ;
  assign n211 = n148 | n210 ;
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  assign n233 = N34 & n215 ;
  assign n234 = n132 & ~n233 ;
  buffer buf_n235( .i (n234), .o (n235) );
  assign n242 = ~N40 & n235 ;
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  assign n243 = N99 & n214 ;
  assign n244 = n171 & ~n243 ;
  buffer buf_n245( .i (n244), .o (n245) );
  assign n254 = ~N105 & n245 ;
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  assign n255 = N21 & n214 ;
  assign n256 = n145 & ~n255 ;
  buffer buf_n257( .i (n256), .o (n257) );
  assign n265 = ~N27 & n257 ;
  assign n266 = n254 | n265 ;
  assign n267 = n242 | n266 ;
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  assign n268 = N8 & n214 ;
  assign n269 = n159 & ~n268 ;
  buffer buf_n270( .i (n269), .o (n270) );
  assign n284 = ~N14 & n270 ;
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n285( .i (n213), .o (n285) );
  assign n286 = N86 & n285 ;
  assign n287 = n118 & ~n286 ;
  buffer buf_n288( .i (n287), .o (n288) );
  assign n297 = ~N92 & n288 ;
  assign n298 = n284 | n297 ;
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  assign n299 = N73 & n213 ;
  assign n300 = n194 & ~n299 ;
  buffer buf_n301( .i (n300), .o (n301) );
  assign n311 = ~N79 & n301 ;
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  assign n312 = N60 & n212 ;
  assign n313 = n182 & ~n312 ;
  buffer buf_n314( .i (n313), .o (n314) );
  assign n324 = ~N66 & n314 ;
  buffer buf_n325( .i (n324), .o (n325) );
  assign n334 = n311 | n325 ;
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  assign n335 = N47 & n213 ;
  assign n336 = n206 & ~n335 ;
  buffer buf_n337( .i (n336), .o (n337) );
  assign n346 = ~N53 & n337 ;
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n347( .i (n212), .o (n347) );
  assign n348 = N112 & n347 ;
  assign n349 = n106 & ~n348 ;
  buffer buf_n350( .i (n349), .o (n350) );
  assign n362 = ~N115 & n350 ;
  assign n363 = n346 | n362 ;
  assign n364 = n334 | n363 ;
  assign n365 = n298 | n364 ;
  assign n366 = n267 | n365 ;
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  assign n378 = N40 & n368 ;
  assign n379 = n241 & ~n378 ;
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  assign n385 = N27 & n368 ;
  assign n386 = n264 & ~n385 ;
  buffer buf_n387( .i (n386), .o (n387) );
  assign n393 = n380 | n387 ;
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  assign n397 = N53 & n368 ;
  assign n398 = n345 & ~n397 ;
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  assign n402 = n323 & ~n369 ;
  assign n403 = n333 | n402 ;
  assign n404 = n399 | n403 ;
  buffer buf_n405( .i (n404), .o (n405) );
  assign n407 = n394 | n405 ;
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  assign n411 = N92 & n369 ;
  assign n412 = n296 & ~n411 ;
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  assign n414 = N79 & n369 ;
  assign n415 = n310 & ~n414 ;
  buffer buf_n416( .i (n415), .o (n416) );
  assign n418 = n413 | n416 ;
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n420( .i (n367), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  assign n422 = N105 & n421 ;
  assign n423 = n253 & ~n422 ;
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  assign n426 = N115 & n371 ;
  assign n427 = n361 & ~n426 ;
  assign n428 = n425 | n427 ;
  assign n429 = n419 | n428 ;
  assign n430 = n408 | n429 ;
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  assign n431 = N14 & n374 ;
  assign n432 = n283 & ~n431 ;
  assign n433 = n430 & ~n432 ;
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n406( .i (n405), .o (n406) );
  assign n434 = ~n406 & n419 ;
  assign n435 = n396 | n434 ;
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n417( .i (n416), .o (n417) );
  assign n437 = ~n405 & n417 ;
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  assign n438 = ~n413 & n424 ;
  assign n439 = n401 | n438 ;
  assign n440 = n437 | n439 ;
  assign n441 = ~n384 & n440 ;
  assign n442 = n392 | n441 ;
  assign N223 = n96 ;
  assign N329 = n232 ;
  assign N370 = n377 ;
  assign N421 = n433 ;
  assign N430 = n410 ;
  assign N431 = n436 ;
  assign N432 = n442 ;
endmodule
