module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( in_0_ , in_1_ , in_2_ , in_3_ , in_4_ , in_5_ , in_6_ , in_7_ , in_8_ , in_9_ , in_10_ , in_11_ , in_12_ , in_13_ , in_14_ , in_15_ , out_0_ , out_1_ , out_2_ , out_3_ , out_4_ );
  input in_0_ , in_1_ , in_2_ , in_3_ , in_4_ , in_5_ , in_6_ , in_7_ , in_8_ , in_9_ , in_10_ , in_11_ , in_12_ , in_13_ , in_14_ , in_15_ ;
  output out_0_ , out_1_ , out_2_ , out_3_ , out_4_ ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 ;
  assign n17 = in_14_ & in_15_ ;
  buffer buf_n18( .i (n17), .o (n18) );
  assign n19 = in_12_ | in_13_ ;
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  assign n23 = in_4_ | in_5_ ;
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  assign n27 = in_0_ | in_1_ ;
  buffer buf_n28( .i (n27), .o (n28) );
  assign n29 = in_2_ & in_3_ ;
  buffer buf_n30( .i (n29), .o (n30) );
  assign n31 = ( n24 & n28 ) | ( n24 & n30 ) | ( n28 & n30 ) ;
  buffer buf_n32( .i (n31), .o (n32) );
  assign n37 = ( ~n24 & n28 ) | ( ~n24 & n30 ) | ( n28 & n30 ) ;
  buffer buf_n38( .i (n37), .o (n38) );
  assign n39 = ( n26 & ~n32 ) | ( n26 & n38 ) | ( ~n32 & n38 ) ;
  buffer buf_n40( .i (n39), .o (n40) );
  assign n41 = in_10_ & in_11_ ;
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  assign n45 = in_6_ & in_7_ ;
  buffer buf_n46( .i (n45), .o (n46) );
  assign n47 = in_8_ | in_9_ ;
  buffer buf_n48( .i (n47), .o (n48) );
  assign n49 = ( n42 & n46 ) | ( n42 & n48 ) | ( n46 & n48 ) ;
  buffer buf_n50( .i (n49), .o (n50) );
  assign n55 = ( ~n42 & n46 ) | ( ~n42 & n48 ) | ( n46 & n48 ) ;
  buffer buf_n56( .i (n55), .o (n56) );
  assign n57 = ( n44 & ~n50 ) | ( n44 & n56 ) | ( ~n50 & n56 ) ;
  buffer buf_n58( .i (n57), .o (n58) );
  assign n59 = ( n20 & n40 ) | ( n20 & n58 ) | ( n40 & n58 ) ;
  buffer buf_n60( .i (n59), .o (n60) );
  assign n63 = ( ~n20 & n40 ) | ( ~n20 & n58 ) | ( n40 & n58 ) ;
  buffer buf_n64( .i (n63), .o (n64) );
  assign n65 = ( n22 & ~n60 ) | ( n22 & n64 ) | ( ~n60 & n64 ) ;
  buffer buf_n66( .i (n65), .o (n66) );
  assign n67 = n18 & n66 ;
  buffer buf_n68( .i (n67), .o (n68) );
  assign n69 = n18 | n66 ;
  buffer buf_n70( .i (n69), .o (n70) );
  assign n71 = ~n68 & n70 ;
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  assign n72 = ( n36 & n54 ) | ( n36 & n60 ) | ( n54 & n60 ) ;
  buffer buf_n73( .i (n72), .o (n73) );
  assign n78 = ( n36 & n54 ) | ( n36 & ~n60 ) | ( n54 & ~n60 ) ;
  buffer buf_n79( .i (n78), .o (n79) );
  assign n80 = ( n62 & ~n73 ) | ( n62 & n79 ) | ( ~n73 & n79 ) ;
  buffer buf_n81( .i (n80), .o (n81) );
  assign n82 = n68 & n81 ;
  buffer buf_n83( .i (n82), .o (n83) );
  assign n84 = n68 | n81 ;
  buffer buf_n85( .i (n84), .o (n85) );
  assign n86 = ~n83 & n85 ;
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  assign n87 = n77 & n83 ;
  buffer buf_n88( .i (n87), .o (n88) );
  assign n89 = n77 | n83 ;
  buffer buf_n90( .i (n89), .o (n90) );
  assign n91 = ~n88 & n90 ;
  assign out_0_ = 1'b0 ;
  assign out_1_ = n71 ;
  assign out_2_ = n86 ;
  assign out_3_ = n91 ;
  assign out_4_ = n88 ;
endmodule
