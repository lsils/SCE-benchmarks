module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 ;
  buffer buf_n125( .i (x5), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n78( .i (x3), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n31( .i (x1), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n145( .i (x6), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  assign n190 = ( n47 & ~n94 ) | ( n47 & n161 ) | ( ~n94 & n161 ) ;
  buffer buf_n54( .i (x2), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  assign n191 = n47 | n70 ;
  assign n192 = ( n95 & n190 ) | ( n95 & n191 ) | ( n190 & n191 ) ;
  assign n193 = n143 & ~n192 ;
  buffer buf_n48( .i (n47), .o (n48) );
  assign n194 = n90 & n157 ;
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  assign n205 = ( n70 & n161 ) | ( n70 & n197 ) | ( n161 & n197 ) ;
  assign n206 = n48 & n205 ;
  assign n207 = n143 | n206 ;
  assign n208 = ~n193 & n207 ;
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n165( .i (x7), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n71( .i (n70), .o (n71) );
  assign n211 = ( n69 & ~n140 ) | ( n69 & n160 ) | ( ~n140 & n160 ) ;
  buffer buf_n212( .i (n211), .o (n212) );
  assign n213 = ( ~n71 & n95 ) | ( ~n71 & n212 ) | ( n95 & n212 ) ;
  buffer buf_n162( .i (n161), .o (n162) );
  assign n214 = ( n95 & n162 ) | ( n95 & ~n212 ) | ( n162 & ~n212 ) ;
  assign n215 = n213 & ~n214 ;
  assign n216 = ( ~n50 & n184 ) | ( ~n50 & n215 ) | ( n184 & n215 ) ;
  assign n217 = ( n69 & n93 ) | ( n69 & n140 ) | ( n93 & n140 ) ;
  buffer buf_n218( .i (n217), .o (n218) );
  assign n219 = ( n71 & n162 ) | ( n71 & ~n218 ) | ( n162 & ~n218 ) ;
  buffer buf_n220( .i (n94), .o (n220) );
  assign n221 = ( n162 & n218 ) | ( n162 & ~n220 ) | ( n218 & ~n220 ) ;
  assign n222 = ~n219 & n221 ;
  assign n223 = ( n50 & n184 ) | ( n50 & n222 ) | ( n184 & n222 ) ;
  assign n224 = n216 & n223 ;
  assign n225 = ~n209 & n224 ;
  buffer buf_n9( .i (x0), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n103( .i (x4), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  assign n226 = n30 & n124 ;
  assign n227 = ( n210 & n225 ) | ( n210 & n226 ) | ( n225 & n226 ) ;
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  assign n230 = ( n42 & n65 ) | ( n42 & n136 ) | ( n65 & n136 ) ;
  buffer buf_n231( .i (n230), .o (n231) );
  assign n236 = ( n67 & n158 ) | ( n67 & ~n231 ) | ( n158 & ~n231 ) ;
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  assign n241 = ( n46 & n140 ) | ( n46 & ~n237 ) | ( n140 & ~n237 ) ;
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  assign n244 = ~n235 & n242 ;
  assign n245 = ( n240 & n243 ) | ( n240 & n244 ) | ( n243 & n244 ) ;
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  assign n248 = ( n29 & n123 ) | ( n29 & ~n246 ) | ( n123 & ~n246 ) ;
  assign n249 = n27 & ~n49 ;
  assign n250 = n49 & n143 ;
  assign n251 = ~n19 & n64 ;
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n142), .o (n259) );
  assign n260 = ~n258 & n259 ;
  assign n261 = ( n249 & n250 ) | ( n249 & ~n260 ) | ( n250 & ~n260 ) ;
  assign n262 = n123 & n261 ;
  assign n263 = ( n247 & n248 ) | ( n247 & n262 ) | ( n248 & n262 ) ;
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  assign n266 = ( ~n20 & n65 ) | ( ~n20 & n156 ) | ( n65 & n156 ) ;
  assign n267 = n19 & ~n155 ;
  assign n268 = ( n65 & n136 ) | ( n65 & ~n267 ) | ( n136 & ~n267 ) ;
  assign n269 = ~n266 & n268 ;
  assign n270 = n91 & ~n269 ;
  assign n271 = ~n135 & n155 ;
  buffer buf_n272( .i (n271), .o (n272) );
  assign n281 = n252 & n272 ;
  assign n282 = n91 | n281 ;
  assign n283 = ~n270 & n282 ;
  assign n284 = n118 & ~n283 ;
  assign n285 = ~n66 & n90 ;
  assign n286 = n136 & ~n156 ;
  buffer buf_n287( .i (n286), .o (n287) );
  assign n292 = ( n67 & n285 ) | ( n67 & n287 ) | ( n285 & n287 ) ;
  assign n293 = n23 & n292 ;
  assign n294 = n118 | n293 ;
  assign n295 = ~n284 & n294 ;
  assign n296 = n182 & n295 ;
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  assign n299 = ( n67 & n158 ) | ( n67 & ~n178 ) | ( n158 & ~n178 ) ;
  buffer buf_n300( .i (n299), .o (n300) );
  assign n301 = ( ~n69 & n93 ) | ( ~n69 & n300 ) | ( n93 & n300 ) ;
  assign n302 = ( n93 & n160 ) | ( n93 & ~n300 ) | ( n160 & ~n300 ) ;
  assign n303 = n301 & ~n302 ;
  assign n304 = ~n142 & n303 ;
  assign n305 = n121 & n304 ;
  assign n306 = n297 | n305 ;
  assign n307 = ( n29 & n298 ) | ( n29 & n306 ) | ( n298 & n306 ) ;
  assign n308 = n52 & ~n307 ;
  assign n309 = ( ~n91 & n116 ) | ( ~n91 & n178 ) | ( n116 & n178 ) ;
  buffer buf_n310( .i (n309), .o (n310) );
  assign n311 = ( n160 & ~n180 ) | ( n160 & n310 ) | ( ~n180 & n310 ) ;
  buffer buf_n312( .i (n159), .o (n312) );
  assign n313 = ( n118 & ~n310 ) | ( n118 & n312 ) | ( ~n310 & n312 ) ;
  assign n314 = n311 & ~n313 ;
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n72( .i (n71), .o (n72) );
  assign n317 = ( n72 & n259 ) | ( n72 & ~n315 ) | ( n259 & ~n315 ) ;
  assign n318 = n157 & ~n177 ;
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n117), .o (n321) );
  assign n322 = n320 & n321 ;
  assign n323 = ( n70 & n94 ) | ( n70 & n322 ) | ( n94 & n322 ) ;
  assign n324 = ~n71 & n323 ;
  assign n325 = n259 & n324 ;
  assign n326 = ( n316 & n317 ) | ( n316 & n325 ) | ( n317 & n325 ) ;
  assign n327 = n29 & n326 ;
  assign n328 = n52 | n327 ;
  assign n329 = ~n308 & n328 ;
  assign n330 = n138 & n158 ;
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  assign n336 = n28 & n335 ;
  assign n337 = ( n51 & n123 ) | ( n51 & n336 ) | ( n123 & n336 ) ;
  assign n338 = ~n124 & n337 ;
  buffer buf_n339( .i (n68), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  assign n341 = ( n141 & ~n161 ) | ( n141 & n340 ) | ( ~n161 & n340 ) ;
  assign n342 = n218 & ~n341 ;
  assign n343 = n49 & n342 ;
  assign n344 = n28 | n343 ;
  buffer buf_n96( .i (n95), .o (n96) );
  assign n345 = ( n38 & n61 ) | ( n38 & n152 ) | ( n61 & n152 ) ;
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  assign n350 = ( ~n137 & n157 ) | ( ~n137 & n349 ) | ( n157 & n349 ) ;
  buffer buf_n351( .i (n350), .o (n351) );
  assign n354 = n159 & ~n351 ;
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  assign n357 = n353 | n355 ;
  buffer buf_n358( .i (n312), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  assign n360 = ( n356 & n357 ) | ( n356 & ~n359 ) | ( n357 & ~n359 ) ;
  assign n361 = ~n96 & n360 ;
  assign n362 = n28 & ~n361 ;
  assign n363 = n344 & ~n362 ;
  assign n364 = ~n45 & n68 ;
  assign n365 = n24 & n364 ;
  assign n366 = n332 & n365 ;
  assign n367 = ( n120 & n220 ) | ( n120 & n366 ) | ( n220 & n366 ) ;
  assign n368 = ~n121 & n367 ;
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n122), .o (n371) );
  assign n372 = n369 | n371 ;
  assign n373 = ( n363 & n370 ) | ( n363 & n372 ) | ( n370 & n372 ) ;
  assign n374 = n338 | n373 ;
  assign n375 = ( ~n264 & n329 ) | ( ~n264 & n374 ) | ( n329 & n374 ) ;
  assign n376 = n265 | n375 ;
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  assign n377 = n155 & n175 ;
  buffer buf_n378( .i (n135), .o (n378) );
  assign n379 = n377 & ~n378 ;
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  assign n385 = ~n86 & n111 ;
  buffer buf_n386( .i (n385), .o (n386) );
  assign n390 = ~n111 & n133 ;
  buffer buf_n391( .i (n390), .o (n391) );
  assign n396 = ( n113 & ~n386 ) | ( n113 & n391 ) | ( ~n386 & n391 ) ;
  assign n397 = ( n156 & ~n176 ) | ( n156 & n396 ) | ( ~n176 & n396 ) ;
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n154), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  assign n404 = n398 & ~n403 ;
  assign n405 = ( n179 & n399 ) | ( n179 & n404 ) | ( n399 & n404 ) ;
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  assign n408 = n119 & ~n406 ;
  assign n409 = ( n384 & n407 ) | ( n384 & ~n408 ) | ( n407 & ~n408 ) ;
  assign n410 = n27 & n409 ;
  assign n411 = n178 & ~n403 ;
  assign n412 = n139 & n411 ;
  assign n413 = ~n321 & n412 ;
  buffer buf_n414( .i (n92), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  assign n416 = n413 & n415 ;
  assign n417 = ~n139 & n319 ;
  assign n418 = ( n321 & n414 ) | ( n321 & n417 ) | ( n414 & n417 ) ;
  assign n419 = ~n415 & n418 ;
  assign n420 = n416 | n419 ;
  assign n421 = ~n27 & n420 ;
  assign n422 = n410 | n421 ;
  assign n423 = ( n51 & ~n74 ) | ( n51 & n422 ) | ( ~n74 & n422 ) ;
  assign n424 = ( ~n21 & n115 ) | ( ~n21 & n177 ) | ( n115 & n177 ) ;
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  assign n427 = ( n312 & n321 ) | ( n312 & n426 ) | ( n321 & n426 ) ;
  assign n428 = ( n23 & ~n179 ) | ( n23 & n425 ) | ( ~n179 & n425 ) ;
  assign n429 = n117 & ~n425 ;
  assign n430 = ( ~n312 & n428 ) | ( ~n312 & n429 ) | ( n428 & n429 ) ;
  assign n431 = ( ~n119 & n427 ) | ( ~n119 & n430 ) | ( n427 & n430 ) ;
  assign n432 = ~n116 & n380 ;
  assign n433 = n23 & n432 ;
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  assign n436 = n141 | n434 ;
  assign n437 = ( n431 & n435 ) | ( n431 & n436 ) | ( n435 & n436 ) ;
  assign n438 = n96 & ~n437 ;
  buffer buf_n439( .i (n117), .o (n439) );
  buffer buf_n440( .i (n159), .o (n440) );
  assign n441 = ( n180 & n439 ) | ( n180 & ~n440 ) | ( n439 & ~n440 ) ;
  buffer buf_n442( .i (n139), .o (n442) );
  assign n443 = ( n180 & n439 ) | ( n180 & ~n442 ) | ( n439 & ~n442 ) ;
  assign n444 = ~n441 & n443 ;
  assign n445 = n26 & n444 ;
  assign n446 = n96 | n445 ;
  assign n447 = ~n438 & n446 ;
  assign n448 = ( n51 & n74 ) | ( n51 & n447 ) | ( n74 & n447 ) ;
  assign n449 = n423 & n448 ;
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n66), .o (n452) );
  assign n453 = n403 & n452 ;
  buffer buf_n454( .i (n453), .o (n454) );
  assign n457 = ( n439 & n442 ) | ( n439 & n454 ) | ( n442 & n454 ) ;
  buffer buf_n458( .i (n457), .o (n458) );
  assign n459 = n120 | n458 ;
  assign n460 = n120 & n458 ;
  assign n461 = n459 & ~n460 ;
  buffer buf_n462( .i (n26), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  assign n464 = n461 | n463 ;
  buffer buf_n465( .i (n116), .o (n465) );
  buffer buf_n466( .i (n138), .o (n466) );
  assign n467 = n465 & ~n466 ;
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  assign n470 = ~n359 & n469 ;
  assign n471 = ~n72 & n470 ;
  assign n472 = n463 & ~n471 ;
  assign n473 = n464 & ~n472 ;
  assign n474 = n52 & ~n473 ;
  buffer buf_n144( .i (n143), .o (n144) );
  assign n475 = n465 & n466 ;
  buffer buf_n476( .i (n475), .o (n476) );
  assign n479 = ( n340 & n358 ) | ( n340 & n476 ) | ( n358 & n476 ) ;
  buffer buf_n480( .i (n479), .o (n480) );
  assign n481 = ~n259 & n480 ;
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  assign n482 = ( ~n121 & n478 ) | ( ~n121 & n480 ) | ( n478 & n480 ) ;
  assign n483 = ( n144 & n481 ) | ( n144 & ~n482 ) | ( n481 & ~n482 ) ;
  buffer buf_n484( .i (n463), .o (n484) );
  assign n485 = n483 & n484 ;
  buffer buf_n486( .i (n50), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  assign n488 = n485 | n487 ;
  assign n489 = ~n474 & n488 ;
  assign n490 = ~n63 & n174 ;
  assign n491 = ( n135 & ~n400 ) | ( n135 & n490 ) | ( ~n400 & n490 ) ;
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  assign n495 = ( n66 & n402 ) | ( n66 & n492 ) | ( n402 & n492 ) ;
  buffer buf_n496( .i (n177), .o (n496) );
  assign n497 = ( n138 & ~n495 ) | ( n138 & n496 ) | ( ~n495 & n496 ) ;
  assign n498 = ~n494 & n497 ;
  assign n499 = n439 & ~n498 ;
  assign n500 = n68 & n381 ;
  buffer buf_n501( .i (n465), .o (n501) );
  assign n502 = n500 | n501 ;
  assign n503 = ~n499 & n502 ;
  assign n504 = n220 & ~n503 ;
  assign n505 = n114 & ~n401 ;
  assign n506 = n114 | n401 ;
  assign n507 = ( ~n115 & n505 ) | ( ~n115 & n506 ) | ( n505 & n506 ) ;
  buffer buf_n508( .i (n507), .o (n508) );
  assign n518 = n466 & n508 ;
  buffer buf_n519( .i (n179), .o (n519) );
  assign n520 = n518 & ~n519 ;
  assign n521 = n340 & n520 ;
  assign n522 = n220 | n521 ;
  assign n523 = ~n504 & n522 ;
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  assign n526 = ( ~n484 & n486 ) | ( ~n484 & n524 ) | ( n486 & n524 ) ;
  assign n527 = n339 & n414 ;
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n119), .o (n531) );
  assign n532 = n384 & n531 ;
  assign n533 = ~n462 & n532 ;
  assign n534 = n530 & n533 ;
  assign n535 = ~n486 & n534 ;
  assign n536 = ( n525 & ~n526 ) | ( n525 & n535 ) | ( ~n526 & n535 ) ;
  buffer buf_n537( .i (n403), .o (n537) );
  assign n538 = n92 | n537 ;
  assign n539 = n442 | n538 ;
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n64), .o (n542) );
  assign n543 = n20 & n542 ;
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  assign n551 = ( n48 & n540 ) | ( n48 & n548 ) | ( n540 & n548 ) ;
  assign n552 = ~n541 & n551 ;
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  assign n555 = ( n21 & ~n90 ) | ( n21 & n402 ) | ( ~n90 & n402 ) ;
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n559( .i (n542), .o (n559) );
  buffer buf_n560( .i (n89), .o (n560) );
  assign n561 = n559 | n560 ;
  buffer buf_n562( .i (n561), .o (n562) );
  assign n566 = ( ~n537 & n556 ) | ( ~n537 & n562 ) | ( n556 & n562 ) ;
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  assign n569 = ( n340 & n558 ) | ( n340 & ~n567 ) | ( n558 & ~n567 ) ;
  assign n570 = ( n359 & n568 ) | ( n359 & ~n569 ) | ( n568 & ~n569 ) ;
  buffer buf_n571( .i (n48), .o (n571) );
  buffer buf_n572( .i (n142), .o (n572) );
  assign n573 = ( n570 & n571 ) | ( n570 & ~n572 ) | ( n571 & ~n572 ) ;
  assign n574 = n25 & ~n415 ;
  buffer buf_n575( .i (n402), .o (n575) );
  assign n576 = ~n452 & n575 ;
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  assign n579 = n25 & ~n578 ;
  assign n580 = ( n528 & n574 ) | ( n528 & ~n579 ) | ( n574 & ~n579 ) ;
  assign n581 = ( n571 & n572 ) | ( n571 & n580 ) | ( n572 & n580 ) ;
  assign n582 = ~n573 & n581 ;
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  assign n583 = ( n92 & n395 ) | ( n92 & ~n537 ) | ( n395 & ~n537 ) ;
  assign n584 = ~n414 & n583 ;
  assign n585 = n25 & n584 ;
  buffer buf_n586( .i (n47), .o (n586) );
  buffer buf_n587( .i (n339), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  assign n589 = ( n585 & n586 ) | ( n585 & n588 ) | ( n586 & n588 ) ;
  assign n590 = ~n72 & n589 ;
  buffer buf_n591( .i (n590), .o (n591) );
  assign n592 = ( ~n553 & n582 ) | ( ~n553 & n591 ) | ( n582 & n591 ) ;
  assign n593 = n371 | n591 ;
  assign n594 = ( n554 & n592 ) | ( n554 & n593 ) | ( n592 & n593 ) ;
  assign n595 = n536 | n594 ;
  assign n596 = ( ~n450 & n489 ) | ( ~n450 & n595 ) | ( n489 & n595 ) ;
  assign n597 = n451 | n596 ;
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n598( .i (n415), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  assign n600 = n278 & ~n599 ;
  assign n601 = ~n122 & n600 ;
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  assign n604 = n44 & n253 ;
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  assign n612 = n602 & ~n611 ;
  buffer buf_n613( .i (n401), .o (n613) );
  assign n614 = n43 & n613 ;
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n560), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  assign n620 = ( n442 & n616 ) | ( n442 & n619 ) | ( n616 & n619 ) ;
  assign n621 = ( n45 & ~n615 ) | ( n45 & n618 ) | ( ~n615 & n618 ) ;
  buffer buf_n622( .i (n466), .o (n622) );
  assign n623 = ( n440 & n621 ) | ( n440 & n622 ) | ( n621 & n622 ) ;
  assign n624 = ~n620 & n623 ;
  assign n625 = n588 & ~n624 ;
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  assign n626 = ~n537 & n618 ;
  buffer buf_n627( .i (n137), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  assign n629 = ~n618 & n628 ;
  assign n630 = ( ~n289 & n626 ) | ( ~n289 & n629 ) | ( n626 & n629 ) ;
  buffer buf_n631( .i (n46), .o (n631) );
  assign n632 = n630 & n631 ;
  assign n633 = n588 | n632 ;
  assign n634 = ~n625 & n633 ;
  assign n635 = ( ~n122 & n463 ) | ( ~n122 & n634 ) | ( n463 & n634 ) ;
  assign n636 = ( n46 & n339 ) | ( n46 & ~n622 ) | ( n339 & ~n622 ) ;
  buffer buf_n637( .i (n636), .o (n637) );
  assign n639 = ( n359 & n588 ) | ( n359 & ~n637 ) | ( n588 & ~n637 ) ;
  buffer buf_n640( .i (n358), .o (n640) );
  assign n641 = ( ~n586 & n637 ) | ( ~n586 & n640 ) | ( n637 & n640 ) ;
  assign n642 = n639 & ~n641 ;
  buffer buf_n643( .i (n462), .o (n643) );
  buffer buf_n644( .i (n531), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  assign n646 = ( n642 & n643 ) | ( n642 & n645 ) | ( n643 & n645 ) ;
  assign n647 = n635 & n646 ;
  assign n648 = ( n196 & n501 ) | ( n196 & n605 ) | ( n501 & n605 ) ;
  buffer buf_n649( .i (n501), .o (n649) );
  assign n650 = n648 & ~n649 ;
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  assign n654 = ( n42 & n89 ) | ( n42 & ~n542 ) | ( n89 & ~n542 ) ;
  assign n655 = ( n43 & ~n613 ) | ( n43 & n654 ) | ( ~n613 & n654 ) ;
  buffer buf_n656( .i (n655), .o (n656) );
  assign n659 = n45 & ~n656 ;
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  assign n662 = n658 | n660 ;
  assign n663 = ( ~n586 & n661 ) | ( ~n586 & n662 ) | ( n661 & n662 ) ;
  assign n664 = ( n462 & n651 ) | ( n462 & n663 ) | ( n651 & n663 ) ;
  assign n665 = n645 & ~n664 ;
  assign n666 = ( n371 & n653 ) | ( n371 & ~n665 ) | ( n653 & ~n665 ) ;
  assign n667 = n647 | n666 ;
  assign n668 = ( n603 & ~n612 ) | ( n603 & n667 ) | ( ~n612 & n667 ) ;
  assign n669 = ( ~n452 & n575 ) | ( ~n452 & n627 ) | ( n575 & n627 ) ;
  buffer buf_n670( .i (n669), .o (n670) );
  assign n671 = ( ~n440 & n501 ) | ( ~n440 & n670 ) | ( n501 & n670 ) ;
  buffer buf_n672( .i (n465), .o (n672) );
  assign n673 = ( n622 & ~n670 ) | ( n622 & n672 ) | ( ~n670 & n672 ) ;
  assign n674 = n671 & ~n673 ;
  assign n675 = ( ~n586 & n598 ) | ( ~n586 & n674 ) | ( n598 & n674 ) ;
  buffer buf_n676( .i (n115), .o (n676) );
  assign n677 = ( n452 & n627 ) | ( n452 & n676 ) | ( n627 & n676 ) ;
  buffer buf_n678( .i (n677), .o (n678) );
  assign n679 = ( n440 & n672 ) | ( n440 & ~n678 ) | ( n672 & ~n678 ) ;
  buffer buf_n680( .i (n575), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  assign n682 = ( ~n622 & n678 ) | ( ~n622 & n681 ) | ( n678 & n681 ) ;
  assign n683 = ~n679 & n682 ;
  buffer buf_n684( .i (n631), .o (n684) );
  assign n685 = ( n598 & n683 ) | ( n598 & n684 ) | ( n683 & n684 ) ;
  assign n686 = n675 & n685 ;
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  assign n689 = n484 & n687 ;
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  assign n690 = ( n20 & n378 ) | ( n20 & n542 ) | ( n378 & n542 ) ;
  assign n691 = ( ~n43 & n137 ) | ( ~n43 & n690 ) | ( n137 & n690 ) ;
  buffer buf_n692( .i (n691), .o (n692) );
  assign n695 = n628 & ~n692 ;
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  assign n698 = n694 | n696 ;
  buffer buf_n699( .i (n141), .o (n699) );
  assign n700 = ( n697 & n698 ) | ( n697 & ~n699 ) | ( n698 & ~n699 ) ;
  assign n701 = ( n512 & n599 ) | ( n512 & ~n700 ) | ( n599 & ~n700 ) ;
  buffer buf_n702( .i (n134), .o (n702) );
  assign n703 = n64 & n702 ;
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n559), .o (n707) );
  assign n708 = ( n676 & n705 ) | ( n676 & n707 ) | ( n705 & n707 ) ;
  buffer buf_n709( .i (n114), .o (n709) );
  buffer buf_n710( .i (n378), .o (n710) );
  assign n711 = ( n21 & ~n709 ) | ( n21 & n710 ) | ( ~n709 & n710 ) ;
  buffer buf_n712( .i (n19), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  assign n714 = ( n704 & ~n710 ) | ( n704 & n713 ) | ( ~n710 & n713 ) ;
  assign n715 = n711 & ~n714 ;
  assign n716 = ( ~n706 & n708 ) | ( ~n706 & n715 ) | ( n708 & n715 ) ;
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  assign n719 = ( n358 & ~n631 ) | ( n358 & n717 ) | ( ~n631 & n717 ) ;
  buffer buf_n720( .i (n22), .o (n720) );
  buffer buf_n721( .i (n676), .o (n721) );
  assign n722 = ~n720 & n721 ;
  assign n723 = n331 & n722 ;
  assign n724 = n631 & n723 ;
  assign n725 = ( n718 & ~n719 ) | ( n718 & n724 ) | ( ~n719 & n724 ) ;
  assign n726 = ~n599 & n725 ;
  assign n727 = ( n513 & ~n701 ) | ( n513 & n726 ) | ( ~n701 & n726 ) ;
  assign n728 = ~n575 & n707 ;
  buffer buf_n729( .i (n728), .o (n729) );
  assign n731 = n672 & n729 ;
  buffer buf_n732( .i (n42), .o (n732) );
  assign n733 = n713 & n732 ;
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n737( .i (n44), .o (n737) );
  assign n738 = ~n734 & n737 ;
  buffer buf_n739( .i (n738), .o (n739) );
  assign n740 = n731 & n739 ;
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  assign n741 = n577 & ~n672 ;
  assign n742 = ( ~n736 & n739 ) | ( ~n736 & n741 ) | ( n739 & n741 ) ;
  assign n743 = ( n26 & n740 ) | ( n26 & n742 ) | ( n740 & n742 ) ;
  assign n744 = n599 & ~n743 ;
  assign n745 = ~n544 & n707 ;
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n721), .o (n747) );
  assign n748 = n746 & n747 ;
  assign n749 = ( ~n546 & n681 ) | ( ~n546 & n746 ) | ( n681 & n746 ) ;
  buffer buf_n750( .i (n24), .o (n750) );
  assign n751 = ( n748 & n749 ) | ( n748 & n750 ) | ( n749 & n750 ) ;
  assign n752 = ~n684 & n751 ;
  buffer buf_n753( .i (n598), .o (n753) );
  assign n754 = n752 | n753 ;
  assign n755 = ~n744 & n754 ;
  assign n756 = n727 | n755 ;
  assign n757 = ( n688 & ~n689 ) | ( n688 & n756 ) | ( ~n689 & n756 ) ;
  buffer buf_n758( .i (n757), .o (n758) );
  assign n759 = ( n188 & n668 ) | ( n188 & n758 ) | ( n668 & n758 ) ;
  buffer buf_n638( .i (n637), .o (n638) );
  assign n760 = n638 | n753 ;
  buffer buf_n761( .i (n587), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  assign n763 = ( n638 & n753 ) | ( n638 & ~n762 ) | ( n753 & ~n762 ) ;
  assign n764 = ( n73 & ~n760 ) | ( n73 & n763 ) | ( ~n760 & n763 ) ;
  assign n765 = n484 & ~n764 ;
  buffer buf_n766( .i (n628), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  assign n768 = ~n587 & n767 ;
  buffer buf_n769( .i (n619), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  assign n771 = n768 & n770 ;
  assign n772 = n571 & n771 ;
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n643), .o (n774) );
  assign n775 = n773 | n774 ;
  assign n776 = ~n765 & n775 ;
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  assign n777 = ( n57 & ~n106 ) | ( n57 & n128 ) | ( ~n106 & n128 ) ;
  buffer buf_n778( .i (n777), .o (n778) );
  assign n783 = ( n83 & ~n130 ) | ( n83 & n778 ) | ( ~n130 & n778 ) ;
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  assign n788 = ( n61 & ~n110 ) | ( n61 & n784 ) | ( ~n110 & n784 ) ;
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  assign n791 = ~n782 & n789 ;
  assign n792 = ( ~n787 & n790 ) | ( ~n787 & n791 ) | ( n790 & n791 ) ;
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  assign n795 = ( n613 & n732 ) | ( n613 & ~n793 ) | ( n732 & ~n793 ) ;
  assign n796 = n88 & n113 ;
  assign n797 = n113 | n702 ;
  assign n798 = n40 & ~n87 ;
  assign n799 = n702 | n798 ;
  assign n800 = ( n796 & ~n797 ) | ( n796 & n799 ) | ( ~n797 & n799 ) ;
  assign n801 = n613 & n800 ;
  assign n802 = ( n794 & n795 ) | ( n794 & n801 ) | ( n795 & n801 ) ;
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  assign n806 = ( n63 & n112 ) | ( n63 & ~n154 ) | ( n112 & ~n154 ) ;
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n112), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  assign n813 = n807 & ~n812 ;
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  assign n816 = ( n617 & ~n707 ) | ( n617 & n814 ) | ( ~n707 & n814 ) ;
  assign n817 = ( n810 & n815 ) | ( n810 & n816 ) | ( n815 & n816 ) ;
  buffer buf_n818( .i (n737), .o (n818) );
  assign n819 = ( n803 & n817 ) | ( n803 & n818 ) | ( n817 & n818 ) ;
  assign n820 = n767 & ~n819 ;
  assign n821 = ( n699 & n805 ) | ( n699 & ~n820 ) | ( n805 & ~n820 ) ;
  buffer buf_n822( .i (n750), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  assign n824 = n821 & n823 ;
  assign n825 = ( n87 & n134 ) | ( n87 & n154 ) | ( n134 & n154 ) ;
  assign n826 = ( n400 & ~n811 ) | ( n400 & n825 ) | ( ~n811 & n825 ) ;
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n830( .i (n400), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  assign n832 = ~n827 & n831 ;
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  assign n835 = n829 | n833 ;
  assign n836 = ( ~n681 & n834 ) | ( ~n681 & n835 ) | ( n834 & n835 ) ;
  buffer buf_n837( .i (n818), .o (n837) );
  assign n838 = ~n836 & n837 ;
  assign n839 = n273 & n676 ;
  buffer buf_n840( .i (n839), .o (n840) );
  assign n844 = n619 & n840 ;
  assign n845 = n837 | n844 ;
  assign n846 = ~n838 & n845 ;
  assign n847 = ( n762 & n823 ) | ( n762 & n846 ) | ( n823 & n846 ) ;
  assign n848 = ( ~n550 & n824 ) | ( ~n550 & n847 ) | ( n824 & n847 ) ;
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  assign n851 = n515 | n849 ;
  assign n852 = ( n776 & n850 ) | ( n776 & n851 ) | ( n850 & n851 ) ;
  assign n853 = ( ~n188 & n758 ) | ( ~n188 & n852 ) | ( n758 & n852 ) ;
  assign n854 = n759 | n853 ;
  assign n855 = ( n44 & n617 ) | ( n44 & n627 ) | ( n617 & n627 ) ;
  buffer buf_n856( .i (n559), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  assign n858 = ( n628 & n855 ) | ( n628 & ~n857 ) | ( n855 & ~n857 ) ;
  buffer buf_n859( .i (n858), .o (n859) );
  assign n862 = n767 & ~n859 ;
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  assign n865 = n861 | n863 ;
  assign n866 = ( ~n144 & n864 ) | ( ~n144 & n865 ) | ( n864 & n865 ) ;
  assign n867 = n774 | n866 ;
  assign n868 = ~n773 & n774 ;
  assign n869 = n867 & ~n868 ;
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  assign n872 = ~n517 & n870 ;
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n873( .i (n710), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  assign n875 = n857 & ~n874 ;
  buffer buf_n876( .i (n875), .o (n876) );
  assign n877 = ( n750 & n769 ) | ( n750 & n876 ) | ( n769 & n876 ) ;
  assign n878 = ~n770 & n877 ;
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  assign n879 = n750 & n769 ;
  buffer buf_n880( .i (n857), .o (n880) );
  assign n881 = ~n747 & n880 ;
  buffer buf_n882( .i (n24), .o (n882) );
  assign n883 = ~n881 & n882 ;
  assign n884 = ( n565 & ~n879 ) | ( n565 & n883 ) | ( ~n879 & n883 ) ;
  assign n885 = ~n878 & n884 ;
  assign n886 = n164 & n885 ;
  assign n887 = ( n378 & ~n712 ) | ( n378 & n812 ) | ( ~n712 & n812 ) ;
  buffer buf_n888( .i (n887), .o (n888) );
  assign n892 = ( n617 & ~n873 ) | ( n617 & n888 ) | ( ~n873 & n888 ) ;
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n896( .i (n720), .o (n896) );
  assign n897 = ( n766 & n893 ) | ( n766 & n896 ) | ( n893 & n896 ) ;
  assign n898 = n891 & ~n897 ;
  assign n899 = ( n770 & ~n895 ) | ( n770 & n898 ) | ( ~n895 & n898 ) ;
  assign n900 = n762 & n899 ;
  assign n901 = n164 | n900 ;
  assign n902 = ~n886 & n901 ;
  assign n903 = n487 & n902 ;
  buffer buf_n904( .i (n709), .o (n904) );
  buffer buf_n905( .i (n831), .o (n905) );
  assign n906 = n904 & n905 ;
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  assign n907 = ( n389 & n856 ) | ( n389 & n904 ) | ( n856 & n904 ) ;
  assign n908 = ( n810 & n906 ) | ( n810 & ~n907 ) | ( n906 & ~n907 ) ;
  assign n909 = n766 & n908 ;
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n730( .i (n729), .o (n730) );
  assign n912 = ( n468 & ~n587 ) | ( n468 & n730 ) | ( ~n587 & n730 ) ;
  assign n913 = n910 | n912 ;
  assign n914 = ( n753 & n911 ) | ( n753 & n913 ) | ( n911 & n913 ) ;
  assign n915 = n643 | n914 ;
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  assign n916 = n529 & n843 ;
  assign n917 = n643 & ~n916 ;
  assign n918 = n915 & ~n917 ;
  assign n919 = n487 | n918 ;
  assign n920 = ( ~n53 & n903 ) | ( ~n53 & n919 ) | ( n903 & n919 ) ;
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  assign n921 = ( n289 & ~n766 ) | ( n289 & n880 ) | ( ~n766 & n880 ) ;
  assign n922 = n837 | n921 ;
  assign n923 = ( n291 & n640 ) | ( n291 & n922 ) | ( n640 & n922 ) ;
  assign n924 = n823 & ~n923 ;
  buffer buf_n925( .i (n41), .o (n925) );
  buffer buf_n926( .i (n702), .o (n926) );
  assign n927 = ( n830 & n925 ) | ( n830 & n926 ) | ( n925 & n926 ) ;
  assign n928 = ( ~n559 & n831 ) | ( ~n559 & n927 ) | ( n831 & n927 ) ;
  buffer buf_n929( .i (n928), .o (n929) );
  assign n932 = n680 & ~n929 ;
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  assign n935 = n931 | n933 ;
  assign n936 = ( ~n640 & n934 ) | ( ~n640 & n935 ) | ( n934 & n935 ) ;
  assign n937 = n823 | n936 ;
  buffer buf_n938( .i (n822), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  assign n940 = ( n924 & n937 ) | ( n924 & ~n939 ) | ( n937 & ~n939 ) ;
  assign n941 = ( n63 & ~n134 ) | ( n63 & n346 ) | ( ~n134 & n346 ) ;
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n945( .i (n62), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  assign n948 = ~n942 & n947 ;
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  assign n951 = n944 | n949 ;
  assign n952 = ( ~n857 & n950 ) | ( ~n857 & n951 ) | ( n950 & n951 ) ;
  assign n953 = n896 & n952 ;
  assign n954 = ( n856 & n873 ) | ( n856 & n905 ) | ( n873 & n905 ) ;
  assign n955 = n737 & n954 ;
  assign n956 = n896 | n955 ;
  assign n957 = ( ~n882 & n953 ) | ( ~n882 & n956 ) | ( n953 & n956 ) ;
  assign n958 = ( ~n182 & n531 ) | ( ~n182 & n957 ) | ( n531 & n957 ) ;
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  assign n961 = ( n184 & ~n645 ) | ( n184 & n959 ) | ( ~n645 & n959 ) ;
  assign n962 = ( n940 & n960 ) | ( n940 & n961 ) | ( n960 & n961 ) ;
  assign n963 = n99 & n962 ;
  buffer buf_n964( .i (n496), .o (n964) );
  assign n965 = ( n680 & n874 ) | ( n680 & n964 ) | ( n874 & n964 ) ;
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n874), .o (n967) );
  assign n968 = ( n519 & n896 ) | ( n519 & n967 ) | ( n896 & n967 ) ;
  buffer buf_n969( .i (n720), .o (n969) );
  assign n970 = n681 & ~n969 ;
  assign n971 = ( ~n966 & n968 ) | ( ~n966 & n970 ) | ( n968 & n970 ) ;
  assign n972 = n761 & ~n971 ;
  assign n973 = n496 | n905 ;
  assign n974 = ( n319 & ~n680 ) | ( n319 & n973 ) | ( ~n680 & n973 ) ;
  buffer buf_n975( .i (n974), .o (n975) );
  assign n976 = n882 & n975 ;
  assign n977 = n761 | n976 ;
  assign n978 = ~n972 & n977 ;
  buffer buf_n979( .i (n571), .o (n979) );
  assign n980 = ~n978 & n979 ;
  buffer buf_n981( .i (n880), .o (n981) );
  assign n982 = ( n181 & n876 ) | ( n181 & n981 ) | ( n876 & n981 ) ;
  assign n983 = ( n181 & n876 ) | ( n181 & ~n981 ) | ( n876 & ~n981 ) ;
  assign n984 = ( n761 & ~n982 ) | ( n761 & n983 ) | ( ~n982 & n983 ) ;
  assign n985 = n938 & n984 ;
  assign n986 = n979 | n985 ;
  assign n987 = ~n980 & n986 ;
  assign n988 = n99 | n987 ;
  assign n989 = ( ~n100 & n963 ) | ( ~n100 & n988 ) | ( n963 & n988 ) ;
  assign n990 = n920 | n989 ;
  assign n991 = ( n871 & ~n872 ) | ( n871 & n990 ) | ( ~n872 & n990 ) ;
  buffer buf_n455( .i (n454), .o (n455) );
  assign n992 = n455 | n769 ;
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n456( .i (n455), .o (n456) );
  assign n995 = ( n456 & ~n699 ) | ( n456 & n770 ) | ( ~n699 & n770 ) ;
  assign n996 = n993 & ~n995 ;
  assign n997 = ( ~n97 & n994 ) | ( ~n97 & n996 ) | ( n994 & n996 ) ;
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  assign n1000 = n487 & n998 ;
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n1001( .i (n684), .o (n1001) );
  buffer buf_n1002( .i (n619), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  assign n1005 = n1001 & n1004 ;
  assign n1006 = ( n73 & ~n279 ) | ( n73 & n1005 ) | ( ~n279 & n1005 ) ;
  assign n1007 = n280 & n1006 ;
  assign n1008 = ( n519 & n818 ) | ( n519 & n967 ) | ( n818 & n967 ) ;
  buffer buf_n1009( .i (n905), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  assign n1011 = ~n818 & n1010 ;
  assign n1012 = ( ~n966 & n1008 ) | ( ~n966 & n1011 ) | ( n1008 & n1011 ) ;
  assign n1013 = n1003 & ~n1012 ;
  assign n1014 = n837 & n975 ;
  assign n1015 = n1003 | n1014 ;
  assign n1016 = ~n1013 & n1015 ;
  assign n1017 = n73 & ~n1016 ;
  buffer buf_n1018( .i (n560), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  assign n1020 = ~n874 & n1019 ;
  buffer buf_n1021( .i (n1020), .o (n1021) );
  assign n1022 = ( n181 & n1002 ) | ( n181 & n1021 ) | ( n1002 & n1021 ) ;
  buffer buf_n1023( .i (n519), .o (n1023) );
  assign n1024 = ( ~n1002 & n1021 ) | ( ~n1002 & n1023 ) | ( n1021 & n1023 ) ;
  assign n1025 = ( n1003 & ~n1022 ) | ( n1003 & n1024 ) | ( ~n1022 & n1024 ) ;
  assign n1026 = n1001 & n1025 ;
  buffer buf_n1027( .i (n762), .o (n1027) );
  assign n1028 = n1026 | n1027 ;
  assign n1029 = ~n1017 & n1028 ;
  assign n1030 = n1007 | n1029 ;
  assign n1031 = ( n999 & ~n1000 ) | ( n999 & n1030 ) | ( ~n1000 & n1030 ) ;
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  assign n1034 = n188 | n204 ;
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  assign n1035 = n77 & ~n204 ;
  buffer buf_n1036( .i (n187), .o (n1036) );
  assign n1037 = ( n77 & ~n204 ) | ( n77 & n1036 ) | ( ~n204 & n1036 ) ;
  assign n1038 = ( n1034 & n1035 ) | ( n1034 & ~n1037 ) | ( n1035 & ~n1037 ) ;
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n189( .i (n188), .o (n189) );
  assign n1039 = n102 & n189 ;
  assign y0 = n229 ;
  assign y1 = n376 ;
  assign y2 = n597 ;
  assign y3 = n854 ;
  assign y4 = n991 ;
  assign y5 = n1033 ;
  assign y6 = n1038 ;
  assign y7 = n1039 ;
endmodule
