module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 ;
  wire n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 ;
  buffer buf_n735( .i (x28), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n685( .i (x26), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n542( .i (x21), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n457( .i (x18), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n485( .i (x19), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  assign n1211 = ~n470 & n498 ;
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  assign n1224 = n562 & n1217 ;
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  assign n1229 = n708 & n1226 ;
  buffer buf_n763( .i (x29), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n793( .i (x30), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  assign n1230 = ~n782 & n812 ;
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  assign n1239 = ( n759 & n1229 ) | ( n759 & n1234 ) | ( n1229 & n1234 ) ;
  assign n1240 = ~n760 & n1239 ;
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n1247( .i (n1246), .o (n1247) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n46( .i (x0), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  assign n1248 = ~n67 & n478 ;
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n512( .i (x20), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  assign n1251 = ~n527 & n557 ;
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  assign n1259 = ( n508 & n1249 ) | ( n508 & n1258 ) | ( n1249 & n1258 ) ;
  assign n1260 = ~n509 & n1259 ;
  assign n1261 = ( n760 & n1235 ) | ( n760 & n1260 ) | ( n1235 & n1260 ) ;
  assign n1262 = ~n761 & n1261 ;
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  assign n1268 = n503 & n560 ;
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  assign n1273 = ( n535 & ~n1249 ) | ( n535 & n1272 ) | ( ~n1249 & n1272 ) ;
  assign n1274 = n1250 & n1273 ;
  buffer buf_n629( .i (x24), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  assign n1275 = n651 & n815 ;
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  assign n1278 = ( n788 & n1274 ) | ( n788 & n1277 ) | ( n1274 & n1277 ) ;
  assign n1279 = ~n789 & n1278 ;
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n292( .i (x10), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  assign n1284 = n312 & n562 ;
  assign n1285 = ( n478 & n506 ) | ( n478 & n1284 ) | ( n506 & n1284 ) ;
  assign n1286 = ~n479 & n1285 ;
  buffer buf_n655( .i (x25), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  assign n1287 = n677 & ~n785 ;
  assign n1288 = ( n758 & n1286 ) | ( n758 & n1287 ) | ( n1286 & n1287 ) ;
  assign n1289 = ~n759 & n1288 ;
  assign n1290 = n818 & n1289 ;
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  assign n1296 = n654 & n1228 ;
  assign n1297 = ( n761 & n1236 ) | ( n761 & n1296 ) | ( n1236 & n1296 ) ;
  assign n1298 = ~n762 & n1297 ;
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  assign n1301 = ~n471 & n526 ;
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  assign n1311 = ( n68 & ~n507 ) | ( n68 & n1308 ) | ( ~n507 & n1308 ) ;
  assign n1312 = ~n69 & n1311 ;
  assign n1313 = n566 & n1312 ;
  assign n1314 = ( n654 & n788 ) | ( n654 & n1313 ) | ( n788 & n1313 ) ;
  assign n1315 = ~n789 & n1314 ;
  assign n1316 = n820 & n1315 ;
  buffer buf_n1317( .i (n1316), .o (n1317) );
  assign n1318 = n1299 | n1317 ;
  assign n1319 = n1294 | n1318 ;
  assign n1320 = n1283 | n1319 ;
  assign n1321 = ( ~n1246 & n1267 ) | ( ~n1246 & n1320 ) | ( n1267 & n1320 ) ;
  assign n1322 = n1247 | n1321 ;
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  assign n1328 = n1281 | n1317 ;
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  assign n1338 = n1241 | n1291 ;
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  assign n1350 = n1242 | n1280 ;
  assign n1351 = n1299 | n1350 ;
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  assign n1361 = ~n498 & n525 ;
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  assign n1373 = ( n65 & n476 ) | ( n65 & n1366 ) | ( n476 & n1366 ) ;
  assign n1374 = ~n477 & n1373 ;
  buffer buf_n1375( .i (n1374), .o (n1375) );
  assign n1376 = n564 & n1375 ;
  buffer buf_n1377( .i (n1376), .o (n1377) );
  assign n1379 = ( n787 & n1276 ) | ( n787 & n1377 ) | ( n1276 & n1377 ) ;
  assign n1380 = ~n788 & n1379 ;
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  assign n1386 = n63 & n502 ;
  buffer buf_n1387( .i (n1386), .o (n1387) );
  assign n1391 = n476 & n1387 ;
  buffer buf_n1392( .i (n1391), .o (n1392) );
  assign n1393 = n533 & n1392 ;
  assign n1394 = n561 & n812 ;
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  assign n1399 = ( n785 & n1393 ) | ( n785 & n1396 ) | ( n1393 & n1396 ) ;
  assign n1400 = ~n786 & n1399 ;
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  assign n1409 = n61 & ~n500 ;
  buffer buf_n1410( .i (n1409), .o (n1410) );
  assign n1416 = n474 & n1410 ;
  assign n1417 = ~n753 & n1416 ;
  assign n1418 = ( n531 & n561 ) | ( n531 & n1417 ) | ( n561 & n1417 ) ;
  assign n1419 = ~n532 & n1418 ;
  assign n1420 = n1231 & n1419 ;
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n480( .i (n479), .o (n480) );
  assign n1429 = n67 & n563 ;
  assign n1430 = ( n479 & n507 ) | ( n479 & n1429 ) | ( n507 & n1429 ) ;
  assign n1431 = ~n480 & n1430 ;
  assign n1432 = n754 & n812 ;
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  assign n1439 = ( n787 & n1431 ) | ( n787 & n1436 ) | ( n1431 & n1436 ) ;
  buffer buf_n1440( .i (n787), .o (n1440) );
  assign n1441 = n1439 & ~n1440 ;
  buffer buf_n1442( .i (n1441), .o (n1442) );
  assign n1449 = n1425 | n1442 ;
  assign n1450 = ( ~n1382 & n1404 ) | ( ~n1382 & n1449 ) | ( n1404 & n1449 ) ;
  assign n1451 = n1383 | n1450 ;
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  buffer buf_n1455( .i (n1454), .o (n1455) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n318( .i (x11), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  assign n1461 = n308 & n473 ;
  buffer buf_n1462( .i (n1461), .o (n1462) );
  assign n1463 = ( n64 & n336 ) | ( n64 & n1462 ) | ( n336 & n1462 ) ;
  assign n1464 = ~n337 & n1463 ;
  assign n1465 = n498 & ~n555 ;
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  assign n1472 = ( n532 & n1464 ) | ( n532 & n1471 ) | ( n1464 & n1471 ) ;
  assign n1473 = ~n533 & n1472 ;
  assign n1474 = n677 & n1473 ;
  assign n1475 = ( n786 & n816 ) | ( n786 & n1474 ) | ( n816 & n1474 ) ;
  assign n1476 = ~n817 & n1475 ;
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n131( .i (x3), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  assign n1488 = n150 & n504 ;
  assign n1489 = ( ~n66 & n477 ) | ( ~n66 & n1488 ) | ( n477 & n1488 ) ;
  assign n1490 = n67 & n1489 ;
  buffer buf_n711( .i (x27), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  assign n1491 = n533 & n732 ;
  assign n1492 = ( n564 & n1490 ) | ( n564 & n1491 ) | ( n1490 & n1491 ) ;
  assign n1493 = ~n565 & n1492 ;
  buffer buf_n1494( .i (n786), .o (n1494) );
  assign n1495 = n1493 & ~n1494 ;
  assign n1496 = ~n818 & n1495 ;
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n180( .i (x5), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  assign n1505 = n57 & ~n191 ;
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  assign n1514 = n505 & n1513 ;
  assign n1515 = n478 & n1514 ;
  assign n1516 = n532 & ~n731 ;
  buffer buf_n1517( .i (n1516), .o (n1517) );
  assign n1518 = ( n564 & n1515 ) | ( n564 & n1517 ) | ( n1515 & n1517 ) ;
  assign n1519 = ~n565 & n1518 ;
  assign n1520 = n817 & n1519 ;
  assign n1521 = ( n760 & n1440 ) | ( n760 & n1520 ) | ( n1440 & n1520 ) ;
  assign n1522 = ~n761 & n1521 ;
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n157( .i (x4), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  assign n1529 = ~n176 & n504 ;
  assign n1530 = ( n66 & n477 ) | ( n66 & n1529 ) | ( n477 & n1529 ) ;
  buffer buf_n1531( .i (n66), .o (n1531) );
  assign n1532 = n1530 & ~n1531 ;
  buffer buf_n1533( .i (n563), .o (n1533) );
  assign n1534 = ( n1517 & n1532 ) | ( n1517 & n1533 ) | ( n1532 & n1533 ) ;
  assign n1535 = ~n565 & n1534 ;
  assign n1536 = n759 & n1535 ;
  assign n1537 = ( n818 & n1440 ) | ( n818 & n1536 ) | ( n1440 & n1536 ) ;
  assign n1538 = ~n819 & n1537 ;
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  assign n1546 = n1528 | n1544 ;
  assign n1547 = n1504 | n1546 ;
  assign n1548 = ~n561 & n704 ;
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1553( .i (n531), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  assign n1555 = ( n1392 & n1549 ) | ( n1392 & n1554 ) | ( n1549 & n1554 ) ;
  assign n1556 = ~n534 & n1555 ;
  assign n1557 = ~n816 & n1556 ;
  buffer buf_n1558( .i (n758), .o (n1558) );
  assign n1559 = ( n1494 & n1557 ) | ( n1494 & n1558 ) | ( n1557 & n1558 ) ;
  buffer buf_n1560( .i (n1558), .o (n1560) );
  assign n1561 = n1559 & ~n1560 ;
  buffer buf_n1562( .i (n1561), .o (n1562) );
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  assign n1571 = n339 & n506 ;
  assign n1572 = ( ~n68 & n479 ) | ( ~n68 & n1571 ) | ( n479 & n1571 ) ;
  assign n1573 = n69 & n1572 ;
  assign n1574 = ( n536 & n1552 ) | ( n536 & n1573 ) | ( n1552 & n1573 ) ;
  assign n1575 = ~n537 & n1574 ;
  assign n1576 = ( n789 & n1438 ) | ( n789 & n1575 ) | ( n1438 & n1575 ) ;
  assign n1577 = ~n790 & n1576 ;
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1585( .i (n476), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  assign n1588 = ( n340 & n1390 ) | ( n340 & n1587 ) | ( n1390 & n1587 ) ;
  assign n1589 = ~n341 & n1588 ;
  assign n1590 = ( n536 & n1552 ) | ( n536 & n1589 ) | ( n1552 & n1589 ) ;
  assign n1591 = ~n537 & n1590 ;
  buffer buf_n1592( .i (n1440), .o (n1592) );
  assign n1593 = ( n1438 & n1591 ) | ( n1438 & n1592 ) | ( n1591 & n1592 ) ;
  assign n1594 = ~n790 & n1593 ;
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  assign n1599 = n1580 | n1597 ;
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  assign n1602 = n1569 | n1601 ;
  assign n1603 = ( ~n1486 & n1547 ) | ( ~n1486 & n1602 ) | ( n1547 & n1602 ) ;
  assign n1604 = n1487 | n1603 ;
  buffer buf_n107( .i (x2), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  assign n1605 = n63 & ~n148 ;
  assign n1606 = ( n125 & ~n475 ) | ( n125 & n1605 ) | ( ~n475 & n1605 ) ;
  assign n1607 = ~n126 & n1606 ;
  assign n1608 = ~n562 & n1607 ;
  assign n1609 = ( n506 & n1554 ) | ( n506 & n1608 ) | ( n1554 & n1608 ) ;
  assign n1610 = ~n507 & n1609 ;
  buffer buf_n1611( .i (n785), .o (n1611) );
  assign n1612 = ( n1435 & n1610 ) | ( n1435 & n1611 ) | ( n1610 & n1611 ) ;
  assign n1613 = ~n1494 & n1612 ;
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n604( .i (x23), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  assign n1622 = ~n757 & n1375 ;
  buffer buf_n1623( .i (n1533), .o (n1623) );
  assign n1624 = ( n627 & n1622 ) | ( n627 & n1623 ) | ( n1622 & n1623 ) ;
  assign n1625 = ~n566 & n1624 ;
  buffer buf_n1626( .i (n817), .o (n1626) );
  assign n1627 = n1625 & ~n1626 ;
  assign n1628 = n1592 & n1627 ;
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  assign n1637 = n124 & ~n474 ;
  assign n1638 = ( n64 & n149 ) | ( n64 & n1637 ) | ( n149 & n1637 ) ;
  assign n1639 = ~n150 & n1638 ;
  assign n1640 = ~n1553 & n1639 ;
  buffer buf_n1641( .i (n505), .o (n1641) );
  assign n1642 = ( ~n563 & n1640 ) | ( ~n563 & n1641 ) | ( n1640 & n1641 ) ;
  buffer buf_n1643( .i (n1641), .o (n1643) );
  assign n1644 = n1642 & ~n1643 ;
  assign n1645 = ( n1435 & n1611 ) | ( n1435 & n1644 ) | ( n1611 & n1644 ) ;
  assign n1646 = ~n1494 & n1645 ;
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n391( .i (x15), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  assign n1656 = ~n410 & n1512 ;
  assign n1657 = n338 & n1656 ;
  assign n1658 = n471 & n526 ;
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  assign n1669 = ( n1641 & n1657 ) | ( n1641 & n1664 ) | ( n1657 & n1664 ) ;
  assign n1670 = ~n1643 & n1669 ;
  assign n1671 = n1623 & n1670 ;
  assign n1672 = ( n709 & n1558 ) | ( n709 & n1671 ) | ( n1558 & n1671 ) ;
  assign n1673 = ~n1560 & n1672 ;
  assign n1674 = n1236 & n1673 ;
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  assign n1681 = ~n331 & n1506 ;
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  assign n1684 = ~n407 & n1683 ;
  assign n1685 = ( n502 & n1660 ) | ( n502 & n1684 ) | ( n1660 & n1684 ) ;
  assign n1686 = ~n503 & n1685 ;
  buffer buf_n1687( .i (n560), .o (n1687) );
  assign n1688 = n1686 & n1687 ;
  assign n1689 = ( n705 & n755 ) | ( n705 & n1688 ) | ( n755 & n1688 ) ;
  assign n1690 = ~n756 & n1689 ;
  assign n1691 = n1232 & n1690 ;
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n411( .i (n410), .o (n411) );
  assign n1704 = n334 & n1509 ;
  assign n1705 = n309 & n1704 ;
  assign n1706 = ~n503 & n1705 ;
  buffer buf_n1707( .i (n475), .o (n1707) );
  assign n1708 = ( n410 & n1706 ) | ( n410 & n1707 ) | ( n1706 & n1707 ) ;
  assign n1709 = ~n411 & n1708 ;
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  assign n1712 = n530 & n673 ;
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  assign n1716 = ( n1533 & ~n1710 ) | ( n1533 & n1715 ) | ( ~n1710 & n1715 ) ;
  assign n1717 = n1711 & n1716 ;
  assign n1718 = ( n1234 & n1558 ) | ( n1234 & n1717 ) | ( n1558 & n1717 ) ;
  assign n1719 = ~n1560 & n1718 ;
  buffer buf_n1720( .i (n1719), .o (n1720) );
  assign n1727 = ( n149 & ~n475 ) | ( n149 & n1511 ) | ( ~n475 & n1511 ) ;
  assign n1728 = ~n150 & n1727 ;
  assign n1729 = ~n1553 & n1728 ;
  buffer buf_n1730( .i (n1687), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  assign n1732 = ( n1641 & n1729 ) | ( n1641 & ~n1731 ) | ( n1729 & ~n1731 ) ;
  assign n1733 = ~n1643 & n1732 ;
  assign n1734 = ~n816 & n1733 ;
  buffer buf_n1735( .i (n758), .o (n1735) );
  buffer buf_n1736( .i (n1611), .o (n1736) );
  assign n1737 = ( n1734 & n1735 ) | ( n1734 & n1736 ) | ( n1735 & n1736 ) ;
  assign n1738 = ~n1560 & n1737 ;
  buffer buf_n1739( .i (n1738), .o (n1739) );
  assign n1746 = n1720 | n1739 ;
  assign n1747 = ( ~n1675 & n1696 ) | ( ~n1675 & n1746 ) | ( n1696 & n1746 ) ;
  assign n1748 = n1676 | n1747 ;
  assign n1749 = n1651 | n1748 ;
  assign n1750 = ( ~n1619 & n1632 ) | ( ~n1619 & n1749 ) | ( n1632 & n1749 ) ;
  assign n1751 = n1620 | n1750 ;
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n573( .i (x22), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  assign n1754 = n593 & n813 ;
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1736), .o (n1759) );
  assign n1760 = ( n1378 & n1758 ) | ( n1378 & n1759 ) | ( n1758 & n1759 ) ;
  assign n1761 = ~n1592 & n1760 ;
  buffer buf_n1762( .i (n1761), .o (n1762) );
  assign n1763 = n311 & ~n1707 ;
  buffer buf_n1764( .i (n65), .o (n1764) );
  assign n1765 = ( n338 & n1763 ) | ( n338 & n1764 ) | ( n1763 & n1764 ) ;
  assign n1766 = ~n339 & n1765 ;
  assign n1767 = n1533 & n1766 ;
  assign n1768 = ( n508 & n535 ) | ( n508 & n1767 ) | ( n535 & n1767 ) ;
  assign n1769 = ~n509 & n1768 ;
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n1770( .i (n815), .o (n1770) );
  assign n1771 = n678 & n1770 ;
  buffer buf_n1772( .i (n1771), .o (n1772) );
  assign n1774 = ( n1759 & n1769 ) | ( n1759 & n1772 ) | ( n1769 & n1772 ) ;
  assign n1775 = ~n1592 & n1774 ;
  buffer buf_n1776( .i (n1775), .o (n1776) );
  assign n1782 = n1762 | n1776 ;
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  assign n1788 = n337 & ~n504 ;
  assign n1789 = ( n1585 & n1764 ) | ( n1585 & n1788 ) | ( n1764 & n1788 ) ;
  assign n1790 = ~n1586 & n1789 ;
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  assign n1793 = n529 & n702 ;
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  assign n1800 = ( n1623 & ~n1791 ) | ( n1623 & n1798 ) | ( ~n1791 & n1798 ) ;
  assign n1801 = n1792 & n1800 ;
  assign n1802 = n1235 & n1801 ;
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n412( .i (n411), .o (n412) );
  assign n1809 = ( n411 & n1217 ) | ( n411 & n1513 ) | ( n1217 & n1513 ) ;
  assign n1810 = ~n412 & n1809 ;
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  assign n1813 = n529 & n590 ;
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  buffer buf_n1818( .i (n1817), .o (n1818) );
  assign n1819 = ( n1623 & ~n1811 ) | ( n1623 & n1818 ) | ( ~n1811 & n1818 ) ;
  assign n1820 = n1812 & n1819 ;
  buffer buf_n1821( .i (n1735), .o (n1821) );
  assign n1822 = ( n1235 & n1820 ) | ( n1235 & n1821 ) | ( n1820 & n1821 ) ;
  buffer buf_n1823( .i (n1821), .o (n1823) );
  assign n1824 = n1822 & ~n1823 ;
  buffer buf_n1825( .i (n1824), .o (n1825) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  assign n1837 = n307 & n1682 ;
  assign n1838 = ~n501 & n1837 ;
  assign n1839 = ( n408 & n474 ) | ( n408 & n1838 ) | ( n474 & n1838 ) ;
  assign n1840 = ~n409 & n1839 ;
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  assign n1843 = ( n1713 & n1730 ) | ( n1713 & ~n1841 ) | ( n1730 & ~n1841 ) ;
  assign n1844 = n1842 & n1843 ;
  assign n1845 = ( n757 & n1232 ) | ( n757 & n1844 ) | ( n1232 & n1844 ) ;
  buffer buf_n1846( .i (n757), .o (n1846) );
  assign n1847 = n1845 & ~n1846 ;
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  buffer buf_n1856( .i (n502), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  assign n1858 = n1512 & ~n1857 ;
  assign n1859 = ( n411 & n1585 ) | ( n411 & n1858 ) | ( n1585 & n1858 ) ;
  assign n1860 = ~n412 & n1859 ;
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1731), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  assign n1865 = ( n1818 & ~n1861 ) | ( n1818 & n1864 ) | ( ~n1861 & n1864 ) ;
  assign n1866 = n1862 & n1865 ;
  buffer buf_n1867( .i (n1234), .o (n1867) );
  assign n1868 = ( n1821 & n1866 ) | ( n1821 & n1867 ) | ( n1866 & n1867 ) ;
  assign n1869 = ~n1823 & n1868 ;
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  assign n1872 = n1852 | n1871 ;
  buffer buf_n1873( .i (n1872), .o (n1873) );
  assign n1875 = n1828 | n1873 ;
  assign n1876 = n1808 | n1875 ;
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n510( .i (n509), .o (n510) );
  assign n1877 = n312 & n1764 ;
  assign n1878 = ( n339 & n1586 ) | ( n339 & n1877 ) | ( n1586 & n1877 ) ;
  assign n1879 = ~n1587 & n1878 ;
  assign n1880 = n1864 & n1879 ;
  assign n1881 = ( n509 & n536 ) | ( n509 & n1880 ) | ( n536 & n1880 ) ;
  assign n1882 = ~n510 & n1881 ;
  buffer buf_n1883( .i (n1759), .o (n1883) );
  assign n1884 = ( n1773 & n1882 ) | ( n1773 & n1883 ) | ( n1882 & n1883 ) ;
  assign n1885 = ~n790 & n1884 ;
  buffer buf_n1886( .i (n1885), .o (n1886) );
  assign n1888 = n65 & ~n1707 ;
  assign n1889 = ( n338 & ~n505 ) | ( n338 & n1888 ) | ( ~n505 & n1888 ) ;
  buffer buf_n1890( .i (n337), .o (n1890) );
  buffer buf_n1891( .i (n1890), .o (n1891) );
  assign n1892 = n1889 & ~n1891 ;
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  assign n1895 = ( n1798 & n1864 ) | ( n1798 & ~n1893 ) | ( n1864 & ~n1893 ) ;
  assign n1896 = n1894 & n1895 ;
  assign n1897 = n1867 & n1896 ;
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  assign n1904 = n1886 | n1900 ;
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1907( .i (n1906), .o (n1907) );
  assign n1908 = n1876 | n1907 ;
  assign n1909 = ( ~n1752 & n1787 ) | ( ~n1752 & n1908 ) | ( n1787 & n1908 ) ;
  assign n1910 = n1753 | n1909 ;
  assign n1911 = ~n559 & n590 ;
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  assign n1915 = ( n1392 & n1554 ) | ( n1392 & n1914 ) | ( n1554 & n1914 ) ;
  assign n1916 = ~n534 & n1915 ;
  assign n1917 = ~n1770 & n1916 ;
  assign n1918 = n1736 & n1917 ;
  buffer buf_n1919( .i (n1918), .o (n1919) );
  buffer buf_n1920( .i (n1919), .o (n1920) );
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  assign n1929 = n62 & n528 ;
  buffer buf_n1930( .i (n473), .o (n1930) );
  buffer buf_n1931( .i (n501), .o (n1931) );
  assign n1932 = ( n1929 & n1930 ) | ( n1929 & n1931 ) | ( n1930 & n1931 ) ;
  buffer buf_n1933( .i (n1930), .o (n1933) );
  assign n1934 = n1932 & ~n1933 ;
  assign n1935 = n1912 & n1934 ;
  assign n1936 = n755 & n1935 ;
  assign n1937 = ( n784 & n814 ) | ( n784 & n1936 ) | ( n814 & n1936 ) ;
  assign n1938 = ~n815 & n1937 ;
  buffer buf_n1939( .i (n1938), .o (n1939) );
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  assign n1949 = n1215 & n1511 ;
  assign n1950 = ( n1687 & n1814 ) | ( n1687 & n1949 ) | ( n1814 & n1949 ) ;
  assign n1951 = ~n1730 & n1950 ;
  assign n1952 = ~n814 & n1951 ;
  buffer buf_n1953( .i (n756), .o (n1953) );
  buffer buf_n1954( .i (n784), .o (n1954) );
  assign n1955 = ( n1952 & n1953 ) | ( n1952 & n1954 ) | ( n1953 & n1954 ) ;
  assign n1956 = ~n1846 & n1955 ;
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  buffer buf_n1960( .i (n1959), .o (n1960) );
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n437( .i (x17), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  assign n1967 = n62 & n453 ;
  assign n1968 = ( n1930 & n1931 ) | ( n1930 & n1967 ) | ( n1931 & n1967 ) ;
  assign n1969 = ~n1856 & n1968 ;
  assign n1970 = ( n1687 & n1794 ) | ( n1687 & n1969 ) | ( n1794 & n1969 ) ;
  assign n1971 = ~n1730 & n1970 ;
  assign n1972 = ~n814 & n1971 ;
  assign n1973 = ( n1953 & n1954 ) | ( n1953 & n1972 ) | ( n1954 & n1972 ) ;
  assign n1974 = ~n1846 & n1973 ;
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  assign n1983 = ( n454 & n1410 ) | ( n454 & n1930 ) | ( n1410 & n1930 ) ;
  assign n1984 = ~n455 & n1983 ;
  buffer buf_n1985( .i (n560), .o (n1985) );
  assign n1986 = ( n1794 & n1984 ) | ( n1794 & n1985 ) | ( n1984 & n1985 ) ;
  buffer buf_n1987( .i (n1985), .o (n1987) );
  assign n1988 = n1986 & ~n1987 ;
  buffer buf_n1989( .i (n813), .o (n1989) );
  assign n1990 = n1988 & ~n1989 ;
  assign n1991 = ( n1953 & n1954 ) | ( n1953 & n1990 ) | ( n1954 & n1990 ) ;
  assign n1992 = ~n1846 & n1991 ;
  buffer buf_n1993( .i (n1992), .o (n1993) );
  assign n2002 = n1975 | n1993 ;
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n2003), .o (n2004) );
  buffer buf_n2005( .i (n2004), .o (n2005) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n2007( .i (n2006), .o (n2007) );
  buffer buf_n2008( .i (n2007), .o (n2008) );
  assign n2009 = n1964 | n2008 ;
  assign n2010 = n1948 | n2009 ;
  assign n2011 = ( ~n64 & n336 ) | ( ~n64 & n1462 ) | ( n336 & n1462 ) ;
  buffer buf_n2012( .i (n63), .o (n2012) );
  buffer buf_n2013( .i (n2012), .o (n2013) );
  assign n2014 = n2011 & n2013 ;
  assign n2015 = ( n1471 & n1553 ) | ( n1471 & n2014 ) | ( n1553 & n2014 ) ;
  assign n2016 = ~n1554 & n2015 ;
  assign n2017 = n677 & n2016 ;
  assign n2018 = ( n1611 & n1770 ) | ( n1611 & n2017 ) | ( n1770 & n2017 ) ;
  buffer buf_n2019( .i (n1770), .o (n2019) );
  assign n2020 = n2018 & ~n2019 ;
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2028( .i (n2027), .o (n2028) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  assign n2029 = ( n340 & n1415 ) | ( n340 & n1587 ) | ( n1415 & n1587 ) ;
  assign n2030 = ~n341 & n2029 ;
  assign n2031 = ( n566 & n1799 ) | ( n566 & n2030 ) | ( n1799 & n2030 ) ;
  assign n2032 = ~n567 & n2031 ;
  assign n2033 = ( n1438 & n1883 ) | ( n1438 & n2032 ) | ( n1883 & n2032 ) ;
  buffer buf_n2034( .i (n1883), .o (n2034) );
  assign n2035 = n2033 & ~n2034 ;
  buffer buf_n2036( .i (n2035), .o (n2036) );
  assign n2040 = n1531 & n1891 ;
  assign n2041 = ( n1587 & n1643 ) | ( n1587 & n2040 ) | ( n1643 & n2040 ) ;
  assign n2042 = ~n508 & n2041 ;
  buffer buf_n2043( .i (n1864), .o (n2043) );
  assign n2044 = ( n1799 & n2042 ) | ( n1799 & n2043 ) | ( n2042 & n2043 ) ;
  assign n2045 = ~n567 & n2044 ;
  assign n2046 = ( n1438 & n1883 ) | ( n1438 & n2045 ) | ( n1883 & n2045 ) ;
  assign n2047 = ~n2034 & n2046 ;
  buffer buf_n2048( .i (n2047), .o (n2048) );
  assign n2053 = n2036 | n2048 ;
  buffer buf_n2054( .i (n2053), .o (n2054) );
  buffer buf_n2055( .i (n2054), .o (n2055) );
  buffer buf_n2056( .i (n2055), .o (n2056) );
  assign n2057 = n2028 | n2056 ;
  assign n2058 = ( ~n1927 & n2010 ) | ( ~n1927 & n2057 ) | ( n2010 & n2057 ) ;
  assign n2059 = n1928 | n2058 ;
  assign n2060 = n1910 | n2059 ;
  assign n2061 = n1604 | n2060 ;
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  assign n2063 = n1852 | n1886 ;
  assign n2064 = n1778 | n2063 ;
  assign n2065 = n1482 | n2064 ;
  assign n2066 = ( ~n1725 & n2027 ) | ( ~n1725 & n2065 ) | ( n2027 & n2065 ) ;
  assign n2067 = n1726 | n2066 ;
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  assign n2073 = n1784 | n1828 ;
  assign n2074 = n1903 | n2073 ;
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1874( .i (n1873), .o (n1874) );
  assign n2075 = n1744 | n1874 ;
  assign n2076 = ( ~n1701 & n2074 ) | ( ~n1701 & n2075 ) | ( n2074 & n2075 ) ;
  assign n2077 = n1702 | n2076 ;
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  assign n2078 = n1617 | n2048 ;
  assign n2079 = ( ~n1923 & n1945 ) | ( ~n1923 & n2078 ) | ( n1945 & n2078 ) ;
  assign n2080 = n1924 | n2079 ;
  assign n2081 = n1598 | n2080 ;
  assign n2082 = ( n1484 & ~n1544 ) | ( n1484 & n2081 ) | ( ~n1544 & n2081 ) ;
  assign n2083 = n1545 | n2082 ;
  assign n2084 = n2077 | n2083 ;
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  assign n2088 = n1499 | n1630 ;
  assign n2089 = n1651 | n2088 ;
  buffer buf_n2090( .i (n2089), .o (n2090) );
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  assign n2098 = ~n496 & n553 ;
  buffer buf_n2099( .i (n2098), .o (n2099) );
  assign n2102 = ( n470 & ~n525 ) | ( n470 & n2099 ) | ( ~n525 & n2099 ) ;
  assign n2103 = ~n471 & n2102 ;
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n2111( .i (n2110), .o (n2111) );
  assign n2113 = n591 & n781 ;
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n1953), .o (n2118) );
  assign n2119 = ( n2111 & n2117 ) | ( n2111 & n2118 ) | ( n2117 & n2118 ) ;
  assign n2120 = ~n1735 & n2119 ;
  assign n2121 = n1626 & n2120 ;
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n1090( .i (x40), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1138( .i (x42), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1111( .i (x41), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1064( .i (x39), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1049( .i (x38), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n274( .i (x9), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  assign n2128 = n461 | n516 ;
  assign n2129 = ( ~n279 & n490 ) | ( ~n279 & n2128 ) | ( n490 & n2128 ) ;
  assign n2130 = n280 | n2129 ;
  assign n2131 = n549 & ~n2130 ;
  assign n2132 = ( n581 & n743 ) | ( n581 & n2131 ) | ( n743 & n2131 ) ;
  assign n2133 = ~n744 & n2132 ;
  buffer buf_n2134( .i (n2133), .o (n2134) );
  assign n2149 = ~n804 & n2134 ;
  assign n2150 = n775 & n2149 ;
  buffer buf_n2151( .i (n2150), .o (n2151) );
  assign n2152 = ~n1063 & n2151 ;
  buffer buf_n2153( .i (n2152), .o (n2153) );
  assign n2163 = ~n1080 & n2153 ;
  buffer buf_n2164( .i (n2163), .o (n2164) );
  assign n2171 = ~n1129 & n2164 ;
  assign n2172 = ( n1109 & ~n1157 ) | ( n1109 & n2171 ) | ( ~n1157 & n2171 ) ;
  assign n2173 = ~n1110 & n2172 ;
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n1163( .i (x43), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1187( .i (x44), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  assign n2175 = ~n1184 & n1208 ;
  assign n2176 = n2174 & n2175 ;
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n2177), .o (n2178) );
  buffer buf_n2179( .i (n2178), .o (n2179) );
  buffer buf_n2180( .i (n2179), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  buffer buf_n2182( .i (n2181), .o (n2182) );
  buffer buf_n2183( .i (n2182), .o (n2183) );
  buffer buf_n2184( .i (n2183), .o (n2184) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n2155( .i (n2154), .o (n2155) );
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n2158( .i (n2157), .o (n2158) );
  buffer buf_n2159( .i (n2158), .o (n2159) );
  buffer buf_n2160( .i (n2159), .o (n2160) );
  buffer buf_n2161( .i (n2160), .o (n2161) );
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  assign n2189 = n1088 & n1162 ;
  assign n2190 = ( n1136 & n2162 ) | ( n1136 & n2189 ) | ( n2162 & n2189 ) ;
  assign n2191 = ~n1137 & n2190 ;
  buffer buf_n2192( .i (n2191), .o (n2192) );
  buffer buf_n2193( .i (n2192), .o (n2193) );
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n2166( .i (n2165), .o (n2166) );
  buffer buf_n2167( .i (n2166), .o (n2167) );
  buffer buf_n2168( .i (n2167), .o (n2168) );
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  assign n2197 = ~n1134 & n1161 ;
  assign n2198 = n2170 & n2197 ;
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n2200( .i (n2199), .o (n2200) );
  buffer buf_n2201( .i (n2200), .o (n2201) );
  assign n2207 = n1087 & ~n1161 ;
  assign n2208 = ( n1135 & n2161 ) | ( n1135 & n2207 ) | ( n2161 & n2207 ) ;
  assign n2209 = ~n1136 & n2208 ;
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n2211( .i (n2210), .o (n2211) );
  assign n2214 = n2201 | n2211 ;
  assign n2215 = n2193 | n2214 ;
  buffer buf_n2216( .i (n2215), .o (n2216) );
  assign n2219 = n2184 | n2216 ;
  assign n2220 = n2127 | n2219 ;
  buffer buf_n2221( .i (n2220), .o (n2221) );
  buffer buf_n2222( .i (n2221), .o (n2222) );
  buffer buf_n456( .i (n455), .o (n456) );
  assign n2226 = ( n456 & n1662 ) | ( n456 & n1857 ) | ( n1662 & n1857 ) ;
  buffer buf_n2227( .i (n1857), .o (n2227) );
  assign n2228 = n2226 & ~n2227 ;
  assign n2229 = n1549 & n2228 ;
  buffer buf_n2230( .i (n2229), .o (n2230) );
  assign n2232 = ~n2118 & n2230 ;
  buffer buf_n2233( .i (n2232), .o (n2233) );
  assign n2234 = ~n1626 & n2233 ;
  buffer buf_n2235( .i (n1759), .o (n2235) );
  assign n2236 = n2234 & n2235 ;
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  assign n2246 = ( n452 & n472 ) | ( n452 & n1362 ) | ( n472 & n1362 ) ;
  assign n2247 = ~n453 & n2246 ;
  assign n2248 = ~n752 & n2247 ;
  buffer buf_n2249( .i (n559), .o (n2249) );
  assign n2250 = ( n703 & n2248 ) | ( n703 & n2249 ) | ( n2248 & n2249 ) ;
  assign n2251 = ~n1985 & n2250 ;
  buffer buf_n2252( .i (n2251), .o (n2252) );
  assign n2256 = n1989 & n2252 ;
  assign n2257 = n1954 & n2256 ;
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  buffer buf_n2265( .i (n2264), .o (n2265) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  assign n2274 = n473 & ~n558 ;
  assign n2275 = ( n529 & n1931 ) | ( n529 & n2274 ) | ( n1931 & n2274 ) ;
  assign n2276 = ~n1856 & n2275 ;
  buffer buf_n2277( .i (n2276), .o (n2277) );
  buffer buf_n2278( .i (n2277), .o (n2278) );
  assign n2279 = n703 & n781 ;
  buffer buf_n2280( .i (n2279), .o (n2280) );
  assign n2281 = ( n755 & ~n2277 ) | ( n755 & n2280 ) | ( ~n2277 & n2280 ) ;
  assign n2282 = n2278 & n2281 ;
  buffer buf_n2283( .i (n1989), .o (n2283) );
  assign n2284 = n2282 & ~n2283 ;
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n2289( .i (n2288), .o (n2289) );
  buffer buf_n2290( .i (n2289), .o (n2290) );
  buffer buf_n2291( .i (n2290), .o (n2291) );
  buffer buf_n2292( .i (n2291), .o (n2292) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  assign n2301 = ~n557 & n1212 ;
  assign n2302 = n528 & n2301 ;
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  assign n2307 = ~n756 & n2306 ;
  assign n2308 = n595 & n2307 ;
  buffer buf_n2309( .i (n2308), .o (n2309) );
  assign n2311 = n2019 & n2309 ;
  buffer buf_n2312( .i (n1736), .o (n2312) );
  assign n2313 = n2311 & n2312 ;
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  assign n2321 = n753 & n2303 ;
  assign n2322 = n592 & n2321 ;
  buffer buf_n2323( .i (n2322), .o (n2323) );
  assign n2328 = n1989 & n2323 ;
  buffer buf_n2329( .i (n784), .o (n2329) );
  assign n2330 = n2328 & n2329 ;
  buffer buf_n2331( .i (n2330), .o (n2331) );
  buffer buf_n2332( .i (n2331), .o (n2332) );
  buffer buf_n2333( .i (n2332), .o (n2333) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n2335( .i (n2334), .o (n2335) );
  buffer buf_n79( .i (x1), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  assign n2342 = n94 & ~n527 ;
  buffer buf_n2343( .i (n472), .o (n2343) );
  assign n2344 = ( n501 & n2342 ) | ( n501 & n2343 ) | ( n2342 & n2343 ) ;
  buffer buf_n2345( .i (n2343), .o (n2345) );
  assign n2346 = n2344 & ~n2345 ;
  buffer buf_n2347( .i (n2346), .o (n2347) );
  buffer buf_n2348( .i (n2347), .o (n2348) );
  buffer buf_n2349( .i (n2348), .o (n2349) );
  assign n2350 = ~n1731 & n2349 ;
  buffer buf_n2351( .i (n2350), .o (n2351) );
  assign n2352 = n627 & n2351 ;
  buffer buf_n2353( .i (n2329), .o (n2353) );
  buffer buf_n2354( .i (n2353), .o (n2354) );
  assign n2355 = ( n2019 & n2352 ) | ( n2019 & n2354 ) | ( n2352 & n2354 ) ;
  assign n2356 = ~n1626 & n2355 ;
  buffer buf_n2357( .i (n2356), .o (n2357) );
  buffer buf_n2358( .i (n2357), .o (n2358) );
  assign n2365 = n2335 | n2358 ;
  assign n2366 = n2316 | n2365 ;
  buffer buf_n2367( .i (n2366), .o (n2367) );
  assign n2371 = n2292 | n2367 ;
  assign n2372 = ( ~n2241 & n2266 ) | ( ~n2241 & n2371 ) | ( n2266 & n2371 ) ;
  assign n2373 = n2242 | n2372 ;
  assign n2374 = n1135 & n2161 ;
  buffer buf_n2375( .i (n2374), .o (n2375) );
  buffer buf_n2376( .i (n2375), .o (n2376) );
  buffer buf_n2377( .i (n2376), .o (n2377) );
  buffer buf_n2378( .i (n2377), .o (n2378) );
  buffer buf_n2379( .i (n2378), .o (n2379) );
  buffer buf_n2380( .i (n2379), .o (n2380) );
  buffer buf_n2381( .i (n2380), .o (n2381) );
  assign n2386 = n1063 & n2151 ;
  buffer buf_n2387( .i (n2386), .o (n2387) );
  buffer buf_n2388( .i (n2387), .o (n2388) );
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2391( .i (n2390), .o (n2391) );
  buffer buf_n2392( .i (n2391), .o (n2392) );
  buffer buf_n2393( .i (n2392), .o (n2393) );
  buffer buf_n2394( .i (n2393), .o (n2394) );
  buffer buf_n2395( .i (n2394), .o (n2395) );
  buffer buf_n2396( .i (n2395), .o (n2396) );
  buffer buf_n2397( .i (n2396), .o (n2397) );
  buffer buf_n2398( .i (n2397), .o (n2398) );
  buffer buf_n2399( .i (n2398), .o (n2399) );
  buffer buf_n2400( .i (n2399), .o (n2400) );
  buffer buf_n2401( .i (n2400), .o (n2401) );
  buffer buf_n2402( .i (n2401), .o (n2402) );
  buffer buf_n823( .i (x31), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  assign n2405 = n291 & ~n1931 ;
  assign n2406 = ( ~n530 & n1933 ) | ( ~n530 & n2405 ) | ( n1933 & n2405 ) ;
  assign n2407 = ~n1707 & n2406 ;
  assign n2408 = n1987 & n2407 ;
  buffer buf_n2409( .i (n754), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  assign n2411 = ( n594 & n2408 ) | ( n594 & n2410 ) | ( n2408 & n2410 ) ;
  buffer buf_n2412( .i (n2410), .o (n2412) );
  assign n2413 = n2411 & ~n2412 ;
  assign n2414 = n1233 & n2413 ;
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n2416( .i (n2415), .o (n2416) );
  buffer buf_n883( .i (x33), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  assign n2424 = ~n908 & n1089 ;
  assign n2425 = ( n849 & n2416 ) | ( n849 & n2424 ) | ( n2416 & n2424 ) ;
  assign n2426 = ~n850 & n2425 ;
  buffer buf_n2427( .i (n2426), .o (n2427) );
  buffer buf_n2428( .i (n2427), .o (n2428) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  assign n2433 = n472 & n500 ;
  assign n2434 = ( n528 & n558 ) | ( n528 & n2433 ) | ( n558 & n2433 ) ;
  assign n2435 = ~n559 & n2434 ;
  buffer buf_n2436( .i (n2435), .o (n2436) );
  buffer buf_n2437( .i (n2436), .o (n2437) );
  buffer buf_n2438( .i (n2437), .o (n2438) );
  buffer buf_n2441( .i (n783), .o (n2441) );
  assign n2442 = n2438 & n2441 ;
  assign n2443 = ( n733 & n2412 ) | ( n733 & n2442 ) | ( n2412 & n2442 ) ;
  assign n2444 = ~n734 & n2443 ;
  assign n2445 = n2019 & n2444 ;
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n2448( .i (n2447), .o (n2448) );
  buffer buf_n2449( .i (n2448), .o (n2449) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  buffer buf_n2137( .i (n2136), .o (n2137) );
  buffer buf_n2138( .i (n2137), .o (n2138) );
  buffer buf_n2139( .i (n2138), .o (n2139) );
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n2143( .i (n2142), .o (n2143) );
  buffer buf_n2144( .i (n2143), .o (n2144) );
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  assign n2457 = n1867 & n2148 ;
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n2439( .i (n2438), .o (n2439) );
  buffer buf_n2440( .i (n2439), .o (n2440) );
  assign n2464 = n733 & n2283 ;
  assign n2465 = ( n2353 & n2440 ) | ( n2353 & n2464 ) | ( n2440 & n2464 ) ;
  assign n2466 = ~n2354 & n2465 ;
  buffer buf_n2467( .i (n2466), .o (n2467) );
  buffer buf_n2468( .i (n2467), .o (n2468) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  assign n2477 = n2459 | n2469 ;
  assign n2478 = n2449 | n2477 ;
  assign n2479 = n2428 | n2478 ;
  assign n2480 = ( ~n2380 & n2402 ) | ( ~n2380 & n2479 ) | ( n2402 & n2479 ) ;
  assign n2481 = n2381 | n2480 ;
  assign n2482 = n2438 & ~n2441 ;
  assign n2483 = ( n733 & n2412 ) | ( n733 & n2482 ) | ( n2412 & n2482 ) ;
  assign n2484 = ~n734 & n2483 ;
  buffer buf_n2485( .i (n2484), .o (n2485) );
  buffer buf_n2488( .i (n2283), .o (n2488) );
  buffer buf_n2489( .i (n2488), .o (n2489) );
  buffer buf_n2490( .i (n2489), .o (n2490) );
  assign n2491 = n2485 & ~n2490 ;
  buffer buf_n2492( .i (n2491), .o (n2492) );
  buffer buf_n2493( .i (n2492), .o (n2493) );
  buffer buf_n2494( .i (n2493), .o (n2494) );
  buffer buf_n2495( .i (n2494), .o (n2495) );
  buffer buf_n2496( .i (n2495), .o (n2496) );
  buffer buf_n2497( .i (n2496), .o (n2497) );
  buffer buf_n2498( .i (n470), .o (n2498) );
  buffer buf_n2499( .i (n2498), .o (n2499) );
  assign n2500 = ( n527 & n1466 ) | ( n527 & n2499 ) | ( n1466 & n2499 ) ;
  buffer buf_n2501( .i (n526), .o (n2501) );
  buffer buf_n2502( .i (n2501), .o (n2502) );
  assign n2503 = n2500 & ~n2502 ;
  buffer buf_n2504( .i (n2503), .o (n2504) );
  assign n2513 = n753 & n2504 ;
  assign n2514 = n704 & n2513 ;
  buffer buf_n2515( .i (n2514), .o (n2515) );
  buffer buf_n2516( .i (n813), .o (n2516) );
  assign n2517 = n2515 & ~n2516 ;
  assign n2518 = n2329 & n2517 ;
  buffer buf_n2519( .i (n2518), .o (n2519) );
  buffer buf_n2520( .i (n2519), .o (n2520) );
  buffer buf_n2521( .i (n2520), .o (n2521) );
  buffer buf_n2522( .i (n2521), .o (n2522) );
  buffer buf_n2523( .i (n2522), .o (n2523) );
  buffer buf_n2524( .i (n2523), .o (n2524) );
  buffer buf_n2525( .i (n2524), .o (n2525) );
  buffer buf_n2526( .i (n2525), .o (n2526) );
  buffer buf_n2505( .i (n2504), .o (n2505) );
  buffer buf_n2506( .i (n2505), .o (n2506) );
  buffer buf_n2507( .i (n2506), .o (n2507) );
  buffer buf_n2508( .i (n2507), .o (n2508) );
  buffer buf_n2509( .i (n2508), .o (n2509) );
  assign n2529 = ( n1755 & n2329 ) | ( n1755 & ~n2508 ) | ( n2329 & ~n2508 ) ;
  assign n2530 = n2509 & n2529 ;
  buffer buf_n2531( .i (n2530), .o (n2531) );
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n2532), .o (n2533) );
  buffer buf_n2534( .i (n2533), .o (n2534) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  buffer buf_n2536( .i (n2535), .o (n2536) );
  assign n2539 = ~n2409 & n2506 ;
  assign n2540 = n706 & n2539 ;
  buffer buf_n2541( .i (n2540), .o (n2541) );
  assign n2543 = n2488 & n2541 ;
  assign n2544 = n2354 & n2543 ;
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2510( .i (n2509), .o (n2510) );
  buffer buf_n2511( .i (n2510), .o (n2511) );
  buffer buf_n2512( .i (n2511), .o (n2512) );
  assign n2554 = ( n1772 & n2312 ) | ( n1772 & ~n2511 ) | ( n2312 & ~n2511 ) ;
  assign n2555 = n2512 & n2554 ;
  buffer buf_n2556( .i (n2555), .o (n2556) );
  buffer buf_n2557( .i (n2556), .o (n2557) );
  assign n2564 = n2548 | n2557 ;
  assign n2565 = n2536 | n2564 ;
  assign n2566 = n2526 | n2565 ;
  assign n2567 = n2497 | n2566 ;
  assign n2568 = n2481 | n2567 ;
  assign n2569 = ( ~n2221 & n2373 ) | ( ~n2221 & n2568 ) | ( n2373 & n2568 ) ;
  assign n2570 = n2222 | n2569 ;
  buffer buf_n2571( .i (n2570), .o (n2571) );
  buffer buf_n2572( .i (n2571), .o (n2572) );
  buffer buf_n2573( .i (n531), .o (n2573) );
  assign n2574 = ( n1269 & ~n1585 ) | ( n1269 & n2573 ) | ( ~n1585 & n2573 ) ;
  assign n2575 = n1586 & n2574 ;
  buffer buf_n2576( .i (n2575), .o (n2576) );
  assign n2577 = ~n2488 & n2576 ;
  assign n2578 = n2354 & n2577 ;
  buffer buf_n2579( .i (n2578), .o (n2579) );
  buffer buf_n2580( .i (n2579), .o (n2580) );
  buffer buf_n2581( .i (n2580), .o (n2581) );
  buffer buf_n2582( .i (n2581), .o (n2582) );
  buffer buf_n2583( .i (n2582), .o (n2583) );
  buffer buf_n2584( .i (n2583), .o (n2584) );
  buffer buf_n2585( .i (n2584), .o (n2585) );
  buffer buf_n2586( .i (n2585), .o (n2586) );
  buffer buf_n2587( .i (n2586), .o (n2587) );
  buffer buf_n2588( .i (n2587), .o (n2588) );
  buffer buf_n2589( .i (n2588), .o (n2589) );
  assign n2590 = n673 & n781 ;
  buffer buf_n2591( .i (n2590), .o (n2591) );
  buffer buf_n2592( .i (n500), .o (n2592) );
  assign n2593 = ( n334 & n1659 ) | ( n334 & n2592 ) | ( n1659 & n2592 ) ;
  buffer buf_n2594( .i (n2592), .o (n2594) );
  assign n2595 = n2593 & ~n2594 ;
  assign n2596 = n2249 & n2595 ;
  buffer buf_n2597( .i (n2596), .o (n2597) );
  assign n2598 = ( n2409 & n2591 ) | ( n2409 & n2597 ) | ( n2591 & n2597 ) ;
  assign n2599 = ~n2410 & n2598 ;
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  buffer buf_n2602( .i (n2601), .o (n2602) );
  buffer buf_n2603( .i (n2602), .o (n2603) );
  buffer buf_n2604( .i (n2603), .o (n2604) );
  buffer buf_n2605( .i (n2604), .o (n2605) );
  buffer buf_n2606( .i (n2605), .o (n2606) );
  buffer buf_n2607( .i (n2606), .o (n2607) );
  buffer buf_n2608( .i (n2607), .o (n2608) );
  buffer buf_n2609( .i (n2608), .o (n2609) );
  buffer buf_n2610( .i (n2609), .o (n2610) );
  buffer buf_n2611( .i (n2610), .o (n2611) );
  assign n2613 = ( n334 & n1363 ) | ( n334 & n2343 ) | ( n1363 & n2343 ) ;
  assign n2614 = ~n335 & n2613 ;
  assign n2615 = n2249 & n2614 ;
  buffer buf_n2616( .i (n2615), .o (n2616) );
  assign n2617 = ( n2280 & n2409 ) | ( n2280 & n2616 ) | ( n2409 & n2616 ) ;
  assign n2618 = ~n2410 & n2617 ;
  buffer buf_n2619( .i (n2618), .o (n2619) );
  buffer buf_n2620( .i (n2619), .o (n2620) );
  buffer buf_n2621( .i (n2620), .o (n2621) );
  buffer buf_n2622( .i (n2621), .o (n2622) );
  buffer buf_n2623( .i (n2622), .o (n2623) );
  buffer buf_n2624( .i (n2623), .o (n2624) );
  buffer buf_n2625( .i (n2624), .o (n2625) );
  buffer buf_n2626( .i (n2625), .o (n2626) );
  buffer buf_n2627( .i (n2626), .o (n2627) );
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  assign n2631 = n820 & ~n2623 ;
  buffer buf_n2632( .i (n2631), .o (n2632) );
  buffer buf_n2633( .i (n2632), .o (n2633) );
  buffer buf_n2634( .i (n2633), .o (n2634) );
  buffer buf_n2635( .i (n2634), .o (n2635) );
  buffer buf_n2636( .i (n2635), .o (n2636) );
  buffer buf_n2637( .i (n2636), .o (n2637) );
  assign n2638 = ( n2611 & n2630 ) | ( n2611 & ~n2637 ) | ( n2630 & ~n2637 ) ;
  buffer buf_n2639( .i (n754), .o (n2639) );
  assign n2640 = ( n2280 & n2597 ) | ( n2280 & n2639 ) | ( n2597 & n2639 ) ;
  buffer buf_n2641( .i (n2639), .o (n2641) );
  assign n2642 = n2640 & ~n2641 ;
  buffer buf_n2643( .i (n2642), .o (n2643) );
  buffer buf_n2644( .i (n2643), .o (n2644) );
  buffer buf_n2645( .i (n2644), .o (n2645) );
  buffer buf_n2646( .i (n2645), .o (n2646) );
  buffer buf_n2647( .i (n2646), .o (n2647) );
  buffer buf_n2648( .i (n2647), .o (n2648) );
  buffer buf_n2649( .i (n2648), .o (n2649) );
  buffer buf_n2650( .i (n2649), .o (n2650) );
  buffer buf_n2651( .i (n2650), .o (n2651) );
  buffer buf_n2652( .i (n2651), .o (n2652) );
  buffer buf_n2653( .i (n2652), .o (n2653) );
  buffer buf_n2654( .i (n2653), .o (n2654) );
  buffer buf_n596( .i (n595), .o (n596) );
  assign n2655 = n596 & n2351 ;
  buffer buf_n2656( .i (n2353), .o (n2656) );
  assign n2657 = ( n2489 & n2655 ) | ( n2489 & n2656 ) | ( n2655 & n2656 ) ;
  assign n2658 = ~n2490 & n2657 ;
  buffer buf_n2659( .i (n2658), .o (n2659) );
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2660), .o (n2661) );
  buffer buf_n2662( .i (n2661), .o (n2662) );
  buffer buf_n2663( .i (n2662), .o (n2663) );
  buffer buf_n2664( .i (n2663), .o (n2664) );
  buffer buf_n2665( .i (n2664), .o (n2665) );
  buffer buf_n2668( .i (n558), .o (n2668) );
  assign n2669 = ( n1364 & n2345 ) | ( n1364 & ~n2668 ) | ( n2345 & ~n2668 ) ;
  assign n2670 = ~n1933 & n2669 ;
  buffer buf_n2671( .i (n2670), .o (n2671) );
  buffer buf_n2672( .i (n2671), .o (n2672) );
  buffer buf_n2673( .i (n2672), .o (n2673) );
  buffer buf_n2674( .i (n2673), .o (n2674) );
  assign n2680 = n2488 & n2674 ;
  assign n2681 = ( n1735 & n2656 ) | ( n1735 & n2680 ) | ( n2656 & n2680 ) ;
  assign n2682 = ~n1821 & n2681 ;
  buffer buf_n2683( .i (n2682), .o (n2683) );
  buffer buf_n2684( .i (n2683), .o (n2684) );
  buffer buf_n2685( .i (n2684), .o (n2685) );
  buffer buf_n2686( .i (n2685), .o (n2686) );
  buffer buf_n2687( .i (n2686), .o (n2687) );
  buffer buf_n2688( .i (n2687), .o (n2688) );
  assign n2693 = n2118 & n2674 ;
  assign n2694 = ( n2489 & n2656 ) | ( n2489 & n2693 ) | ( n2656 & n2693 ) ;
  assign n2695 = ~n2490 & n2694 ;
  buffer buf_n2696( .i (n2695), .o (n2696) );
  buffer buf_n2697( .i (n2696), .o (n2697) );
  buffer buf_n2698( .i (n2697), .o (n2698) );
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n2700( .i (n2699), .o (n2700) );
  assign n2705 = n1856 | n2249 ;
  buffer buf_n2706( .i (n1933), .o (n2706) );
  buffer buf_n2707( .i (n530), .o (n2707) );
  assign n2708 = ( n2705 & ~n2706 ) | ( n2705 & n2707 ) | ( ~n2706 & n2707 ) ;
  buffer buf_n2709( .i (n2706), .o (n2709) );
  assign n2710 = n2708 | n2709 ;
  buffer buf_n2711( .i (n2710), .o (n2711) );
  buffer buf_n2712( .i (n2711), .o (n2712) );
  buffer buf_n2714( .i (n2283), .o (n2714) );
  assign n2715 = ~n2712 & n2714 ;
  buffer buf_n2716( .i (n2118), .o (n2716) );
  assign n2717 = ( n2656 & n2715 ) | ( n2656 & n2716 ) | ( n2715 & n2716 ) ;
  buffer buf_n2718( .i (n2716), .o (n2718) );
  assign n2719 = n2717 & ~n2718 ;
  buffer buf_n2720( .i (n2719), .o (n2720) );
  buffer buf_n2721( .i (n2720), .o (n2721) );
  buffer buf_n2727( .i (n2412), .o (n2727) );
  assign n2728 = ~n2712 & n2727 ;
  buffer buf_n2729( .i (n2353), .o (n2729) );
  assign n2730 = ( n2489 & n2728 ) | ( n2489 & n2729 ) | ( n2728 & n2729 ) ;
  assign n2731 = ~n2490 & n2730 ;
  buffer buf_n2732( .i (n2731), .o (n2732) );
  buffer buf_n2733( .i (n2732), .o (n2733) );
  assign n2740 = n2721 | n2733 ;
  buffer buf_n2741( .i (n2740), .o (n2741) );
  buffer buf_n2742( .i (n2741), .o (n2742) );
  assign n2743 = n2700 | n2742 ;
  assign n2744 = ( ~n2664 & n2688 ) | ( ~n2664 & n2743 ) | ( n2688 & n2743 ) ;
  assign n2745 = n2665 | n2744 ;
  assign n2746 = n2654 | n2745 ;
  assign n2747 = ( ~n2588 & n2638 ) | ( ~n2588 & n2746 ) | ( n2638 & n2746 ) ;
  assign n2748 = n2589 | n2747 ;
  assign n2749 = n534 & n1225 ;
  assign n2750 = ( n2117 & n2727 ) | ( n2117 & n2749 ) | ( n2727 & n2749 ) ;
  assign n2751 = ~n2716 & n2750 ;
  buffer buf_n2752( .i (n2751), .o (n2752) );
  assign n2755 = ~n819 & n2752 ;
  buffer buf_n2756( .i (n2755), .o (n2756) );
  buffer buf_n2757( .i (n2756), .o (n2757) );
  buffer buf_n2758( .i (n2757), .o (n2758) );
  buffer buf_n2759( .i (n2758), .o (n2759) );
  buffer buf_n2760( .i (n2759), .o (n2760) );
  buffer buf_n2761( .i (n2760), .o (n2761) );
  buffer buf_n2762( .i (n2761), .o (n2762) );
  buffer buf_n2763( .i (n2762), .o (n2763) );
  assign n2764 = ( n1252 & n2345 ) | ( n1252 & n2594 ) | ( n2345 & n2594 ) ;
  buffer buf_n2765( .i (n2594), .o (n2765) );
  assign n2766 = n2764 & ~n2765 ;
  buffer buf_n2767( .i (n2766), .o (n2767) );
  buffer buf_n2772( .i (n811), .o (n2772) );
  buffer buf_n2773( .i (n2772), .o (n2773) );
  assign n2774 = n2767 & ~n2773 ;
  assign n2775 = ( n2441 & n2641 ) | ( n2441 & n2774 ) | ( n2641 & n2774 ) ;
  buffer buf_n2776( .i (n2641), .o (n2776) );
  assign n2777 = n2775 & ~n2776 ;
  buffer buf_n2778( .i (n2777), .o (n2778) );
  buffer buf_n2779( .i (n2778), .o (n2779) );
  buffer buf_n2780( .i (n2779), .o (n2780) );
  buffer buf_n2781( .i (n2780), .o (n2781) );
  buffer buf_n2782( .i (n2781), .o (n2782) );
  buffer buf_n2783( .i (n2782), .o (n2783) );
  buffer buf_n2784( .i (n2783), .o (n2784) );
  buffer buf_n2785( .i (n2784), .o (n2785) );
  buffer buf_n2786( .i (n2785), .o (n2786) );
  buffer buf_n2787( .i (n2786), .o (n2787) );
  buffer buf_n2788( .i (n2787), .o (n2788) );
  assign n2789 = n1225 & n2776 ;
  buffer buf_n2790( .i (n2441), .o (n2790) );
  buffer buf_n2791( .i (n2790), .o (n2791) );
  assign n2792 = ( n2714 & n2789 ) | ( n2714 & n2791 ) | ( n2789 & n2791 ) ;
  buffer buf_n2793( .i (n2714), .o (n2793) );
  assign n2794 = n2792 & ~n2793 ;
  buffer buf_n2795( .i (n2794), .o (n2795) );
  buffer buf_n2796( .i (n2795), .o (n2796) );
  buffer buf_n2797( .i (n2796), .o (n2797) );
  buffer buf_n2798( .i (n2797), .o (n2798) );
  buffer buf_n2799( .i (n2798), .o (n2799) );
  buffer buf_n2800( .i (n2799), .o (n2800) );
  buffer buf_n2801( .i (n2800), .o (n2801) );
  buffer buf_n2802( .i (n2801), .o (n2802) );
  assign n2803 = ( n2591 & n2616 ) | ( n2591 & n2639 ) | ( n2616 & n2639 ) ;
  assign n2804 = ~n2641 & n2803 ;
  buffer buf_n2805( .i (n2804), .o (n2805) );
  assign n2811 = ~n2714 & n2805 ;
  buffer buf_n2812( .i (n2811), .o (n2812) );
  buffer buf_n2813( .i (n2812), .o (n2813) );
  buffer buf_n2814( .i (n2813), .o (n2814) );
  buffer buf_n2815( .i (n2814), .o (n2815) );
  buffer buf_n2816( .i (n2815), .o (n2816) );
  assign n2819 = n2345 & n2668 ;
  buffer buf_n2820( .i (n2502), .o (n2820) );
  buffer buf_n2821( .i (n2820), .o (n2821) );
  assign n2822 = ( n2765 & n2819 ) | ( n2765 & n2821 ) | ( n2819 & n2821 ) ;
  assign n2823 = ~n1857 & n2822 ;
  assign n2824 = ( n2114 & n2639 ) | ( n2114 & n2823 ) | ( n2639 & n2823 ) ;
  buffer buf_n2825( .i (n752), .o (n2825) );
  buffer buf_n2826( .i (n2825), .o (n2826) );
  buffer buf_n2827( .i (n2826), .o (n2827) );
  buffer buf_n2828( .i (n2827), .o (n2828) );
  assign n2829 = n2824 & ~n2828 ;
  buffer buf_n2830( .i (n2829), .o (n2830) );
  buffer buf_n2831( .i (n2830), .o (n2831) );
  buffer buf_n2832( .i (n2831), .o (n2832) );
  buffer buf_n2836( .i (n2793), .o (n2836) );
  assign n2837 = n2832 & ~n2836 ;
  buffer buf_n2838( .i (n2837), .o (n2838) );
  buffer buf_n2839( .i (n2838), .o (n2839) );
  buffer buf_n2840( .i (n2839), .o (n2840) );
  assign n2845 = n2816 | n2840 ;
  buffer buf_n2846( .i (n2845), .o (n2846) );
  buffer buf_n2847( .i (n2846), .o (n2847) );
  buffer buf_n2848( .i (n2847), .o (n2848) );
  assign n2849 = n2802 | n2848 ;
  assign n2850 = ( ~n2762 & n2788 ) | ( ~n2762 & n2849 ) | ( n2788 & n2849 ) ;
  assign n2851 = n2763 | n2850 ;
  assign n2852 = n1985 & n2347 ;
  buffer buf_n2853( .i (n2852), .o (n2853) );
  assign n2854 = ( n625 & n2828 ) | ( n625 & n2853 ) | ( n2828 & n2853 ) ;
  assign n2855 = ~n2776 & n2854 ;
  assign n2856 = n1233 & n2855 ;
  buffer buf_n2857( .i (n2856), .o (n2857) );
  buffer buf_n2858( .i (n2857), .o (n2858) );
  buffer buf_n2859( .i (n2858), .o (n2859) );
  buffer buf_n2860( .i (n2859), .o (n2860) );
  buffer buf_n2861( .i (n2860), .o (n2861) );
  buffer buf_n2862( .i (n2861), .o (n2862) );
  buffer buf_n2863( .i (n2862), .o (n2863) );
  buffer buf_n2864( .i (n2863), .o (n2864) );
  buffer buf_n2865( .i (n2864), .o (n2865) );
  buffer buf_n2866( .i (n2865), .o (n2866) );
  buffer buf_n2867( .i (n2866), .o (n2867) );
  buffer buf_n2100( .i (n2099), .o (n2100) );
  buffer buf_n2101( .i (n2100), .o (n2101) );
  assign n2868 = ( n2101 & n2499 ) | ( n2101 & n2501 ) | ( n2499 & n2501 ) ;
  assign n2869 = ~n2343 & n2868 ;
  buffer buf_n2870( .i (n2869), .o (n2870) );
  buffer buf_n2871( .i (n2870), .o (n2871) );
  buffer buf_n2872( .i (n2871), .o (n2872) );
  buffer buf_n2873( .i (n2872), .o (n2873) );
  assign n2882 = ~n2516 & n2873 ;
  assign n2883 = ( n707 & n2790 ) | ( n707 & n2882 ) | ( n2790 & n2882 ) ;
  assign n2884 = ~n708 & n2883 ;
  buffer buf_n2885( .i (n2884), .o (n2885) );
  assign n2894 = n706 & n2873 ;
  buffer buf_n2895( .i (n2516), .o (n2895) );
  assign n2896 = ( n2790 & n2894 ) | ( n2790 & n2895 ) | ( n2894 & n2895 ) ;
  buffer buf_n2897( .i (n2895), .o (n2897) );
  assign n2898 = n2896 & ~n2897 ;
  buffer buf_n2899( .i (n2898), .o (n2899) );
  assign n2907 = n2885 | n2899 ;
  buffer buf_n2908( .i (n2907), .o (n2908) );
  buffer buf_n2909( .i (n2908), .o (n2909) );
  buffer buf_n2910( .i (n2909), .o (n2910) );
  buffer buf_n2911( .i (n2910), .o (n2911) );
  buffer buf_n2912( .i (n2911), .o (n2912) );
  buffer buf_n2913( .i (n2912), .o (n2913) );
  buffer buf_n2914( .i (n2913), .o (n2914) );
  buffer buf_n2915( .i (n2914), .o (n2915) );
  buffer buf_n2874( .i (n2873), .o (n2874) );
  buffer buf_n2875( .i (n2874), .o (n2875) );
  buffer buf_n2876( .i (n2875), .o (n2876) );
  assign n2917 = n705 & n2773 ;
  buffer buf_n2918( .i (n2917), .o (n2918) );
  buffer buf_n2919( .i (n2918), .o (n2919) );
  assign n2920 = ( n2791 & ~n2875 ) | ( n2791 & n2919 ) | ( ~n2875 & n2919 ) ;
  assign n2921 = n2876 & n2920 ;
  buffer buf_n2922( .i (n2921), .o (n2922) );
  buffer buf_n2923( .i (n2922), .o (n2923) );
  buffer buf_n2924( .i (n2923), .o (n2924) );
  buffer buf_n2925( .i (n2924), .o (n2925) );
  buffer buf_n2926( .i (n2925), .o (n2926) );
  buffer buf_n2927( .i (n2926), .o (n2927) );
  buffer buf_n2928( .i (n2927), .o (n2928) );
  buffer buf_n2929( .i (n2928), .o (n2929) );
  assign n2934 = ( n594 & n2828 ) | ( n594 & n2853 ) | ( n2828 & n2853 ) ;
  assign n2935 = ~n2776 & n2934 ;
  assign n2936 = n1233 & n2935 ;
  buffer buf_n2937( .i (n2936), .o (n2937) );
  assign n2946 = n650 & n2873 ;
  assign n2947 = ( n2790 & n2895 ) | ( n2790 & n2946 ) | ( n2895 & n2946 ) ;
  assign n2948 = ~n2897 & n2947 ;
  buffer buf_n2949( .i (n2948), .o (n2949) );
  assign n2961 = n2937 | n2949 ;
  buffer buf_n2962( .i (n2961), .o (n2962) );
  buffer buf_n2963( .i (n2962), .o (n2963) );
  buffer buf_n2964( .i (n2963), .o (n2964) );
  buffer buf_n2965( .i (n2964), .o (n2965) );
  buffer buf_n2966( .i (n2965), .o (n2966) );
  buffer buf_n2967( .i (n2966), .o (n2967) );
  buffer buf_n2968( .i (n2967), .o (n2968) );
  assign n2969 = n2929 | n2968 ;
  assign n2970 = ( ~n2866 & n2915 ) | ( ~n2866 & n2969 ) | ( n2915 & n2969 ) ;
  assign n2971 = n2867 | n2970 ;
  assign n2972 = n2851 | n2971 ;
  assign n2973 = ( ~n2571 & n2748 ) | ( ~n2571 & n2972 ) | ( n2748 & n2972 ) ;
  assign n2974 = n2572 | n2973 ;
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  assign n2975 = ~n1209 & n2174 ;
  assign n2976 = n1186 & n2975 ;
  buffer buf_n2977( .i (n2976), .o (n2977) );
  buffer buf_n2978( .i (n2977), .o (n2978) );
  buffer buf_n2979( .i (n2978), .o (n2979) );
  buffer buf_n2980( .i (n2979), .o (n2980) );
  buffer buf_n2981( .i (n2980), .o (n2981) );
  buffer buf_n2982( .i (n2981), .o (n2982) );
  buffer buf_n2983( .i (n2982), .o (n2983) );
  buffer buf_n2984( .i (n2983), .o (n2984) );
  buffer buf_n2985( .i (n2984), .o (n2985) );
  buffer buf_n2986( .i (n2985), .o (n2986) );
  buffer buf_n2987( .i (n2986), .o (n2987) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n2988( .i (n149), .o (n2988) );
  buffer buf_n2989( .i (n2765), .o (n2989) );
  assign n2990 = ( n1662 & n2988 ) | ( n1662 & n2989 ) | ( n2988 & n2989 ) ;
  assign n2991 = ~n151 & n2990 ;
  buffer buf_n2992( .i (n783), .o (n2992) );
  assign n2993 = n2991 & ~n2992 ;
  buffer buf_n2994( .i (n732), .o (n2994) );
  assign n2995 = ( n1863 & n2993 ) | ( n1863 & n2994 ) | ( n2993 & n2994 ) ;
  buffer buf_n2996( .i (n1863), .o (n2996) );
  assign n2997 = n2995 & ~n2996 ;
  assign n2998 = ~n2793 & n2997 ;
  buffer buf_n2999( .i (n2998), .o (n2999) );
  buffer buf_n3000( .i (n2999), .o (n3000) );
  buffer buf_n3001( .i (n3000), .o (n3001) );
  buffer buf_n3002( .i (n3001), .o (n3002) );
  buffer buf_n3003( .i (n3002), .o (n3003) );
  assign n3009 = n2495 | n3003 ;
  buffer buf_n3010( .i (n3009), .o (n3010) );
  buffer buf_n3011( .i (n3010), .o (n3011) );
  buffer buf_n3012( .i (n3011), .o (n3012) );
  buffer buf_n2470( .i (n2469), .o (n2470) );
  buffer buf_n2471( .i (n2470), .o (n2471) );
  buffer buf_n2472( .i (n2471), .o (n2472) );
  buffer buf_n2473( .i (n2472), .o (n2473) );
  buffer buf_n2474( .i (n2473), .o (n2474) );
  buffer buf_n2231( .i (n2230), .o (n2231) );
  assign n3013 = ~n2773 & n2827 ;
  buffer buf_n3014( .i (n3013), .o (n3014) );
  buffer buf_n3015( .i (n3014), .o (n3015) );
  buffer buf_n3016( .i (n3015), .o (n3016) );
  assign n3021 = ( n2231 & n2729 ) | ( n2231 & n3016 ) | ( n2729 & n3016 ) ;
  assign n3022 = ~n2312 & n3021 ;
  buffer buf_n3023( .i (n3022), .o (n3023) );
  buffer buf_n3024( .i (n3023), .o (n3024) );
  buffer buf_n3025( .i (n3024), .o (n3025) );
  buffer buf_n3026( .i (n3025), .o (n3026) );
  buffer buf_n3027( .i (n3026), .o (n3027) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  assign n3032 = n2515 & ~n2992 ;
  assign n3033 = ~n2895 & n3032 ;
  buffer buf_n3034( .i (n3033), .o (n3034) );
  buffer buf_n3035( .i (n3034), .o (n3035) );
  buffer buf_n3036( .i (n3035), .o (n3036) );
  buffer buf_n3037( .i (n3036), .o (n3037) );
  buffer buf_n3038( .i (n3037), .o (n3038) );
  assign n3044 = n2547 | n3038 ;
  buffer buf_n3045( .i (n3044), .o (n3045) );
  assign n3049 = n2317 | n3045 ;
  assign n3050 = ( ~n2240 & n3027 ) | ( ~n2240 & n3049 ) | ( n3027 & n3049 ) ;
  assign n3051 = n2241 | n3050 ;
  assign n3052 = n2474 | n3051 ;
  assign n3053 = ( ~n2986 & n3012 ) | ( ~n2986 & n3052 ) | ( n3012 & n3052 ) ;
  assign n3054 = n2987 | n3053 ;
  buffer buf_n3055( .i (n3054), .o (n3055) );
  buffer buf_n3056( .i (n3055), .o (n3056) );
  buffer buf_n2689( .i (n2688), .o (n2689) );
  buffer buf_n2690( .i (n2689), .o (n2690) );
  buffer buf_n2691( .i (n2690), .o (n2691) );
  buffer buf_n2692( .i (n2691), .o (n2692) );
  buffer buf_n2701( .i (n2700), .o (n2701) );
  buffer buf_n2702( .i (n2701), .o (n2702) );
  buffer buf_n2703( .i (n2702), .o (n2703) );
  buffer buf_n2704( .i (n2703), .o (n2704) );
  buffer buf_n2734( .i (n2733), .o (n2734) );
  buffer buf_n2735( .i (n2734), .o (n2735) );
  buffer buf_n2736( .i (n2735), .o (n2736) );
  buffer buf_n2737( .i (n2736), .o (n2737) );
  buffer buf_n2738( .i (n2737), .o (n2738) );
  buffer buf_n2739( .i (n2738), .o (n2739) );
  buffer buf_n2722( .i (n2721), .o (n2722) );
  buffer buf_n2723( .i (n2722), .o (n2723) );
  buffer buf_n2724( .i (n2723), .o (n2724) );
  buffer buf_n2725( .i (n2724), .o (n2725) );
  buffer buf_n2726( .i (n2725), .o (n2726) );
  assign n3057 = n2586 | n2726 ;
  assign n3058 = n2739 | n3057 ;
  assign n3059 = n2704 | n3058 ;
  assign n3060 = n2692 | n3059 ;
  assign n3061 = n819 & n2752 ;
  buffer buf_n3062( .i (n3061), .o (n3062) );
  buffer buf_n3063( .i (n3062), .o (n3063) );
  buffer buf_n3064( .i (n3063), .o (n3064) );
  buffer buf_n3065( .i (n3064), .o (n3065) );
  buffer buf_n3066( .i (n3065), .o (n3066) );
  assign n3069 = ( ~n1227 & n1436 ) | ( ~n1227 & n2729 ) | ( n1436 & n2729 ) ;
  assign n3070 = n1228 & n3069 ;
  buffer buf_n3071( .i (n3070), .o (n3071) );
  buffer buf_n3072( .i (n3071), .o (n3072) );
  buffer buf_n3073( .i (n3072), .o (n3073) );
  assign n3076 = n2757 | n3073 ;
  assign n3077 = n2799 | n3076 ;
  buffer buf_n2768( .i (n2767), .o (n2768) );
  assign n3078 = n2516 & n2768 ;
  buffer buf_n3079( .i (n2828), .o (n3079) );
  buffer buf_n3080( .i (n2992), .o (n3080) );
  assign n3081 = ( n3078 & n3079 ) | ( n3078 & n3080 ) | ( n3079 & n3080 ) ;
  assign n3082 = ~n2727 & n3081 ;
  buffer buf_n3083( .i (n3082), .o (n3083) );
  buffer buf_n3084( .i (n3083), .o (n3084) );
  buffer buf_n3085( .i (n3084), .o (n3085) );
  buffer buf_n3086( .i (n3085), .o (n3086) );
  buffer buf_n3087( .i (n3086), .o (n3087) );
  buffer buf_n2806( .i (n2805), .o (n2806) );
  buffer buf_n2807( .i (n2806), .o (n2807) );
  buffer buf_n2808( .i (n2807), .o (n2808) );
  buffer buf_n2809( .i (n2808), .o (n2809) );
  buffer buf_n2810( .i (n2809), .o (n2810) );
  buffer buf_n2833( .i (n2832), .o (n2833) );
  buffer buf_n2834( .i (n2833), .o (n2834) );
  buffer buf_n2835( .i (n2834), .o (n2835) );
  assign n3088 = n2810 | n2835 ;
  assign n3089 = n3087 | n3088 ;
  assign n3090 = n2784 | n3089 ;
  assign n3091 = ( ~n3065 & n3077 ) | ( ~n3065 & n3090 ) | ( n3077 & n3090 ) ;
  assign n3092 = n3066 | n3091 ;
  buffer buf_n3093( .i (n3092), .o (n3093) );
  buffer buf_n3094( .i (n3093), .o (n3094) );
  buffer buf_n2950( .i (n2949), .o (n2950) );
  buffer buf_n2951( .i (n2950), .o (n2951) );
  assign n3095 = n2923 | n2951 ;
  buffer buf_n3096( .i (n3095), .o (n3096) );
  buffer buf_n3097( .i (n3096), .o (n3097) );
  buffer buf_n3098( .i (n3097), .o (n3098) );
  buffer buf_n3099( .i (n3098), .o (n3099) );
  buffer buf_n3100( .i (n3099), .o (n3100) );
  buffer buf_n3101( .i (n3100), .o (n3101) );
  assign n3102 = n624 & n1217 ;
  buffer buf_n3103( .i (n2573), .o (n3103) );
  assign n3104 = ( n1731 & n3102 ) | ( n1731 & n3103 ) | ( n3102 & n3103 ) ;
  buffer buf_n3105( .i (n3103), .o (n3105) );
  assign n3106 = n3104 & ~n3105 ;
  assign n3107 = ~n2897 & n3106 ;
  assign n3108 = ( n2716 & n2729 ) | ( n2716 & n3107 ) | ( n2729 & n3107 ) ;
  assign n3109 = ~n2718 & n3108 ;
  buffer buf_n3110( .i (n3109), .o (n3110) );
  buffer buf_n3111( .i (n3110), .o (n3111) );
  buffer buf_n3112( .i (n3111), .o (n3112) );
  buffer buf_n3113( .i (n3112), .o (n3113) );
  buffer buf_n3114( .i (n3113), .o (n3114) );
  assign n3116 = n592 & n1216 ;
  assign n3117 = ( n1987 & n2573 ) | ( n1987 & n3116 ) | ( n2573 & n3116 ) ;
  assign n3118 = ~n3103 & n3117 ;
  buffer buf_n3119( .i (n2773), .o (n3119) );
  buffer buf_n3120( .i (n3119), .o (n3120) );
  assign n3121 = n3118 & ~n3120 ;
  assign n3122 = ( n2727 & n2791 ) | ( n2727 & n3121 ) | ( n2791 & n3121 ) ;
  buffer buf_n3123( .i (n3079), .o (n3123) );
  buffer buf_n3124( .i (n3123), .o (n3124) );
  assign n3125 = n3122 & ~n3124 ;
  buffer buf_n3126( .i (n3125), .o (n3126) );
  buffer buf_n3127( .i (n3126), .o (n3127) );
  buffer buf_n3128( .i (n3127), .o (n3128) );
  buffer buf_n3129( .i (n3128), .o (n3129) );
  buffer buf_n3130( .i (n3129), .o (n3130) );
  buffer buf_n2938( .i (n2937), .o (n2938) );
  buffer buf_n2939( .i (n2938), .o (n2939) );
  buffer buf_n2877( .i (n2876), .o (n2877) );
  buffer buf_n3134( .i (n2791), .o (n3134) );
  assign n3135 = ( n1276 & ~n2876 ) | ( n1276 & n3134 ) | ( ~n2876 & n3134 ) ;
  assign n3136 = n2877 & n3135 ;
  buffer buf_n3137( .i (n3136), .o (n3137) );
  assign n3144 = n2939 | n3137 ;
  buffer buf_n3145( .i (n3144), .o (n3145) );
  buffer buf_n3146( .i (n3145), .o (n3146) );
  assign n3147 = n3130 | n3146 ;
  assign n3148 = ( ~n2863 & n3114 ) | ( ~n2863 & n3147 ) | ( n3114 & n3147 ) ;
  assign n3149 = n2864 | n3148 ;
  buffer buf_n2900( .i (n2899), .o (n2900) );
  buffer buf_n2901( .i (n2900), .o (n2901) );
  buffer buf_n2902( .i (n2901), .o (n2902) );
  buffer buf_n2903( .i (n2902), .o (n2903) );
  buffer buf_n2904( .i (n2903), .o (n2904) );
  buffer buf_n2905( .i (n2904), .o (n2905) );
  buffer buf_n2906( .i (n2905), .o (n2906) );
  buffer buf_n2886( .i (n2885), .o (n2886) );
  buffer buf_n2887( .i (n2886), .o (n2887) );
  buffer buf_n2888( .i (n2887), .o (n2888) );
  buffer buf_n2889( .i (n2888), .o (n2889) );
  buffer buf_n2890( .i (n2889), .o (n2890) );
  buffer buf_n2891( .i (n2890), .o (n2891) );
  buffer buf_n710( .i (n709), .o (n710) );
  assign n3150 = n2875 & n2897 ;
  assign n3151 = ( n709 & n3134 ) | ( n709 & n3150 ) | ( n3134 & n3150 ) ;
  assign n3152 = ~n710 & n3151 ;
  buffer buf_n3153( .i (n3152), .o (n3153) );
  buffer buf_n3154( .i (n3153), .o (n3154) );
  buffer buf_n3155( .i (n3154), .o (n3155) );
  buffer buf_n3156( .i (n3155), .o (n3156) );
  buffer buf_n3157( .i (n3156), .o (n3157) );
  assign n3159 = n2891 | n3157 ;
  assign n3160 = n2906 | n3159 ;
  assign n3161 = n3149 | n3160 ;
  assign n3162 = ( ~n3093 & n3101 ) | ( ~n3093 & n3161 ) | ( n3101 & n3161 ) ;
  assign n3163 = n3094 | n3162 ;
  buffer buf_n2612( .i (n2611), .o (n2612) );
  assign n3164 = n2602 & ~n2836 ;
  buffer buf_n3165( .i (n3164), .o (n3165) );
  buffer buf_n3166( .i (n3165), .o (n3166) );
  buffer buf_n3167( .i (n3166), .o (n3167) );
  buffer buf_n3168( .i (n3167), .o (n3168) );
  buffer buf_n3169( .i (n3168), .o (n3169) );
  buffer buf_n3170( .i (n3169), .o (n3170) );
  buffer buf_n3171( .i (n3170), .o (n3171) );
  buffer buf_n3172( .i (n3171), .o (n3172) );
  buffer buf_n3173( .i (n3172), .o (n3173) );
  assign n3174 = n2630 | n2654 ;
  assign n3175 = ( n2612 & ~n3173 ) | ( n2612 & n3174 ) | ( ~n3173 & n3174 ) ;
  assign n3176 = n3163 | n3175 ;
  assign n3177 = ( ~n3055 & n3060 ) | ( ~n3055 & n3176 ) | ( n3060 & n3176 ) ;
  assign n3178 = n3056 | n3177 ;
  buffer buf_n2475( .i (n2474), .o (n2475) );
  buffer buf_n2476( .i (n2475), .o (n2476) );
  assign n3179 = n2446 | n2999 ;
  buffer buf_n3180( .i (n3179), .o (n3180) );
  buffer buf_n3181( .i (n3180), .o (n3181) );
  buffer buf_n3182( .i (n3181), .o (n3182) );
  buffer buf_n3183( .i (n3182), .o (n3183) );
  buffer buf_n3184( .i (n3183), .o (n3184) );
  buffer buf_n3185( .i (n3184), .o (n3185) );
  buffer buf_n3186( .i (n3185), .o (n3186) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  assign n3187 = n2290 | n2557 ;
  assign n3188 = ( n2536 & ~n2549 ) | ( n2536 & n3187 ) | ( ~n2549 & n3187 ) ;
  assign n3189 = n2550 | n3188 ;
  assign n3190 = n2519 | n3034 ;
  buffer buf_n3191( .i (n3190), .o (n3191) );
  buffer buf_n3192( .i (n3191), .o (n3192) );
  buffer buf_n3193( .i (n3192), .o (n3193) );
  buffer buf_n3194( .i (n3193), .o (n3194) );
  buffer buf_n3195( .i (n3194), .o (n3195) );
  buffer buf_n3196( .i (n3195), .o (n3196) );
  assign n3201 = n2496 | n3196 ;
  assign n3202 = n3189 | n3201 ;
  buffer buf_n1210( .i (n1209), .o (n1210) );
  assign n3203 = ~n1185 & n2174 ;
  assign n3204 = ~n1210 & n3203 ;
  buffer buf_n3205( .i (n3204), .o (n3205) );
  buffer buf_n3206( .i (n3205), .o (n3206) );
  buffer buf_n3207( .i (n3206), .o (n3207) );
  buffer buf_n3208( .i (n3207), .o (n3208) );
  buffer buf_n3209( .i (n3208), .o (n3209) );
  buffer buf_n3210( .i (n3209), .o (n3210) );
  buffer buf_n3211( .i (n3210), .o (n3211) );
  buffer buf_n3212( .i (n3211), .o (n3212) );
  buffer buf_n2460( .i (n2459), .o (n2460) );
  buffer buf_n2461( .i (n2460), .o (n2461) );
  buffer buf_n2462( .i (n2461), .o (n2462) );
  assign n3213 = n2184 | n2462 ;
  assign n3214 = n3212 | n3213 ;
  assign n3215 = n3202 | n3214 ;
  assign n3216 = ( ~n2475 & n3186 ) | ( ~n2475 & n3215 ) | ( n3186 & n3215 ) ;
  assign n3217 = n2476 | n3216 ;
  buffer buf_n3218( .i (n3217), .o (n3218) );
  buffer buf_n3219( .i (n3218), .o (n3219) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n3028( .i (n3027), .o (n3028) );
  buffer buf_n3029( .i (n3028), .o (n3029) );
  buffer buf_n3030( .i (n3029), .o (n3030) );
  buffer buf_n3031( .i (n3030), .o (n3031) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  buffer buf_n2368( .i (n2367), .o (n2368) );
  buffer buf_n2369( .i (n2368), .o (n2369) );
  buffer buf_n2370( .i (n2369), .o (n2370) );
  assign n3220 = n2268 | n2370 ;
  assign n3221 = ( ~n2244 & n3031 ) | ( ~n2244 & n3220 ) | ( n3031 & n3220 ) ;
  assign n3222 = n2245 | n3221 ;
  buffer buf_n3223( .i (n3120), .o (n3223) );
  assign n3224 = n2600 & n3223 ;
  buffer buf_n3225( .i (n3224), .o (n3225) );
  buffer buf_n3226( .i (n3225), .o (n3226) );
  buffer buf_n3227( .i (n3226), .o (n3227) );
  buffer buf_n3228( .i (n3227), .o (n3228) );
  buffer buf_n3229( .i (n3228), .o (n3229) );
  buffer buf_n3230( .i (n3229), .o (n3230) );
  buffer buf_n3231( .i (n3230), .o (n3231) );
  buffer buf_n3232( .i (n3231), .o (n3232) );
  buffer buf_n3234( .i (n2836), .o (n3234) );
  assign n3235 = n2808 & n3234 ;
  buffer buf_n3236( .i (n3235), .o (n3236) );
  assign n3242 = n3166 | n3236 ;
  buffer buf_n3243( .i (n3242), .o (n3243) );
  buffer buf_n3244( .i (n3243), .o (n3244) );
  assign n3247 = n2830 & n3223 ;
  buffer buf_n3248( .i (n3247), .o (n3248) );
  buffer buf_n3249( .i (n3248), .o (n3249) );
  assign n3260 = n2813 | n3249 ;
  buffer buf_n3261( .i (n3260), .o (n3261) );
  buffer buf_n3262( .i (n3261), .o (n3262) );
  buffer buf_n3263( .i (n3262), .o (n3263) );
  assign n3264 = n2840 | n3087 ;
  assign n3265 = n3263 | n3264 ;
  assign n3266 = ( ~n3231 & n3244 ) | ( ~n3231 & n3265 ) | ( n3244 & n3265 ) ;
  assign n3267 = n3232 | n3266 ;
  buffer buf_n3268( .i (n3267), .o (n3268) );
  buffer buf_n3269( .i (n3268), .o (n3269) );
  assign n3270 = n2796 | n3110 ;
  buffer buf_n3271( .i (n3270), .o (n3271) );
  assign n3272 = n3073 | n3271 ;
  buffer buf_n3273( .i (n3272), .o (n3273) );
  assign n3277 = n3065 | n3273 ;
  assign n3278 = ( ~n2760 & n2786 ) | ( ~n2760 & n3277 ) | ( n2786 & n3277 ) ;
  assign n3279 = n2761 | n3278 ;
  assign n3280 = n2643 & n3223 ;
  buffer buf_n3281( .i (n3280), .o (n3281) );
  buffer buf_n3282( .i (n3281), .o (n3282) );
  buffer buf_n3283( .i (n3282), .o (n3283) );
  buffer buf_n3284( .i (n3283), .o (n3284) );
  buffer buf_n3285( .i (n3284), .o (n3285) );
  buffer buf_n3286( .i (n3285), .o (n3286) );
  buffer buf_n3287( .i (n3286), .o (n3287) );
  buffer buf_n3288( .i (n3287), .o (n3288) );
  assign n3289 = ( n1462 & n2765 ) | ( n1462 & n2821 ) | ( n2765 & n2821 ) ;
  assign n3290 = ~n2707 & n3289 ;
  buffer buf_n3291( .i (n3290), .o (n3291) );
  buffer buf_n3292( .i (n3291), .o (n3292) );
  assign n3294 = ( n676 & n1395 ) | ( n676 & ~n3291 ) | ( n1395 & ~n3291 ) ;
  assign n3295 = n3292 & n3294 ;
  buffer buf_n3296( .i (n3295), .o (n3296) );
  buffer buf_n3297( .i (n3296), .o (n3297) );
  buffer buf_n3298( .i (n3297), .o (n3298) );
  buffer buf_n3299( .i (n3298), .o (n3299) );
  buffer buf_n3300( .i (n3299), .o (n3300) );
  buffer buf_n3301( .i (n3300), .o (n3301) );
  buffer buf_n3302( .i (n3301), .o (n3302) );
  buffer buf_n3303( .i (n3302), .o (n3303) );
  assign n3306 = ( n1269 & n2573 ) | ( n1269 & n2709 ) | ( n2573 & n2709 ) ;
  assign n3307 = ~n3103 & n3306 ;
  buffer buf_n3308( .i (n3307), .o (n3308) );
  assign n3312 = n3223 & n3308 ;
  assign n3313 = n709 & n3312 ;
  buffer buf_n3314( .i (n3313), .o (n3314) );
  buffer buf_n3315( .i (n3314), .o (n3315) );
  buffer buf_n3316( .i (n3315), .o (n3316) );
  buffer buf_n3317( .i (n3316), .o (n3317) );
  buffer buf_n3318( .i (n3317), .o (n3318) );
  assign n3321 = ( n2625 & ~n2632 ) | ( n2625 & n2649 ) | ( ~n2632 & n2649 ) ;
  assign n3322 = n3318 | n3321 ;
  assign n3323 = ( ~n3287 & n3303 ) | ( ~n3287 & n3322 ) | ( n3303 & n3322 ) ;
  assign n3324 = n3288 | n3323 ;
  buffer buf_n3131( .i (n3130), .o (n3131) );
  buffer buf_n3132( .i (n3131), .o (n3132) );
  buffer buf_n3138( .i (n3137), .o (n3138) );
  buffer buf_n3139( .i (n3138), .o (n3139) );
  buffer buf_n3140( .i (n3139), .o (n3140) );
  buffer buf_n3141( .i (n3140), .o (n3141) );
  buffer buf_n2952( .i (n2951), .o (n2952) );
  buffer buf_n2953( .i (n2952), .o (n2953) );
  buffer buf_n2954( .i (n2953), .o (n2954) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n2878( .i (n2877), .o (n2878) );
  buffer buf_n2879( .i (n2878), .o (n2879) );
  buffer buf_n2880( .i (n2879), .o (n2880) );
  buffer buf_n2881( .i (n2880), .o (n2881) );
  assign n3325 = n792 & n2881 ;
  assign n3326 = n2954 | n3325 ;
  assign n3327 = ( ~n3131 & n3141 ) | ( ~n3131 & n3326 ) | ( n3141 & n3326 ) ;
  assign n3328 = n3132 | n3327 ;
  assign n3329 = n3324 | n3328 ;
  assign n3330 = ( ~n3268 & n3279 ) | ( ~n3268 & n3329 ) | ( n3279 & n3329 ) ;
  assign n3331 = n3269 | n3330 ;
  buffer buf_n2666( .i (n2665), .o (n2666) );
  buffer buf_n2667( .i (n2666), .o (n2667) );
  buffer buf_n3332( .i (n3120), .o (n3332) );
  assign n3333 = n2576 & n3332 ;
  buffer buf_n3334( .i (n3333), .o (n3334) );
  assign n3339 = n2312 & n3334 ;
  buffer buf_n3340( .i (n3339), .o (n3340) );
  buffer buf_n3341( .i (n3340), .o (n3341) );
  buffer buf_n3342( .i (n3341), .o (n3342) );
  buffer buf_n3343( .i (n3342), .o (n3343) );
  buffer buf_n3344( .i (n3343), .o (n3344) );
  assign n3345 = n2583 | n2741 ;
  assign n3346 = n3344 | n3345 ;
  buffer buf_n3347( .i (n3346), .o (n3347) );
  assign n3348 = n2702 | n3347 ;
  assign n3349 = ( ~n2666 & n2690 ) | ( ~n2666 & n3348 ) | ( n2690 & n3348 ) ;
  assign n3350 = n2667 | n3349 ;
  assign n3351 = n3331 | n3350 ;
  assign n3352 = ( ~n3218 & n3222 ) | ( ~n3218 & n3351 ) | ( n3222 & n3351 ) ;
  assign n3353 = n3219 | n3352 ;
  buffer buf_n2223( .i (n2222), .o (n2223) );
  buffer buf_n2224( .i (n2223), .o (n2224) );
  buffer buf_n2225( .i (n2224), .o (n2225) );
  buffer buf_n3354( .i (n3134), .o (n3354) );
  assign n3355 = ( n1758 & n2511 ) | ( n1758 & n3354 ) | ( n2511 & n3354 ) ;
  assign n3356 = ~n2235 & n3355 ;
  buffer buf_n3357( .i (n3356), .o (n3357) );
  buffer buf_n3358( .i (n3357), .o (n3358) );
  buffer buf_n3359( .i (n3358), .o (n3359) );
  buffer buf_n3360( .i (n3359), .o (n3360) );
  buffer buf_n3361( .i (n3360), .o (n3361) );
  buffer buf_n3362( .i (n3361), .o (n3362) );
  buffer buf_n3363( .i (n3362), .o (n3363) );
  buffer buf_n3364( .i (n3363), .o (n3364) );
  buffer buf_n3365( .i (n3364), .o (n3365) );
  assign n3366 = n2258 | n2285 ;
  buffer buf_n3367( .i (n3366), .o (n3367) );
  buffer buf_n3368( .i (n3367), .o (n3368) );
  buffer buf_n3369( .i (n3368), .o (n3369) );
  buffer buf_n3370( .i (n3369), .o (n3370) );
  buffer buf_n3371( .i (n3370), .o (n3371) );
  buffer buf_n3372( .i (n3371), .o (n3372) );
  buffer buf_n3373( .i (n3372), .o (n3373) );
  buffer buf_n3374( .i (n3373), .o (n3374) );
  buffer buf_n3375( .i (n3374), .o (n3375) );
  buffer buf_n3376( .i (n3375), .o (n3376) );
  assign n3377 = n1867 & n2233 ;
  buffer buf_n3378( .i (n3377), .o (n3378) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n3385( .i (n1232), .o (n3385) );
  buffer buf_n3386( .i (n3385), .o (n3386) );
  assign n3387 = n2255 & n3386 ;
  buffer buf_n3388( .i (n3387), .o (n3388) );
  buffer buf_n3389( .i (n3388), .o (n3389) );
  assign n3399 = n3378 | n3389 ;
  assign n3400 = n3024 | n3399 ;
  buffer buf_n3401( .i (n3400), .o (n3401) );
  buffer buf_n3402( .i (n3401), .o (n3402) );
  buffer buf_n3403( .i (n3402), .o (n3403) );
  buffer buf_n3404( .i (n3403), .o (n3404) );
  buffer buf_n3405( .i (n3404), .o (n3405) );
  buffer buf_n2542( .i (n2541), .o (n2542) );
  assign n3406 = n2542 & n3386 ;
  buffer buf_n3407( .i (n3406), .o (n3407) );
  buffer buf_n3408( .i (n3407), .o (n3408) );
  buffer buf_n3409( .i (n3408), .o (n3409) );
  buffer buf_n3410( .i (n3409), .o (n3410) );
  buffer buf_n3411( .i (n3410), .o (n3411) );
  buffer buf_n3412( .i (n3411), .o (n3412) );
  buffer buf_n3413( .i (n3412), .o (n3413) );
  buffer buf_n3414( .i (n3413), .o (n3414) );
  buffer buf_n3039( .i (n3038), .o (n3039) );
  buffer buf_n3040( .i (n3039), .o (n3040) );
  buffer buf_n3041( .i (n3040), .o (n3041) );
  buffer buf_n3042( .i (n3041), .o (n3042) );
  buffer buf_n2537( .i (n2536), .o (n2537) );
  buffer buf_n2558( .i (n2557), .o (n2558) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n3293( .i (n3292), .o (n3293) );
  buffer buf_n3418( .i (n3080), .o (n3418) );
  assign n3419 = n3293 & ~n3418 ;
  assign n3420 = ( n679 & n2043 ) | ( n679 & n3419 ) | ( n2043 & n3419 ) ;
  assign n3421 = ~n567 & n3420 ;
  buffer buf_n3422( .i (n3421), .o (n3422) );
  assign n3425 = n820 & n3422 ;
  buffer buf_n3426( .i (n3425), .o (n3426) );
  buffer buf_n3427( .i (n3426), .o (n3427) );
  assign n3432 = n2558 | n3427 ;
  assign n3433 = n2537 | n3432 ;
  assign n3434 = n3042 | n3433 ;
  assign n3435 = n3414 | n3434 ;
  assign n3436 = n3405 | n3435 ;
  assign n3437 = ( ~n3364 & n3376 ) | ( ~n3364 & n3436 ) | ( n3376 & n3436 ) ;
  assign n3438 = n3365 | n3437 ;
  buffer buf_n2336( .i (n2335), .o (n2336) );
  buffer buf_n2337( .i (n2336), .o (n2337) );
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  buffer buf_n2340( .i (n2339), .o (n2340) );
  buffer buf_n2341( .i (n2340), .o (n2341) );
  assign n3439 = n146 & n2501 ;
  buffer buf_n3440( .i (n2499), .o (n3440) );
  assign n3441 = ( n2592 & n3439 ) | ( n2592 & n3440 ) | ( n3439 & n3440 ) ;
  buffer buf_n3442( .i (n3440), .o (n3442) );
  assign n3443 = n3441 & ~n3442 ;
  assign n3444 = n2825 & n3443 ;
  buffer buf_n3445( .i (n2668), .o (n3445) );
  buffer buf_n3446( .i (n3445), .o (n3446) );
  assign n3447 = ( n592 & n3444 ) | ( n592 & n3446 ) | ( n3444 & n3446 ) ;
  assign n3448 = ~n1987 & n3447 ;
  assign n3449 = n1231 & n3448 ;
  buffer buf_n3450( .i (n3449), .o (n3450) );
  buffer buf_n3451( .i (n3450), .o (n3451) );
  buffer buf_n3452( .i (n3451), .o (n3452) );
  buffer buf_n3453( .i (n3452), .o (n3453) );
  buffer buf_n3454( .i (n3453), .o (n3454) );
  buffer buf_n3455( .i (n3454), .o (n3455) );
  buffer buf_n3456( .i (n3455), .o (n3456) );
  buffer buf_n3457( .i (n3456), .o (n3457) );
  buffer buf_n3458( .i (n3457), .o (n3458) );
  buffer buf_n3459( .i (n3458), .o (n3459) );
  buffer buf_n3460( .i (n3459), .o (n3460) );
  assign n3461 = ~n147 & n2592 ;
  assign n3462 = ( n124 & ~n3442 ) | ( n124 & n3461 ) | ( ~n3442 & n3461 ) ;
  assign n3463 = ~n125 & n3462 ;
  assign n3464 = ( n1814 & n3446 ) | ( n1814 & n3463 ) | ( n3446 & n3463 ) ;
  buffer buf_n3465( .i (n3446), .o (n3465) );
  assign n3466 = n3464 & ~n3465 ;
  assign n3467 = ( n1433 & n2992 ) | ( n1433 & n3466 ) | ( n2992 & n3466 ) ;
  assign n3468 = ~n3080 & n3467 ;
  buffer buf_n3469( .i (n3468), .o (n3469) );
  buffer buf_n3470( .i (n3469), .o (n3470) );
  buffer buf_n3471( .i (n3470), .o (n3471) );
  buffer buf_n3472( .i (n3471), .o (n3472) );
  buffer buf_n3473( .i (n3472), .o (n3473) );
  buffer buf_n3474( .i (n3473), .o (n3474) );
  buffer buf_n3475( .i (n3474), .o (n3475) );
  buffer buf_n3476( .i (n3475), .o (n3476) );
  buffer buf_n3477( .i (n3476), .o (n3477) );
  assign n3479 = n2278 & n3119 ;
  buffer buf_n3480( .i (n3479), .o (n3480) );
  assign n3482 = n596 & n3480 ;
  buffer buf_n3483( .i (n3482), .o (n3483) );
  buffer buf_n3484( .i (n3483), .o (n3484) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n3481( .i (n3480), .o (n3481) );
  assign n3493 = n628 & n3481 ;
  buffer buf_n3494( .i (n3493), .o (n3494) );
  assign n3500 = n3484 | n3494 ;
  buffer buf_n3501( .i (n3500), .o (n3501) );
  buffer buf_n3502( .i (n3501), .o (n3502) );
  buffer buf_n3503( .i (n3502), .o (n3503) );
  buffer buf_n3504( .i (n3503), .o (n3504) );
  buffer buf_n3505( .i (n3504), .o (n3505) );
  assign n3506 = n3477 | n3505 ;
  assign n3507 = ( ~n2340 & n3460 ) | ( ~n2340 & n3506 ) | ( n3460 & n3506 ) ;
  assign n3508 = n2341 | n3507 ;
  buffer buf_n2940( .i (n2939), .o (n2940) );
  buffer buf_n2941( .i (n2940), .o (n2941) );
  buffer buf_n2942( .i (n2941), .o (n2942) );
  buffer buf_n2943( .i (n2942), .o (n2943) );
  buffer buf_n2944( .i (n2943), .o (n2944) );
  buffer buf_n2945( .i (n2944), .o (n2945) );
  assign n3509 = n3168 | n3302 ;
  assign n3510 = n2863 | n3509 ;
  buffer buf_n3511( .i (n2707), .o (n3511) );
  buffer buf_n3512( .i (n1216), .o (n3512) );
  assign n3513 = ~n3511 & n3512 ;
  buffer buf_n3514( .i (n3465), .o (n3514) );
  assign n3515 = n3513 & ~n3514 ;
  buffer buf_n3516( .i (n3515), .o (n3516) );
  assign n3517 = ( n1756 & n3418 ) | ( n1756 & n3516 ) | ( n3418 & n3516 ) ;
  assign n3518 = ~n3134 & n3517 ;
  buffer buf_n3519( .i (n3518), .o (n3519) );
  buffer buf_n3520( .i (n3519), .o (n3520) );
  buffer buf_n3521( .i (n3520), .o (n3521) );
  buffer buf_n3522( .i (n3521), .o (n3522) );
  buffer buf_n3523( .i (n3522), .o (n3523) );
  assign n3529 = n623 & ~n782 ;
  buffer buf_n3530( .i (n3529), .o (n3530) );
  buffer buf_n3531( .i (n3530), .o (n3531) );
  assign n3532 = ( n2673 & n3079 ) | ( n2673 & n3531 ) | ( n3079 & n3531 ) ;
  assign n3533 = ~n3123 & n3532 ;
  assign n3534 = n2793 & n3533 ;
  buffer buf_n3535( .i (n3534), .o (n3535) );
  buffer buf_n3536( .i (n3535), .o (n3536) );
  buffer buf_n3537( .i (n3536), .o (n3537) );
  buffer buf_n3538( .i (n3537), .o (n3538) );
  buffer buf_n3542( .i (n1231), .o (n3542) );
  assign n3543 = ( ~n2711 & n3079 ) | ( ~n2711 & n3542 ) | ( n3079 & n3542 ) ;
  assign n3544 = ~n3123 & n3543 ;
  buffer buf_n3545( .i (n3544), .o (n3545) );
  buffer buf_n3546( .i (n3545), .o (n3546) );
  buffer buf_n3547( .i (n3546), .o (n3547) );
  assign n3554 = n3340 | n3547 ;
  assign n3555 = n3316 | n3554 ;
  assign n3556 = n3538 | n3555 ;
  assign n3557 = n3523 | n3556 ;
  buffer buf_n367( .i (x14), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  assign n3558 = n386 & ~n2826 ;
  assign n3559 = ( n731 & ~n783 ) | ( n731 & n3558 ) | ( ~n783 & n3558 ) ;
  assign n3560 = ~n732 & n3559 ;
  assign n3561 = ~n3120 & n3560 ;
  buffer buf_n3562( .i (n3561), .o (n3562) );
  buffer buf_n345( .i (x13), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  assign n3570 = n362 & ~n728 ;
  assign n3571 = ( n385 & n3445 ) | ( n385 & n3570 ) | ( n3445 & n3570 ) ;
  assign n3572 = ~n386 & n3571 ;
  buffer buf_n3573( .i (n782), .o (n3573) );
  assign n3574 = n3572 & ~n3573 ;
  buffer buf_n3575( .i (n2827), .o (n3575) );
  assign n3576 = ( ~n3119 & n3574 ) | ( ~n3119 & n3575 ) | ( n3574 & n3575 ) ;
  buffer buf_n3577( .i (n3575), .o (n3577) );
  assign n3578 = n3576 & ~n3577 ;
  buffer buf_n3579( .i (n3578), .o (n3579) );
  assign n3590 = n3562 | n3579 ;
  buffer buf_n3591( .i (n3590), .o (n3591) );
  buffer buf_n3592( .i (n3591), .o (n3592) );
  buffer buf_n3593( .i (n3592), .o (n3593) );
  buffer buf_n3594( .i (n3593), .o (n3594) );
  buffer buf_n3595( .i (n3594), .o (n3595) );
  buffer buf_n3596( .i (n3595), .o (n3596) );
  assign n3597 = n3557 | n3596 ;
  assign n3598 = ( ~n2944 & n3510 ) | ( ~n2944 & n3597 ) | ( n3510 & n3597 ) ;
  assign n3599 = n2945 | n3598 ;
  assign n3600 = n705 & ~n3573 ;
  assign n3601 = ( n2306 & n3575 ) | ( n2306 & n3600 ) | ( n3575 & n3600 ) ;
  assign n3602 = ~n3577 & n3601 ;
  assign n3603 = n3332 & n3602 ;
  buffer buf_n3604( .i (n3603), .o (n3604) );
  buffer buf_n3605( .i (n3604), .o (n3605) );
  buffer buf_n3606( .i (n3605), .o (n3606) );
  buffer buf_n3607( .i (n3606), .o (n3607) );
  buffer buf_n3608( .i (n3607), .o (n3608) );
  buffer buf_n3609( .i (n3608), .o (n3609) );
  buffer buf_n3610( .i (n3609), .o (n3610) );
  buffer buf_n3611( .i (n3610), .o (n3611) );
  assign n3612 = ( n2306 & n3530 ) | ( n2306 & n3575 ) | ( n3530 & n3575 ) ;
  assign n3613 = ~n3577 & n3612 ;
  assign n3614 = n3332 & n3613 ;
  buffer buf_n3615( .i (n3614), .o (n3615) );
  buffer buf_n3616( .i (n3615), .o (n3616) );
  buffer buf_n3617( .i (n3616), .o (n3617) );
  buffer buf_n3618( .i (n3617), .o (n3618) );
  buffer buf_n3619( .i (n3618), .o (n3619) );
  buffer buf_n3620( .i (n3619), .o (n3620) );
  buffer buf_n3621( .i (n3620), .o (n3621) );
  buffer buf_n2310( .i (n2309), .o (n2310) );
  buffer buf_n3624( .i (n3386), .o (n3624) );
  assign n3625 = n2310 & n3624 ;
  buffer buf_n3626( .i (n3625), .o (n3626) );
  buffer buf_n3627( .i (n3626), .o (n3627) );
  buffer buf_n3628( .i (n3627), .o (n3628) );
  buffer buf_n3629( .i (n3628), .o (n3629) );
  buffer buf_n3636( .i (n2772), .o (n3636) );
  assign n3637 = n624 & n3636 ;
  buffer buf_n3638( .i (n3637), .o (n3638) );
  buffer buf_n3639( .i (n3638), .o (n3639) );
  assign n3640 = ( n3418 & n3516 ) | ( n3418 & n3639 ) | ( n3516 & n3639 ) ;
  buffer buf_n3641( .i (n3418), .o (n3641) );
  assign n3642 = n3640 & ~n3641 ;
  buffer buf_n3643( .i (n3642), .o (n3643) );
  buffer buf_n3644( .i (n3643), .o (n3644) );
  buffer buf_n3645( .i (n3644), .o (n3645) );
  assign n3652 = n2358 | n3645 ;
  assign n3653 = n2661 | n3652 ;
  assign n3654 = n3629 | n3653 ;
  assign n3655 = ( ~n3610 & n3621 ) | ( ~n3610 & n3654 ) | ( n3621 & n3654 ) ;
  assign n3656 = n3611 | n3655 ;
  buffer buf_n3657( .i (n3656), .o (n3657) );
  assign n3660 = n3599 | n3657 ;
  assign n3661 = n3508 | n3660 ;
  buffer buf_n3004( .i (n3003), .o (n3004) );
  buffer buf_n3005( .i (n3004), .o (n3005) );
  buffer buf_n3006( .i (n3005), .o (n3006) );
  buffer buf_n3007( .i (n3006), .o (n3007) );
  buffer buf_n3008( .i (n3007), .o (n3008) );
  buffer buf_n2429( .i (n2428), .o (n2429) );
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  buffer buf_n2432( .i (n2431), .o (n2432) );
  buffer buf_n2527( .i (n2526), .o (n2527) );
  buffer buf_n2528( .i (n2527), .o (n2528) );
  buffer buf_n2450( .i (n2449), .o (n2450) );
  buffer buf_n2451( .i (n2450), .o (n2451) );
  buffer buf_n2452( .i (n2451), .o (n2452) );
  assign n3662 = ~n730 & n2436 ;
  assign n3663 = ~n2827 & n3662 ;
  buffer buf_n3664( .i (n3663), .o (n3664) );
  buffer buf_n3665( .i (n3664), .o (n3665) );
  assign n3666 = n3385 & n3665 ;
  buffer buf_n3667( .i (n3666), .o (n3667) );
  buffer buf_n3668( .i (n3667), .o (n3668) );
  buffer buf_n3669( .i (n3668), .o (n3669) );
  buffer buf_n3670( .i (n3669), .o (n3670) );
  buffer buf_n3671( .i (n3670), .o (n3671) );
  buffer buf_n3672( .i (n3671), .o (n3672) );
  buffer buf_n3673( .i (n3672), .o (n3673) );
  buffer buf_n3674( .i (n3673), .o (n3674) );
  assign n3676 = n2452 | n3674 ;
  assign n3677 = n2528 | n3676 ;
  assign n3678 = n2432 | n3677 ;
  assign n3679 = n3008 | n3678 ;
  assign n3680 = n3661 | n3679 ;
  assign n3681 = ( ~n2224 & n3438 ) | ( ~n2224 & n3680 ) | ( n3438 & n3680 ) ;
  assign n3682 = n2225 | n3681 ;
  buffer buf_n2212( .i (n2211), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  assign n3683 = n1110 & ~n1158 ;
  assign n3684 = ( n1132 & n2167 ) | ( n1132 & n3683 ) | ( n2167 & n3683 ) ;
  assign n3685 = ~n1133 & n3684 ;
  buffer buf_n3686( .i (n3685), .o (n3686) );
  buffer buf_n3687( .i (n3686), .o (n3687) );
  buffer buf_n3688( .i (n3687), .o (n3688) );
  buffer buf_n3689( .i (n3688), .o (n3689) );
  buffer buf_n3690( .i (n3689), .o (n3690) );
  buffer buf_n3691( .i (n3690), .o (n3691) );
  assign n3695 = n2124 | n3691 ;
  assign n3696 = n2213 | n3695 ;
  buffer buf_n3697( .i (n3696), .o (n3697) );
  buffer buf_n3698( .i (n3697), .o (n3698) );
  buffer buf_n3699( .i (n3698), .o (n3699) );
  buffer buf_n3700( .i (n3699), .o (n3700) );
  buffer buf_n3701( .i (n3700), .o (n3701) );
  buffer buf_n3702( .i (n3701), .o (n3702) );
  buffer buf_n3703( .i (n3702), .o (n3703) );
  buffer buf_n2382( .i (n2381), .o (n2382) );
  buffer buf_n2383( .i (n2382), .o (n2383) );
  buffer buf_n2384( .i (n2383), .o (n2384) );
  buffer buf_n2385( .i (n2384), .o (n2385) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n2417( .i (n2416), .o (n2417) );
  buffer buf_n2418( .i (n2417), .o (n2418) );
  assign n3704 = n911 & n2418 ;
  buffer buf_n3705( .i (n3704), .o (n3705) );
  buffer buf_n3706( .i (n3705), .o (n3706) );
  buffer buf_n3707( .i (n3706), .o (n3707) );
  buffer buf_n3708( .i (n3707), .o (n3708) );
  buffer buf_n3709( .i (n3708), .o (n3709) );
  buffer buf_n3710( .i (n3709), .o (n3710) );
  assign n3711 = n2432 | n3007 ;
  assign n3712 = ( ~n2384 & n3710 ) | ( ~n2384 & n3711 ) | ( n3710 & n3711 ) ;
  assign n3713 = n2385 | n3712 ;
  buffer buf_n2359( .i (n2358), .o (n2359) );
  buffer buf_n2360( .i (n2359), .o (n2360) );
  buffer buf_n2361( .i (n2360), .o (n2361) );
  buffer buf_n2362( .i (n2361), .o (n2362) );
  buffer buf_n2363( .i (n2362), .o (n2363) );
  buffer buf_n3319( .i (n3318), .o (n3319) );
  assign n3714 = n2663 | n3319 ;
  assign n3715 = ( ~n2362 & n3459 ) | ( ~n2362 & n3714 ) | ( n3459 & n3714 ) ;
  assign n3716 = n2363 | n3715 ;
  assign n3717 = n2335 | n3473 ;
  buffer buf_n3718( .i (n3717), .o (n3718) );
  buffer buf_n3719( .i (n3718), .o (n3719) );
  buffer buf_n3720( .i (n3719), .o (n3720) );
  buffer buf_n3721( .i (n3720), .o (n3721) );
  assign n3724 = n2622 & n3234 ;
  buffer buf_n3725( .i (n3724), .o (n3725) );
  buffer buf_n3726( .i (n3725), .o (n3726) );
  buffer buf_n3727( .i (n3726), .o (n3727) );
  assign n3730 = n2859 | n2923 ;
  assign n3731 = ( ~n3062 & n3072 ) | ( ~n3062 & n3730 ) | ( n3072 & n3730 ) ;
  assign n3732 = n3063 | n3731 ;
  assign n3733 = n3727 | n3732 ;
  assign n3734 = ( n3169 & ~n3287 ) | ( n3169 & n3733 ) | ( ~n3287 & n3733 ) ;
  assign n3735 = n3288 | n3734 ;
  assign n3736 = n3721 | n3735 ;
  assign n3737 = ( ~n3030 & n3716 ) | ( ~n3030 & n3736 ) | ( n3716 & n3736 ) ;
  assign n3738 = n3031 | n3737 ;
  buffer buf_n3197( .i (n3196), .o (n3197) );
  buffer buf_n3198( .i (n3197), .o (n3198) );
  buffer buf_n3199( .i (n3198), .o (n3199) );
  buffer buf_n3200( .i (n3199), .o (n3200) );
  buffer buf_n2453( .i (n2452), .o (n2453) );
  buffer buf_n2454( .i (n2453), .o (n2454) );
  assign n3739 = n2532 | n3367 ;
  buffer buf_n3740( .i (n3739), .o (n3740) );
  buffer buf_n3741( .i (n3740), .o (n3741) );
  assign n3742 = n2557 | n3741 ;
  buffer buf_n3743( .i (n3742), .o (n3743) );
  buffer buf_n3744( .i (n3743), .o (n3744) );
  buffer buf_n3745( .i (n3744), .o (n3745) );
  buffer buf_n3746( .i (n3745), .o (n3746) );
  assign n3747 = n2454 | n3746 ;
  assign n3748 = n3200 | n3747 ;
  assign n3749 = n3738 | n3748 ;
  assign n3750 = ( ~n3702 & n3713 ) | ( ~n3702 & n3749 ) | ( n3713 & n3749 ) ;
  assign n3751 = n3703 | n3750 ;
  buffer buf_n852( .i (x32), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  assign n3752 = n620 & n2104 ;
  assign n3753 = ( n780 & n810 ) | ( n780 & n3752 ) | ( n810 & n3752 ) ;
  assign n3754 = ~n811 & n3753 ;
  buffer buf_n3755( .i (n3754), .o (n3755) );
  buffer buf_n3756( .i (n3755), .o (n3756) );
  buffer buf_n3757( .i (n3756), .o (n3757) );
  buffer buf_n3758( .i (n3757), .o (n3758) );
  buffer buf_n3759( .i (n3758), .o (n3759) );
  buffer buf_n3760( .i (n3759), .o (n3760) );
  buffer buf_n3761( .i (n3760), .o (n3761) );
  buffer buf_n3762( .i (n3761), .o (n3762) );
  buffer buf_n3763( .i (n3762), .o (n3763) );
  assign n3769 = n850 & n3762 ;
  assign n3770 = ( n880 & n3763 ) | ( n880 & n3769 ) | ( n3763 & n3769 ) ;
  buffer buf_n3771( .i (n3770), .o (n3771) );
  buffer buf_n3772( .i (n3771), .o (n3772) );
  assign n3773 = ( n2110 & n3080 ) | ( n2110 & n3638 ) | ( n3080 & n3638 ) ;
  buffer buf_n3774( .i (n3573), .o (n3774) );
  buffer buf_n3775( .i (n3774), .o (n3775) );
  buffer buf_n3776( .i (n3775), .o (n3776) );
  assign n3777 = n3773 & ~n3776 ;
  buffer buf_n3778( .i (n3777), .o (n3778) );
  buffer buf_n3779( .i (n3778), .o (n3779) );
  buffer buf_n3780( .i (n3779), .o (n3780) );
  buffer buf_n3781( .i (n3780), .o (n3781) );
  buffer buf_n3782( .i (n3781), .o (n3782) );
  buffer buf_n3783( .i (n3782), .o (n3783) );
  buffer buf_n1016( .i (x37), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n951( .i (x35), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  assign n3787 = ~n872 & n3755 ;
  assign n3788 = ( n844 & ~n904 ) | ( n844 & n3787 ) | ( ~n904 & n3787 ) ;
  assign n3789 = ~n845 & n3788 ;
  buffer buf_n3790( .i (n3789), .o (n3790) );
  buffer buf_n3791( .i (n3790), .o (n3791) );
  buffer buf_n917( .i (x34), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  assign n3799 = n941 & n3790 ;
  assign n3800 = ( n976 & n3791 ) | ( n976 & n3799 ) | ( n3791 & n3799 ) ;
  buffer buf_n3801( .i (n3800), .o (n3801) );
  buffer buf_n3802( .i (n3801), .o (n3802) );
  buffer buf_n3803( .i (n3802), .o (n3803) );
  buffer buf_n984( .i (x36), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  assign n3804 = ~n941 & n3790 ;
  assign n3805 = ~n976 & n3804 ;
  buffer buf_n3806( .i (n3805), .o (n3806) );
  assign n3812 = ( ~n1011 & n3801 ) | ( ~n1011 & n3806 ) | ( n3801 & n3806 ) ;
  assign n3813 = n1044 & ~n3812 ;
  assign n3814 = ( n1045 & n3803 ) | ( n1045 & ~n3813 ) | ( n3803 & ~n3813 ) ;
  assign n3815 = n3783 | n3814 ;
  assign n3816 = ( ~n2983 & n3772 ) | ( ~n2983 & n3815 ) | ( n3772 & n3815 ) ;
  assign n3817 = n2984 | n3816 ;
  buffer buf_n3818( .i (n3817), .o (n3818) );
  buffer buf_n3819( .i (n3818), .o (n3819) );
  buffer buf_n3820( .i (n731), .o (n3820) );
  assign n3821 = n3774 & n3820 ;
  assign n3822 = ( n2439 & n3577 ) | ( n2439 & n3821 ) | ( n3577 & n3821 ) ;
  assign n3823 = ~n3123 & n3822 ;
  buffer buf_n3824( .i (n3332), .o (n3824) );
  assign n3825 = n3823 & ~n3824 ;
  buffer buf_n3826( .i (n3825), .o (n3826) );
  buffer buf_n3827( .i (n3826), .o (n3827) );
  buffer buf_n3828( .i (n3827), .o (n3828) );
  buffer buf_n3829( .i (n3828), .o (n3829) );
  buffer buf_n3830( .i (n3829), .o (n3830) );
  buffer buf_n3831( .i (n3830), .o (n3831) );
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n3833( .i (n2826), .o (n3833) );
  buffer buf_n3834( .i (n3833), .o (n3834) );
  buffer buf_n3835( .i (n3834), .o (n3835) );
  buffer buf_n3836( .i (n3835), .o (n3836) );
  assign n3837 = ( n1756 & ~n2111 ) | ( n1756 & n3836 ) | ( ~n2111 & n3836 ) ;
  assign n3838 = n2112 & n3837 ;
  buffer buf_n3839( .i (n3838), .o (n3839) );
  buffer buf_n3840( .i (n3839), .o (n3840) );
  buffer buf_n3841( .i (n3840), .o (n3841) );
  buffer buf_n3842( .i (n3841), .o (n3842) );
  buffer buf_n3843( .i (n3842), .o (n3843) );
  buffer buf_n3844( .i (n3843), .o (n3844) );
  assign n3846 = n3831 | n3844 ;
  buffer buf_n3847( .i (n3846), .o (n3847) );
  buffer buf_n3848( .i (n3847), .o (n3848) );
  assign n3849 = n1498 | n2469 ;
  buffer buf_n3850( .i (n3849), .o (n3850) );
  buffer buf_n3851( .i (n3850), .o (n3851) );
  buffer buf_n3852( .i (n3851), .o (n3852) );
  buffer buf_n3853( .i (n3852), .o (n3853) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n3854( .i (n2227), .o (n3854) );
  assign n3855 = ( ~n178 & n1664 ) | ( ~n178 & n3854 ) | ( n1664 & n3854 ) ;
  assign n3856 = n179 & n3855 ;
  assign n3857 = ~n2994 & n3835 ;
  assign n3858 = ( n2996 & n3856 ) | ( n2996 & n3857 ) | ( n3856 & n3857 ) ;
  assign n3859 = ~n2043 & n3858 ;
  assign n3860 = ~n2836 & n3859 ;
  assign n3861 = n2235 & n3860 ;
  buffer buf_n3862( .i (n3861), .o (n3862) );
  buffer buf_n3863( .i (n3862), .o (n3863) );
  buffer buf_n3864( .i (n3863), .o (n3864) );
  buffer buf_n3865( .i (n3864), .o (n3865) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  assign n3869 = ( ~n199 & n1662 ) | ( ~n199 & n2989 ) | ( n1662 & n2989 ) ;
  assign n3870 = n200 & n3869 ;
  assign n3871 = ~n3820 & n3870 ;
  assign n3872 = ( n1863 & ~n3835 ) | ( n1863 & n3871 ) | ( ~n3835 & n3871 ) ;
  assign n3873 = ~n2996 & n3872 ;
  assign n3874 = n3824 & n3873 ;
  assign n3875 = n3354 & n3874 ;
  buffer buf_n3876( .i (n3875), .o (n3876) );
  buffer buf_n3877( .i (n3876), .o (n3877) );
  buffer buf_n3878( .i (n3877), .o (n3878) );
  assign n3882 = n2494 | n3878 ;
  buffer buf_n3883( .i (n3882), .o (n3883) );
  assign n3887 = ( ~n2451 & n3865 ) | ( ~n2451 & n3883 ) | ( n3865 & n3883 ) ;
  assign n3888 = n2452 | n3887 ;
  assign n3889 = n3853 | n3888 ;
  assign n3890 = ( ~n3818 & n3848 ) | ( ~n3818 & n3889 ) | ( n3848 & n3889 ) ;
  assign n3891 = n3819 | n3890 ;
  buffer buf_n3892( .i (n3891), .o (n3892) );
  buffer buf_n3893( .i (n3892), .o (n3893) );
  assign n3894 = n2646 & ~n3234 ;
  buffer buf_n3895( .i (n3894), .o (n3895) );
  buffer buf_n3896( .i (n3895), .o (n3896) );
  buffer buf_n3897( .i (n3896), .o (n3897) );
  buffer buf_n3898( .i (n3897), .o (n3898) );
  buffer buf_n3899( .i (n3898), .o (n3899) );
  buffer buf_n3900( .i (n3899), .o (n3900) );
  buffer buf_n3901( .i (n3900), .o (n3901) );
  buffer buf_n3902( .i (n3901), .o (n3902) );
  buffer buf_n3903( .i (n148), .o (n3903) );
  buffer buf_n3904( .i (n3442), .o (n3904) );
  assign n3905 = n3903 & ~n3904 ;
  buffer buf_n3906( .i (n3905), .o (n3906) );
  assign n3911 = ~n2227 & n3906 ;
  assign n3912 = ~n3514 & n3911 ;
  assign n3913 = ( n3105 & ~n3835 ) | ( n3105 & n3912 ) | ( ~n3835 & n3912 ) ;
  assign n3914 = ~n535 & n3913 ;
  assign n3915 = ~n3824 & n3914 ;
  assign n3916 = n3354 & n3915 ;
  buffer buf_n3917( .i (n3916), .o (n3917) );
  buffer buf_n3918( .i (n3917), .o (n3918) );
  buffer buf_n3919( .i (n3918), .o (n3919) );
  buffer buf_n3920( .i (n3919), .o (n3920) );
  buffer buf_n3921( .i (n3920), .o (n3921) );
  buffer buf_n3922( .i (n3921), .o (n3922) );
  buffer buf_n3923( .i (n3922), .o (n3923) );
  buffer buf_n3924( .i (n3923), .o (n3924) );
  buffer buf_n3925( .i (n3119), .o (n3925) );
  buffer buf_n3926( .i (n3925), .o (n3926) );
  assign n3927 = n2619 & ~n3926 ;
  buffer buf_n3928( .i (n3927), .o (n3928) );
  buffer buf_n3929( .i (n3928), .o (n3929) );
  buffer buf_n3930( .i (n3929), .o (n3930) );
  buffer buf_n3931( .i (n3930), .o (n3931) );
  buffer buf_n3932( .i (n3931), .o (n3932) );
  buffer buf_n3933( .i (n3932), .o (n3933) );
  buffer buf_n3934( .i (n3933), .o (n3934) );
  buffer buf_n3935( .i (n3934), .o (n3935) );
  buffer buf_n3936( .i (n3935), .o (n3936) );
  assign n3939 = n2586 | n3936 ;
  assign n3940 = ( ~n3901 & n3924 ) | ( ~n3901 & n3939 ) | ( n3924 & n3939 ) ;
  assign n3941 = n3902 | n3940 ;
  buffer buf_n3524( .i (n3523), .o (n3524) );
  buffer buf_n3525( .i (n3524), .o (n3525) );
  assign n3942 = n1619 | n2700 ;
  assign n3943 = n3525 | n3942 ;
  buffer buf_n2675( .i (n2674), .o (n2675) );
  assign n3944 = ( n1276 & n2675 ) | ( n1276 & n3641 ) | ( n2675 & n3641 ) ;
  assign n3945 = ~n3354 & n3944 ;
  buffer buf_n3946( .i (n3945), .o (n3946) );
  buffer buf_n3947( .i (n3946), .o (n3947) );
  buffer buf_n3948( .i (n3947), .o (n3948) );
  buffer buf_n3949( .i (n3948), .o (n3949) );
  buffer buf_n3950( .i (n3949), .o (n3950) );
  buffer buf_n3951( .i (n3950), .o (n3951) );
  buffer buf_n205( .i (x6), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  assign n3952 = n224 & ~n2989 ;
  assign n3953 = ( n151 & n2709 ) | ( n151 & n3952 ) | ( n2709 & n3952 ) ;
  buffer buf_n3954( .i (n2709), .o (n3954) );
  assign n3955 = n3953 & ~n3954 ;
  assign n3956 = n3511 & n3833 ;
  buffer buf_n3957( .i (n3956), .o (n3957) );
  buffer buf_n3962( .i (n3514), .o (n3962) );
  assign n3963 = ( n3955 & n3957 ) | ( n3955 & n3962 ) | ( n3957 & n3962 ) ;
  assign n3964 = ~n2996 & n3963 ;
  assign n3965 = n3386 & n3964 ;
  buffer buf_n3966( .i (n3965), .o (n3966) );
  assign n3973 = ~n148 & n222 ;
  assign n3974 = ( n125 & ~n3904 ) | ( n125 & n3973 ) | ( ~n3904 & n3973 ) ;
  assign n3975 = ~n126 & n3974 ;
  assign n3976 = ~n3465 & n3975 ;
  buffer buf_n3977( .i (n3511), .o (n3977) );
  assign n3978 = ( n3854 & n3976 ) | ( n3854 & n3977 ) | ( n3976 & n3977 ) ;
  buffer buf_n3979( .i (n3854), .o (n3979) );
  assign n3980 = n3978 & ~n3979 ;
  assign n3981 = ( n1435 & n3776 ) | ( n1435 & n3980 ) | ( n3776 & n3980 ) ;
  assign n3982 = ~n3641 & n3981 ;
  buffer buf_n3983( .i (n3982), .o (n3983) );
  assign n3988 = n3966 | n3983 ;
  buffer buf_n3989( .i (n3988), .o (n3989) );
  buffer buf_n3990( .i (n3989), .o (n3990) );
  buffer buf_n3991( .i (n3990), .o (n3991) );
  buffer buf_n3992( .i (n3991), .o (n3992) );
  buffer buf_n3993( .i (n3992), .o (n3993) );
  assign n3994 = n3951 | n3993 ;
  assign n3995 = ( ~n2689 & n3943 ) | ( ~n2689 & n3994 ) | ( n3943 & n3994 ) ;
  assign n3996 = n2690 | n3995 ;
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n3997( .i (n2706), .o (n3997) );
  assign n3998 = n200 & ~n3997 ;
  assign n3999 = ( n152 & ~n3854 ) | ( n152 & n3998 ) | ( ~n3854 & n3998 ) ;
  assign n4000 = ~n153 & n3999 ;
  buffer buf_n4001( .i (n3962), .o (n4001) );
  assign n4002 = n4000 & ~n4001 ;
  buffer buf_n4003( .i (n3105), .o (n4003) );
  buffer buf_n4004( .i (n4003), .o (n4004) );
  assign n4005 = ( ~n3124 & n4002 ) | ( ~n3124 & n4004 ) | ( n4002 & n4004 ) ;
  assign n4006 = ~n537 & n4005 ;
  assign n4007 = ~n3234 & n4006 ;
  assign n4008 = n2034 & n4007 ;
  buffer buf_n4009( .i (n4008), .o (n4009) );
  buffer buf_n4010( .i (n4009), .o (n4010) );
  buffer buf_n4011( .i (n4010), .o (n4011) );
  buffer buf_n4012( .i (n4011), .o (n4012) );
  assign n4015 = n2737 | n4012 ;
  assign n4016 = ( ~n1654 & n2726 ) | ( ~n1654 & n4015 ) | ( n2726 & n4015 ) ;
  assign n4017 = n1655 | n4016 ;
  assign n4018 = n3996 | n4017 ;
  assign n4019 = n3941 | n4018 ;
  buffer buf_n3379( .i (n3378), .o (n3379) );
  buffer buf_n3380( .i (n3379), .o (n3380) );
  buffer buf_n3381( .i (n3380), .o (n3381) );
  buffer buf_n3382( .i (n3381), .o (n3382) );
  buffer buf_n3383( .i (n3382), .o (n3383) );
  buffer buf_n3384( .i (n3383), .o (n3384) );
  buffer buf_n4020( .i (n147), .o (n4020) );
  assign n4021 = ( n124 & n1214 ) | ( n124 & n4020 ) | ( n1214 & n4020 ) ;
  assign n4022 = ~n3903 & n4021 ;
  assign n4023 = ( n1814 & n3446 ) | ( n1814 & n4022 ) | ( n3446 & n4022 ) ;
  assign n4024 = ~n3465 & n4023 ;
  assign n4025 = ( n1433 & n3774 ) | ( n1433 & n4024 ) | ( n3774 & n4024 ) ;
  assign n4026 = ~n3775 & n4025 ;
  buffer buf_n4027( .i (n4026), .o (n4027) );
  buffer buf_n4028( .i (n4027), .o (n4028) );
  buffer buf_n4029( .i (n4028), .o (n4029) );
  buffer buf_n4030( .i (n4029), .o (n4030) );
  buffer buf_n4031( .i (n4030), .o (n4031) );
  buffer buf_n4032( .i (n4031), .o (n4032) );
  buffer buf_n4033( .i (n4032), .o (n4033) );
  buffer buf_n4034( .i (n4033), .o (n4034) );
  buffer buf_n4035( .i (n4034), .o (n4035) );
  assign n4036 = n2339 | n4035 ;
  assign n4037 = ( ~n2242 & n3384 ) | ( ~n2242 & n4036 ) | ( n3384 & n4036 ) ;
  assign n4038 = n2243 | n4037 ;
  assign n4039 = n2550 | n3743 ;
  assign n4040 = ( ~n2527 & n3413 ) | ( ~n2527 & n4039 ) | ( n3413 & n4039 ) ;
  assign n4041 = n2528 | n4040 ;
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  assign n4042 = n195 & n2501 ;
  buffer buf_n4043( .i (n499), .o (n4043) );
  buffer buf_n4044( .i (n4043), .o (n4044) );
  assign n4045 = ( n3440 & n4042 ) | ( n3440 & n4044 ) | ( n4042 & n4044 ) ;
  assign n4046 = ~n3442 & n4045 ;
  buffer buf_n4047( .i (n4046), .o (n4047) );
  assign n4053 = ~n2826 & n4047 ;
  buffer buf_n4054( .i (n3445), .o (n4054) );
  buffer buf_n4055( .i (n4054), .o (n4055) );
  assign n4056 = ( n593 & n4053 ) | ( n593 & n4055 ) | ( n4053 & n4055 ) ;
  assign n4057 = ~n3514 & n4056 ;
  assign n4058 = ~n3925 & n4057 ;
  assign n4059 = n3776 & n4058 ;
  buffer buf_n4060( .i (n4059), .o (n4060) );
  buffer buf_n4061( .i (n4060), .o (n4061) );
  buffer buf_n4062( .i (n4061), .o (n4062) );
  buffer buf_n4063( .i (n4062), .o (n4063) );
  buffer buf_n4064( .i (n4063), .o (n4064) );
  buffer buf_n4065( .i (n4064), .o (n4065) );
  buffer buf_n4066( .i (n4065), .o (n4066) );
  assign n4069 = n2361 | n4066 ;
  assign n4070 = ( ~n2319 & n2664 ) | ( ~n2319 & n4069 ) | ( n2664 & n4069 ) ;
  assign n4071 = n2320 | n4070 ;
  assign n4072 = n4041 | n4071 ;
  assign n4073 = n4038 | n4072 ;
  assign n4074 = n2795 | n2858 ;
  buffer buf_n4075( .i (n4074), .o (n4075) );
  buffer buf_n4076( .i (n4075), .o (n4076) );
  buffer buf_n4077( .i (n4076), .o (n4077) );
  buffer buf_n4078( .i (n4077), .o (n4078) );
  assign n4079 = n3596 | n4078 ;
  assign n4080 = ( n2913 & ~n2967 ) | ( n2913 & n4079 ) | ( ~n2967 & n4079 ) ;
  assign n4081 = n2968 | n4080 ;
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n2769( .i (n2768), .o (n2769) );
  assign n4082 = ( n2769 & n3014 ) | ( n2769 & n3775 ) | ( n3014 & n3775 ) ;
  assign n4083 = ~n3776 & n4082 ;
  buffer buf_n4084( .i (n4083), .o (n4084) );
  buffer buf_n4085( .i (n4084), .o (n4085) );
  buffer buf_n4086( .i (n4085), .o (n4086) );
  buffer buf_n4087( .i (n4086), .o (n4087) );
  buffer buf_n4088( .i (n4087), .o (n4088) );
  buffer buf_n4089( .i (n4088), .o (n4089) );
  assign n4092 = n1428 | n4089 ;
  assign n4093 = ( ~n2759 & n2785 ) | ( ~n2759 & n4092 ) | ( n2785 & n4092 ) ;
  assign n4094 = n2760 | n4093 ;
  assign n4095 = n2848 | n4094 ;
  assign n4096 = ( ~n3172 & n4081 ) | ( ~n3172 & n4095 ) | ( n4081 & n4095 ) ;
  assign n4097 = n3173 | n4096 ;
  assign n4098 = n4073 | n4097 ;
  assign n4099 = ( ~n3892 & n4019 ) | ( ~n3892 & n4098 ) | ( n4019 & n4098 ) ;
  assign n4100 = n3893 | n4099 ;
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  buffer buf_n2187( .i (n2186), .o (n2187) );
  buffer buf_n2188( .i (n2187), .o (n2188) );
  assign n4101 = n2124 | n2193 ;
  buffer buf_n4102( .i (n4101), .o (n4102) );
  buffer buf_n4103( .i (n4102), .o (n4103) );
  buffer buf_n4104( .i (n4103), .o (n4104) );
  buffer buf_n4105( .i (n4104), .o (n4105) );
  assign n4106 = n2199 | n2375 ;
  assign n4107 = n2210 | n4106 ;
  buffer buf_n4108( .i (n4107), .o (n4108) );
  buffer buf_n4109( .i (n4108), .o (n4109) );
  buffer buf_n4110( .i (n4109), .o (n4110) );
  buffer buf_n4111( .i (n4110), .o (n4111) );
  buffer buf_n4112( .i (n4111), .o (n4112) );
  assign n4113 = n1498 | n3180 ;
  assign n4114 = n3829 | n4113 ;
  assign n4115 = n2401 | n4114 ;
  assign n4116 = ( ~n2429 & n2462 ) | ( ~n2429 & n4115 ) | ( n2462 & n4115 ) ;
  assign n4117 = n2430 | n4116 ;
  assign n4118 = n4112 | n4117 ;
  assign n4119 = ( ~n2187 & n4105 ) | ( ~n2187 & n4118 ) | ( n4105 & n4118 ) ;
  assign n4120 = n2188 | n4119 ;
  buffer buf_n4121( .i (n4120), .o (n4121) );
  buffer buf_n4122( .i (n4121), .o (n4122) );
  buffer buf_n3415( .i (n3414), .o (n3415) );
  buffer buf_n3416( .i (n3415), .o (n3416) );
  buffer buf_n3417( .i (n3416), .o (n3417) );
  buffer buf_n2559( .i (n2558), .o (n2559) );
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  buffer buf_n2563( .i (n2562), .o (n2563) );
  buffer buf_n3428( .i (n3427), .o (n3428) );
  buffer buf_n3429( .i (n3428), .o (n3429) );
  buffer buf_n3430( .i (n3429), .o (n3430) );
  buffer buf_n3431( .i (n3430), .o (n3431) );
  assign n4123 = n3357 | n3740 ;
  buffer buf_n4124( .i (n4123), .o (n4124) );
  buffer buf_n4125( .i (n4124), .o (n4125) );
  buffer buf_n4126( .i (n4125), .o (n4126) );
  buffer buf_n4127( .i (n4126), .o (n4127) );
  buffer buf_n4128( .i (n4127), .o (n4128) );
  assign n4129 = n3431 | n4128 ;
  assign n4130 = ( n2563 & ~n3416 ) | ( n2563 & n4129 ) | ( ~n3416 & n4129 ) ;
  assign n4131 = n3417 | n4130 ;
  buffer buf_n3485( .i (n3484), .o (n3485) );
  buffer buf_n3486( .i (n3485), .o (n3486) );
  buffer buf_n3487( .i (n3486), .o (n3487) );
  buffer buf_n3488( .i (n3487), .o (n3488) );
  buffer buf_n3489( .i (n3488), .o (n3489) );
  buffer buf_n3490( .i (n3489), .o (n3490) );
  assign n4132 = n3469 | n4027 ;
  buffer buf_n4133( .i (n4132), .o (n4133) );
  buffer buf_n4134( .i (n4133), .o (n4134) );
  buffer buf_n4135( .i (n4134), .o (n4135) );
  buffer buf_n4136( .i (n4135), .o (n4136) );
  buffer buf_n4137( .i (n4136), .o (n4137) );
  buffer buf_n4138( .i (n4137), .o (n4138) );
  assign n4139 = n2333 | n4061 ;
  assign n4140 = n3454 | n4139 ;
  assign n4141 = n3604 | n3615 ;
  buffer buf_n4142( .i (n4141), .o (n4142) );
  assign n4151 = n2659 | n4142 ;
  assign n4152 = ( ~n2358 & n4140 ) | ( ~n2358 & n4151 ) | ( n4140 & n4151 ) ;
  assign n4153 = n2359 | n4152 ;
  assign n4154 = n3401 | n4153 ;
  assign n4155 = ( ~n3489 & n4138 ) | ( ~n3489 & n4154 ) | ( n4138 & n4154 ) ;
  assign n4156 = n3490 | n4155 ;
  buffer buf_n4157( .i (n4156), .o (n4157) );
  buffer buf_n4158( .i (n4157), .o (n4158) );
  assign n4159 = n1616 | n3989 ;
  buffer buf_n4160( .i (n4159), .o (n4160) );
  buffer buf_n4161( .i (n4160), .o (n4161) );
  buffer buf_n4162( .i (n4161), .o (n4162) );
  buffer buf_n4163( .i (n4162), .o (n4163) );
  buffer buf_n4164( .i (n4163), .o (n4164) );
  assign n4165 = n3895 | n3918 ;
  assign n4166 = n3932 | n4165 ;
  assign n4167 = n2904 | n4166 ;
  assign n4168 = ( ~n3169 & n3596 ) | ( ~n3169 & n4167 ) | ( n3596 & n4167 ) ;
  assign n4169 = n3170 | n4168 ;
  buffer buf_n4170( .i (n3775), .o (n4170) );
  assign n4171 = ( n1756 & n2674 ) | ( n1756 & n4170 ) | ( n2674 & n4170 ) ;
  assign n4172 = ~n3641 & n4171 ;
  buffer buf_n4173( .i (n4172), .o (n4173) );
  buffer buf_n4174( .i (n4173), .o (n4174) );
  buffer buf_n4175( .i (n4174), .o (n4175) );
  buffer buf_n4176( .i (n4175), .o (n4176) );
  buffer buf_n4177( .i (n4176), .o (n4177) );
  buffer buf_n4178( .i (n4177), .o (n4178) );
  assign n4187 = n650 & n2672 ;
  buffer buf_n4188( .i (n3774), .o (n4188) );
  assign n4189 = ( n3925 & n4187 ) | ( n3925 & n4188 ) | ( n4187 & n4188 ) ;
  assign n4190 = ~n3926 & n4189 ;
  buffer buf_n4191( .i (n4190), .o (n4191) );
  buffer buf_n4192( .i (n4191), .o (n4192) );
  buffer buf_n4193( .i (n4192), .o (n4193) );
  buffer buf_n4194( .i (n4193), .o (n4194) );
  buffer buf_n4195( .i (n4194), .o (n4195) );
  buffer buf_n4196( .i (n4195), .o (n4196) );
  assign n4198 = n4010 | n4196 ;
  assign n4199 = ( ~n1652 & n4178 ) | ( ~n1652 & n4198 ) | ( n4178 & n4198 ) ;
  assign n4200 = n1653 | n4199 ;
  assign n4201 = n4169 | n4200 ;
  assign n4202 = ( ~n4157 & n4164 ) | ( ~n4157 & n4201 ) | ( n4164 & n4201 ) ;
  assign n4203 = n4158 | n4202 ;
  buffer buf_n3866( .i (n3865), .o (n3866) );
  buffer buf_n3867( .i (n3866), .o (n3867) );
  buffer buf_n3868( .i (n3867), .o (n3868) );
  buffer buf_n3884( .i (n3883), .o (n3884) );
  buffer buf_n3885( .i (n3884), .o (n3885) );
  buffer buf_n3886( .i (n3885), .o (n3886) );
  assign n4204 = n3868 | n3886 ;
  assign n4205 = n3664 & ~n3925 ;
  assign n4206 = n4170 & n4205 ;
  buffer buf_n4207( .i (n4206), .o (n4207) );
  buffer buf_n4208( .i (n4207), .o (n4208) );
  buffer buf_n4209( .i (n4208), .o (n4209) );
  assign n4217 = n3669 | n4209 ;
  buffer buf_n4218( .i (n4217), .o (n4218) );
  buffer buf_n4219( .i (n4218), .o (n4219) );
  buffer buf_n4220( .i (n4219), .o (n4220) );
  buffer buf_n4221( .i (n4220), .o (n4221) );
  buffer buf_n4222( .i (n4221), .o (n4222) );
  buffer buf_n4223( .i (n4222), .o (n4223) );
  assign n4224 = n3199 | n4223 ;
  assign n4225 = n4204 | n4224 ;
  assign n4226 = n4203 | n4225 ;
  assign n4227 = ( ~n4121 & n4131 ) | ( ~n4121 & n4226 ) | ( n4131 & n4226 ) ;
  assign n4228 = n4122 | n4227 ;
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n3807( .i (n3806), .o (n3807) );
  buffer buf_n3808( .i (n3807), .o (n3808) );
  buffer buf_n3809( .i (n3808), .o (n3809) );
  buffer buf_n3810( .i (n3809), .o (n3810) );
  buffer buf_n3811( .i (n3810), .o (n3811) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  assign n4229 = n1015 & n3810 ;
  assign n4230 = ( n1048 & n3811 ) | ( n1048 & n4229 ) | ( n3811 & n4229 ) ;
  buffer buf_n4231( .i (n4230), .o (n4231) );
  buffer buf_n3784( .i (n3783), .o (n3784) );
  buffer buf_n3785( .i (n3784), .o (n3785) );
  buffer buf_n3786( .i (n3785), .o (n3786) );
  buffer buf_n3692( .i (n3691), .o (n3692) );
  assign n4232 = n3692 | n3843 ;
  assign n4233 = ( ~n3211 & n3706 ) | ( ~n3211 & n4232 ) | ( n3706 & n4232 ) ;
  assign n4234 = n3212 | n4233 ;
  assign n4235 = n3786 | n4234 ;
  assign n4236 = ( ~n2986 & n4231 ) | ( ~n2986 & n4235 ) | ( n4231 & n4235 ) ;
  assign n4237 = n2987 | n4236 ;
  buffer buf_n4238( .i (n4237), .o (n4238) );
  buffer buf_n4239( .i (n4238), .o (n4239) );
  buffer buf_n2455( .i (n2454), .o (n2455) );
  buffer buf_n2456( .i (n2455), .o (n2456) );
  buffer buf_n2551( .i (n2550), .o (n2551) );
  buffer buf_n2552( .i (n2551), .o (n2552) );
  buffer buf_n2553( .i (n2552), .o (n2553) );
  assign n4240 = n3197 | n3413 ;
  assign n4241 = ( ~n2552 & n2561 ) | ( ~n2552 & n4240 ) | ( n2561 & n4240 ) ;
  assign n4242 = n2553 | n4241 ;
  buffer buf_n4210( .i (n4209), .o (n4210) );
  buffer buf_n4211( .i (n4210), .o (n4211) );
  buffer buf_n4212( .i (n4211), .o (n4212) );
  buffer buf_n4213( .i (n4212), .o (n4213) );
  buffer buf_n4214( .i (n4213), .o (n4214) );
  buffer buf_n4215( .i (n4214), .o (n4215) );
  buffer buf_n4216( .i (n4215), .o (n4216) );
  assign n4243 = n2468 | n3827 ;
  buffer buf_n4244( .i (n4243), .o (n4244) );
  buffer buf_n4245( .i (n4244), .o (n4245) );
  buffer buf_n4246( .i (n4245), .o (n4246) );
  buffer buf_n4247( .i (n4246), .o (n4247) );
  buffer buf_n4248( .i (n4247), .o (n4248) );
  buffer buf_n4249( .i (n4248), .o (n4249) );
  assign n4250 = n4216 | n4249 ;
  assign n4251 = ( ~n2455 & n4242 ) | ( ~n2455 & n4250 ) | ( n4242 & n4250 ) ;
  assign n4252 = n2456 | n4251 ;
  buffer buf_n3728( .i (n3727), .o (n3728) );
  buffer buf_n3729( .i (n3728), .o (n3729) );
  buffer buf_n2841( .i (n2840), .o (n2841) );
  buffer buf_n2770( .i (n2769), .o (n2770) );
  buffer buf_n2771( .i (n2770), .o (n2771) );
  buffer buf_n4253( .i (n4170), .o (n4253) );
  assign n4254 = ( n1436 & n2771 ) | ( n1436 & n4253 ) | ( n2771 & n4253 ) ;
  buffer buf_n4255( .i (n4253), .o (n4255) );
  assign n4256 = n4254 & ~n4255 ;
  buffer buf_n4257( .i (n4256), .o (n4257) );
  buffer buf_n4258( .i (n4257), .o (n4258) );
  buffer buf_n4259( .i (n4258), .o (n4259) );
  assign n4264 = n3086 | n3261 ;
  assign n4265 = ( ~n2840 & n4259 ) | ( ~n2840 & n4264 ) | ( n4259 & n4264 ) ;
  assign n4266 = n2841 | n4265 ;
  assign n4267 = n3230 | n3243 ;
  assign n4268 = ( ~n3728 & n4266 ) | ( ~n3728 & n4267 ) | ( n4266 & n4267 ) ;
  assign n4269 = n3729 | n4268 ;
  buffer buf_n4270( .i (n4269), .o (n4270) );
  buffer buf_n4271( .i (n4270), .o (n4271) );
  buffer buf_n3304( .i (n3303), .o (n3304) );
  buffer buf_n3305( .i (n3304), .o (n3305) );
  buffer buf_n3320( .i (n3319), .o (n3320) );
  buffer buf_n3309( .i (n3308), .o (n3309) );
  buffer buf_n3310( .i (n3309), .o (n3310) );
  buffer buf_n3311( .i (n3310), .o (n3311) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n4272( .i (n3824), .o (n4272) );
  assign n4273 = ( n598 & ~n3310 ) | ( n598 & n4272 ) | ( ~n3310 & n4272 ) ;
  assign n4274 = ( n3282 & n3311 ) | ( n3282 & n4273 ) | ( n3311 & n4273 ) ;
  buffer buf_n4275( .i (n4274), .o (n4275) );
  buffer buf_n4276( .i (n4275), .o (n4276) );
  buffer buf_n4277( .i (n4276), .o (n4277) );
  buffer buf_n4278( .i (n4277), .o (n4278) );
  buffer buf_n4279( .i (n4278), .o (n4279) );
  assign n4280 = n3320 | n4279 ;
  assign n4281 = n3305 | n4280 ;
  assign n4282 = n3096 | n3145 ;
  buffer buf_n4283( .i (n4282), .o (n4283) );
  buffer buf_n4284( .i (n4283), .o (n4284) );
  assign n4285 = ( ~n2861 & n3129 ) | ( ~n2861 & n3271 ) | ( n3129 & n3271 ) ;
  assign n4286 = n2862 | n4285 ;
  buffer buf_n2753( .i (n2752), .o (n2753) );
  buffer buf_n2754( .i (n2753), .o (n2754) );
  assign n4287 = n2754 | n3072 ;
  assign n4288 = n2783 | n4287 ;
  assign n4289 = n2901 | n3592 ;
  assign n4290 = ( ~n2888 & n3154 ) | ( ~n2888 & n4289 ) | ( n3154 & n4289 ) ;
  assign n4291 = n2889 | n4290 ;
  assign n4292 = n4288 | n4291 ;
  assign n4293 = ( ~n4283 & n4286 ) | ( ~n4283 & n4292 ) | ( n4286 & n4292 ) ;
  assign n4294 = n4284 | n4293 ;
  assign n4295 = n3347 | n4294 ;
  assign n4296 = ( ~n4270 & n4281 ) | ( ~n4270 & n4295 ) | ( n4281 & n4295 ) ;
  assign n4297 = n4271 | n4296 ;
  buffer buf_n3722( .i (n3721), .o (n3722) );
  buffer buf_n3723( .i (n3722), .o (n3723) );
  assign n4298 = n2314 | n3454 ;
  buffer buf_n4299( .i (n4298), .o (n4299) );
  buffer buf_n4300( .i (n4299), .o (n4300) );
  buffer buf_n4301( .i (n4300), .o (n4301) );
  buffer buf_n4302( .i (n4301), .o (n4302) );
  buffer buf_n4303( .i (n4302), .o (n4303) );
  buffer buf_n4304( .i (n4303), .o (n4304) );
  assign n4305 = n2262 | n2534 ;
  assign n4306 = ( ~n2290 & n3025 ) | ( ~n2290 & n4305 ) | ( n3025 & n4305 ) ;
  assign n4307 = n2291 | n4306 ;
  assign n4308 = n3381 | n3503 ;
  assign n4309 = ( ~n2240 & n4307 ) | ( ~n2240 & n4308 ) | ( n4307 & n4308 ) ;
  assign n4310 = n2241 | n4309 ;
  assign n4311 = n2698 | n3948 ;
  assign n4312 = n2686 | n4311 ;
  assign n4313 = n3621 | n4312 ;
  assign n4314 = n3525 | n4313 ;
  assign n4315 = n4310 | n4314 ;
  assign n4316 = ( ~n3722 & n4304 ) | ( ~n3722 & n4315 ) | ( n4304 & n4315 ) ;
  assign n4317 = n3723 | n4316 ;
  assign n4318 = n4297 | n4317 ;
  assign n4319 = ( ~n4238 & n4252 ) | ( ~n4238 & n4318 ) | ( n4252 & n4318 ) ;
  assign n4320 = n4239 | n4319 ;
  buffer buf_n3548( .i (n3547), .o (n3548) );
  buffer buf_n3549( .i (n3548), .o (n3549) );
  buffer buf_n3550( .i (n3549), .o (n3550) );
  assign n4321 = n2723 | n3550 ;
  assign n4322 = n2736 | n4321 ;
  assign n4323 = n2584 | n2846 ;
  assign n4324 = n4322 | n4323 ;
  buffer buf_n4325( .i (n4324), .o (n4325) );
  buffer buf_n4326( .i (n4325), .o (n4326) );
  buffer buf_n3526( .i (n3525), .o (n3526) );
  assign n4327 = n3538 | n3948 ;
  buffer buf_n4328( .i (n4327), .o (n4328) );
  assign n4332 = n2700 | n4328 ;
  assign n4333 = ( n2688 & ~n3525 ) | ( n2688 & n4332 ) | ( ~n3525 & n4332 ) ;
  assign n4334 = n3526 | n4333 ;
  buffer buf_n4260( .i (n4259), .o (n4260) );
  buffer buf_n4261( .i (n4260), .o (n4261) );
  buffer buf_n4262( .i (n4261), .o (n4262) );
  assign n4335 = n2757 | n2798 ;
  assign n4336 = n1428 | n4335 ;
  assign n4337 = n2785 | n4336 ;
  assign n4338 = n4262 | n4337 ;
  assign n4339 = n2890 | n2965 ;
  assign n4340 = ( ~n2863 & n3596 ) | ( ~n2863 & n4339 ) | ( n3596 & n4339 ) ;
  assign n4341 = n2864 | n4340 ;
  assign n4342 = n4338 | n4341 ;
  assign n4343 = ( ~n4325 & n4334 ) | ( ~n4325 & n4342 ) | ( n4334 & n4342 ) ;
  assign n4344 = n4326 | n4343 ;
  buffer buf_n4345( .i (n4344), .o (n4345) );
  buffer buf_n4346( .i (n4345), .o (n4346) );
  buffer buf_n3390( .i (n3389), .o (n3390) );
  buffer buf_n3391( .i (n3390), .o (n3391) );
  buffer buf_n3392( .i (n3391), .o (n3392) );
  buffer buf_n3393( .i (n3392), .o (n3393) );
  buffer buf_n3394( .i (n3393), .o (n3394) );
  buffer buf_n3395( .i (n3394), .o (n3395) );
  buffer buf_n3396( .i (n3395), .o (n3396) );
  buffer buf_n3397( .i (n3396), .o (n3397) );
  buffer buf_n3398( .i (n3397), .o (n3398) );
  buffer buf_n3491( .i (n3490), .o (n3491) );
  buffer buf_n3492( .i (n3491), .o (n3492) );
  buffer buf_n4347( .i (n3440), .o (n4347) );
  assign n4348 = ~n2820 & n4347 ;
  buffer buf_n4349( .i (n4348), .o (n4349) );
  assign n4353 = ( n311 & n2989 ) | ( n311 & n4349 ) | ( n2989 & n4349 ) ;
  buffer buf_n4354( .i (n4353), .o (n4354) );
  buffer buf_n4356( .i (n2227), .o (n4356) );
  assign n4357 = n4354 & ~n4356 ;
  buffer buf_n4358( .i (n3636), .o (n4358) );
  buffer buf_n4359( .i (n4358), .o (n4359) );
  assign n4360 = n4357 & n4359 ;
  assign n4361 = ( n678 & n4001 ) | ( n678 & n4360 ) | ( n4001 & n4360 ) ;
  assign n4362 = ~n2043 & n4361 ;
  buffer buf_n4363( .i (n4362), .o (n4363) );
  buffer buf_n4364( .i (n4363), .o (n4364) );
  buffer buf_n4365( .i (n4364), .o (n4365) );
  buffer buf_n4366( .i (n4365), .o (n4366) );
  buffer buf_n4367( .i (n4366), .o (n4367) );
  buffer buf_n4368( .i (n4367), .o (n4368) );
  buffer buf_n4369( .i (n4368), .o (n4369) );
  buffer buf_n4370( .i (n4369), .o (n4370) );
  assign n4371 = n2320 | n4370 ;
  assign n4372 = n3492 | n4371 ;
  assign n4373 = n2244 | n4372 ;
  assign n4374 = n3398 | n4373 ;
  buffer buf_n3658( .i (n3657), .o (n3658) );
  buffer buf_n3659( .i (n3658), .o (n3659) );
  assign n4375 = n2549 | n3359 ;
  assign n4376 = n3428 | n4375 ;
  assign n4377 = n3674 | n4376 ;
  assign n4378 = ( n2474 & ~n3006 ) | ( n2474 & n4377 ) | ( ~n3006 & n4377 ) ;
  assign n4379 = n3007 | n4378 ;
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n3832( .i (n3831), .o (n3832) );
  assign n4380 = ( ~n949 & n983 ) | ( ~n949 & n3832 ) | ( n983 & n3832 ) ;
  buffer buf_n3792( .i (n3791), .o (n3792) );
  buffer buf_n3793( .i (n3792), .o (n3793) );
  buffer buf_n3794( .i (n3793), .o (n3794) );
  buffer buf_n3795( .i (n3794), .o (n3795) );
  buffer buf_n3796( .i (n3795), .o (n3796) );
  buffer buf_n3797( .i (n3796), .o (n3797) );
  buffer buf_n3798( .i (n3797), .o (n3798) );
  assign n4381 = n3798 | n3832 ;
  assign n4382 = ( n950 & n4380 ) | ( n950 & n4381 ) | ( n4380 & n4381 ) ;
  assign n4383 = n4231 | n4382 ;
  assign n4384 = n4379 | n4383 ;
  assign n4385 = n3659 | n4384 ;
  assign n4386 = ( ~n4345 & n4374 ) | ( ~n4345 & n4385 ) | ( n4374 & n4385 ) ;
  assign n4387 = n4346 | n4386 ;
  buffer buf_n3675( .i (n3674), .o (n3675) );
  buffer buf_n3046( .i (n3045), .o (n3046) );
  assign n4388 = n2472 | n3046 ;
  assign n4389 = ( n3010 & ~n3674 ) | ( n3010 & n4388 ) | ( ~n3674 & n4388 ) ;
  assign n4390 = n3675 | n4389 ;
  assign n4391 = ~n942 & n976 ;
  assign n4392 = n3792 & n4391 ;
  buffer buf_n4393( .i (n4392), .o (n4393) );
  buffer buf_n4394( .i (n4393), .o (n4394) );
  buffer buf_n4395( .i (n4394), .o (n4395) );
  buffer buf_n4396( .i (n4395), .o (n4396) );
  buffer buf_n4397( .i (n4396), .o (n4397) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  assign n4398 = ~n876 & n907 ;
  buffer buf_n4399( .i (n4398), .o (n4399) );
  buffer buf_n4400( .i (n4399), .o (n4400) );
  buffer buf_n4401( .i (n4400), .o (n4401) );
  buffer buf_n4402( .i (n4401), .o (n4402) );
  buffer buf_n4403( .i (n4402), .o (n4403) );
  buffer buf_n851( .i (n850), .o (n851) );
  assign n4404 = ~n851 & n3763 ;
  buffer buf_n4405( .i (n4404), .o (n4405) );
  assign n4409 = ( n882 & n4403 ) | ( n882 & n4405 ) | ( n4403 & n4405 ) ;
  buffer buf_n4410( .i (n4409), .o (n4410) );
  assign n4413 = n4397 | n4410 ;
  assign n4414 = n3847 | n4413 ;
  assign n4415 = ( ~n2986 & n4390 ) | ( ~n2986 & n4414 ) | ( n4390 & n4414 ) ;
  assign n4416 = n2987 | n4415 ;
  buffer buf_n4417( .i (n4416), .o (n4417) );
  buffer buf_n4418( .i (n4417), .o (n4418) );
  assign n4419 = n2237 | n3390 ;
  buffer buf_n4420( .i (n4419), .o (n4420) );
  buffer buf_n4421( .i (n4420), .o (n4421) );
  buffer buf_n4422( .i (n4421), .o (n4422) );
  assign n4423 = n3028 | n4422 ;
  buffer buf_n4424( .i (n4423), .o (n4424) );
  assign n4425 = n3431 | n4424 ;
  assign n4426 = ( n3364 & ~n3416 ) | ( n3364 & n4425 ) | ( ~n3416 & n4425 ) ;
  assign n4427 = n3417 | n4426 ;
  buffer buf_n2364( .i (n2363), .o (n2364) );
  buffer buf_n3646( .i (n3645), .o (n3646) );
  buffer buf_n3647( .i (n3646), .o (n3647) );
  buffer buf_n3648( .i (n3647), .o (n3648) );
  buffer buf_n3649( .i (n3648), .o (n3649) );
  buffer buf_n3539( .i (n3538), .o (n3539) );
  assign n4428 = n2686 | n3539 ;
  buffer buf_n4429( .i (n2699), .o (n4429) );
  assign n4430 = n4428 | n4429 ;
  assign n4431 = n3649 | n4430 ;
  assign n4432 = ( ~n2363 & n3526 ) | ( ~n2363 & n4431 ) | ( n3526 & n4431 ) ;
  assign n4433 = n2364 | n4432 ;
  buffer buf_n2842( .i (n2841), .o (n2842) );
  buffer buf_n2843( .i (n2842), .o (n2843) );
  buffer buf_n2844( .i (n2843), .o (n2844) );
  assign n4434 = n1422 | n2778 ;
  buffer buf_n4435( .i (n4434), .o (n4435) );
  buffer buf_n4436( .i (n4435), .o (n4436) );
  buffer buf_n4437( .i (n4436), .o (n4437) );
  buffer buf_n4438( .i (n4437), .o (n4438) );
  buffer buf_n4439( .i (n4438), .o (n4439) );
  buffer buf_n4440( .i (n4439), .o (n4440) );
  buffer buf_n4441( .i (n4440), .o (n4441) );
  assign n4444 = n2908 | n2962 ;
  assign n4445 = ( ~n2756 & n4075 ) | ( ~n2756 & n4444 ) | ( n4075 & n4444 ) ;
  assign n4446 = n2757 | n4445 ;
  buffer buf_n4447( .i (n4446), .o (n4447) );
  assign n4452 = n2816 | n3896 ;
  assign n4453 = n3933 | n4452 ;
  assign n4454 = n4447 | n4453 ;
  assign n4455 = ( ~n2843 & n4441 ) | ( ~n2843 & n4454 ) | ( n4441 & n4454 ) ;
  assign n4456 = n2844 | n4455 ;
  assign n4457 = n2734 | n4176 ;
  buffer buf_n4458( .i (n4457), .o (n4458) );
  buffer buf_n4459( .i (n4458), .o (n4459) );
  buffer buf_n4197( .i (n4196), .o (n4197) );
  assign n4460 = n2579 | n3546 ;
  buffer buf_n4461( .i (n4460), .o (n4461) );
  buffer buf_n4462( .i (n4461), .o (n4462) );
  buffer buf_n4463( .i (n4462), .o (n4463) );
  buffer buf_n4464( .i (n4463), .o (n4464) );
  assign n4465 = n4197 | n4464 ;
  assign n4466 = ( ~n2725 & n4459 ) | ( ~n2725 & n4465 ) | ( n4459 & n4465 ) ;
  assign n4467 = n2726 | n4466 ;
  assign n4468 = n4456 | n4467 ;
  assign n4469 = n4433 | n4468 ;
  buffer buf_n3630( .i (n3629), .o (n3630) );
  buffer buf_n3631( .i (n3630), .o (n3631) );
  buffer buf_n3632( .i (n3631), .o (n3632) );
  buffer buf_n3633( .i (n3632), .o (n3633) );
  buffer buf_n3634( .i (n3633), .o (n3634) );
  buffer buf_n3622( .i (n3621), .o (n3622) );
  buffer buf_n3623( .i (n3622), .o (n3623) );
  buffer buf_n3495( .i (n3494), .o (n3495) );
  buffer buf_n3496( .i (n3495), .o (n3496) );
  buffer buf_n3497( .i (n3496), .o (n3497) );
  buffer buf_n3498( .i (n3497), .o (n3498) );
  buffer buf_n3499( .i (n3498), .o (n3499) );
  assign n4470 = n3382 | n3499 ;
  assign n4471 = n3477 | n4470 ;
  assign n4472 = n3623 | n4471 ;
  assign n4473 = ( ~n3633 & n4304 ) | ( ~n3633 & n4472 ) | ( n4304 & n4472 ) ;
  assign n4474 = n3634 | n4473 ;
  assign n4475 = n4469 | n4474 ;
  assign n4476 = ( ~n4417 & n4427 ) | ( ~n4417 & n4475 ) | ( n4427 & n4475 ) ;
  assign n4477 = n4418 | n4476 ;
  buffer buf_n2269( .i (n2268), .o (n2269) );
  buffer buf_n2270( .i (n2269), .o (n2270) );
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2273( .i (n2272), .o (n2273) );
  buffer buf_n2293( .i (n2292), .o (n2293) );
  buffer buf_n2294( .i (n2293), .o (n2294) );
  buffer buf_n2295( .i (n2294), .o (n2295) );
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n2297( .i (n2296), .o (n2297) );
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  assign n4478 = n2977 | n3778 ;
  assign n4479 = n3206 | n4478 ;
  buffer buf_n4480( .i (n4479), .o (n4480) );
  assign n4483 = n2178 | n3687 ;
  buffer buf_n4484( .i (n4483), .o (n4484) );
  assign n4488 = n3840 | n4484 ;
  assign n4489 = ( ~n2123 & n4480 ) | ( ~n2123 & n4488 ) | ( n4480 & n4488 ) ;
  assign n4490 = n2124 | n4489 ;
  buffer buf_n4491( .i (n4490), .o (n4491) );
  buffer buf_n4492( .i (n4491), .o (n4492) );
  assign n4493 = ( n849 & n3761 ) | ( n849 & n4399 ) | ( n3761 & n4399 ) ;
  assign n4494 = ~n850 & n4493 ;
  buffer buf_n4495( .i (n4494), .o (n4495) );
  buffer buf_n4496( .i (n4495), .o (n4496) );
  assign n4499 = n946 | n4495 ;
  assign n4500 = ( n3796 & n4496 ) | ( n3796 & n4499 ) | ( n4496 & n4499 ) ;
  assign n4501 = ( ~n1012 & n1044 ) | ( ~n1012 & n4393 ) | ( n1044 & n4393 ) ;
  assign n4502 = n3807 | n4393 ;
  assign n4503 = ( n1013 & n4501 ) | ( n1013 & n4502 ) | ( n4501 & n4502 ) ;
  assign n4504 = n3771 | n4503 ;
  assign n4505 = ( ~n4491 & n4500 ) | ( ~n4491 & n4504 ) | ( n4500 & n4504 ) ;
  assign n4506 = n4492 | n4505 ;
  buffer buf_n4507( .i (n4506), .o (n4507) );
  buffer buf_n4508( .i (n4507), .o (n4508) );
  buffer buf_n2403( .i (n2402), .o (n2403) );
  assign n4509 = n2429 | n3706 ;
  assign n4510 = ( ~n2381 & n2403 ) | ( ~n2381 & n4509 ) | ( n2403 & n4509 ) ;
  assign n4511 = n2382 | n4510 ;
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2463( .i (n2462), .o (n2463) );
  assign n4512 = n2494 | n3181 ;
  assign n4513 = n3864 | n4512 ;
  assign n4514 = n3830 | n3850 ;
  assign n4515 = ( ~n2462 & n4513 ) | ( ~n2462 & n4514 ) | ( n4513 & n4514 ) ;
  assign n4516 = n2463 | n4515 ;
  assign n4517 = n2218 | n4516 ;
  assign n4518 = ( ~n4507 & n4511 ) | ( ~n4507 & n4517 ) | ( n4511 & n4517 ) ;
  assign n4519 = n4508 | n4518 ;
  buffer buf_n4520( .i (n4519), .o (n4520) );
  buffer buf_n4521( .i (n4520), .o (n4521) );
  buffer buf_n3233( .i (n3232), .o (n3233) );
  assign n4522 = n3083 | n4084 ;
  buffer buf_n4523( .i (n4522), .o (n4523) );
  assign n4531 = n2838 | n4523 ;
  assign n4532 = n4258 | n4531 ;
  assign n4533 = n3063 | n4532 ;
  assign n4534 = ( ~n2758 & n4439 ) | ( ~n2758 & n4533 ) | ( n4439 & n4533 ) ;
  assign n4535 = n2759 | n4534 ;
  assign n4536 = ~n310 & n1511 ;
  assign n4537 = ~n410 & n4536 ;
  buffer buf_n4538( .i (n2594), .o (n4538) );
  buffer buf_n4539( .i (n4538), .o (n4539) );
  buffer buf_n4540( .i (n4539), .o (n4540) );
  assign n4541 = ( n1663 & n4537 ) | ( n1663 & n4540 ) | ( n4537 & n4540 ) ;
  assign n4542 = ~n4356 & n4541 ;
  assign n4543 = n3962 & n4542 ;
  assign n4544 = ( n678 & n3836 ) | ( n678 & n4543 ) | ( n3836 & n4543 ) ;
  assign n4545 = ~n3124 & n4544 ;
  assign n4546 = n3624 & n4545 ;
  buffer buf_n4547( .i (n4546), .o (n4547) );
  buffer buf_n4548( .i (n4547), .o (n4548) );
  buffer buf_n4549( .i (n4548), .o (n4549) );
  buffer buf_n4550( .i (n4549), .o (n4550) );
  buffer buf_n3250( .i (n3249), .o (n3250) );
  buffer buf_n3251( .i (n3250), .o (n3251) );
  buffer buf_n3252( .i (n3251), .o (n3252) );
  assign n4557 = n198 & ~n4538 ;
  assign n4558 = ( n311 & n2706 ) | ( n311 & n4557 ) | ( n2706 & n4557 ) ;
  assign n4559 = ~n312 & n4558 ;
  buffer buf_n4560( .i (n4559), .o (n4560) );
  buffer buf_n4561( .i (n4560), .o (n4561) );
  assign n4562 = ( n1715 & n3962 ) | ( n1715 & ~n4560 ) | ( n3962 & ~n4560 ) ;
  assign n4563 = n4561 & n4562 ;
  buffer buf_n4564( .i (n3385), .o (n4564) );
  assign n4565 = ( n3124 & n4563 ) | ( n3124 & n4564 ) | ( n4563 & n4564 ) ;
  assign n4566 = ~n2718 & n4565 ;
  buffer buf_n4567( .i (n4566), .o (n4567) );
  buffer buf_n4568( .i (n4567), .o (n4568) );
  assign n4576 = n2815 | n4568 ;
  assign n4577 = ( n3252 & ~n4549 ) | ( n3252 & n4576 ) | ( ~n4549 & n4576 ) ;
  assign n4578 = n4550 | n4577 ;
  assign n4579 = n3244 | n4578 ;
  assign n4580 = ( ~n3232 & n4535 ) | ( ~n3232 & n4579 ) | ( n4535 & n4579 ) ;
  assign n4581 = n3233 | n4580 ;
  buffer buf_n4582( .i (n4581), .o (n4582) );
  buffer buf_n4583( .i (n4582), .o (n4583) );
  buffer buf_n3133( .i (n3132), .o (n3133) );
  assign n4584 = ~n310 & n4538 ;
  buffer buf_n4585( .i (n3904), .o (n4585) );
  assign n4586 = n4584 & ~n4585 ;
  assign n4587 = n4055 & n4586 ;
  assign n4588 = ( n676 & n3834 ) | ( n676 & n4587 ) | ( n3834 & n4587 ) ;
  buffer buf_n4589( .i (n3834), .o (n4589) );
  assign n4590 = n4588 & ~n4589 ;
  assign n4591 = n3385 & n4590 ;
  buffer buf_n4592( .i (n4591), .o (n4592) );
  buffer buf_n4593( .i (n4592), .o (n4593) );
  buffer buf_n4594( .i (n4593), .o (n4594) );
  buffer buf_n4595( .i (n4594), .o (n4595) );
  buffer buf_n4596( .i (n4595), .o (n4596) );
  buffer buf_n4597( .i (n4596), .o (n4597) );
  buffer buf_n4598( .i (n4597), .o (n4598) );
  buffer buf_n4599( .i (n4598), .o (n4599) );
  assign n4602 = n2944 | n4599 ;
  assign n4603 = ( ~n2865 & n3133 ) | ( ~n2865 & n4602 ) | ( n3133 & n4602 ) ;
  assign n4604 = n2866 | n4603 ;
  buffer buf_n3274( .i (n3273), .o (n3274) );
  buffer buf_n3275( .i (n3274), .o (n3275) );
  buffer buf_n3276( .i (n3275), .o (n3276) );
  buffer buf_n2892( .i (n2891), .o (n2892) );
  buffer buf_n2893( .i (n2892), .o (n2893) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n4605( .i (n3979), .o (n4605) );
  buffer buf_n4606( .i (n4605), .o (n4606) );
  assign n4607 = ( n316 & n1310 ) | ( n316 & ~n4606 ) | ( n1310 & ~n4606 ) ;
  assign n4608 = ~n317 & n4607 ;
  assign n4609 = n681 & n4608 ;
  assign n4610 = n569 & n4609 ;
  buffer buf_n4611( .i (n4610), .o (n4611) );
  buffer buf_n4612( .i (n4611), .o (n4612) );
  assign n4616 = n3156 | n4612 ;
  buffer buf_n4617( .i (n4616), .o (n4617) );
  buffer buf_n3563( .i (n3562), .o (n3563) );
  buffer buf_n3564( .i (n3563), .o (n3564) );
  buffer buf_n3565( .i (n3564), .o (n3565) );
  buffer buf_n3566( .i (n3565), .o (n3566) );
  buffer buf_n3567( .i (n3566), .o (n3567) );
  buffer buf_n3568( .i (n3567), .o (n3568) );
  buffer buf_n3569( .i (n3568), .o (n3569) );
  assign n4622 = n2924 | n3138 ;
  assign n4623 = ( n2903 & ~n2953 ) | ( n2903 & n4622 ) | ( ~n2953 & n4622 ) ;
  assign n4624 = n2954 | n4623 ;
  assign n4625 = n3569 | n4624 ;
  assign n4626 = ( ~n2892 & n4617 ) | ( ~n2892 & n4625 ) | ( n4617 & n4625 ) ;
  assign n4627 = n2893 | n4626 ;
  assign n4628 = n3276 | n4627 ;
  assign n4629 = ( ~n4582 & n4604 ) | ( ~n4582 & n4628 ) | ( n4604 & n4628 ) ;
  assign n4630 = n4583 | n4629 ;
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n3423( .i (n3422), .o (n3423) );
  buffer buf_n3424( .i (n3423), .o (n3424) );
  buffer buf_n4355( .i (n4354), .o (n4355) );
  assign n4631 = ~n314 & n4355 ;
  buffer buf_n4632( .i (n4631), .o (n4632) );
  buffer buf_n4633( .i (n4632), .o (n4633) );
  assign n4634 = ~n4255 & n4633 ;
  assign n4635 = ( n568 & n681 ) | ( n568 & n4634 ) | ( n681 & n4634 ) ;
  assign n4636 = ~n569 & n4635 ;
  assign n4637 = n821 & n4636 ;
  assign n4638 = ( n822 & n3424 ) | ( n822 & n4637 ) | ( n3424 & n4637 ) ;
  buffer buf_n4639( .i (n4638), .o (n4639) );
  assign n4641 = n2545 | n3191 ;
  assign n4642 = n3408 | n4641 ;
  assign n4643 = n3877 | n4642 ;
  assign n4644 = n4218 | n4643 ;
  assign n4645 = n4124 | n4644 ;
  assign n4646 = ( ~n2559 & n4639 ) | ( ~n2559 & n4645 ) | ( n4639 & n4645 ) ;
  assign n4647 = n2560 | n4646 ;
  buffer buf_n4648( .i (n4647), .o (n4648) );
  buffer buf_n4649( .i (n4648), .o (n4649) );
  assign n4650 = n3608 | n4299 ;
  assign n4651 = n4065 | n4650 ;
  assign n4652 = n3718 | n4367 ;
  assign n4653 = ( ~n4034 & n4651 ) | ( ~n4034 & n4652 ) | ( n4651 & n4652 ) ;
  assign n4654 = n4035 | n4653 ;
  buffer buf_n4655( .i (n4044), .o (n4655) );
  assign n4656 = n4347 & ~n4655 ;
  buffer buf_n4657( .i (n4656), .o (n4657) );
  buffer buf_n4658( .i (n4657), .o (n4658) );
  buffer buf_n4659( .i (n4658), .o (n4659) );
  buffer buf_n4660( .i (n4659), .o (n4660) );
  assign n4661 = ( n314 & ~n3105 ) | ( n314 & n4660 ) | ( ~n3105 & n4660 ) ;
  assign n4662 = ~n315 & n4661 ;
  buffer buf_n4663( .i (n3926), .o (n4663) );
  assign n4664 = n4662 & n4663 ;
  buffer buf_n4665( .i (n4001), .o (n4665) );
  buffer buf_n4666( .i (n4665), .o (n4666) );
  assign n4667 = ( n680 & n4664 ) | ( n680 & n4666 ) | ( n4664 & n4666 ) ;
  assign n4668 = ~n568 & n4667 ;
  buffer buf_n4669( .i (n4668), .o (n4669) );
  buffer buf_n4670( .i (n4669), .o (n4670) );
  assign n4671 = n3487 | n4670 ;
  assign n4672 = ( ~n3381 & n3498 ) | ( ~n3381 & n4671 ) | ( n3498 & n4671 ) ;
  assign n4673 = n3382 | n4672 ;
  buffer buf_n4674( .i (n4673), .o (n4674) );
  assign n4675 = n4654 | n4674 ;
  assign n4676 = ( n4424 & ~n4648 ) | ( n4424 & n4675 ) | ( ~n4648 & n4675 ) ;
  assign n4677 = n4649 | n4676 ;
  assign n4678 = ( n3341 & ~n3918 ) | ( n3341 & n4461 ) | ( ~n3918 & n4461 ) ;
  assign n4679 = n3919 | n4678 ;
  assign n4680 = n4010 | n4679 ;
  assign n4681 = ( ~n1652 & n2724 ) | ( ~n1652 & n4680 ) | ( n2724 & n4680 ) ;
  assign n4682 = n1653 | n4681 ;
  buffer buf_n4683( .i (n4682), .o (n4683) );
  buffer buf_n4684( .i (n4683), .o (n4684) );
  assign n4685 = n2660 | n3521 ;
  assign n4686 = ( ~n1617 & n3646 ) | ( ~n1617 & n4685 ) | ( n3646 & n4685 ) ;
  assign n4687 = n1618 | n4686 ;
  assign n4688 = n3621 | n4687 ;
  assign n4689 = ( n2362 & ~n3631 ) | ( n2362 & n4688 ) | ( ~n3631 & n4688 ) ;
  assign n4690 = n3632 | n4689 ;
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  assign n4691 = ( n679 & n1398 ) | ( n679 & ~n4632 ) | ( n1398 & ~n4632 ) ;
  assign n4692 = n4633 & n4691 ;
  buffer buf_n4693( .i (n4692), .o (n4693) );
  buffer buf_n4694( .i (n4693), .o (n4694) );
  buffer buf_n4695( .i (n4694), .o (n4695) );
  assign n4701 = ( n598 & n3297 ) | ( n598 & n3310 ) | ( n3297 & n3310 ) ;
  buffer buf_n4702( .i (n4272), .o (n4702) );
  assign n4703 = ~n4701 & n4702 ;
  buffer buf_n4704( .i (n4702), .o (n4704) );
  assign n4705 = ( n3299 & ~n4703 ) | ( n3299 & n4704 ) | ( ~n4703 & n4704 ) ;
  assign n4706 = n3316 | n4705 ;
  assign n4707 = n4695 | n4706 ;
  assign n4708 = n3933 | n4707 ;
  assign n4709 = ( n2651 & ~n3728 ) | ( n2651 & n4708 ) | ( ~n3728 & n4708 ) ;
  assign n4710 = n3729 | n4709 ;
  buffer buf_n3967( .i (n3966), .o (n3967) );
  buffer buf_n3968( .i (n3967), .o (n3968) );
  buffer buf_n3969( .i (n3968), .o (n3969) );
  buffer buf_n3970( .i (n3969), .o (n3970) );
  buffer buf_n3971( .i (n3970), .o (n3971) );
  buffer buf_n3972( .i (n3971), .o (n3972) );
  buffer buf_n3984( .i (n3983), .o (n3984) );
  buffer buf_n3985( .i (n3984), .o (n3985) );
  buffer buf_n3986( .i (n3985), .o (n3986) );
  buffer buf_n3987( .i (n3986), .o (n3987) );
  assign n4711 = n3946 | n4174 ;
  buffer buf_n4712( .i (n4711), .o (n4712) );
  assign n4723 = n3537 | n4194 ;
  assign n4724 = n4712 | n4723 ;
  assign n4725 = n3987 | n4724 ;
  assign n4726 = ( n2687 & ~n3971 ) | ( n2687 & n4725 ) | ( ~n3971 & n4725 ) ;
  assign n4727 = n3972 | n4726 ;
  assign n4728 = n4710 | n4727 ;
  assign n4729 = ( ~n4683 & n4690 ) | ( ~n4683 & n4728 ) | ( n4690 & n4728 ) ;
  assign n4730 = n4684 | n4729 ;
  assign n4731 = n4677 | n4730 ;
  assign n4732 = ( ~n4520 & n4630 ) | ( ~n4520 & n4731 ) | ( n4630 & n4731 ) ;
  assign n4733 = n4521 | n4732 ;
  assign n4734 = n2903 | n3896 ;
  assign n4735 = n3933 | n4734 ;
  buffer buf_n4736( .i (n4735), .o (n4736) );
  buffer buf_n4737( .i (n4736), .o (n4737) );
  buffer buf_n4738( .i (n4737), .o (n4738) );
  buffer buf_n4739( .i (n4738), .o (n4739) );
  buffer buf_n4740( .i (n4739), .o (n4740) );
  buffer buf_n4741( .i (n4740), .o (n4741) );
  buffer buf_n4742( .i (n4741), .o (n4742) );
  buffer buf_n4743( .i (n4742), .o (n4743) );
  buffer buf_n4179( .i (n4178), .o (n4179) );
  buffer buf_n4180( .i (n4179), .o (n4180) );
  buffer buf_n4181( .i (n4180), .o (n4181) );
  buffer buf_n4182( .i (n4181), .o (n4182) );
  buffer buf_n4183( .i (n4182), .o (n4183) );
  buffer buf_n4184( .i (n4183), .o (n4184) );
  buffer buf_n4185( .i (n4184), .o (n4185) );
  buffer buf_n4186( .i (n4185), .o (n4186) );
  buffer buf_n4143( .i (n4142), .o (n4143) );
  buffer buf_n4144( .i (n4143), .o (n4144) );
  buffer buf_n4145( .i (n4144), .o (n4145) );
  buffer buf_n4146( .i (n4145), .o (n4146) );
  buffer buf_n4147( .i (n4146), .o (n4147) );
  buffer buf_n4148( .i (n4147), .o (n4148) );
  buffer buf_n4149( .i (n4148), .o (n4149) );
  buffer buf_n4150( .i (n4149), .o (n4150) );
  buffer buf_n4640( .i (n4639), .o (n4640) );
  assign n4744 = n3410 | n3782 ;
  assign n4745 = n3672 | n4744 ;
  assign n4746 = n3360 | n4745 ;
  assign n4747 = ( ~n3394 & n4640 ) | ( ~n3394 & n4746 ) | ( n4640 & n4746 ) ;
  assign n4748 = n3395 | n4747 ;
  buffer buf_n4350( .i (n4349), .o (n4350) );
  buffer buf_n4351( .i (n4350), .o (n4351) );
  buffer buf_n4352( .i (n4351), .o (n4352) );
  buffer buf_n4749( .i (n4055), .o (n4749) );
  buffer buf_n4750( .i (n4749), .o (n4750) );
  assign n4751 = ( n3979 & n4352 ) | ( n3979 & ~n4750 ) | ( n4352 & ~n4750 ) ;
  assign n4752 = ~n4605 & n4751 ;
  assign n4753 = n4663 & n4752 ;
  assign n4754 = n598 & n4753 ;
  buffer buf_n4755( .i (n4754), .o (n4755) );
  assign n4759 = n4364 | n4755 ;
  buffer buf_n4760( .i (n4759), .o (n4760) );
  buffer buf_n4761( .i (n4760), .o (n4761) );
  buffer buf_n4762( .i (n4761), .o (n4762) );
  buffer buf_n4763( .i (n4762), .o (n4763) );
  buffer buf_n4764( .i (n4763), .o (n4764) );
  assign n4765 = n4674 | n4764 ;
  assign n4766 = ( ~n4149 & n4748 ) | ( ~n4149 & n4765 ) | ( n4748 & n4765 ) ;
  assign n4767 = n4150 | n4766 ;
  buffer buf_n4768( .i (n4767), .o (n4768) );
  buffer buf_n4769( .i (n4768), .o (n4769) );
  buffer buf_n3635( .i (n3634), .o (n3635) );
  buffer buf_n3527( .i (n3526), .o (n3527) );
  buffer buf_n3528( .i (n3527), .o (n3528) );
  buffer buf_n3650( .i (n3649), .o (n3650) );
  buffer buf_n3651( .i (n3650), .o (n3651) );
  buffer buf_n4713( .i (n4712), .o (n4713) );
  buffer buf_n4714( .i (n4713), .o (n4714) );
  buffer buf_n4715( .i (n4714), .o (n4715) );
  buffer buf_n4716( .i (n4715), .o (n4716) );
  buffer buf_n3540( .i (n3539), .o (n3540) );
  buffer buf_n3541( .i (n3540), .o (n3541) );
  assign n4770 = ( n2673 & n2918 ) | ( n2673 & n4188 ) | ( n2918 & n4188 ) ;
  assign n4771 = ~n4170 & n4770 ;
  buffer buf_n4772( .i (n4771), .o (n4772) );
  buffer buf_n4773( .i (n4772), .o (n4773) );
  buffer buf_n4774( .i (n4773), .o (n4774) );
  buffer buf_n4775( .i (n4774), .o (n4775) );
  buffer buf_n4776( .i (n4775), .o (n4776) );
  buffer buf_n4777( .i (n4776), .o (n4777) );
  buffer buf_n4778( .i (n4777), .o (n4778) );
  buffer buf_n4779( .i (n4778), .o (n4779) );
  assign n4780 = n3541 | n4779 ;
  assign n4781 = n4716 | n4780 ;
  assign n4782 = n3651 | n4781 ;
  assign n4783 = ( n3528 & ~n3634 ) | ( n3528 & n4782 ) | ( ~n3634 & n4782 ) ;
  assign n4784 = n3635 | n4783 ;
  buffer buf_n4551( .i (n4550), .o (n4551) );
  buffer buf_n4552( .i (n4551), .o (n4552) );
  buffer buf_n4553( .i (n4552), .o (n4553) );
  buffer buf_n4554( .i (n4553), .o (n4554) );
  buffer buf_n4555( .i (n4554), .o (n4555) );
  buffer buf_n4696( .i (n4695), .o (n4696) );
  buffer buf_n4697( .i (n4696), .o (n4697) );
  buffer buf_n4698( .i (n4697), .o (n4698) );
  buffer buf_n4699( .i (n4698), .o (n4699) );
  buffer buf_n4700( .i (n4699), .o (n4700) );
  buffer buf_n3551( .i (n3550), .o (n3551) );
  buffer buf_n3552( .i (n3551), .o (n3552) );
  buffer buf_n3553( .i (n3552), .o (n3553) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n3335( .i (n3334), .o (n3335) );
  buffer buf_n3336( .i (n3335), .o (n3336) );
  buffer buf_n3337( .i (n3336), .o (n3337) );
  buffer buf_n3338( .i (n3337), .o (n3338) );
  assign n4785 = n602 & n3338 ;
  buffer buf_n4786( .i (n4785), .o (n4786) );
  buffer buf_n4787( .i (n4786), .o (n4787) );
  buffer buf_n4788( .i (n4787), .o (n4788) );
  assign n4789 = n3553 | n4788 ;
  assign n4790 = ( ~n4554 & n4700 ) | ( ~n4554 & n4789 ) | ( n4700 & n4789 ) ;
  assign n4791 = n4555 | n4790 ;
  buffer buf_n4569( .i (n4568), .o (n4569) );
  buffer buf_n4570( .i (n4569), .o (n4570) );
  buffer buf_n4571( .i (n4570), .o (n4571) );
  buffer buf_n4572( .i (n4571), .o (n4572) );
  buffer buf_n4573( .i (n4572), .o (n4573) );
  buffer buf_n4574( .i (n4573), .o (n4574) );
  buffer buf_n4575( .i (n4574), .o (n4575) );
  buffer buf_n3580( .i (n3579), .o (n3580) );
  buffer buf_n3581( .i (n3580), .o (n3581) );
  buffer buf_n3582( .i (n3581), .o (n3582) );
  buffer buf_n3583( .i (n3582), .o (n3583) );
  buffer buf_n3584( .i (n3583), .o (n3584) );
  buffer buf_n3585( .i (n3584), .o (n3585) );
  buffer buf_n3586( .i (n3585), .o (n3586) );
  buffer buf_n3587( .i (n3586), .o (n3587) );
  buffer buf_n3588( .i (n3587), .o (n3588) );
  buffer buf_n3589( .i (n3588), .o (n3589) );
  buffer buf_n4600( .i (n4599), .o (n4600) );
  buffer buf_n4613( .i (n4612), .o (n4613) );
  buffer buf_n4614( .i (n4613), .o (n4614) );
  buffer buf_n4615( .i (n4614), .o (n4615) );
  assign n4792 = n4600 | n4615 ;
  assign n4793 = ( n3589 & ~n4574 ) | ( n3589 & n4792 ) | ( ~n4574 & n4792 ) ;
  assign n4794 = n4575 | n4793 ;
  assign n4795 = n4791 | n4794 ;
  assign n4796 = ( ~n4768 & n4784 ) | ( ~n4768 & n4795 ) | ( n4784 & n4795 ) ;
  assign n4797 = n4769 | n4796 ;
  assign n4798 = n3535 | n3546 ;
  assign n4799 = ( ~n3626 & n3669 ) | ( ~n3626 & n4798 ) | ( n3669 & n4798 ) ;
  assign n4800 = n3627 | n4799 ;
  buffer buf_n4801( .i (n4800), .o (n4801) );
  buffer buf_n4802( .i (n4801), .o (n4802) );
  buffer buf_n4803( .i (n4802), .o (n4803) );
  buffer buf_n4804( .i (n4803), .o (n4804) );
  buffer buf_n4805( .i (n4804), .o (n4805) );
  buffer buf_n4806( .i (n4805), .o (n4806) );
  buffer buf_n4807( .i (n4806), .o (n4807) );
  buffer buf_n4808( .i (n4807), .o (n4808) );
  buffer buf_n4809( .i (n4808), .o (n4809) );
  buffer buf_n4810( .i (n4809), .o (n4810) );
  assign n4811 = n4010 | n4160 ;
  assign n4812 = ( ~n1652 & n3921 ) | ( ~n1652 & n4811 ) | ( n3921 & n4811 ) ;
  assign n4813 = n1653 | n4812 ;
  buffer buf_n3879( .i (n3878), .o (n3879) );
  assign n4814 = n3879 | n4065 ;
  assign n4815 = n4034 | n4814 ;
  assign n4816 = n3866 | n4815 ;
  assign n4817 = ( ~n1503 & n4813 ) | ( ~n1503 & n4816 ) | ( n4813 & n4816 ) ;
  assign n4818 = n1504 | n4817 ;
  buffer buf_n4819( .i (n4818), .o (n4819) );
  buffer buf_n4820( .i (n4819), .o (n4820) );
  buffer buf_n4821( .i (n4820), .o (n4821) );
  buffer buf_n4822( .i (n4821), .o (n4822) );
  buffer buf_n2930( .i (n2929), .o (n2930) );
  buffer buf_n2931( .i (n2930), .o (n2931) );
  buffer buf_n2932( .i (n2931), .o (n2932) );
  buffer buf_n2933( .i (n2932), .o (n2933) );
  buffer buf_n4618( .i (n4617), .o (n4618) );
  buffer buf_n4619( .i (n4618), .o (n4619) );
  buffer buf_n4620( .i (n4619), .o (n4620) );
  buffer buf_n4621( .i (n4620), .o (n4621) );
  buffer buf_n4601( .i (n4600), .o (n4601) );
  buffer buf_n3142( .i (n3141), .o (n3142) );
  buffer buf_n3143( .i (n3142), .o (n3143) );
  assign n4823 = n3133 | n3143 ;
  assign n4824 = n4601 | n4823 ;
  buffer buf_n413( .i (x16), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n231( .i (x7), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  assign n4825 = ( n249 & n431 ) | ( n249 & n1215 ) | ( n431 & n1215 ) ;
  assign n4826 = ~n432 & n4825 ;
  buffer buf_n4827( .i (n4826), .o (n4827) );
  buffer buf_n4828( .i (n4827), .o (n4828) );
  assign n4829 = ( n1816 & n4749 ) | ( n1816 & ~n4827 ) | ( n4749 & ~n4827 ) ;
  assign n4830 = n4828 & n4829 ;
  buffer buf_n4831( .i (n4188), .o (n4831) );
  assign n4832 = ( n3015 & n4830 ) | ( n3015 & n4831 ) | ( n4830 & n4831 ) ;
  assign n4833 = ~n4253 & n4832 ;
  buffer buf_n4834( .i (n4833), .o (n4834) );
  buffer buf_n4835( .i (n4834), .o (n4835) );
  buffer buf_n4836( .i (n4835), .o (n4836) );
  buffer buf_n4837( .i (n4836), .o (n4837) );
  buffer buf_n4838( .i (n4837), .o (n4838) );
  buffer buf_n4839( .i (n4838), .o (n4839) );
  buffer buf_n4840( .i (n4839), .o (n4840) );
  buffer buf_n4841( .i (n4840), .o (n4841) );
  buffer buf_n4842( .i (n4841), .o (n4842) );
  buffer buf_n3017( .i (n3016), .o (n3017) );
  buffer buf_n253( .i (x8), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  assign n4843 = n432 & n4539 ;
  assign n4844 = ( n273 & n3997 ) | ( n273 & n4843 ) | ( n3997 & n4843 ) ;
  assign n4845 = ~n3954 & n4844 ;
  buffer buf_n4846( .i (n4845), .o (n4846) );
  buffer buf_n4847( .i (n4846), .o (n4847) );
  assign n4848 = ( n1818 & n4001 ) | ( n1818 & ~n4846 ) | ( n4001 & ~n4846 ) ;
  assign n4849 = n4847 & n4848 ;
  assign n4850 = ( n3017 & n4255 ) | ( n3017 & n4849 ) | ( n4255 & n4849 ) ;
  assign n4851 = ~n2235 & n4850 ;
  buffer buf_n4852( .i (n4851), .o (n4852) );
  buffer buf_n4853( .i (n4852), .o (n4853) );
  buffer buf_n4854( .i (n4853), .o (n4854) );
  buffer buf_n4855( .i (n4854), .o (n4855) );
  buffer buf_n4856( .i (n4855), .o (n4856) );
  buffer buf_n4857( .i (n4856), .o (n4857) );
  buffer buf_n3115( .i (n3114), .o (n3115) );
  buffer buf_n3074( .i (n3073), .o (n3074) );
  buffer buf_n3075( .i (n3074), .o (n3075) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n4048( .i (n4047), .o (n4048) );
  buffer buf_n4049( .i (n4048), .o (n4049) );
  buffer buf_n4050( .i (n4049), .o (n4050) );
  buffer buf_n4051( .i (n4050), .o (n4051) );
  buffer buf_n4052( .i (n4051), .o (n4052) );
  assign n4858 = n4052 & n4665 ;
  buffer buf_n4859( .i (n597), .o (n4859) );
  assign n4860 = ( n2718 & n4858 ) | ( n2718 & n4859 ) | ( n4858 & n4859 ) ;
  assign n4861 = ~n1823 & n4860 ;
  assign n4862 = n1237 & n4861 ;
  buffer buf_n4863( .i (n4862), .o (n4863) );
  buffer buf_n4864( .i (n4863), .o (n4864) );
  buffer buf_n4865( .i (n4864), .o (n4865) );
  assign n4866 = n3075 | n4865 ;
  assign n4867 = n3115 | n4866 ;
  assign n4868 = n4857 | n4867 ;
  assign n4869 = n4842 | n4868 ;
  assign n4870 = n4824 | n4869 ;
  assign n4871 = ( ~n2932 & n4621 ) | ( ~n2932 & n4870 ) | ( n4621 & n4870 ) ;
  assign n4872 = n2933 | n4871 ;
  buffer buf_n3764( .i (n3763), .o (n3764) );
  buffer buf_n3765( .i (n3764), .o (n3765) );
  buffer buf_n3766( .i (n3765), .o (n3766) );
  buffer buf_n3767( .i (n3766), .o (n3767) );
  buffer buf_n3768( .i (n3767), .o (n3768) );
  buffer buf_n4406( .i (n4405), .o (n4406) );
  buffer buf_n4407( .i (n4406), .o (n4407) );
  buffer buf_n4408( .i (n4407), .o (n4408) );
  buffer buf_n3845( .i (n3844), .o (n3845) );
  assign n4873 = n3212 | n3845 ;
  assign n4874 = ( n3768 & ~n4408 ) | ( n3768 & n4873 ) | ( ~n4408 & n4873 ) ;
  buffer buf_n4875( .i (n4874), .o (n4875) );
  buffer buf_n4876( .i (n4875), .o (n4876) );
  assign n4877 = n3315 | n4693 ;
  assign n4878 = n3300 | n4877 ;
  buffer buf_n4879( .i (n4878), .o (n4879) );
  buffer buf_n4880( .i (n4879), .o (n4880) );
  buffer buf_n4881( .i (n4880), .o (n4881) );
  buffer buf_n4882( .i (n4881), .o (n4882) );
  assign n4883 = n3344 | n4786 ;
  buffer buf_n4756( .i (n4755), .o (n4756) );
  buffer buf_n4757( .i (n4756), .o (n4757) );
  buffer buf_n4758( .i (n4757), .o (n4758) );
  assign n4884 = n4191 | n4772 ;
  buffer buf_n4885( .i (n4884), .o (n4885) );
  buffer buf_n4886( .i (n4885), .o (n4886) );
  buffer buf_n4887( .i (n4886), .o (n4887) );
  assign n4888 = n4670 | n4887 ;
  assign n4889 = ( ~n4367 & n4758 ) | ( ~n4367 & n4888 ) | ( n4758 & n4888 ) ;
  assign n4890 = n4368 | n4889 ;
  assign n4891 = n4883 | n4890 ;
  assign n4892 = ( ~n4180 & n4882 ) | ( ~n4180 & n4891 ) | ( n4882 & n4891 ) ;
  assign n4893 = n4181 | n4892 ;
  buffer buf_n4411( .i (n4410), .o (n4411) );
  buffer buf_n4412( .i (n4411), .o (n4412) );
  assign n4894 = n3802 | n3807 ;
  buffer buf_n4895( .i (n4894), .o (n4895) );
  buffer buf_n4896( .i (n4895), .o (n4896) );
  buffer buf_n4897( .i (n4896), .o (n4897) );
  buffer buf_n4898( .i (n4897), .o (n4898) );
  buffer buf_n4899( .i (n4898), .o (n4899) );
  assign n4900 = n4412 | n4899 ;
  assign n4901 = ( ~n4875 & n4893 ) | ( ~n4875 & n4900 ) | ( n4893 & n4900 ) ;
  assign n4902 = n4876 | n4901 ;
  buffer buf_n4556( .i (n4555), .o (n4556) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  assign n4903 = ( n202 & n1665 ) | ( n202 & n3979 ) | ( n1665 & n3979 ) ;
  assign n4904 = ~n4605 & n4903 ;
  buffer buf_n4905( .i (n4750), .o (n4905) );
  assign n4906 = ~n3836 & n4905 ;
  assign n4907 = ( n679 & n4904 ) | ( n679 & n4906 ) | ( n4904 & n4906 ) ;
  assign n4908 = ~n680 & n4907 ;
  assign n4909 = n1236 & n4908 ;
  buffer buf_n4910( .i (n4909), .o (n4910) );
  buffer buf_n4911( .i (n4910), .o (n4911) );
  buffer buf_n4912( .i (n4911), .o (n4912) );
  buffer buf_n4913( .i (n4912), .o (n4913) );
  buffer buf_n4914( .i (n4913), .o (n4914) );
  buffer buf_n4915( .i (n4914), .o (n4915) );
  buffer buf_n4916( .i (n4915), .o (n4916) );
  buffer buf_n4263( .i (n4262), .o (n4263) );
  assign n4917 = n198 & n310 ;
  assign n4918 = ( n4539 & n4585 ) | ( n4539 & n4917 ) | ( n4585 & n4917 ) ;
  assign n4919 = ~n4540 & n4918 ;
  buffer buf_n4920( .i (n4919), .o (n4920) );
  buffer buf_n4921( .i (n4920), .o (n4921) );
  assign n4922 = ( n1715 & n4750 ) | ( n1715 & ~n4920 ) | ( n4750 & ~n4920 ) ;
  assign n4923 = n4921 & n4922 ;
  buffer buf_n4924( .i (n3836), .o (n4924) );
  assign n4925 = ( n4564 & n4923 ) | ( n4564 & n4924 ) | ( n4923 & n4924 ) ;
  buffer buf_n4926( .i (n4924), .o (n4926) );
  assign n4927 = n4925 & ~n4926 ;
  buffer buf_n4928( .i (n4927), .o (n4928) );
  buffer buf_n4929( .i (n4928), .o (n4929) );
  buffer buf_n4930( .i (n4929), .o (n4930) );
  buffer buf_n4931( .i (n4930), .o (n4931) );
  buffer buf_n4932( .i (n4931), .o (n4932) );
  buffer buf_n4933( .i (n4932), .o (n4933) );
  buffer buf_n4934( .i (n4933), .o (n4934) );
  assign n4935 = n4263 | n4934 ;
  assign n4936 = n4916 | n4935 ;
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  assign n4937 = n252 & ~n4356 ;
  buffer buf_n4938( .i (n3954), .o (n4938) );
  assign n4939 = ( n435 & n4937 ) | ( n435 & n4938 ) | ( n4937 & n4938 ) ;
  assign n4940 = ~n436 & n4939 ;
  buffer buf_n4941( .i (n4940), .o (n4941) );
  buffer buf_n4942( .i (n4941), .o (n4942) );
  buffer buf_n3958( .i (n3957), .o (n3958) );
  buffer buf_n3959( .i (n3958), .o (n3959) );
  buffer buf_n3960( .i (n3959), .o (n3960) );
  assign n4943 = ( n3960 & n4666 ) | ( n3960 & ~n4941 ) | ( n4666 & ~n4941 ) ;
  assign n4944 = n4942 & n4943 ;
  buffer buf_n4945( .i (n4944), .o (n4945) );
  buffer buf_n4946( .i (n4945), .o (n4946) );
  buffer buf_n4947( .i (n4946), .o (n4947) );
  buffer buf_n4948( .i (n4947), .o (n4948) );
  buffer buf_n4949( .i (n4948), .o (n4949) );
  assign n4950 = n273 & n433 ;
  assign n4951 = ( n3954 & n4356 ) | ( n3954 & n4950 ) | ( n4356 & n4950 ) ;
  buffer buf_n4952( .i (n4540), .o (n4952) );
  buffer buf_n4953( .i (n4952), .o (n4953) );
  assign n4954 = n4951 & ~n4953 ;
  buffer buf_n4955( .i (n4954), .o (n4955) );
  buffer buf_n4956( .i (n4955), .o (n4956) );
  assign n4957 = ( n3959 & n4665 ) | ( n3959 & ~n4955 ) | ( n4665 & ~n4955 ) ;
  assign n4958 = n4956 & n4957 ;
  buffer buf_n4959( .i (n4958), .o (n4959) );
  buffer buf_n4960( .i (n4959), .o (n4960) );
  buffer buf_n4961( .i (n4960), .o (n4961) );
  buffer buf_n4962( .i (n4961), .o (n4962) );
  buffer buf_n4963( .i (n4962), .o (n4963) );
  assign n4964 = n4278 | n4963 ;
  assign n4965 = ( ~n3232 & n4949 ) | ( ~n3232 & n4964 ) | ( n4949 & n4964 ) ;
  assign n4966 = n3233 | n4965 ;
  assign n4967 = n4574 | n4966 ;
  assign n4968 = ( ~n4555 & n4936 ) | ( ~n4555 & n4967 ) | ( n4936 & n4967 ) ;
  assign n4969 = n4556 | n4968 ;
  assign n4970 = n4902 | n4969 ;
  assign n4971 = n4872 | n4970 ;
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  assign n4972 = n1525 | n1565 ;
  assign n4973 = n1501 | n4972 ;
  assign n4974 = n1982 | n4973 ;
  assign n4975 = ( n1621 & ~n1965 ) | ( n1621 & n4974 ) | ( ~n1965 & n4974 ) ;
  assign n4976 = n1966 | n4975 ;
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  assign n4977 = n1803 | n1898 ;
  buffer buf_n4978( .i (n4977), .o (n4978) );
  assign n4979 = n1886 | n4978 ;
  assign n4980 = ( ~n1384 & n1783 ) | ( ~n1384 & n4979 ) | ( n1783 & n4979 ) ;
  assign n4981 = n1385 | n4980 ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  assign n4982 = n1444 | n1826 ;
  assign n4983 = n1428 | n4982 ;
  assign n4984 = n1873 | n4983 ;
  assign n4985 = ( ~n1725 & n4981 ) | ( ~n1725 & n4984 ) | ( n4981 & n4984 ) ;
  assign n4986 = n1726 | n4985 ;
  buffer buf_n1677( .i (n1676), .o (n1677) );
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  assign n4987 = n1650 | n1741 ;
  assign n4988 = n1631 | n4987 ;
  assign n4989 = n1699 | n4988 ;
  assign n4990 = ( n1408 & ~n1679 ) | ( n1408 & n4989 ) | ( ~n1679 & n4989 ) ;
  assign n4991 = n1680 | n4990 ;
  assign n4992 = n4986 | n4991 ;
  assign n4993 = n4976 | n4992 ;
  buffer buf_n4994( .i (n4993), .o (n4994) );
  buffer buf_n4995( .i (n4994), .o (n4995) );
  buffer buf_n4996( .i (n4995), .o (n4996) );
  buffer buf_n1994( .i (n1993), .o (n1994) );
  buffer buf_n1995( .i (n1994), .o (n1995) );
  buffer buf_n1996( .i (n1995), .o (n1996) );
  buffer buf_n1997( .i (n1996), .o (n1997) );
  buffer buf_n1998( .i (n1997), .o (n1998) );
  buffer buf_n1999( .i (n1998), .o (n1999) );
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n2001( .i (n2000), .o (n2001) );
  assign n4997 = n1925 | n1947 ;
  assign n4998 = n2001 | n4997 ;
  assign n4999 = n1482 | n2026 ;
  buffer buf_n5000( .i (n4999), .o (n5000) );
  assign n5001 = n1544 | n5000 ;
  assign n5002 = n4998 | n5001 ;
  buffer buf_n5003( .i (n5002), .o (n5003) );
  buffer buf_n5004( .i (n5003), .o (n5004) );
  buffer buf_n5005( .i (n5004), .o (n5005) );
  buffer buf_n5006( .i (n5005), .o (n5006) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n2037( .i (n2036), .o (n2037) );
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  assign n5007 = n1947 | n2039 ;
  assign n5008 = n2052 | n5007 ;
  buffer buf_n5009( .i (n1543), .o (n5009) );
  assign n5010 = n1600 | n5009 ;
  assign n5011 = n5008 | n5010 ;
  buffer buf_n5012( .i (n5011), .o (n5012) );
  buffer buf_n5013( .i (n5012), .o (n5013) );
  buffer buf_n5014( .i (n5013), .o (n5014) );
  buffer buf_n5015( .i (n5014), .o (n5015) );
  buffer buf_n342( .i (x12), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  assign n5016 = ~n345 & n542 ;
  assign n5017 = ( n343 & ~n368 ) | ( n343 & n5016 ) | ( ~n368 & n5016 ) ;
  assign n5018 = ~n344 & n5017 ;
  assign n5019 = ~n738 & n5018 ;
  assign n5020 = ( n715 & ~n767 ) | ( n715 & n5019 ) | ( ~n767 & n5019 ) ;
  assign n5021 = ~n716 & n5020 ;
  assign n5022 = ~n799 & n5021 ;
  buffer buf_n5023( .i (n5022), .o (n5023) );
  buffer buf_n5024( .i (n5023), .o (n5024) );
  buffer buf_n5025( .i (n5024), .o (n5025) );
  buffer buf_n5026( .i (n5025), .o (n5026) );
  buffer buf_n5027( .i (n5026), .o (n5027) );
  buffer buf_n5028( .i (n5027), .o (n5028) );
  buffer buf_n5029( .i (n5028), .o (n5029) );
  buffer buf_n5030( .i (n5029), .o (n5030) );
  buffer buf_n5031( .i (n5030), .o (n5031) );
  buffer buf_n5032( .i (n5031), .o (n5032) );
  buffer buf_n5033( .i (n5032), .o (n5033) );
  buffer buf_n5034( .i (n5033), .o (n5034) );
  buffer buf_n5035( .i (n5034), .o (n5035) );
  buffer buf_n5036( .i (n5035), .o (n5036) );
  buffer buf_n5037( .i (n5036), .o (n5037) );
  buffer buf_n5038( .i (n5037), .o (n5038) );
  buffer buf_n5039( .i (n5038), .o (n5039) );
  buffer buf_n5040( .i (n5039), .o (n5040) );
  buffer buf_n5041( .i (n5040), .o (n5041) );
  buffer buf_n5042( .i (n5041), .o (n5042) );
  buffer buf_n5043( .i (n5042), .o (n5043) );
  buffer buf_n5044( .i (n5043), .o (n5044) );
  buffer buf_n5045( .i (n5044), .o (n5045) );
  buffer buf_n5046( .i (n5045), .o (n5046) );
  buffer buf_n5047( .i (n5046), .o (n5047) );
  buffer buf_n5048( .i (n5047), .o (n5048) );
  buffer buf_n5049( .i (n5048), .o (n5049) );
  buffer buf_n5050( .i (n5049), .o (n5050) );
  buffer buf_n5051( .i (n5050), .o (n5051) );
  buffer buf_n5052( .i (n5051), .o (n5052) );
  buffer buf_n5053( .i (n5052), .o (n5053) );
  buffer buf_n5054( .i (n5053), .o (n5054) );
  buffer buf_n3880( .i (n3879), .o (n3880) );
  assign n5055 = n3850 | n3864 ;
  assign n5056 = ( ~n2451 & n3880 ) | ( ~n2451 & n5055 ) | ( n3880 & n5055 ) ;
  assign n5057 = n2452 | n5056 ;
  buffer buf_n5058( .i (n5057), .o (n5058) );
  buffer buf_n5059( .i (n5058), .o (n5059) );
  buffer buf_n5060( .i (n5059), .o (n5060) );
  buffer buf_n5061( .i (n5060), .o (n5061) );
  buffer buf_n5062( .i (n5061), .o (n5062) );
  buffer buf_n5063( .i (n5062), .o (n5063) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  buffer buf_n2203( .i (n2202), .o (n2203) );
  buffer buf_n2204( .i (n2203), .o (n2204) );
  buffer buf_n2205( .i (n2204), .o (n2205) );
  buffer buf_n2206( .i (n2205), .o (n2206) );
  buffer buf_n2404( .i (n2403), .o (n2404) );
  assign n5064 = n2206 | n2404 ;
  assign n5065 = n2383 | n5064 ;
  assign n5066 = n2185 | n3697 ;
  assign n5067 = n2985 | n5066 ;
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n2419( .i (n2418), .o (n2419) );
  buffer buf_n2420( .i (n2419), .o (n2420) );
  buffer buf_n2421( .i (n2420), .o (n2421) );
  buffer buf_n2422( .i (n2421), .o (n2422) );
  buffer buf_n2423( .i (n2422), .o (n2423) );
  buffer buf_n5068( .i (n849), .o (n5068) );
  assign n5069 = n2417 & n5068 ;
  buffer buf_n5070( .i (n5069), .o (n5070) );
  buffer buf_n5071( .i (n5070), .o (n5071) );
  buffer buf_n5072( .i (n5071), .o (n5072) );
  buffer buf_n5073( .i (n5072), .o (n5073) );
  buffer buf_n5074( .i (n5073), .o (n5074) );
  assign n5075 = ( ~n916 & n2423 ) | ( ~n916 & n5074 ) | ( n2423 & n5074 ) ;
  assign n5076 = n5067 | n5075 ;
  assign n5077 = n5065 | n5076 ;
  buffer buf_n5078( .i (n5077), .o (n5078) );
  buffer buf_n5079( .i (n5078), .o (n5079) );
  buffer buf_n3253( .i (n3252), .o (n3253) );
  buffer buf_n3254( .i (n3253), .o (n3254) );
  buffer buf_n3255( .i (n3254), .o (n3255) );
  buffer buf_n3256( .i (n3255), .o (n3256) );
  buffer buf_n3257( .i (n3256), .o (n3257) );
  buffer buf_n3258( .i (n3257), .o (n3258) );
  buffer buf_n3259( .i (n3258), .o (n3259) );
  buffer buf_n3067( .i (n3066), .o (n3067) );
  buffer buf_n3068( .i (n3067), .o (n3068) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  assign n5080 = n1299 | n1339 ;
  assign n5081 = n2799 | n5080 ;
  buffer buf_n5082( .i (n5081), .o (n5082) );
  buffer buf_n5083( .i (n5082), .o (n5083) );
  assign n5084 = ( n1448 & ~n3067 ) | ( n1448 & n5083 ) | ( ~n3067 & n5083 ) ;
  assign n5085 = n3068 | n5084 ;
  buffer buf_n4524( .i (n4523), .o (n4524) );
  buffer buf_n4525( .i (n4524), .o (n4525) );
  buffer buf_n4526( .i (n4525), .o (n4526) );
  buffer buf_n4527( .i (n4526), .o (n4527) );
  buffer buf_n4528( .i (n4527), .o (n4528) );
  buffer buf_n4529( .i (n4528), .o (n4529) );
  buffer buf_n4530( .i (n4529), .o (n4530) );
  buffer buf_n3237( .i (n3236), .o (n3237) );
  buffer buf_n3238( .i (n3237), .o (n3238) );
  buffer buf_n3239( .i (n3238), .o (n3239) );
  buffer buf_n3240( .i (n3239), .o (n3240) );
  buffer buf_n3241( .i (n3240), .o (n3241) );
  assign n5086 = n2725 | n3729 ;
  assign n5087 = n3241 | n5086 ;
  assign n5088 = n4530 | n5087 ;
  assign n5089 = ( ~n3258 & n5085 ) | ( ~n3258 & n5088 ) | ( n5085 & n5088 ) ;
  assign n5090 = n3259 | n5089 ;
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  buffer buf_n1584( .i (n1583), .o (n1584) );
  assign n5091 = n2039 | n3028 ;
  assign n5092 = n2052 | n5091 ;
  buffer buf_n3047( .i (n3046), .o (n3047) );
  buffer buf_n3048( .i (n3047), .o (n3048) );
  buffer buf_n2486( .i (n2485), .o (n2486) );
  buffer buf_n2487( .i (n2486), .o (n2487) );
  assign n5093 = n2487 & n4704 ;
  buffer buf_n5094( .i (n5093), .o (n5094) );
  buffer buf_n5095( .i (n5094), .o (n5095) );
  buffer buf_n5096( .i (n5095), .o (n5096) );
  assign n5097 = n1523 | n2493 ;
  assign n5098 = n1595 | n5097 ;
  assign n5099 = n1541 | n5098 ;
  assign n5100 = ( ~n3706 & n5096 ) | ( ~n3706 & n5099 ) | ( n5096 & n5099 ) ;
  assign n5101 = n3707 | n5100 ;
  assign n5102 = n3048 | n5101 ;
  assign n5103 = ( ~n1583 & n5092 ) | ( ~n1583 & n5102 ) | ( n5092 & n5102 ) ;
  assign n5104 = n1584 | n5103 ;
  buffer buf_n2676( .i (n2675), .o (n2676) );
  buffer buf_n2677( .i (n2676), .o (n2677) );
  buffer buf_n2678( .i (n2677), .o (n2678) );
  buffer buf_n2679( .i (n2678), .o (n2679) );
  buffer buf_n3018( .i (n3017), .o (n3018) );
  buffer buf_n3019( .i (n3018), .o (n3019) );
  buffer buf_n3020( .i (n3019), .o (n3020) );
  assign n5105 = ( n791 & n2679 ) | ( n791 & n3020 ) | ( n2679 & n3020 ) ;
  assign n5106 = ~n792 & n5105 ;
  buffer buf_n5107( .i (n5106), .o (n5107) );
  buffer buf_n5108( .i (n5107), .o (n5108) );
  buffer buf_n2713( .i (n2712), .o (n2713) );
  assign n5109 = ( ~n2713 & n3016 ) | ( ~n2713 & n4253 ) | ( n3016 & n4253 ) ;
  assign n5110 = ~n4255 & n5109 ;
  buffer buf_n5111( .i (n5110), .o (n5111) );
  assign n5112 = n1648 | n5111 ;
  buffer buf_n5113( .i (n5112), .o (n5113) );
  buffer buf_n5114( .i (n5113), .o (n5114) );
  assign n5115 = n2686 | n5114 ;
  assign n5116 = n1619 | n5115 ;
  assign n5117 = ( ~n2319 & n5108 ) | ( ~n2319 & n5116 ) | ( n5108 & n5116 ) ;
  assign n5118 = n2320 | n5117 ;
  buffer buf_n3478( .i (n3477), .o (n3478) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2325( .i (n2324), .o (n2325) );
  buffer buf_n2326( .i (n2325), .o (n2326) );
  buffer buf_n2327( .i (n2326), .o (n2327) );
  buffer buf_n5119( .i (n4831), .o (n5119) );
  buffer buf_n5120( .i (n5119), .o (n5120) );
  assign n5121 = n2327 & ~n5120 ;
  assign n5122 = ~n4702 & n5121 ;
  buffer buf_n5123( .i (n5122), .o (n5123) );
  buffer buf_n5124( .i (n5123), .o (n5124) );
  buffer buf_n5125( .i (n5124), .o (n5125) );
  buffer buf_n5126( .i (n5125), .o (n5126) );
  assign n5127 = n3458 | n5126 ;
  assign n5128 = n1947 | n5127 ;
  assign n5129 = n3478 | n5128 ;
  assign n5130 = ( ~n2243 & n5118 ) | ( ~n2243 & n5129 ) | ( n5118 & n5129 ) ;
  assign n5131 = n2244 | n5130 ;
  assign n5132 = n5104 | n5131 ;
  assign n5133 = ( ~n5078 & n5090 ) | ( ~n5078 & n5132 ) | ( n5090 & n5132 ) ;
  assign n5134 = n5079 | n5133 ;
  assign n5135 = n4020 | n4347 ;
  buffer buf_n5136( .i (n123), .o (n5136) );
  buffer buf_n5137( .i (n5136), .o (n5137) );
  assign n5138 = ( n223 & n5135 ) | ( n223 & ~n5137 ) | ( n5135 & ~n5137 ) ;
  assign n5139 = n126 | n5138 ;
  assign n5140 = n4055 | n5139 ;
  assign n5141 = ( n3977 & n4952 ) | ( n3977 & ~n5140 ) | ( n4952 & ~n5140 ) ;
  assign n5142 = ~n4953 & n5141 ;
  buffer buf_n5143( .i (n1434), .o (n5143) );
  assign n5144 = ( n4831 & n5142 ) | ( n4831 & n5143 ) | ( n5142 & n5143 ) ;
  assign n5145 = ~n5119 & n5144 ;
  buffer buf_n5146( .i (n5145), .o (n5146) );
  assign n5153 = n1614 | n5146 ;
  assign n5154 = n3520 | n5153 ;
  assign n5155 = n2331 | n3451 ;
  assign n5156 = ( n1940 & ~n1957 ) | ( n1940 & n5155 ) | ( ~n1957 & n5155 ) ;
  assign n5157 = n1958 | n5156 ;
  assign n5158 = n3644 | n5157 ;
  assign n5159 = ( ~n3627 & n5154 ) | ( ~n3627 & n5158 ) | ( n5154 & n5158 ) ;
  assign n5160 = n3628 | n5159 ;
  buffer buf_n5161( .i (n5160), .o (n5161) );
  buffer buf_n5162( .i (n5161), .o (n5162) );
  assign n5163 = n2003 | n3472 ;
  assign n5164 = ( ~n3379 & n3390 ) | ( ~n3379 & n5163 ) | ( n3390 & n5163 ) ;
  assign n5165 = n3380 | n5164 ;
  assign n5166 = n1921 | n3357 ;
  buffer buf_n5167( .i (n5166), .o (n5167) );
  assign n5170 = n5165 | n5167 ;
  assign n5171 = ( n2054 & ~n5161 ) | ( n2054 & n5170 ) | ( ~n5161 & n5170 ) ;
  assign n5172 = n5162 | n5171 ;
  buffer buf_n5173( .i (n5172), .o (n5173) );
  buffer buf_n5174( .i (n5173), .o (n5174) );
  assign n5175 = n1562 | n3408 ;
  buffer buf_n5176( .i (n5175), .o (n5176) );
  assign n5178 = n2024 | n5176 ;
  assign n5179 = ( ~n1481 & n3427 ) | ( ~n1481 & n5178 ) | ( n3427 & n5178 ) ;
  assign n5180 = n1482 | n5179 ;
  assign n5181 = n4221 | n5180 ;
  assign n5182 = n1600 | n5181 ;
  buffer buf_n2194( .i (n2193), .o (n2194) );
  buffer buf_n2195( .i (n2194), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  assign n5183 = n2461 | n3783 ;
  assign n5184 = ( ~n2195 & n2472 ) | ( ~n2195 & n5183 ) | ( n2472 & n5183 ) ;
  assign n5185 = n2196 | n5184 ;
  assign n5186 = n3863 | n5094 ;
  assign n5187 = n3879 | n5186 ;
  assign n5188 = n1542 | n5187 ;
  assign n5189 = n3005 | n5188 ;
  assign n5190 = n5185 | n5189 ;
  assign n5191 = ( ~n5173 & n5182 ) | ( ~n5173 & n5190 ) | ( n5182 & n5190 ) ;
  assign n5192 = n5174 | n5191 ;
  buffer buf_n5193( .i (n5192), .o (n5193) );
  buffer buf_n5194( .i (n5193), .o (n5194) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  assign n5195 = n1762 | n2888 ;
  buffer buf_n5196( .i (n5195), .o (n5196) );
  buffer buf_n5197( .i (n5196), .o (n5197) );
  buffer buf_n5198( .i (n5197), .o (n5198) );
  assign n5199 = n1804 | n2963 ;
  assign n5200 = ( ~n1383 & n2903 ) | ( ~n1383 & n5199 ) | ( n2903 & n5199 ) ;
  assign n5201 = n1384 | n5200 ;
  assign n5202 = n1905 | n5201 ;
  assign n5203 = ( ~n1780 & n5198 ) | ( ~n1780 & n5202 ) | ( n5198 & n5202 ) ;
  assign n5204 = n1781 | n5203 ;
  buffer buf_n5205( .i (n5204), .o (n5205) );
  buffer buf_n5206( .i (n5205), .o (n5206) );
  assign n5207 = n1870 | n2839 ;
  buffer buf_n5208( .i (n5207), .o (n5208) );
  buffer buf_n5209( .i (n5208), .o (n5209) );
  buffer buf_n5210( .i (n5209), .o (n5210) );
  buffer buf_n5211( .i (n5210), .o (n5211) );
  buffer buf_n5212( .i (n5211), .o (n5212) );
  buffer buf_n5213( .i (n5212), .o (n5213) );
  buffer buf_n4442( .i (n4441), .o (n4442) );
  buffer buf_n4443( .i (n4442), .o (n4443) );
  buffer buf_n5214( .i (n2756), .o (n5214) );
  assign n5215 = n1826 | n5214 ;
  buffer buf_n5216( .i (n5215), .o (n5216) );
  assign n5217 = n2800 | n5216 ;
  assign n5218 = ( n1447 & ~n2864 ) | ( n1447 & n5217 ) | ( ~n2864 & n5217 ) ;
  assign n5219 = n2865 | n5218 ;
  assign n5220 = n4443 | n5219 ;
  assign n5221 = ( ~n5205 & n5213 ) | ( ~n5205 & n5220 ) | ( n5213 & n5220 ) ;
  assign n5222 = n5206 | n5221 ;
  buffer buf_n1703( .i (n1702), .o (n1703) );
  assign n5223 = n1407 | n3898 ;
  assign n5224 = ( ~n1679 & n3935 ) | ( ~n1679 & n5223 ) | ( n3935 & n5223 ) ;
  assign n5225 = n1680 | n5224 ;
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n2817( .i (n2816), .o (n2817) );
  buffer buf_n2818( .i (n2817), .o (n2818) );
  assign n5226 = n1724 | n2818 ;
  assign n5227 = n1855 | n5226 ;
  assign n5228 = n3171 | n5227 ;
  assign n5229 = ( ~n1702 & n5225 ) | ( ~n1702 & n5228 ) | ( n5225 & n5228 ) ;
  assign n5230 = n1703 | n5229 ;
  buffer buf_n1633( .i (n1632), .o (n1633) );
  buffer buf_n1634( .i (n1633), .o (n1634) );
  buffer buf_n1635( .i (n1634), .o (n1635) );
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n4329( .i (n4328), .o (n4329) );
  buffer buf_n4330( .i (n4329), .o (n4330) );
  buffer buf_n4331( .i (n4330), .o (n4331) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n3961( .i (n3960), .o (n3961) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n3907( .i (n3906), .o (n3907) );
  buffer buf_n3908( .i (n3907), .o (n3908) );
  buffer buf_n3909( .i (n3908), .o (n3909) );
  buffer buf_n3910( .i (n3909), .o (n3910) );
  assign n5231 = ( n229 & n3910 ) | ( n229 & ~n4606 ) | ( n3910 & ~n4606 ) ;
  assign n5232 = ~n230 & n5231 ;
  assign n5233 = ( n568 & n3961 ) | ( n568 & n5232 ) | ( n3961 & n5232 ) ;
  assign n5234 = ~n569 & n5233 ;
  assign n5235 = n1238 & n5234 ;
  buffer buf_n5236( .i (n5235), .o (n5236) );
  buffer buf_n5237( .i (n5236), .o (n5237) );
  buffer buf_n5238( .i (n5237), .o (n5238) );
  buffer buf_n5239( .i (n5238), .o (n5239) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  assign n5240 = n152 | n4952 ;
  assign n5241 = ( ~n129 & n4938 ) | ( ~n129 & n5240 ) | ( n4938 & n5240 ) ;
  assign n5242 = n130 | n5241 ;
  assign n5243 = n4004 | n5242 ;
  assign n5244 = n4666 | n5243 ;
  buffer buf_n5245( .i (n5120), .o (n5245) );
  buffer buf_n5246( .i (n1437), .o (n5246) );
  assign n5247 = ( ~n5244 & n5245 ) | ( ~n5244 & n5246 ) | ( n5245 & n5246 ) ;
  assign n5248 = ~n2034 & n5247 ;
  buffer buf_n5249( .i (n5248), .o (n5249) );
  buffer buf_n5250( .i (n5249), .o (n5250) );
  buffer buf_n5251( .i (n5250), .o (n5251) );
  assign n5252 = n1742 | n4463 ;
  buffer buf_n5253( .i (n1651), .o (n5253) );
  assign n5254 = ( n5251 & n5252 ) | ( n5251 & ~n5253 ) | ( n5252 & ~n5253 ) ;
  buffer buf_n5255( .i (n5253), .o (n5255) );
  assign n5256 = n5254 | n5255 ;
  assign n5257 = n5239 | n5256 ;
  assign n5258 = ( ~n1635 & n4331 ) | ( ~n1635 & n5257 ) | ( n4331 & n5257 ) ;
  assign n5259 = n1636 | n5258 ;
  assign n5260 = n5230 | n5259 ;
  assign n5261 = ( ~n5193 & n5222 ) | ( ~n5193 & n5260 ) | ( n5222 & n5260 ) ;
  assign n5262 = n5194 | n5261 ;
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n3043( .i (n3042), .o (n3043) );
  assign n5263 = n2497 | n4214 ;
  assign n5264 = n3043 | n5263 ;
  buffer buf_n3693( .i (n3692), .o (n3693) );
  buffer buf_n3694( .i (n3693), .o (n3694) );
  assign n5265 = n1498 | n3001 ;
  assign n5266 = n1540 | n5265 ;
  assign n5267 = n2194 | n5266 ;
  buffer buf_n5268( .i (n3705), .o (n5268) );
  assign n5269 = ( ~n3693 & n5267 ) | ( ~n3693 & n5268 ) | ( n5267 & n5268 ) ;
  assign n5270 = n3694 | n5269 ;
  assign n5271 = n5000 | n5270 ;
  assign n5272 = ( ~n1569 & n5264 ) | ( ~n1569 & n5271 ) | ( n5264 & n5271 ) ;
  assign n5273 = n1570 | n5272 ;
  buffer buf_n5274( .i (n5273), .o (n5274) );
  buffer buf_n5275( .i (n5274), .o (n5275) );
  buffer buf_n2955( .i (n2954), .o (n2955) );
  buffer buf_n2956( .i (n2955), .o (n2956) );
  buffer buf_n2957( .i (n2956), .o (n2957) );
  buffer buf_n2958( .i (n2957), .o (n2958) );
  buffer buf_n2959( .i (n2958), .o (n2959) );
  buffer buf_n2960( .i (n2959), .o (n2960) );
  buffer buf_n2916( .i (n2915), .o (n2916) );
  buffer buf_n387( .i (n386), .o (n387) );
  assign n5276 = ( n386 & ~n2707 ) | ( n386 & n4657 ) | ( ~n2707 & n4657 ) ;
  assign n5277 = ~n387 & n5276 ;
  assign n5278 = ~n3820 & n5277 ;
  assign n5279 = ( ~n4589 & n4750 ) | ( ~n4589 & n5278 ) | ( n4750 & n5278 ) ;
  assign n5280 = ~n4905 & n5279 ;
  assign n5281 = ~n5119 & n5280 ;
  assign n5282 = ~n4272 & n5281 ;
  buffer buf_n5283( .i (n5282), .o (n5283) );
  buffer buf_n5284( .i (n5283), .o (n5284) );
  buffer buf_n5285( .i (n5284), .o (n5285) );
  buffer buf_n5286( .i (n5285), .o (n5286) );
  buffer buf_n5287( .i (n5286), .o (n5287) );
  buffer buf_n5288( .i (n5287), .o (n5288) );
  assign n5289 = ( n383 & n1302 ) | ( n383 & ~n4044 ) | ( n1302 & ~n4044 ) ;
  assign n5290 = ~n384 & n5289 ;
  assign n5291 = ~n622 & n5290 ;
  assign n5292 = ( ~n730 & n4054 ) | ( ~n730 & n5291 ) | ( n4054 & n5291 ) ;
  buffer buf_n5293( .i (n4054), .o (n5293) );
  assign n5294 = n5292 & ~n5293 ;
  buffer buf_n5295( .i (n3573), .o (n5295) );
  assign n5296 = n5294 & ~n5295 ;
  assign n5297 = ( ~n4359 & n4589 ) | ( ~n4359 & n5296 ) | ( n4589 & n5296 ) ;
  buffer buf_n5298( .i (n4589), .o (n5298) );
  assign n5299 = n5297 & ~n5298 ;
  buffer buf_n5300( .i (n5299), .o (n5300) );
  buffer buf_n5301( .i (n5300), .o (n5301) );
  buffer buf_n5302( .i (n5301), .o (n5302) );
  buffer buf_n5303( .i (n5302), .o (n5303) );
  buffer buf_n5304( .i (n5303), .o (n5304) );
  buffer buf_n5305( .i (n5304), .o (n5305) );
  buffer buf_n5306( .i (n5305), .o (n5306) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  assign n5307 = n366 & ~n4749 ;
  assign n5308 = ( n389 & ~n2994 ) | ( n389 & n5307 ) | ( ~n2994 & n5307 ) ;
  assign n5309 = ~n390 & n5308 ;
  assign n5310 = ~n5119 & n5309 ;
  assign n5311 = ( ~n4272 & n4926 ) | ( ~n4272 & n5310 ) | ( n4926 & n5310 ) ;
  assign n5312 = ~n1823 & n5311 ;
  buffer buf_n5313( .i (n5312), .o (n5313) );
  buffer buf_n5314( .i (n5313), .o (n5314) );
  buffer buf_n5315( .i (n5314), .o (n5315) );
  buffer buf_n5316( .i (n5315), .o (n5316) );
  assign n5317 = n5306 | n5316 ;
  assign n5318 = ( ~n5047 & n5288 ) | ( ~n5047 & n5317 ) | ( n5288 & n5317 ) ;
  assign n5319 = n5048 | n5318 ;
  buffer buf_n5320( .i (n409), .o (n5320) );
  buffer buf_n5321( .i (n5320), .o (n5321) );
  assign n5322 = ( n200 & n3512 ) | ( n200 & n5321 ) | ( n3512 & n5321 ) ;
  assign n5323 = ~n201 & n5322 ;
  buffer buf_n5324( .i (n5323), .o (n5324) );
  buffer buf_n5325( .i (n5324), .o (n5325) );
  assign n5326 = ( n1818 & n4905 ) | ( n1818 & ~n5324 ) | ( n4905 & ~n5324 ) ;
  assign n5327 = n5325 & n5326 ;
  assign n5328 = ( n3624 & n4926 ) | ( n3624 & n5327 ) | ( n4926 & n5327 ) ;
  buffer buf_n5329( .i (n4926), .o (n5329) );
  assign n5330 = n5328 & ~n5329 ;
  buffer buf_n5331( .i (n5330), .o (n5331) );
  buffer buf_n5332( .i (n5331), .o (n5332) );
  buffer buf_n5333( .i (n5332), .o (n5333) );
  buffer buf_n5334( .i (n5333), .o (n5334) );
  buffer buf_n5335( .i (n5334), .o (n5335) );
  assign n5336 = ( ~n2760 & n5082 ) | ( ~n2760 & n5335 ) | ( n5082 & n5335 ) ;
  assign n5337 = n2761 | n5336 ;
  assign n5338 = n5319 | n5337 ;
  assign n5339 = ( n2916 & ~n2959 ) | ( n2916 & n5338 ) | ( ~n2959 & n5338 ) ;
  assign n5340 = n2960 | n5339 ;
  assign n5341 = n1998 | n3026 ;
  buffer buf_n5342( .i (n5341), .o (n5342) );
  buffer buf_n5343( .i (n5342), .o (n5343) );
  buffer buf_n5344( .i (n5343), .o (n5344) );
  assign n5345 = n1946 | n5126 ;
  assign n5346 = n1982 | n5345 ;
  assign n5347 = n1739 | n5111 ;
  assign n5348 = ( n2581 & ~n3895 ) | ( n2581 & n5347 ) | ( ~n3895 & n5347 ) ;
  assign n5349 = n3896 | n5348 ;
  assign n5350 = n1631 | n5349 ;
  assign n5351 = ( ~n1963 & n5107 ) | ( ~n1963 & n5350 ) | ( n5107 & n5350 ) ;
  assign n5352 = n1964 | n5351 ;
  assign n5353 = n5346 | n5352 ;
  assign n5354 = ( ~n1927 & n5344 ) | ( ~n1927 & n5353 ) | ( n5344 & n5353 ) ;
  assign n5355 = n1928 | n5354 ;
  buffer buf_n3937( .i (n3936), .o (n3937) );
  buffer buf_n3938( .i (n3937), .o (n3938) );
  buffer buf_n4090( .i (n4089), .o (n4090) );
  buffer buf_n4091( .i (n4090), .o (n4091) );
  assign n5356 = n409 & ~n4538 ;
  assign n5357 = ( n199 & n4585 ) | ( n199 & n5356 ) | ( n4585 & n5356 ) ;
  buffer buf_n5358( .i (n199), .o (n5358) );
  assign n5359 = n5357 & ~n5358 ;
  assign n5360 = n3977 & n5359 ;
  buffer buf_n5361( .i (n4749), .o (n5361) );
  buffer buf_n5362( .i (n3834), .o (n5362) );
  assign n5363 = ( n5360 & n5361 ) | ( n5360 & n5362 ) | ( n5361 & n5362 ) ;
  assign n5364 = ~n5298 & n5363 ;
  assign n5365 = n4564 & n5364 ;
  buffer buf_n5366( .i (n5365), .o (n5366) );
  buffer buf_n5367( .i (n5366), .o (n5367) );
  buffer buf_n5368( .i (n5367), .o (n5368) );
  buffer buf_n5369( .i (n5368), .o (n5369) );
  buffer buf_n5370( .i (n5369), .o (n5370) );
  buffer buf_n5371( .i (n5370), .o (n5371) );
  assign n5372 = ~n432 & n4539 ;
  assign n5373 = ( n251 & ~n3997 ) | ( n251 & n5372 ) | ( ~n3997 & n5372 ) ;
  assign n5374 = ~n252 & n5373 ;
  buffer buf_n5375( .i (n5374), .o (n5375) );
  buffer buf_n5376( .i (n5375), .o (n5376) );
  buffer buf_n5377( .i (n1817), .o (n5377) );
  assign n5378 = ( n4905 & ~n5375 ) | ( n4905 & n5377 ) | ( ~n5375 & n5377 ) ;
  assign n5379 = n5376 & n5378 ;
  assign n5380 = ( n3017 & n5120 ) | ( n3017 & n5379 ) | ( n5120 & n5379 ) ;
  assign n5381 = ~n5245 & n5380 ;
  buffer buf_n5382( .i (n5381), .o (n5382) );
  buffer buf_n5383( .i (n5382), .o (n5383) );
  buffer buf_n5384( .i (n5383), .o (n5384) );
  buffer buf_n5385( .i (n431), .o (n5385) );
  assign n5386 = ( n272 & n1216 ) | ( n272 & n5385 ) | ( n1216 & n5385 ) ;
  assign n5387 = ~n273 & n5386 ;
  buffer buf_n5388( .i (n5387), .o (n5388) );
  buffer buf_n5389( .i (n5388), .o (n5389) );
  assign n5390 = ( n1817 & n5361 ) | ( n1817 & ~n5388 ) | ( n5361 & ~n5388 ) ;
  assign n5391 = n5389 & n5390 ;
  buffer buf_n5392( .i (n4831), .o (n5392) );
  assign n5393 = ( n3016 & n5391 ) | ( n3016 & n5392 ) | ( n5391 & n5392 ) ;
  assign n5394 = ~n5120 & n5393 ;
  buffer buf_n5395( .i (n5394), .o (n5395) );
  buffer buf_n5396( .i (n5395), .o (n5396) );
  buffer buf_n5397( .i (n5396), .o (n5397) );
  assign n5398 = n2783 | n5397 ;
  assign n5399 = n5384 | n5398 ;
  assign n5400 = n5371 | n5399 ;
  assign n5401 = ( ~n2843 & n4091 ) | ( ~n2843 & n5400 ) | ( n4091 & n5400 ) ;
  assign n5402 = n2844 | n5401 ;
  buffer buf_n3245( .i (n3244), .o (n3245) );
  buffer buf_n3246( .i (n3245), .o (n3246) );
  assign n5403 = ~n431 & n3904 ;
  buffer buf_n5404( .i (n4655), .o (n5404) );
  buffer buf_n5405( .i (n5404), .o (n5405) );
  assign n5406 = ( n250 & n5403 ) | ( n250 & ~n5405 ) | ( n5403 & ~n5405 ) ;
  assign n5407 = ~n251 & n5406 ;
  buffer buf_n5408( .i (n5407), .o (n5408) );
  buffer buf_n5409( .i (n5408), .o (n5409) );
  assign n5410 = ( n3957 & n5361 ) | ( n3957 & ~n5408 ) | ( n5361 & ~n5408 ) ;
  assign n5411 = n5409 & n5410 ;
  buffer buf_n5412( .i (n5411), .o (n5412) );
  buffer buf_n5413( .i (n5412), .o (n5413) );
  buffer buf_n5414( .i (n5413), .o (n5414) );
  buffer buf_n5415( .i (n5414), .o (n5415) );
  buffer buf_n5416( .i (n5415), .o (n5416) );
  buffer buf_n5417( .i (n5416), .o (n5417) );
  buffer buf_n5418( .i (n5417), .o (n5418) );
  buffer buf_n5419( .i (n5418), .o (n5419) );
  buffer buf_n5420( .i (n430), .o (n5420) );
  assign n5421 = ~n5404 & n5420 ;
  assign n5422 = ( n272 & n4585 ) | ( n272 & n5421 ) | ( n4585 & n5421 ) ;
  assign n5423 = ~n273 & n5422 ;
  buffer buf_n5424( .i (n5423), .o (n5424) );
  buffer buf_n5425( .i (n5424), .o (n5425) );
  assign n5426 = ( n3957 & n5361 ) | ( n3957 & ~n5424 ) | ( n5361 & ~n5424 ) ;
  assign n5427 = n5425 & n5426 ;
  buffer buf_n5428( .i (n5427), .o (n5428) );
  buffer buf_n5429( .i (n5428), .o (n5429) );
  buffer buf_n5430( .i (n5429), .o (n5430) );
  buffer buf_n5431( .i (n5430), .o (n5431) );
  buffer buf_n5432( .i (n5431), .o (n5432) );
  buffer buf_n5433( .i (n5432), .o (n5433) );
  buffer buf_n5434( .i (n5433), .o (n5434) );
  assign n5435 = n2818 | n5434 ;
  assign n5436 = n5419 | n5435 ;
  assign n5437 = n3246 | n5436 ;
  assign n5438 = ( ~n3937 & n5402 ) | ( ~n3937 & n5437 ) | ( n5402 & n5437 ) ;
  assign n5439 = n3938 | n5438 ;
  assign n5440 = n5355 | n5439 ;
  assign n5441 = ( ~n5274 & n5340 ) | ( ~n5274 & n5440 ) | ( n5340 & n5440 ) ;
  assign n5442 = n5275 | n5441 ;
  buffer buf_n4497( .i (n4496), .o (n4497) );
  buffer buf_n4498( .i (n4497), .o (n4498) );
  buffer buf_n4481( .i (n4480), .o (n4481) );
  buffer buf_n4482( .i (n4481), .o (n4482) );
  assign n5443 = n4482 | n4895 ;
  assign n5444 = ( n3772 & ~n4497 ) | ( n3772 & n5443 ) | ( ~n4497 & n5443 ) ;
  assign n5445 = n4498 | n5444 ;
  buffer buf_n5446( .i (n5445), .o (n5446) );
  buffer buf_n5447( .i (n5446), .o (n5447) );
  assign n5448 = n1541 | n5095 ;
  assign n5449 = n3865 | n5448 ;
  assign n5450 = ( n912 & n2419 ) | ( n912 & n5070 ) | ( n2419 & n5070 ) ;
  assign n5451 = n2460 | n4244 ;
  assign n5452 = n5450 | n5451 ;
  assign n5453 = n3183 | n5452 ;
  assign n5454 = ( ~n1502 & n5449 ) | ( ~n1502 & n5453 ) | ( n5449 & n5453 ) ;
  assign n5455 = n1503 | n5454 ;
  buffer buf_n4485( .i (n4484), .o (n4485) );
  buffer buf_n4486( .i (n4485), .o (n4486) );
  buffer buf_n4487( .i (n4486), .o (n4487) );
  buffer buf_n5456( .i (n848), .o (n5456) );
  assign n5457 = n2416 & ~n5456 ;
  assign n5458 = ~n910 & n5457 ;
  assign n5459 = n2399 | n5458 ;
  assign n5460 = n4108 | n5459 ;
  assign n5461 = n4487 | n5460 ;
  assign n5462 = ( ~n3844 & n4102 ) | ( ~n3844 & n5461 ) | ( n4102 & n5461 ) ;
  assign n5463 = n3845 | n5462 ;
  assign n5464 = n1578 | n3039 ;
  assign n5465 = n1596 | n5464 ;
  buffer buf_n5177( .i (n5176), .o (n5177) );
  assign n5466 = n2520 | n4207 ;
  assign n5467 = n3668 | n5466 ;
  assign n5468 = n2492 | n5467 ;
  assign n5469 = ( ~n1523 & n3877 ) | ( ~n1523 & n5468 ) | ( n3877 & n5468 ) ;
  assign n5470 = n1524 | n5469 ;
  assign n5471 = n5177 | n5470 ;
  assign n5472 = ( ~n2550 & n5465 ) | ( ~n2550 & n5471 ) | ( n5465 & n5471 ) ;
  assign n5473 = n2551 | n5472 ;
  assign n5474 = n5463 | n5473 ;
  assign n5475 = ( ~n5446 & n5455 ) | ( ~n5446 & n5474 ) | ( n5455 & n5474 ) ;
  assign n5476 = n5447 | n5475 ;
  buffer buf_n5477( .i (n5476), .o (n5477) );
  buffer buf_n5478( .i (n5477), .o (n5478) );
  buffer buf_n5147( .i (n5146), .o (n5147) );
  buffer buf_n5148( .i (n5147), .o (n5148) );
  buffer buf_n5149( .i (n5148), .o (n5149) );
  buffer buf_n5150( .i (n5149), .o (n5150) );
  buffer buf_n5151( .i (n5150), .o (n5151) );
  buffer buf_n5152( .i (n5151), .o (n5152) );
  assign n5479 = n4160 | n5236 ;
  assign n5480 = ( n5107 & ~n5151 ) | ( n5107 & n5479 ) | ( ~n5151 & n5479 ) ;
  assign n5481 = n5152 | n5480 ;
  assign n5482 = n1960 | n5123 ;
  assign n5483 = n2316 | n5482 ;
  assign n5484 = n1941 | n4133 ;
  assign n5485 = ( ~n2334 & n3454 ) | ( ~n2334 & n5484 ) | ( n3454 & n5484 ) ;
  assign n5486 = n2335 | n5485 ;
  assign n5487 = n4144 | n5486 ;
  assign n5488 = ( ~n4065 & n5483 ) | ( ~n4065 & n5487 ) | ( n5483 & n5487 ) ;
  assign n5489 = n4066 | n5488 ;
  assign n5490 = n2659 | n2696 ;
  assign n5491 = n3521 | n5490 ;
  assign n5492 = n2359 | n5491 ;
  assign n5493 = ( ~n3629 & n3647 ) | ( ~n3629 & n5492 ) | ( n3647 & n5492 ) ;
  assign n5494 = n3630 | n5493 ;
  assign n5495 = n5489 | n5494 ;
  assign n5496 = n5481 | n5495 ;
  buffer buf_n5497( .i (n5496), .o (n5497) );
  buffer buf_n5498( .i (n5497), .o (n5498) );
  buffer buf_n2538( .i (n2537), .o (n2538) );
  buffer buf_n5168( .i (n5167), .o (n5168) );
  buffer buf_n5169( .i (n5168), .o (n5169) );
  assign n5499 = n2538 | n5169 ;
  assign n5500 = ( n2056 & ~n2294 ) | ( n2056 & n5499 ) | ( ~n2294 & n5499 ) ;
  assign n5501 = n2295 | n5500 ;
  assign n5502 = n3501 | n4669 ;
  assign n5503 = ( ~n3380 & n4760 ) | ( ~n3380 & n5502 ) | ( n4760 & n5502 ) ;
  assign n5504 = n3381 | n5503 ;
  assign n5505 = n1980 | n4420 ;
  assign n5506 = n5504 | n5505 ;
  assign n5507 = ( ~n2266 & n5342 ) | ( ~n2266 & n5506 ) | ( n5342 & n5506 ) ;
  assign n5508 = n2267 | n5507 ;
  assign n5509 = n2026 | n4639 ;
  assign n5510 = ( ~n1483 & n2560 ) | ( ~n1483 & n5509 ) | ( n2560 & n5509 ) ;
  assign n5511 = n1484 | n5510 ;
  assign n5512 = n5508 | n5511 ;
  assign n5513 = ( ~n5497 & n5501 ) | ( ~n5497 & n5512 ) | ( n5501 & n5512 ) ;
  assign n5514 = n5498 | n5513 ;
  assign n5515 = n1693 | n3225 ;
  assign n5516 = n3929 | n5515 ;
  assign n5517 = n3165 | n5516 ;
  assign n5518 = ( ~n1721 & n3236 ) | ( ~n1721 & n5517 ) | ( n3236 & n5517 ) ;
  assign n5519 = n1722 | n5518 ;
  buffer buf_n5520( .i (n5519), .o (n5520) );
  buffer buf_n5521( .i (n5520), .o (n5521) );
  assign n5522 = n3895 | n4275 ;
  assign n5523 = ( ~n1676 & n3726 ) | ( ~n1676 & n5522 ) | ( n3726 & n5522 ) ;
  assign n5524 = n1677 | n5523 ;
  assign n5525 = n1848 | n5428 ;
  assign n5526 = n2813 | n5525 ;
  assign n5527 = n4959 | n5526 ;
  assign n5528 = ( ~n4548 & n4945 ) | ( ~n4548 & n5527 ) | ( n4945 & n5527 ) ;
  assign n5529 = n4549 | n5528 ;
  assign n5530 = n3248 | n5412 ;
  assign n5531 = n5366 | n5530 ;
  assign n5532 = n4928 | n5531 ;
  assign n5533 = ( ~n4568 & n4910 ) | ( ~n4568 & n5532 ) | ( n4910 & n5532 ) ;
  assign n5534 = n4569 | n5533 ;
  assign n5535 = n5529 | n5534 ;
  assign n5536 = ( ~n5520 & n5524 ) | ( ~n5520 & n5535 ) | ( n5524 & n5535 ) ;
  assign n5537 = n5521 | n5536 ;
  buffer buf_n5538( .i (n5537), .o (n5538) );
  buffer buf_n5539( .i (n5538), .o (n5539) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  assign n5540 = n3549 | n3919 ;
  assign n5541 = n3343 | n5540 ;
  assign n5542 = n4011 | n5541 ;
  assign n5543 = ( ~n1744 & n2725 ) | ( ~n1744 & n5542 ) | ( n2725 & n5542 ) ;
  assign n5544 = n1745 | n5543 ;
  assign n5545 = n5113 | n5249 ;
  assign n5546 = n3536 | n4885 ;
  assign n5547 = ( ~n1629 & n2684 ) | ( ~n1629 & n5546 ) | ( n2684 & n5546 ) ;
  assign n5548 = n1630 | n5547 ;
  assign n5549 = n5545 | n5548 ;
  assign n5550 = ( ~n3950 & n4458 ) | ( ~n3950 & n5549 ) | ( n4458 & n5549 ) ;
  assign n5551 = n3951 | n5550 ;
  assign n5552 = n2583 | n4879 ;
  assign n5553 = ( ~n1407 & n4786 ) | ( ~n1407 & n5552 ) | ( n4786 & n5552 ) ;
  assign n5554 = n1408 | n5553 ;
  assign n5555 = n5551 | n5554 ;
  assign n5556 = ( ~n5538 & n5544 ) | ( ~n5538 & n5555 ) | ( n5544 & n5555 ) ;
  assign n5557 = n5539 | n5556 ;
  assign n5558 = n4435 | n4834 ;
  assign n5559 = n5395 | n5558 ;
  assign n5560 = ( ~n4852 & n5382 ) | ( ~n4852 & n5559 ) | ( n5382 & n5559 ) ;
  assign n5561 = n4853 | n5560 ;
  assign n5562 = n5208 | n5561 ;
  assign n5563 = ( ~n4261 & n4527 ) | ( ~n4261 & n5562 ) | ( n4527 & n5562 ) ;
  assign n5564 = n4262 | n5563 ;
  buffer buf_n5565( .i (n5564), .o (n5565) );
  buffer buf_n5566( .i (n5565), .o (n5566) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  assign n5567 = n1300 | n3140 ;
  assign n5568 = n1295 | n5567 ;
  assign n5569 = n1382 | n2924 ;
  assign n5570 = n2953 | n5569 ;
  buffer buf_n5571( .i (n2902), .o (n5571) );
  assign n5572 = n4978 | n5571 ;
  assign n5573 = n5570 | n5572 ;
  assign n5574 = n2943 | n5573 ;
  assign n5575 = ( ~n1246 & n5568 ) | ( ~n1246 & n5574 ) | ( n5568 & n5574 ) ;
  assign n5576 = n1247 | n5575 ;
  assign n5577 = n2857 | n4592 ;
  assign n5578 = n3126 | n5577 ;
  assign n5579 = n3110 | n5578 ;
  assign n5580 = ( n1443 & ~n2797 ) | ( n1443 & n5579 ) | ( ~n2797 & n5579 ) ;
  assign n5581 = n2798 | n5580 ;
  assign n5582 = n3072 | n5331 ;
  assign n5583 = n4863 | n5582 ;
  assign n5584 = n5581 | n5583 ;
  assign n5585 = ( ~n3065 & n5216 ) | ( ~n3065 & n5584 ) | ( n5216 & n5584 ) ;
  assign n5586 = n3066 | n5585 ;
  buffer buf_n3158( .i (n3157), .o (n3158) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  assign n5587 = n1777 | n4611 ;
  assign n5588 = n1887 | n5587 ;
  assign n5589 = n706 & n1395 ;
  buffer buf_n5590( .i (n5589), .o (n5590) );
  buffer buf_n5591( .i (n5590), .o (n5591) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  assign n5592 = ( n1666 & n4605 ) | ( n1666 & ~n5590 ) | ( n4605 & ~n5590 ) ;
  assign n5593 = n5591 & n5592 ;
  assign n5594 = n5300 | n5593 ;
  assign n5595 = n3564 | n5594 ;
  assign n5596 = n5283 | n5595 ;
  assign n5597 = ( ~n5043 & n5313 ) | ( ~n5043 & n5596 ) | ( n5313 & n5596 ) ;
  assign n5598 = n5044 | n5597 ;
  assign n5599 = n5196 | n5598 ;
  assign n5600 = ( ~n3157 & n5588 ) | ( ~n3157 & n5599 ) | ( n5588 & n5599 ) ;
  assign n5601 = n3158 | n5600 ;
  assign n5602 = n5586 | n5601 ;
  assign n5603 = ( ~n5565 & n5576 ) | ( ~n5565 & n5602 ) | ( n5576 & n5602 ) ;
  assign n5604 = n5566 | n5603 ;
  assign n5605 = n5557 | n5604 ;
  assign n5606 = ( ~n5477 & n5514 ) | ( ~n5477 & n5605 ) | ( n5514 & n5605 ) ;
  assign n5607 = n5478 | n5606 ;
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  assign n5608 = n4564 & n4665 ;
  assign n5609 = ( n482 & n1372 ) | ( n482 & n5608 ) | ( n1372 & n5608 ) ;
  assign n5610 = ~n483 & n5609 ;
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n5611( .i (n5293), .o (n5611) );
  assign n5612 = n5295 & ~n5611 ;
  buffer buf_n5613( .i (n5612), .o (n5613) );
  assign n5614 = ~n3926 & n5613 ;
  assign n5615 = n481 & n5614 ;
  buffer buf_n5616( .i (n4004), .o (n5616) );
  assign n5617 = ( n510 & n5615 ) | ( n510 & n5616 ) | ( n5615 & n5616 ) ;
  assign n5618 = ~n538 & n5617 ;
  assign n5619 = n5610 | n5618 ;
  buffer buf_n5620( .i (n5619), .o (n5620) );
  buffer buf_n5621( .i (n5620), .o (n5621) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  assign n5622 = n684 & n5620 ;
  assign n5623 = ( n603 & n5621 ) | ( n603 & n5622 ) | ( n5621 & n5622 ) ;
  buffer buf_n5624( .i (n5623), .o (n5624) );
  buffer buf_n5625( .i (n5624), .o (n5625) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  assign n5626 = n751 & ~n4044 ;
  buffer buf_n5627( .i (n5626), .o (n5627) );
  buffer buf_n5628( .i (n5627), .o (n5628) );
  assign n5633 = n335 & n810 ;
  assign n5634 = ( n703 & ~n5627 ) | ( n703 & n5633 ) | ( ~n5627 & n5633 ) ;
  assign n5635 = n5628 & n5634 ;
  buffer buf_n5636( .i (n5635), .o (n5636) );
  buffer buf_n5637( .i (n5636), .o (n5637) );
  buffer buf_n5638( .i (n5637), .o (n5638) );
  assign n5639 = ( n152 & n4952 ) | ( n152 & n5636 ) | ( n4952 & n5636 ) ;
  assign n5640 = n2994 & ~n5639 ;
  assign n5641 = ( n734 & n5638 ) | ( n734 & ~n5640 ) | ( n5638 & ~n5640 ) ;
  assign n5642 = n481 & ~n5641 ;
  buffer buf_n5629( .i (n5628), .o (n5629) );
  buffer buf_n5630( .i (n5629), .o (n5630) );
  buffer buf_n5631( .i (n5630), .o (n5631) );
  buffer buf_n5632( .i (n5631), .o (n5632) );
  buffer buf_n5643( .i (n151), .o (n5643) );
  assign n5644 = n4358 & ~n5643 ;
  assign n5645 = n129 & n5644 ;
  assign n5646 = n5632 & n5645 ;
  assign n5647 = n481 | n5646 ;
  assign n5648 = ~n5642 & n5647 ;
  assign n5649 = ~n5245 & n5648 ;
  buffer buf_n5650( .i (n591), .o (n5650) );
  buffer buf_n5651( .i (n2825), .o (n5651) );
  assign n5652 = n5650 & n5651 ;
  assign n5653 = ( n593 & ~n5358 ) | ( n593 & n5652 ) | ( ~n5358 & n5652 ) ;
  buffer buf_n5654( .i (n4540), .o (n5654) );
  assign n5655 = ~n5653 & n5654 ;
  assign n5656 = n624 & ~n3833 ;
  assign n5657 = n5654 | n5656 ;
  assign n5658 = ~n5655 & n5657 ;
  buffer buf_n5659( .i (n4359), .o (n5659) );
  assign n5660 = ( n480 & n5658 ) | ( n480 & ~n5659 ) | ( n5658 & ~n5659 ) ;
  buffer buf_n5661( .i (n730), .o (n5661) );
  assign n5662 = n177 | n5661 ;
  assign n5663 = ~n752 & n4655 ;
  buffer buf_n5664( .i (n5663), .o (n5664) );
  assign n5667 = n5405 & ~n5664 ;
  buffer buf_n5668( .i (n5667), .o (n5668) );
  assign n5669 = ~n5662 & n5668 ;
  buffer buf_n5665( .i (n5664), .o (n5665) );
  buffer buf_n5666( .i (n5665), .o (n5666) );
  buffer buf_n5670( .i (n704), .o (n5670) );
  buffer buf_n5671( .i (n5670), .o (n5671) );
  assign n5672 = ( ~n5666 & n5668 ) | ( ~n5666 & n5671 ) | ( n5668 & n5671 ) ;
  assign n5673 = ( ~n5362 & n5669 ) | ( ~n5362 & n5672 ) | ( n5669 & n5672 ) ;
  assign n5674 = ( n480 & n5659 ) | ( n480 & ~n5673 ) | ( n5659 & ~n5673 ) ;
  assign n5675 = n5660 & ~n5674 ;
  assign n5676 = n3636 & ~n5358 ;
  assign n5677 = ~n3820 & n5676 ;
  assign n5678 = n4938 & n5677 ;
  buffer buf_n5679( .i (n4953), .o (n5679) );
  assign n5680 = ( n5298 & n5678 ) | ( n5298 & n5679 ) | ( n5678 & n5679 ) ;
  assign n5681 = ~n4924 & n5680 ;
  assign n5682 = n5675 | n5681 ;
  assign n5683 = n5245 & n5682 ;
  assign n5684 = n5649 | n5683 ;
  assign n5685 = n540 & n5684 ;
  buffer buf_n484( .i (n483), .o (n484) );
  assign n5686 = ( ~n707 & n4188 ) | ( ~n707 & n5362 ) | ( n4188 & n5362 ) ;
  buffer buf_n5687( .i (n5686), .o (n5687) );
  assign n5688 = ( n4663 & n5392 ) | ( n4663 & ~n5687 ) | ( n5392 & ~n5687 ) ;
  assign n5689 = ( n4663 & ~n4924 ) | ( n4663 & n5687 ) | ( ~n4924 & n5687 ) ;
  assign n5690 = n5688 & ~n5689 ;
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  assign n5691 = ~n1221 & n4606 ;
  buffer buf_n5692( .i (n5691), .o (n5692) );
  assign n5693 = n5690 & n5692 ;
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n5694( .i (n5295), .o (n5694) );
  assign n5695 = ~n5362 & n5694 ;
  assign n5696 = ( n203 & ~n5659 ) | ( n203 & n5695 ) | ( ~n5659 & n5695 ) ;
  assign n5697 = ~n204 & n5696 ;
  buffer buf_n5698( .i (n3833), .o (n5698) );
  buffer buf_n5699( .i (n5698), .o (n5699) );
  assign n5700 = ( n129 & n3542 ) | ( n129 & n5699 ) | ( n3542 & n5699 ) ;
  assign n5701 = ~n130 & n5700 ;
  assign n5702 = ~n155 & n5701 ;
  assign n5703 = ( ~n156 & n5697 ) | ( ~n156 & n5702 ) | ( n5697 & n5702 ) ;
  assign n5704 = ( ~n1223 & n5692 ) | ( ~n1223 & n5703 ) | ( n5692 & n5703 ) ;
  assign n5705 = ( ~n484 & n5693 ) | ( ~n484 & n5704 ) | ( n5693 & n5704 ) ;
  assign n5706 = n540 | n5705 ;
  assign n5707 = ( ~n541 & n5685 ) | ( ~n541 & n5706 ) | ( n5685 & n5706 ) ;
  assign n5708 = n572 | n5707 ;
  buffer buf_n5709( .i (n198), .o (n5709) );
  assign n5710 = n5651 | n5709 ;
  assign n5711 = n5321 | n5710 ;
  buffer buf_n5712( .i (n5711), .o (n5712) );
  buffer buf_n5713( .i (n5712), .o (n5713) );
  assign n5716 = ( n594 & n3977 ) | ( n594 & n5698 ) | ( n3977 & n5698 ) ;
  assign n5717 = n5712 | n5716 ;
  assign n5718 = ( n5298 & ~n5713 ) | ( n5298 & n5717 ) | ( ~n5713 & n5717 ) ;
  assign n5719 = n4606 & ~n5718 ;
  buffer buf_n5720( .i (n5679), .o (n5720) );
  assign n5721 = n1799 | n5720 ;
  assign n5722 = ~n5719 & n5721 ;
  buffer buf_n5723( .i (n5722), .o (n5723) );
  buffer buf_n5724( .i (n5723), .o (n5724) );
  assign n5725 = ( n484 & ~n4704 ) | ( n484 & n5723 ) | ( ~n4704 & n5723 ) ;
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n5714( .i (n5713), .o (n5714) );
  buffer buf_n5715( .i (n5714), .o (n5715) );
  assign n5726 = ( n510 & n1668 ) | ( n510 & ~n5715 ) | ( n1668 & ~n5715 ) ;
  assign n5727 = ~n511 & n5726 ;
  assign n5728 = n4704 & n5727 ;
  assign n5729 = ( n5724 & ~n5725 ) | ( n5724 & n5728 ) | ( ~n5725 & n5728 ) ;
  assign n5730 = ~n792 & n5729 ;
  assign n5731 = n572 & ~n5730 ;
  assign n5732 = n5708 & ~n5731 ;
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  assign n5733 = ~n597 & n628 ;
  assign n5734 = n5295 | n5698 ;
  assign n5735 = n4359 & n5734 ;
  assign n5736 = ( n1397 & n5613 ) | ( n1397 & ~n5735 ) | ( n5613 & ~n5735 ) ;
  assign n5737 = ~n4004 & n5736 ;
  assign n5738 = ( n4859 & n5733 ) | ( n4859 & n5737 ) | ( n5733 & n5737 ) ;
  assign n5739 = ( n105 & n1223 ) | ( n105 & n5738 ) | ( n1223 & n5738 ) ;
  assign n5740 = ~n106 & n5739 ;
  assign n5741 = n1263 | n5740 ;
  assign n5742 = ( ~n1281 & n1317 ) | ( ~n1281 & n5741 ) | ( n1317 & n5741 ) ;
  assign n5743 = n1282 | n5742 ;
  buffer buf_n5744( .i (n5743), .o (n5744) );
  assign n5745 = ( ~n5624 & n5732 ) | ( ~n5624 & n5744 ) | ( n5732 & n5744 ) ;
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  assign n5746 = n78 & ~n5744 ;
  assign n5747 = ( n5625 & n5745 ) | ( n5625 & ~n5746 ) | ( n5745 & ~n5746 ) ;
  buffer buf_n5748( .i (n5747), .o (n5748) );
  buffer buf_n5749( .i (n5748), .o (n5749) );
  buffer buf_n5750( .i (n5749), .o (n5750) );
  buffer buf_n5751( .i (n5750), .o (n5751) );
  buffer buf_n5752( .i (n5751), .o (n5752) );
  assign n5753 = n3743 | n3865 ;
  assign n5754 = ( n2473 & ~n2527 ) | ( n2473 & n5753 ) | ( ~n2527 & n5753 ) ;
  assign n5755 = n2528 | n5754 ;
  buffer buf_n5756( .i (n5755), .o (n5756) );
  buffer buf_n5757( .i (n5756), .o (n5757) );
  buffer buf_n4448( .i (n4447), .o (n4448) );
  buffer buf_n4449( .i (n4448), .o (n4449) );
  buffer buf_n4450( .i (n4449), .o (n4450) );
  buffer buf_n4451( .i (n4450), .o (n4451) );
  assign n5758 = n2782 | n2815 ;
  buffer buf_n5759( .i (n2839), .o (n5759) );
  assign n5760 = ( ~n3167 & n5758 ) | ( ~n3167 & n5759 ) | ( n5758 & n5759 ) ;
  assign n5761 = n3168 | n5760 ;
  assign n5762 = n3934 | n5761 ;
  assign n5763 = ( n2585 & ~n3899 ) | ( n2585 & n5762 ) | ( ~n3899 & n5762 ) ;
  assign n5764 = n3900 | n5763 ;
  buffer buf_n4067( .i (n4066), .o (n4067) );
  assign n5765 = n2697 | n2733 ;
  assign n5766 = ( ~n2661 & n2685 ) | ( ~n2661 & n5765 ) | ( n2685 & n5765 ) ;
  assign n5767 = n2662 | n5766 ;
  assign n5768 = n4034 | n5767 ;
  assign n5769 = ( ~n2362 & n4067 ) | ( ~n2362 & n5768 ) | ( n4067 & n5768 ) ;
  assign n5770 = n2363 | n5769 ;
  assign n5771 = n5764 | n5770 ;
  assign n5772 = ( n4451 & ~n5756 ) | ( n4451 & n5771 ) | ( ~n5756 & n5771 ) ;
  assign n5773 = n5757 | n5772 ;
  buffer buf_n5774( .i (n5773), .o (n5774) );
  buffer buf_n5775( .i (n5774), .o (n5775) );
  buffer buf_n4013( .i (n4012), .o (n4013) );
  buffer buf_n4014( .i (n4013), .o (n4014) );
  buffer buf_n4068( .i (n4067), .o (n4068) );
  buffer buf_n3881( .i (n3880), .o (n3881) );
  assign n5776 = n4863 | n4911 ;
  assign n5777 = ( ~n3920 & n4931 ) | ( ~n3920 & n5776 ) | ( n4931 & n5776 ) ;
  assign n5778 = n3921 | n5777 ;
  assign n5779 = n3881 | n5778 ;
  assign n5780 = ( ~n4013 & n4068 ) | ( ~n4013 & n5779 ) | ( n4068 & n5779 ) ;
  assign n5781 = n4014 | n5780 ;
  buffer buf_n5782( .i (n5781), .o (n5782) );
  buffer buf_n5783( .i (n5782), .o (n5783) );
  buffer buf_n5784( .i (n5783), .o (n5784) );
  buffer buf_n5785( .i (n5784), .o (n5785) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n4717( .i (n4716), .o (n4717) );
  buffer buf_n4718( .i (n4717), .o (n4718) );
  buffer buf_n4719( .i (n4718), .o (n4719) );
  buffer buf_n4720( .i (n4719), .o (n4720) );
  buffer buf_n4721( .i (n4720), .o (n4721) );
  buffer buf_n4722( .i (n4721), .o (n4722) );
  assign y0 = n1327 ;
  assign y1 = n1337 ;
  assign y2 = 1'b0 ;
  assign y3 = n1349 ;
  assign y4 = n1360 ;
  assign y5 = n1460 ;
  assign y6 = n2062 ;
  assign y7 = n2072 ;
  assign y8 = n2087 ;
  assign y9 = n2097 ;
  assign y10 = n2974 ;
  assign y11 = n3178 ;
  assign y12 = n3353 ;
  assign y13 = n3682 ;
  assign y14 = n3751 ;
  assign y15 = n4100 ;
  assign y16 = n4228 ;
  assign y17 = n4320 ;
  assign y18 = n4387 ;
  assign y19 = n4477 ;
  assign y20 = n2273 ;
  assign y21 = n2300 ;
  assign y22 = n4733 ;
  assign y23 = n4743 ;
  assign y24 = n4186 ;
  assign y25 = n4797 ;
  assign y26 = n4810 ;
  assign y27 = n4822 ;
  assign y28 = n4971 ;
  assign y29 = n4996 ;
  assign y30 = n5006 ;
  assign y31 = n5015 ;
  assign y32 = n5054 ;
  assign y33 = n5063 ;
  assign y34 = n5134 ;
  assign y35 = n5262 ;
  assign y36 = n5442 ;
  assign y37 = n5607 ;
  assign y38 = n5752 ;
  assign y39 = n5775 ;
  assign y40 = n5785 ;
  assign y41 = n1836 ;
  assign y42 = 1'b0 ;
  assign y43 = n4722 ;
  assign y44 = n4186 ;
endmodule
