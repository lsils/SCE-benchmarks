module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 ;
  buffer buf_n4239( .i (x67), .o (n4239) );
  buffer buf_n4240( .i (n4239), .o (n4240) );
  buffer buf_n4241( .i (n4240), .o (n4241) );
  buffer buf_n4242( .i (n4241), .o (n4242) );
  buffer buf_n4243( .i (n4242), .o (n4243) );
  buffer buf_n4244( .i (n4243), .o (n4244) );
  buffer buf_n4245( .i (n4244), .o (n4245) );
  buffer buf_n4246( .i (n4245), .o (n4246) );
  buffer buf_n4247( .i (n4246), .o (n4247) );
  buffer buf_n4248( .i (n4247), .o (n4248) );
  buffer buf_n4249( .i (n4248), .o (n4249) );
  buffer buf_n4250( .i (n4249), .o (n4250) );
  buffer buf_n4251( .i (n4250), .o (n4251) );
  buffer buf_n4252( .i (n4251), .o (n4252) );
  buffer buf_n4253( .i (n4252), .o (n4253) );
  buffer buf_n4254( .i (n4253), .o (n4254) );
  buffer buf_n4255( .i (n4254), .o (n4255) );
  buffer buf_n4256( .i (n4255), .o (n4256) );
  buffer buf_n4257( .i (n4256), .o (n4257) );
  buffer buf_n4258( .i (n4257), .o (n4258) );
  buffer buf_n4259( .i (n4258), .o (n4259) );
  buffer buf_n4260( .i (n4259), .o (n4260) );
  buffer buf_n4261( .i (n4260), .o (n4261) );
  buffer buf_n4262( .i (n4261), .o (n4262) );
  buffer buf_n4263( .i (n4262), .o (n4263) );
  buffer buf_n4264( .i (n4263), .o (n4264) );
  buffer buf_n4265( .i (n4264), .o (n4265) );
  buffer buf_n4266( .i (n4265), .o (n4266) );
  buffer buf_n4267( .i (n4266), .o (n4267) );
  buffer buf_n4268( .i (n4267), .o (n4268) );
  buffer buf_n4269( .i (n4268), .o (n4269) );
  buffer buf_n4270( .i (n4269), .o (n4270) );
  buffer buf_n4271( .i (n4270), .o (n4271) );
  buffer buf_n4272( .i (n4271), .o (n4272) );
  buffer buf_n4273( .i (n4272), .o (n4273) );
  buffer buf_n4274( .i (n4273), .o (n4274) );
  buffer buf_n4275( .i (n4274), .o (n4275) );
  buffer buf_n4276( .i (n4275), .o (n4276) );
  buffer buf_n4277( .i (n4276), .o (n4277) );
  buffer buf_n4278( .i (n4277), .o (n4278) );
  buffer buf_n4279( .i (n4278), .o (n4279) );
  buffer buf_n4280( .i (n4279), .o (n4280) );
  buffer buf_n4281( .i (n4280), .o (n4281) );
  buffer buf_n4282( .i (n4281), .o (n4282) );
  buffer buf_n4283( .i (n4282), .o (n4283) );
  buffer buf_n4284( .i (n4283), .o (n4284) );
  buffer buf_n4285( .i (n4284), .o (n4285) );
  buffer buf_n4286( .i (n4285), .o (n4286) );
  buffer buf_n4287( .i (n4286), .o (n4287) );
  buffer buf_n4288( .i (n4287), .o (n4288) );
  buffer buf_n4289( .i (n4288), .o (n4289) );
  buffer buf_n4290( .i (n4289), .o (n4290) );
  buffer buf_n4291( .i (n4290), .o (n4291) );
  buffer buf_n4292( .i (n4291), .o (n4292) );
  buffer buf_n4293( .i (n4292), .o (n4293) );
  buffer buf_n4294( .i (n4293), .o (n4294) );
  buffer buf_n4295( .i (n4294), .o (n4295) );
  buffer buf_n4296( .i (n4295), .o (n4296) );
  buffer buf_n4297( .i (n4296), .o (n4297) );
  buffer buf_n4298( .i (n4297), .o (n4298) );
  buffer buf_n4299( .i (n4298), .o (n4299) );
  buffer buf_n4300( .i (n4299), .o (n4300) );
  buffer buf_n4301( .i (n4300), .o (n4301) );
  buffer buf_n4302( .i (n4301), .o (n4302) );
  buffer buf_n4303( .i (n4302), .o (n4303) );
  buffer buf_n4304( .i (n4303), .o (n4304) );
  buffer buf_n4305( .i (n4304), .o (n4305) );
  buffer buf_n4306( .i (n4305), .o (n4306) );
  buffer buf_n4307( .i (n4306), .o (n4307) );
  buffer buf_n4308( .i (n4307), .o (n4308) );
  buffer buf_n4309( .i (n4308), .o (n4309) );
  buffer buf_n4310( .i (n4309), .o (n4310) );
  buffer buf_n4311( .i (n4310), .o (n4311) );
  buffer buf_n4312( .i (n4311), .o (n4312) );
  buffer buf_n4313( .i (n4312), .o (n4313) );
  buffer buf_n4314( .i (n4313), .o (n4314) );
  buffer buf_n4315( .i (n4314), .o (n4315) );
  buffer buf_n4316( .i (n4315), .o (n4316) );
  buffer buf_n4317( .i (n4316), .o (n4317) );
  buffer buf_n4318( .i (n4317), .o (n4318) );
  buffer buf_n4319( .i (n4318), .o (n4319) );
  buffer buf_n4320( .i (n4319), .o (n4320) );
  buffer buf_n4321( .i (n4320), .o (n4321) );
  buffer buf_n4322( .i (n4321), .o (n4322) );
  buffer buf_n4323( .i (n4322), .o (n4323) );
  buffer buf_n4324( .i (n4323), .o (n4324) );
  buffer buf_n4325( .i (n4324), .o (n4325) );
  buffer buf_n4326( .i (n4325), .o (n4326) );
  buffer buf_n4327( .i (n4326), .o (n4327) );
  buffer buf_n4328( .i (n4327), .o (n4328) );
  buffer buf_n4329( .i (n4328), .o (n4329) );
  buffer buf_n4330( .i (n4329), .o (n4330) );
  buffer buf_n4331( .i (n4330), .o (n4331) );
  buffer buf_n4332( .i (n4331), .o (n4332) );
  buffer buf_n4333( .i (n4332), .o (n4333) );
  buffer buf_n4334( .i (n4333), .o (n4334) );
  buffer buf_n4335( .i (n4334), .o (n4335) );
  buffer buf_n4336( .i (n4335), .o (n4336) );
  buffer buf_n4337( .i (n4336), .o (n4337) );
  buffer buf_n4338( .i (n4337), .o (n4338) );
  buffer buf_n4339( .i (n4338), .o (n4339) );
  buffer buf_n4340( .i (n4339), .o (n4340) );
  buffer buf_n4341( .i (n4340), .o (n4341) );
  buffer buf_n4342( .i (n4341), .o (n4342) );
  buffer buf_n4343( .i (n4342), .o (n4343) );
  buffer buf_n4344( .i (n4343), .o (n4344) );
  buffer buf_n4345( .i (n4344), .o (n4345) );
  buffer buf_n4346( .i (n4345), .o (n4346) );
  buffer buf_n4347( .i (n4346), .o (n4347) );
  buffer buf_n4348( .i (n4347), .o (n4348) );
  buffer buf_n4349( .i (n4348), .o (n4349) );
  buffer buf_n4350( .i (n4349), .o (n4350) );
  buffer buf_n4351( .i (n4350), .o (n4351) );
  buffer buf_n365( .i (x8), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n3868( .i (x61), .o (n3868) );
  buffer buf_n3869( .i (n3868), .o (n3869) );
  buffer buf_n3870( .i (n3869), .o (n3870) );
  buffer buf_n3871( .i (n3870), .o (n3871) );
  buffer buf_n3872( .i (n3871), .o (n3872) );
  buffer buf_n3873( .i (n3872), .o (n3873) );
  buffer buf_n3874( .i (n3873), .o (n3874) );
  buffer buf_n3875( .i (n3874), .o (n3875) );
  buffer buf_n3876( .i (n3875), .o (n3876) );
  buffer buf_n3877( .i (n3876), .o (n3877) );
  buffer buf_n3878( .i (n3877), .o (n3878) );
  buffer buf_n3879( .i (n3878), .o (n3879) );
  buffer buf_n3880( .i (n3879), .o (n3880) );
  buffer buf_n3881( .i (n3880), .o (n3881) );
  buffer buf_n3882( .i (n3881), .o (n3882) );
  buffer buf_n3883( .i (n3882), .o (n3883) );
  buffer buf_n3884( .i (n3883), .o (n3884) );
  buffer buf_n3885( .i (n3884), .o (n3885) );
  buffer buf_n3886( .i (n3885), .o (n3886) );
  buffer buf_n3887( .i (n3886), .o (n3887) );
  buffer buf_n3888( .i (n3887), .o (n3888) );
  buffer buf_n3889( .i (n3888), .o (n3889) );
  buffer buf_n3890( .i (n3889), .o (n3890) );
  buffer buf_n3891( .i (n3890), .o (n3891) );
  buffer buf_n3892( .i (n3891), .o (n3892) );
  buffer buf_n3893( .i (n3892), .o (n3893) );
  buffer buf_n3894( .i (n3893), .o (n3894) );
  buffer buf_n3895( .i (n3894), .o (n3895) );
  buffer buf_n3896( .i (n3895), .o (n3896) );
  buffer buf_n3897( .i (n3896), .o (n3897) );
  buffer buf_n3898( .i (n3897), .o (n3898) );
  buffer buf_n3899( .i (n3898), .o (n3899) );
  buffer buf_n3900( .i (n3899), .o (n3900) );
  buffer buf_n3901( .i (n3900), .o (n3901) );
  buffer buf_n3902( .i (n3901), .o (n3902) );
  buffer buf_n3903( .i (n3902), .o (n3903) );
  buffer buf_n3904( .i (n3903), .o (n3904) );
  buffer buf_n3905( .i (n3904), .o (n3905) );
  buffer buf_n3906( .i (n3905), .o (n3906) );
  buffer buf_n3907( .i (n3906), .o (n3907) );
  buffer buf_n3908( .i (n3907), .o (n3908) );
  buffer buf_n3909( .i (n3908), .o (n3909) );
  buffer buf_n3910( .i (n3909), .o (n3910) );
  buffer buf_n3911( .i (n3910), .o (n3911) );
  buffer buf_n3912( .i (n3911), .o (n3912) );
  buffer buf_n2573( .i (x43), .o (n2573) );
  buffer buf_n2574( .i (n2573), .o (n2574) );
  buffer buf_n2575( .i (n2574), .o (n2575) );
  buffer buf_n2576( .i (n2575), .o (n2576) );
  buffer buf_n2577( .i (n2576), .o (n2577) );
  buffer buf_n2578( .i (n2577), .o (n2578) );
  buffer buf_n2579( .i (n2578), .o (n2579) );
  buffer buf_n2580( .i (n2579), .o (n2580) );
  buffer buf_n2581( .i (n2580), .o (n2581) );
  buffer buf_n2582( .i (n2581), .o (n2582) );
  buffer buf_n2583( .i (n2582), .o (n2583) );
  buffer buf_n2584( .i (n2583), .o (n2584) );
  buffer buf_n2585( .i (n2584), .o (n2585) );
  buffer buf_n2586( .i (n2585), .o (n2586) );
  buffer buf_n2587( .i (n2586), .o (n2587) );
  buffer buf_n2588( .i (n2587), .o (n2588) );
  buffer buf_n2589( .i (n2588), .o (n2589) );
  buffer buf_n2590( .i (n2589), .o (n2590) );
  buffer buf_n2591( .i (n2590), .o (n2591) );
  buffer buf_n2592( .i (n2591), .o (n2592) );
  buffer buf_n2593( .i (n2592), .o (n2593) );
  buffer buf_n2594( .i (n2593), .o (n2594) );
  buffer buf_n2595( .i (n2594), .o (n2595) );
  buffer buf_n2596( .i (n2595), .o (n2596) );
  buffer buf_n2597( .i (n2596), .o (n2597) );
  buffer buf_n2598( .i (n2597), .o (n2598) );
  buffer buf_n2599( .i (n2598), .o (n2599) );
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  buffer buf_n2602( .i (n2601), .o (n2602) );
  buffer buf_n2603( .i (n2602), .o (n2603) );
  buffer buf_n2604( .i (n2603), .o (n2604) );
  buffer buf_n2605( .i (n2604), .o (n2605) );
  buffer buf_n2606( .i (n2605), .o (n2606) );
  buffer buf_n2607( .i (n2606), .o (n2607) );
  buffer buf_n2608( .i (n2607), .o (n2608) );
  buffer buf_n2609( .i (n2608), .o (n2609) );
  buffer buf_n2610( .i (n2609), .o (n2610) );
  buffer buf_n2611( .i (n2610), .o (n2611) );
  buffer buf_n2612( .i (n2611), .o (n2612) );
  buffer buf_n2613( .i (n2612), .o (n2613) );
  buffer buf_n2614( .i (n2613), .o (n2614) );
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n3436( .i (x55), .o (n3436) );
  buffer buf_n3437( .i (n3436), .o (n3437) );
  buffer buf_n3438( .i (n3437), .o (n3438) );
  buffer buf_n3439( .i (n3438), .o (n3439) );
  buffer buf_n3440( .i (n3439), .o (n3440) );
  buffer buf_n3441( .i (n3440), .o (n3441) );
  buffer buf_n3442( .i (n3441), .o (n3442) );
  buffer buf_n3443( .i (n3442), .o (n3443) );
  buffer buf_n3444( .i (n3443), .o (n3444) );
  buffer buf_n3445( .i (n3444), .o (n3445) );
  buffer buf_n3446( .i (n3445), .o (n3446) );
  buffer buf_n3447( .i (n3446), .o (n3447) );
  buffer buf_n3448( .i (n3447), .o (n3448) );
  buffer buf_n3449( .i (n3448), .o (n3449) );
  buffer buf_n3450( .i (n3449), .o (n3450) );
  buffer buf_n3451( .i (n3450), .o (n3451) );
  buffer buf_n3452( .i (n3451), .o (n3452) );
  buffer buf_n3453( .i (n3452), .o (n3453) );
  buffer buf_n3454( .i (n3453), .o (n3454) );
  buffer buf_n3455( .i (n3454), .o (n3455) );
  buffer buf_n3456( .i (n3455), .o (n3456) );
  buffer buf_n3457( .i (n3456), .o (n3457) );
  buffer buf_n3458( .i (n3457), .o (n3458) );
  buffer buf_n3459( .i (n3458), .o (n3459) );
  buffer buf_n3460( .i (n3459), .o (n3460) );
  buffer buf_n3461( .i (n3460), .o (n3461) );
  buffer buf_n3462( .i (n3461), .o (n3462) );
  buffer buf_n3463( .i (n3462), .o (n3463) );
  buffer buf_n3464( .i (n3463), .o (n3464) );
  buffer buf_n3465( .i (n3464), .o (n3465) );
  buffer buf_n3466( .i (n3465), .o (n3466) );
  buffer buf_n3467( .i (n3466), .o (n3467) );
  buffer buf_n3468( .i (n3467), .o (n3468) );
  buffer buf_n3469( .i (n3468), .o (n3469) );
  buffer buf_n3470( .i (n3469), .o (n3470) );
  buffer buf_n3471( .i (n3470), .o (n3471) );
  buffer buf_n3472( .i (n3471), .o (n3472) );
  buffer buf_n3473( .i (n3472), .o (n3473) );
  buffer buf_n3474( .i (n3473), .o (n3474) );
  buffer buf_n3475( .i (n3474), .o (n3475) );
  buffer buf_n3476( .i (n3475), .o (n3476) );
  buffer buf_n2793( .i (x47), .o (n2793) );
  buffer buf_n2794( .i (n2793), .o (n2794) );
  buffer buf_n2795( .i (n2794), .o (n2795) );
  buffer buf_n2796( .i (n2795), .o (n2796) );
  buffer buf_n2797( .i (n2796), .o (n2797) );
  buffer buf_n2798( .i (n2797), .o (n2798) );
  buffer buf_n2799( .i (n2798), .o (n2799) );
  buffer buf_n2800( .i (n2799), .o (n2800) );
  buffer buf_n2801( .i (n2800), .o (n2801) );
  buffer buf_n2802( .i (n2801), .o (n2802) );
  buffer buf_n2803( .i (n2802), .o (n2803) );
  buffer buf_n2804( .i (n2803), .o (n2804) );
  buffer buf_n2805( .i (n2804), .o (n2805) );
  buffer buf_n2806( .i (n2805), .o (n2806) );
  buffer buf_n2807( .i (n2806), .o (n2807) );
  buffer buf_n2808( .i (n2807), .o (n2808) );
  buffer buf_n2809( .i (n2808), .o (n2809) );
  buffer buf_n2810( .i (n2809), .o (n2810) );
  buffer buf_n2811( .i (n2810), .o (n2811) );
  buffer buf_n2812( .i (n2811), .o (n2812) );
  buffer buf_n2813( .i (n2812), .o (n2813) );
  buffer buf_n2814( .i (n2813), .o (n2814) );
  buffer buf_n2815( .i (n2814), .o (n2815) );
  buffer buf_n2816( .i (n2815), .o (n2816) );
  buffer buf_n2817( .i (n2816), .o (n2817) );
  buffer buf_n2818( .i (n2817), .o (n2818) );
  buffer buf_n2819( .i (n2818), .o (n2819) );
  buffer buf_n2820( .i (n2819), .o (n2820) );
  buffer buf_n2821( .i (n2820), .o (n2821) );
  buffer buf_n2822( .i (n2821), .o (n2822) );
  buffer buf_n2823( .i (n2822), .o (n2823) );
  buffer buf_n2824( .i (n2823), .o (n2824) );
  buffer buf_n2825( .i (n2824), .o (n2825) );
  buffer buf_n2826( .i (n2825), .o (n2826) );
  buffer buf_n2827( .i (n2826), .o (n2827) );
  buffer buf_n2828( .i (n2827), .o (n2828) );
  buffer buf_n2829( .i (n2828), .o (n2829) );
  buffer buf_n2830( .i (n2829), .o (n2830) );
  buffer buf_n2831( .i (n2830), .o (n2831) );
  buffer buf_n1103( .i (x20), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n137( .i (x3), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n2198( .i (x37), .o (n2198) );
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n2200( .i (n2199), .o (n2200) );
  buffer buf_n2201( .i (n2200), .o (n2201) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  buffer buf_n2203( .i (n2202), .o (n2203) );
  buffer buf_n2204( .i (n2203), .o (n2204) );
  buffer buf_n2205( .i (n2204), .o (n2205) );
  buffer buf_n2206( .i (n2205), .o (n2206) );
  buffer buf_n2207( .i (n2206), .o (n2207) );
  buffer buf_n2208( .i (n2207), .o (n2208) );
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n2211( .i (n2210), .o (n2211) );
  buffer buf_n2212( .i (n2211), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  buffer buf_n2214( .i (n2213), .o (n2214) );
  buffer buf_n2215( .i (n2214), .o (n2215) );
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n2221( .i (n2220), .o (n2221) );
  buffer buf_n2222( .i (n2221), .o (n2222) );
  buffer buf_n2223( .i (n2222), .o (n2223) );
  buffer buf_n2224( .i (n2223), .o (n2224) );
  buffer buf_n2225( .i (n2224), .o (n2225) );
  buffer buf_n2226( .i (n2225), .o (n2226) );
  buffer buf_n2227( .i (n2226), .o (n2227) );
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  buffer buf_n413( .i (x9), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n2054( .i (x34), .o (n2054) );
  buffer buf_n2055( .i (n2054), .o (n2055) );
  buffer buf_n2056( .i (n2055), .o (n2056) );
  buffer buf_n2057( .i (n2056), .o (n2057) );
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  buffer buf_n2064( .i (n2063), .o (n2064) );
  buffer buf_n2065( .i (n2064), .o (n2065) );
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n2073( .i (n2072), .o (n2073) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n2075( .i (n2074), .o (n2075) );
  buffer buf_n2076( .i (n2075), .o (n2076) );
  buffer buf_n2077( .i (n2076), .o (n2077) );
  buffer buf_n2078( .i (n2077), .o (n2078) );
  buffer buf_n2079( .i (n2078), .o (n2079) );
  buffer buf_n2080( .i (n2079), .o (n2080) );
  buffer buf_n2081( .i (n2080), .o (n2081) );
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n326( .i (x7), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n3705( .i (x59), .o (n3705) );
  buffer buf_n3706( .i (n3705), .o (n3706) );
  buffer buf_n3707( .i (n3706), .o (n3707) );
  buffer buf_n3708( .i (n3707), .o (n3708) );
  buffer buf_n3709( .i (n3708), .o (n3709) );
  buffer buf_n3710( .i (n3709), .o (n3710) );
  buffer buf_n3711( .i (n3710), .o (n3711) );
  buffer buf_n3712( .i (n3711), .o (n3712) );
  buffer buf_n3713( .i (n3712), .o (n3713) );
  buffer buf_n3714( .i (n3713), .o (n3714) );
  buffer buf_n3715( .i (n3714), .o (n3715) );
  buffer buf_n3716( .i (n3715), .o (n3716) );
  buffer buf_n3717( .i (n3716), .o (n3717) );
  buffer buf_n3718( .i (n3717), .o (n3718) );
  buffer buf_n3719( .i (n3718), .o (n3719) );
  buffer buf_n3720( .i (n3719), .o (n3720) );
  buffer buf_n3721( .i (n3720), .o (n3721) );
  buffer buf_n3722( .i (n3721), .o (n3722) );
  buffer buf_n3723( .i (n3722), .o (n3723) );
  buffer buf_n3724( .i (n3723), .o (n3724) );
  buffer buf_n3725( .i (n3724), .o (n3725) );
  buffer buf_n3726( .i (n3725), .o (n3726) );
  buffer buf_n3727( .i (n3726), .o (n3727) );
  buffer buf_n3728( .i (n3727), .o (n3728) );
  buffer buf_n3729( .i (n3728), .o (n3729) );
  buffer buf_n3936( .i (x62), .o (n3936) );
  buffer buf_n3937( .i (n3936), .o (n3937) );
  buffer buf_n3938( .i (n3937), .o (n3938) );
  buffer buf_n3939( .i (n3938), .o (n3939) );
  buffer buf_n3940( .i (n3939), .o (n3940) );
  buffer buf_n3941( .i (n3940), .o (n3941) );
  buffer buf_n3942( .i (n3941), .o (n3942) );
  buffer buf_n3943( .i (n3942), .o (n3943) );
  buffer buf_n3944( .i (n3943), .o (n3944) );
  buffer buf_n3945( .i (n3944), .o (n3945) );
  buffer buf_n3946( .i (n3945), .o (n3946) );
  buffer buf_n3947( .i (n3946), .o (n3947) );
  buffer buf_n3948( .i (n3947), .o (n3948) );
  buffer buf_n3949( .i (n3948), .o (n3949) );
  buffer buf_n3950( .i (n3949), .o (n3950) );
  buffer buf_n3951( .i (n3950), .o (n3951) );
  buffer buf_n3952( .i (n3951), .o (n3952) );
  buffer buf_n3953( .i (n3952), .o (n3953) );
  buffer buf_n3954( .i (n3953), .o (n3954) );
  buffer buf_n3955( .i (n3954), .o (n3955) );
  buffer buf_n3956( .i (n3955), .o (n3956) );
  buffer buf_n3957( .i (n3956), .o (n3957) );
  buffer buf_n3958( .i (n3957), .o (n3958) );
  buffer buf_n1780( .i (x30), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n2418( .i (x40), .o (n2418) );
  buffer buf_n2419( .i (n2418), .o (n2419) );
  buffer buf_n2420( .i (n2419), .o (n2420) );
  buffer buf_n2421( .i (n2420), .o (n2421) );
  buffer buf_n2422( .i (n2421), .o (n2422) );
  buffer buf_n2423( .i (n2422), .o (n2423) );
  buffer buf_n2424( .i (n2423), .o (n2424) );
  buffer buf_n2425( .i (n2424), .o (n2425) );
  buffer buf_n2426( .i (n2425), .o (n2426) );
  buffer buf_n2427( .i (n2426), .o (n2427) );
  buffer buf_n2428( .i (n2427), .o (n2428) );
  buffer buf_n2429( .i (n2428), .o (n2429) );
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  buffer buf_n2432( .i (n2431), .o (n2432) );
  buffer buf_n2433( .i (n2432), .o (n2433) );
  buffer buf_n2434( .i (n2433), .o (n2434) );
  buffer buf_n2435( .i (n2434), .o (n2435) );
  buffer buf_n2436( .i (n2435), .o (n2436) );
  buffer buf_n3480( .i (x56), .o (n3480) );
  buffer buf_n3481( .i (n3480), .o (n3481) );
  buffer buf_n3482( .i (n3481), .o (n3482) );
  buffer buf_n3483( .i (n3482), .o (n3483) );
  buffer buf_n3484( .i (n3483), .o (n3484) );
  buffer buf_n3485( .i (n3484), .o (n3485) );
  buffer buf_n3486( .i (n3485), .o (n3486) );
  buffer buf_n3487( .i (n3486), .o (n3487) );
  buffer buf_n3488( .i (n3487), .o (n3488) );
  buffer buf_n3489( .i (n3488), .o (n3489) );
  buffer buf_n3490( .i (n3489), .o (n3490) );
  buffer buf_n3491( .i (n3490), .o (n3491) );
  buffer buf_n3492( .i (n3491), .o (n3492) );
  buffer buf_n3493( .i (n3492), .o (n3493) );
  buffer buf_n3494( .i (n3493), .o (n3494) );
  buffer buf_n3495( .i (n3494), .o (n3495) );
  buffer buf_n3496( .i (n3495), .o (n3496) );
  buffer buf_n1743( .i (x29), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n2619( .i (x44), .o (n2619) );
  buffer buf_n2620( .i (n2619), .o (n2620) );
  buffer buf_n2621( .i (n2620), .o (n2621) );
  buffer buf_n2622( .i (n2621), .o (n2622) );
  buffer buf_n2623( .i (n2622), .o (n2623) );
  buffer buf_n2624( .i (n2623), .o (n2624) );
  buffer buf_n2625( .i (n2624), .o (n2625) );
  buffer buf_n2626( .i (n2625), .o (n2626) );
  buffer buf_n2627( .i (n2626), .o (n2627) );
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  buffer buf_n2631( .i (n2630), .o (n2631) );
  buffer buf_n85( .i (x2), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n1818( .i (x31), .o (n1818) );
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  buffer buf_n1821( .i (n1820), .o (n1821) );
  buffer buf_n1822( .i (n1821), .o (n1822) );
  buffer buf_n1823( .i (n1822), .o (n1823) );
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1825( .i (n1824), .o (n1825) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n3519( .i (x57), .o (n3519) );
  buffer buf_n3520( .i (n3519), .o (n3520) );
  buffer buf_n3521( .i (n3520), .o (n3521) );
  buffer buf_n3522( .i (n3521), .o (n3522) );
  buffer buf_n3523( .i (n3522), .o (n3523) );
  buffer buf_n3524( .i (n3523), .o (n3524) );
  buffer buf_n3525( .i (n3524), .o (n3525) );
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n2531( .i (x42), .o (n2531) );
  assign n4352 = n2 | n2531 ;
  buffer buf_n4353( .i (n4352), .o (n4353) );
  buffer buf_n4354( .i (n4353), .o (n4354) );
  buffer buf_n4355( .i (n4354), .o (n4355) );
  buffer buf_n4356( .i (n4355), .o (n4356) );
  buffer buf_n4357( .i (n4356), .o (n4357) );
  assign n4393 = n3525 | n4357 ;
  buffer buf_n4394( .i (n4393), .o (n4394) );
  assign n4421 = n1826 | n4394 ;
  buffer buf_n4422( .i (n4421), .o (n4422) );
  assign n4448 = n95 | n4422 ;
  buffer buf_n4449( .i (n4448), .o (n4449) );
  assign n4473 = n2631 | n4449 ;
  buffer buf_n4474( .i (n4473), .o (n4474) );
  assign n4476 = n1757 | n4474 ;
  buffer buf_n4477( .i (n4476), .o (n4477) );
  assign n4479 = n3496 | n4477 ;
  buffer buf_n4480( .i (n4479), .o (n4480) );
  assign n4482 = n2436 | n4480 ;
  buffer buf_n4483( .i (n4482), .o (n4483) );
  assign n4485 = n1800 | n4483 ;
  buffer buf_n4486( .i (n4485), .o (n4486) );
  assign n4488 = n3958 | n4486 ;
  buffer buf_n4489( .i (n4488), .o (n4489) );
  assign n4491 = n3729 | n4489 ;
  buffer buf_n4492( .i (n4491), .o (n4492) );
  assign n4494 = n352 | n4492 ;
  buffer buf_n4495( .i (n4494), .o (n4495) );
  assign n4497 = n2082 | n4495 ;
  buffer buf_n4498( .i (n4497), .o (n4498) );
  assign n4500 = n443 | n4498 ;
  buffer buf_n4501( .i (n4500), .o (n4501) );
  assign n4503 = n2230 | n4501 ;
  buffer buf_n4504( .i (n4503), .o (n4504) );
  assign n4506 = n171 | n4504 ;
  buffer buf_n4507( .i (n4506), .o (n4507) );
  assign n4508 = n1139 | n4507 ;
  buffer buf_n4509( .i (n4508), .o (n4509) );
  assign n4510 = n2831 | n4509 ;
  buffer buf_n4511( .i (n4510), .o (n4511) );
  assign n4512 = n3476 | n4511 ;
  buffer buf_n4513( .i (n4512), .o (n4513) );
  assign n4514 = n2615 | n4513 ;
  buffer buf_n4515( .i (n4514), .o (n4515) );
  assign n4516 = n3912 & n4515 ;
  buffer buf_n4517( .i (n4516), .o (n4517) );
  assign n4518 = n411 & n4517 ;
  assign n4519 = n411 | n4517 ;
  assign n4520 = ~n4518 & n4519 ;
  buffer buf_n4521( .i (n4520), .o (n4521) );
  buffer buf_n4522( .i (n4521), .o (n4522) );
  buffer buf_n4523( .i (n4522), .o (n4523) );
  buffer buf_n4524( .i (n4523), .o (n4524) );
  buffer buf_n4525( .i (n4524), .o (n4525) );
  buffer buf_n4526( .i (n4525), .o (n4526) );
  buffer buf_n4527( .i (n4526), .o (n4527) );
  buffer buf_n4528( .i (n4527), .o (n4528) );
  buffer buf_n4529( .i (n4528), .o (n4529) );
  buffer buf_n4530( .i (n4529), .o (n4530) );
  buffer buf_n4531( .i (n4530), .o (n4531) );
  buffer buf_n4532( .i (n4531), .o (n4532) );
  buffer buf_n4533( .i (n4532), .o (n4533) );
  buffer buf_n4534( .i (n4533), .o (n4534) );
  buffer buf_n4535( .i (n4534), .o (n4535) );
  buffer buf_n4536( .i (n4535), .o (n4536) );
  buffer buf_n4537( .i (n4536), .o (n4537) );
  buffer buf_n4538( .i (n4537), .o (n4538) );
  buffer buf_n4539( .i (n4538), .o (n4539) );
  buffer buf_n4540( .i (n4539), .o (n4540) );
  buffer buf_n4541( .i (n4540), .o (n4541) );
  buffer buf_n4542( .i (n4541), .o (n4542) );
  buffer buf_n4543( .i (n4542), .o (n4543) );
  buffer buf_n4544( .i (n4543), .o (n4544) );
  buffer buf_n4545( .i (n4544), .o (n4545) );
  buffer buf_n4546( .i (n4545), .o (n4546) );
  buffer buf_n4547( .i (n4546), .o (n4547) );
  buffer buf_n4548( .i (n4547), .o (n4548) );
  buffer buf_n4549( .i (n4548), .o (n4549) );
  buffer buf_n4550( .i (n4549), .o (n4550) );
  buffer buf_n4551( .i (n4550), .o (n4551) );
  buffer buf_n4552( .i (n4551), .o (n4552) );
  buffer buf_n4553( .i (n4552), .o (n4553) );
  buffer buf_n4554( .i (n4553), .o (n4554) );
  buffer buf_n4555( .i (n4554), .o (n4555) );
  buffer buf_n4556( .i (n4555), .o (n4556) );
  buffer buf_n4557( .i (n4556), .o (n4557) );
  buffer buf_n4558( .i (n4557), .o (n4558) );
  buffer buf_n4559( .i (n4558), .o (n4559) );
  buffer buf_n4560( .i (n4559), .o (n4560) );
  buffer buf_n4561( .i (n4560), .o (n4561) );
  buffer buf_n4562( .i (n4561), .o (n4562) );
  buffer buf_n4563( .i (n4562), .o (n4563) );
  buffer buf_n4564( .i (n4563), .o (n4564) );
  buffer buf_n4565( .i (n4564), .o (n4565) );
  buffer buf_n4566( .i (n4565), .o (n4566) );
  buffer buf_n4567( .i (n4566), .o (n4567) );
  buffer buf_n4568( .i (n4567), .o (n4568) );
  buffer buf_n4569( .i (n4568), .o (n4569) );
  buffer buf_n4570( .i (n4569), .o (n4570) );
  buffer buf_n4571( .i (n4570), .o (n4571) );
  buffer buf_n4572( .i (n4571), .o (n4572) );
  buffer buf_n4573( .i (n4572), .o (n4573) );
  buffer buf_n4574( .i (n4573), .o (n4574) );
  buffer buf_n4575( .i (n4574), .o (n4575) );
  buffer buf_n4576( .i (n4575), .o (n4576) );
  buffer buf_n4577( .i (n4576), .o (n4577) );
  buffer buf_n4578( .i (n4577), .o (n4578) );
  buffer buf_n4579( .i (n4578), .o (n4579) );
  buffer buf_n4580( .i (n4579), .o (n4580) );
  buffer buf_n4581( .i (n4580), .o (n4581) );
  buffer buf_n1483( .i (x26), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n1488( .i (n1487), .o (n1488) );
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n1522( .i (n1521), .o (n1522) );
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  buffer buf_n1534( .i (n1533), .o (n1534) );
  buffer buf_n1535( .i (n1534), .o (n1535) );
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n1556( .i (n1555), .o (n1556) );
  buffer buf_n1557( .i (n1556), .o (n1557) );
  buffer buf_n1558( .i (n1557), .o (n1558) );
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  buffer buf_n2617( .i (n2616), .o (n2617) );
  assign n4584 = n3910 & n4513 ;
  buffer buf_n4585( .i (n4584), .o (n4585) );
  assign n4586 = ~n2617 & n4585 ;
  assign n4587 = n2617 & ~n4585 ;
  assign n4588 = n4586 | n4587 ;
  buffer buf_n4589( .i (n4588), .o (n4589) );
  buffer buf_n4590( .i (n4589), .o (n4590) );
  buffer buf_n4591( .i (n4590), .o (n4591) );
  buffer buf_n4592( .i (n4591), .o (n4592) );
  buffer buf_n4593( .i (n4592), .o (n4593) );
  buffer buf_n4594( .i (n4593), .o (n4594) );
  buffer buf_n4595( .i (n4594), .o (n4595) );
  buffer buf_n4596( .i (n4595), .o (n4596) );
  buffer buf_n4597( .i (n4596), .o (n4597) );
  buffer buf_n4598( .i (n4597), .o (n4598) );
  buffer buf_n4599( .i (n4598), .o (n4599) );
  buffer buf_n4600( .i (n4599), .o (n4600) );
  buffer buf_n4601( .i (n4600), .o (n4601) );
  buffer buf_n4602( .i (n4601), .o (n4602) );
  buffer buf_n4603( .i (n4602), .o (n4603) );
  buffer buf_n4604( .i (n4603), .o (n4604) );
  buffer buf_n4605( .i (n4604), .o (n4605) );
  buffer buf_n4606( .i (n4605), .o (n4606) );
  buffer buf_n4607( .i (n4606), .o (n4607) );
  buffer buf_n4608( .i (n4607), .o (n4608) );
  buffer buf_n4609( .i (n4608), .o (n4609) );
  buffer buf_n4610( .i (n4609), .o (n4610) );
  buffer buf_n4611( .i (n4610), .o (n4611) );
  buffer buf_n4612( .i (n4611), .o (n4612) );
  buffer buf_n4613( .i (n4612), .o (n4613) );
  buffer buf_n4614( .i (n4613), .o (n4614) );
  buffer buf_n4615( .i (n4614), .o (n4615) );
  buffer buf_n4616( .i (n4615), .o (n4616) );
  buffer buf_n4617( .i (n4616), .o (n4617) );
  buffer buf_n4618( .i (n4617), .o (n4618) );
  buffer buf_n4619( .i (n4618), .o (n4619) );
  buffer buf_n4620( .i (n4619), .o (n4620) );
  buffer buf_n4621( .i (n4620), .o (n4621) );
  buffer buf_n4622( .i (n4621), .o (n4622) );
  buffer buf_n4623( .i (n4622), .o (n4623) );
  buffer buf_n4624( .i (n4623), .o (n4624) );
  buffer buf_n4625( .i (n4624), .o (n4625) );
  buffer buf_n4626( .i (n4625), .o (n4626) );
  buffer buf_n4627( .i (n4626), .o (n4627) );
  buffer buf_n4628( .i (n4627), .o (n4628) );
  buffer buf_n4629( .i (n4628), .o (n4629) );
  buffer buf_n4630( .i (n4629), .o (n4630) );
  buffer buf_n4631( .i (n4630), .o (n4631) );
  buffer buf_n4632( .i (n4631), .o (n4632) );
  buffer buf_n4633( .i (n4632), .o (n4633) );
  buffer buf_n4634( .i (n4633), .o (n4634) );
  buffer buf_n4635( .i (n4634), .o (n4635) );
  buffer buf_n4636( .i (n4635), .o (n4636) );
  buffer buf_n4637( .i (n4636), .o (n4637) );
  buffer buf_n4638( .i (n4637), .o (n4638) );
  buffer buf_n4639( .i (n4638), .o (n4639) );
  buffer buf_n4640( .i (n4639), .o (n4640) );
  buffer buf_n4641( .i (n4640), .o (n4641) );
  buffer buf_n4642( .i (n4641), .o (n4642) );
  buffer buf_n4643( .i (n4642), .o (n4643) );
  buffer buf_n4644( .i (n4643), .o (n4644) );
  buffer buf_n4645( .i (n4644), .o (n4645) );
  buffer buf_n4646( .i (n4645), .o (n4646) );
  buffer buf_n578( .i (x12), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n3477( .i (n3476), .o (n3477) );
  buffer buf_n3478( .i (n3477), .o (n3478) );
  assign n4649 = n3908 & n4511 ;
  buffer buf_n4650( .i (n4649), .o (n4650) );
  assign n4651 = n3478 & n4650 ;
  assign n4652 = n3478 | n4650 ;
  assign n4653 = ~n4651 & n4652 ;
  buffer buf_n4654( .i (n4653), .o (n4654) );
  buffer buf_n4655( .i (n4654), .o (n4655) );
  buffer buf_n4656( .i (n4655), .o (n4656) );
  buffer buf_n4657( .i (n4656), .o (n4657) );
  buffer buf_n4658( .i (n4657), .o (n4658) );
  buffer buf_n4659( .i (n4658), .o (n4659) );
  buffer buf_n4660( .i (n4659), .o (n4660) );
  buffer buf_n4661( .i (n4660), .o (n4661) );
  buffer buf_n4662( .i (n4661), .o (n4662) );
  buffer buf_n4663( .i (n4662), .o (n4663) );
  buffer buf_n4664( .i (n4663), .o (n4664) );
  buffer buf_n4665( .i (n4664), .o (n4665) );
  buffer buf_n4666( .i (n4665), .o (n4666) );
  buffer buf_n4667( .i (n4666), .o (n4667) );
  buffer buf_n4668( .i (n4667), .o (n4668) );
  buffer buf_n4669( .i (n4668), .o (n4669) );
  buffer buf_n4670( .i (n4669), .o (n4670) );
  buffer buf_n4671( .i (n4670), .o (n4671) );
  buffer buf_n4672( .i (n4671), .o (n4672) );
  buffer buf_n4673( .i (n4672), .o (n4673) );
  buffer buf_n4674( .i (n4673), .o (n4674) );
  buffer buf_n4675( .i (n4674), .o (n4675) );
  buffer buf_n4676( .i (n4675), .o (n4676) );
  buffer buf_n4677( .i (n4676), .o (n4677) );
  buffer buf_n4678( .i (n4677), .o (n4678) );
  buffer buf_n4679( .i (n4678), .o (n4679) );
  buffer buf_n4680( .i (n4679), .o (n4680) );
  buffer buf_n4681( .i (n4680), .o (n4681) );
  buffer buf_n4682( .i (n4681), .o (n4682) );
  buffer buf_n4683( .i (n4682), .o (n4683) );
  buffer buf_n4684( .i (n4683), .o (n4684) );
  buffer buf_n4685( .i (n4684), .o (n4685) );
  buffer buf_n4686( .i (n4685), .o (n4686) );
  buffer buf_n4687( .i (n4686), .o (n4687) );
  buffer buf_n4688( .i (n4687), .o (n4688) );
  buffer buf_n4689( .i (n4688), .o (n4689) );
  buffer buf_n4690( .i (n4689), .o (n4690) );
  buffer buf_n4691( .i (n4690), .o (n4691) );
  buffer buf_n4692( .i (n4691), .o (n4692) );
  buffer buf_n4693( .i (n4692), .o (n4693) );
  buffer buf_n4694( .i (n4693), .o (n4694) );
  buffer buf_n4695( .i (n4694), .o (n4695) );
  buffer buf_n4696( .i (n4695), .o (n4696) );
  buffer buf_n4697( .i (n4696), .o (n4697) );
  buffer buf_n4698( .i (n4697), .o (n4698) );
  buffer buf_n4699( .i (n4698), .o (n4699) );
  buffer buf_n4700( .i (n4699), .o (n4700) );
  buffer buf_n4701( .i (n4700), .o (n4701) );
  buffer buf_n4702( .i (n4701), .o (n4702) );
  buffer buf_n4703( .i (n4702), .o (n4703) );
  buffer buf_n4704( .i (n4703), .o (n4704) );
  buffer buf_n4705( .i (n4704), .o (n4705) );
  buffer buf_n4706( .i (n4705), .o (n4706) );
  buffer buf_n4707( .i (n4706), .o (n4707) );
  buffer buf_n4708( .i (n4707), .o (n4708) );
  buffer buf_n1644( .i (x28), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  buffer buf_n1658( .i (n1657), .o (n1658) );
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n758( .i (x15), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n489( .i (x11), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n2835( .i (x48), .o (n2835) );
  buffer buf_n2836( .i (n2835), .o (n2836) );
  buffer buf_n2837( .i (n2836), .o (n2837) );
  buffer buf_n2838( .i (n2837), .o (n2838) );
  buffer buf_n2839( .i (n2838), .o (n2839) );
  buffer buf_n2840( .i (n2839), .o (n2840) );
  buffer buf_n2841( .i (n2840), .o (n2841) );
  buffer buf_n2842( .i (n2841), .o (n2842) );
  buffer buf_n2843( .i (n2842), .o (n2843) );
  buffer buf_n2844( .i (n2843), .o (n2844) );
  buffer buf_n2845( .i (n2844), .o (n2845) );
  buffer buf_n2846( .i (n2845), .o (n2846) );
  buffer buf_n2847( .i (n2846), .o (n2847) );
  buffer buf_n2848( .i (n2847), .o (n2848) );
  buffer buf_n2849( .i (n2848), .o (n2849) );
  buffer buf_n2850( .i (n2849), .o (n2850) );
  buffer buf_n2851( .i (n2850), .o (n2851) );
  buffer buf_n2852( .i (n2851), .o (n2852) );
  buffer buf_n2853( .i (n2852), .o (n2853) );
  buffer buf_n2854( .i (n2853), .o (n2854) );
  buffer buf_n2855( .i (n2854), .o (n2855) );
  buffer buf_n2856( .i (n2855), .o (n2856) );
  buffer buf_n2857( .i (n2856), .o (n2857) );
  buffer buf_n2858( .i (n2857), .o (n2858) );
  buffer buf_n2859( .i (n2858), .o (n2859) );
  buffer buf_n2860( .i (n2859), .o (n2860) );
  buffer buf_n2861( .i (n2860), .o (n2861) );
  buffer buf_n2862( .i (n2861), .o (n2862) );
  buffer buf_n2863( .i (n2862), .o (n2863) );
  buffer buf_n2864( .i (n2863), .o (n2864) );
  buffer buf_n2865( .i (n2864), .o (n2865) );
  buffer buf_n2866( .i (n2865), .o (n2866) );
  buffer buf_n2867( .i (n2866), .o (n2867) );
  buffer buf_n2868( .i (n2867), .o (n2868) );
  buffer buf_n2869( .i (n2868), .o (n2869) );
  buffer buf_n2870( .i (n2869), .o (n2870) );
  buffer buf_n2871( .i (n2870), .o (n2871) );
  buffer buf_n2872( .i (n2871), .o (n2872) );
  buffer buf_n2873( .i (n2872), .o (n2873) );
  buffer buf_n2874( .i (n2873), .o (n2874) );
  buffer buf_n2875( .i (n2874), .o (n2875) );
  buffer buf_n2876( .i (n2875), .o (n2876) );
  buffer buf_n2877( .i (n2876), .o (n2877) );
  buffer buf_n2878( .i (n2877), .o (n2878) );
  buffer buf_n2879( .i (n2878), .o (n2879) );
  buffer buf_n2880( .i (n2879), .o (n2880) );
  buffer buf_n2881( .i (n2880), .o (n2881) );
  buffer buf_n2882( .i (n2881), .o (n2882) );
  buffer buf_n2883( .i (n2882), .o (n2883) );
  buffer buf_n2884( .i (n2883), .o (n2884) );
  buffer buf_n2885( .i (n2884), .o (n2885) );
  buffer buf_n2886( .i (n2885), .o (n2886) );
  buffer buf_n2887( .i (n2886), .o (n2887) );
  buffer buf_n2888( .i (n2887), .o (n2888) );
  buffer buf_n2889( .i (n2888), .o (n2889) );
  buffer buf_n2890( .i (n2889), .o (n2890) );
  buffer buf_n2891( .i (n2890), .o (n2891) );
  buffer buf_n2892( .i (n2891), .o (n2892) );
  buffer buf_n2893( .i (n2892), .o (n2893) );
  buffer buf_n2894( .i (n2893), .o (n2894) );
  buffer buf_n2895( .i (n2894), .o (n2895) );
  buffer buf_n2896( .i (n2895), .o (n2896) );
  buffer buf_n2897( .i (n2896), .o (n2897) );
  buffer buf_n2898( .i (n2897), .o (n2898) );
  buffer buf_n2899( .i (n2898), .o (n2899) );
  buffer buf_n2900( .i (n2899), .o (n2900) );
  buffer buf_n2901( .i (n2900), .o (n2901) );
  buffer buf_n2902( .i (n2901), .o (n2902) );
  buffer buf_n2903( .i (n2902), .o (n2903) );
  buffer buf_n2904( .i (n2903), .o (n2904) );
  buffer buf_n2905( .i (n2904), .o (n2905) );
  buffer buf_n2906( .i (n2905), .o (n2906) );
  buffer buf_n2907( .i (n2906), .o (n2907) );
  buffer buf_n2908( .i (n2907), .o (n2908) );
  buffer buf_n2909( .i (n2908), .o (n2909) );
  buffer buf_n2910( .i (n2909), .o (n2910) );
  buffer buf_n2911( .i (n2910), .o (n2911) );
  buffer buf_n2912( .i (n2911), .o (n2912) );
  buffer buf_n2913( .i (n2912), .o (n2913) );
  buffer buf_n2914( .i (n2913), .o (n2914) );
  buffer buf_n2915( .i (n2914), .o (n2915) );
  buffer buf_n2916( .i (n2915), .o (n2916) );
  buffer buf_n2917( .i (n2916), .o (n2917) );
  buffer buf_n1312( .i (x23), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n4499( .i (n4498), .o (n4499) );
  assign n4711 = n3899 & n4499 ;
  buffer buf_n4712( .i (n4711), .o (n4712) );
  assign n4713 = ~n446 & n4712 ;
  assign n4714 = n446 & ~n4712 ;
  assign n4715 = n4713 | n4714 ;
  buffer buf_n4716( .i (n4715), .o (n4716) );
  buffer buf_n4717( .i (n4716), .o (n4717) );
  buffer buf_n4718( .i (n4717), .o (n4718) );
  buffer buf_n4719( .i (n4718), .o (n4719) );
  buffer buf_n4720( .i (n4719), .o (n4720) );
  buffer buf_n4721( .i (n4720), .o (n4721) );
  buffer buf_n4722( .i (n4721), .o (n4722) );
  buffer buf_n4723( .i (n4722), .o (n4723) );
  buffer buf_n4724( .i (n4723), .o (n4724) );
  buffer buf_n4725( .i (n4724), .o (n4725) );
  buffer buf_n4726( .i (n4725), .o (n4726) );
  buffer buf_n4727( .i (n4726), .o (n4727) );
  buffer buf_n4728( .i (n4727), .o (n4728) );
  buffer buf_n4729( .i (n4728), .o (n4729) );
  buffer buf_n4730( .i (n4729), .o (n4730) );
  buffer buf_n4731( .i (n4730), .o (n4731) );
  buffer buf_n4732( .i (n4731), .o (n4732) );
  buffer buf_n4733( .i (n4732), .o (n4733) );
  buffer buf_n4734( .i (n4733), .o (n4734) );
  buffer buf_n4735( .i (n4734), .o (n4735) );
  buffer buf_n4736( .i (n4735), .o (n4736) );
  buffer buf_n4737( .i (n4736), .o (n4737) );
  buffer buf_n4738( .i (n4737), .o (n4738) );
  buffer buf_n4739( .i (n4738), .o (n4739) );
  buffer buf_n4740( .i (n4739), .o (n4740) );
  buffer buf_n4741( .i (n4740), .o (n4741) );
  buffer buf_n4742( .i (n4741), .o (n4742) );
  buffer buf_n4743( .i (n4742), .o (n4743) );
  buffer buf_n4744( .i (n4743), .o (n4744) );
  buffer buf_n4745( .i (n4744), .o (n4745) );
  buffer buf_n4746( .i (n4745), .o (n4746) );
  buffer buf_n4747( .i (n4746), .o (n4747) );
  buffer buf_n4748( .i (n4747), .o (n4748) );
  buffer buf_n4749( .i (n4748), .o (n4749) );
  buffer buf_n4750( .i (n4749), .o (n4750) );
  buffer buf_n4751( .i (n4750), .o (n4751) );
  buffer buf_n4752( .i (n4751), .o (n4752) );
  buffer buf_n4753( .i (n4752), .o (n4753) );
  buffer buf_n4754( .i (n4753), .o (n4754) );
  buffer buf_n1029( .i (x19), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1867( .i (x32), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  buffer buf_n1872( .i (n1871), .o (n1872) );
  buffer buf_n1873( .i (n1872), .o (n1873) );
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  buffer buf_n1879( .i (n1878), .o (n1879) );
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n1888( .i (n1887), .o (n1888) );
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1907( .i (n1906), .o (n1907) );
  buffer buf_n1908( .i (n1907), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n1915( .i (n1914), .o (n1915) );
  buffer buf_n1916( .i (n1915), .o (n1916) );
  buffer buf_n1917( .i (n1916), .o (n1917) );
  buffer buf_n1918( .i (n1917), .o (n1918) );
  buffer buf_n1919( .i (n1918), .o (n1919) );
  buffer buf_n1920( .i (n1919), .o (n1920) );
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  buffer buf_n1930( .i (n1929), .o (n1930) );
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n2093( .i (x35), .o (n2093) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n2099( .i (n2098), .o (n2099) );
  buffer buf_n2100( .i (n2099), .o (n2100) );
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n2102( .i (n2101), .o (n2102) );
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n2111( .i (n2110), .o (n2111) );
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  buffer buf_n2119( .i (n2118), .o (n2119) );
  buffer buf_n2120( .i (n2119), .o (n2120) );
  buffer buf_n2121( .i (n2120), .o (n2121) );
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  buffer buf_n2129( .i (n2128), .o (n2129) );
  buffer buf_n2130( .i (n2129), .o (n2130) );
  buffer buf_n2131( .i (n2130), .o (n2131) );
  buffer buf_n2132( .i (n2131), .o (n2132) );
  buffer buf_n2133( .i (n2132), .o (n2133) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  buffer buf_n2137( .i (n2136), .o (n2137) );
  buffer buf_n2138( .i (n2137), .o (n2138) );
  buffer buf_n2139( .i (n2138), .o (n2139) );
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n2143( .i (n2142), .o (n2143) );
  buffer buf_n2144( .i (n2143), .o (n2144) );
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  buffer buf_n2152( .i (n2151), .o (n2152) );
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n176( .i (x4), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n3959( .i (n3958), .o (n3959) );
  buffer buf_n3960( .i (n3959), .o (n3960) );
  buffer buf_n3961( .i (n3960), .o (n3961) );
  buffer buf_n4487( .i (n4486), .o (n4487) );
  assign n4757 = n3891 & n4487 ;
  buffer buf_n4758( .i (n4757), .o (n4758) );
  assign n4759 = ~n3961 & n4758 ;
  assign n4760 = n3961 & ~n4758 ;
  assign n4761 = n4759 | n4760 ;
  buffer buf_n4762( .i (n4761), .o (n4762) );
  buffer buf_n4763( .i (n4762), .o (n4763) );
  buffer buf_n4764( .i (n4763), .o (n4764) );
  buffer buf_n4765( .i (n4764), .o (n4765) );
  buffer buf_n4766( .i (n4765), .o (n4766) );
  buffer buf_n4767( .i (n4766), .o (n4767) );
  buffer buf_n4768( .i (n4767), .o (n4768) );
  buffer buf_n4769( .i (n4768), .o (n4769) );
  buffer buf_n4770( .i (n4769), .o (n4770) );
  buffer buf_n4771( .i (n4770), .o (n4771) );
  buffer buf_n4772( .i (n4771), .o (n4772) );
  buffer buf_n4773( .i (n4772), .o (n4773) );
  buffer buf_n4774( .i (n4773), .o (n4774) );
  buffer buf_n4775( .i (n4774), .o (n4775) );
  buffer buf_n4776( .i (n4775), .o (n4776) );
  buffer buf_n4777( .i (n4776), .o (n4777) );
  buffer buf_n4778( .i (n4777), .o (n4778) );
  buffer buf_n4779( .i (n4778), .o (n4779) );
  buffer buf_n4780( .i (n4779), .o (n4780) );
  buffer buf_n4781( .i (n4780), .o (n4781) );
  buffer buf_n4782( .i (n4781), .o (n4782) );
  buffer buf_n4783( .i (n4782), .o (n4783) );
  buffer buf_n4784( .i (n4783), .o (n4784) );
  buffer buf_n4785( .i (n4784), .o (n4785) );
  buffer buf_n4786( .i (n4785), .o (n4786) );
  buffer buf_n4187( .i (x66), .o (n4187) );
  buffer buf_n4188( .i (n4187), .o (n4188) );
  buffer buf_n4189( .i (n4188), .o (n4189) );
  buffer buf_n4190( .i (n4189), .o (n4190) );
  buffer buf_n4191( .i (n4190), .o (n4191) );
  buffer buf_n4192( .i (n4191), .o (n4192) );
  buffer buf_n4193( .i (n4192), .o (n4193) );
  buffer buf_n4194( .i (n4193), .o (n4194) );
  buffer buf_n4195( .i (n4194), .o (n4195) );
  buffer buf_n4196( .i (n4195), .o (n4196) );
  buffer buf_n4197( .i (n4196), .o (n4197) );
  buffer buf_n4198( .i (n4197), .o (n4198) );
  buffer buf_n4199( .i (n4198), .o (n4199) );
  buffer buf_n4200( .i (n4199), .o (n4200) );
  buffer buf_n4201( .i (n4200), .o (n4201) );
  buffer buf_n4202( .i (n4201), .o (n4202) );
  buffer buf_n4203( .i (n4202), .o (n4203) );
  buffer buf_n4204( .i (n4203), .o (n4204) );
  buffer buf_n4205( .i (n4204), .o (n4205) );
  buffer buf_n4206( .i (n4205), .o (n4206) );
  buffer buf_n4207( .i (n4206), .o (n4207) );
  buffer buf_n4208( .i (n4207), .o (n4208) );
  buffer buf_n4209( .i (n4208), .o (n4209) );
  buffer buf_n4210( .i (n4209), .o (n4210) );
  buffer buf_n4211( .i (n4210), .o (n4211) );
  buffer buf_n4212( .i (n4211), .o (n4212) );
  buffer buf_n4213( .i (n4212), .o (n4213) );
  buffer buf_n4214( .i (n4213), .o (n4214) );
  buffer buf_n4215( .i (n4214), .o (n4215) );
  buffer buf_n4216( .i (n4215), .o (n4216) );
  buffer buf_n4217( .i (n4216), .o (n4217) );
  buffer buf_n4218( .i (n4217), .o (n4218) );
  buffer buf_n4219( .i (n4218), .o (n4219) );
  buffer buf_n4220( .i (n4219), .o (n4220) );
  buffer buf_n4221( .i (n4220), .o (n4221) );
  buffer buf_n4222( .i (n4221), .o (n4222) );
  buffer buf_n4223( .i (n4222), .o (n4223) );
  buffer buf_n4224( .i (n4223), .o (n4224) );
  buffer buf_n4225( .i (n4224), .o (n4225) );
  buffer buf_n4226( .i (n4225), .o (n4226) );
  buffer buf_n4227( .i (n4226), .o (n4227) );
  buffer buf_n4228( .i (n4227), .o (n4228) );
  buffer buf_n4229( .i (n4228), .o (n4229) );
  buffer buf_n4230( .i (n4229), .o (n4230) );
  buffer buf_n4231( .i (n4230), .o (n4231) );
  buffer buf_n4232( .i (n4231), .o (n4232) );
  buffer buf_n4233( .i (n4232), .o (n4233) );
  buffer buf_n4234( .i (n4233), .o (n4234) );
  buffer buf_n4235( .i (n4234), .o (n4235) );
  buffer buf_n4236( .i (n4235), .o (n4236) );
  buffer buf_n4237( .i (n4236), .o (n4237) );
  buffer buf_n3233( .i (x53), .o (n3233) );
  buffer buf_n3234( .i (n3233), .o (n3234) );
  buffer buf_n3235( .i (n3234), .o (n3235) );
  buffer buf_n3236( .i (n3235), .o (n3236) );
  buffer buf_n3237( .i (n3236), .o (n3237) );
  buffer buf_n3238( .i (n3237), .o (n3238) );
  buffer buf_n3239( .i (n3238), .o (n3239) );
  buffer buf_n3240( .i (n3239), .o (n3240) );
  buffer buf_n3241( .i (n3240), .o (n3241) );
  buffer buf_n3242( .i (n3241), .o (n3242) );
  buffer buf_n3243( .i (n3242), .o (n3243) );
  buffer buf_n3244( .i (n3243), .o (n3244) );
  buffer buf_n3245( .i (n3244), .o (n3245) );
  buffer buf_n3246( .i (n3245), .o (n3246) );
  buffer buf_n3247( .i (n3246), .o (n3247) );
  buffer buf_n3248( .i (n3247), .o (n3248) );
  buffer buf_n3249( .i (n3248), .o (n3249) );
  buffer buf_n3250( .i (n3249), .o (n3250) );
  buffer buf_n3251( .i (n3250), .o (n3251) );
  buffer buf_n3252( .i (n3251), .o (n3252) );
  buffer buf_n3253( .i (n3252), .o (n3253) );
  buffer buf_n3254( .i (n3253), .o (n3254) );
  buffer buf_n3255( .i (n3254), .o (n3255) );
  buffer buf_n3256( .i (n3255), .o (n3256) );
  buffer buf_n3257( .i (n3256), .o (n3257) );
  buffer buf_n3258( .i (n3257), .o (n3258) );
  buffer buf_n3259( .i (n3258), .o (n3259) );
  buffer buf_n3260( .i (n3259), .o (n3260) );
  buffer buf_n3261( .i (n3260), .o (n3261) );
  buffer buf_n3262( .i (n3261), .o (n3262) );
  buffer buf_n3263( .i (n3262), .o (n3263) );
  buffer buf_n3264( .i (n3263), .o (n3264) );
  buffer buf_n3265( .i (n3264), .o (n3265) );
  buffer buf_n3266( .i (n3265), .o (n3266) );
  buffer buf_n3267( .i (n3266), .o (n3267) );
  buffer buf_n3268( .i (n3267), .o (n3268) );
  buffer buf_n3269( .i (n3268), .o (n3269) );
  buffer buf_n3270( .i (n3269), .o (n3270) );
  buffer buf_n3271( .i (n3270), .o (n3271) );
  buffer buf_n3272( .i (n3271), .o (n3272) );
  buffer buf_n3273( .i (n3272), .o (n3273) );
  buffer buf_n3274( .i (n3273), .o (n3274) );
  buffer buf_n3275( .i (n3274), .o (n3275) );
  buffer buf_n3276( .i (n3275), .o (n3276) );
  buffer buf_n3277( .i (n3276), .o (n3277) );
  buffer buf_n3278( .i (n3277), .o (n3278) );
  buffer buf_n1441( .i (x25), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  buffer buf_n1455( .i (n1454), .o (n1455) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n47( .i (x1), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n682( .i (x13), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n720( .i (x14), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n4013( .i (x64), .o (n4013) );
  buffer buf_n4014( .i (n4013), .o (n4014) );
  buffer buf_n4015( .i (n4014), .o (n4015) );
  buffer buf_n4016( .i (n4015), .o (n4016) );
  buffer buf_n4017( .i (n4016), .o (n4017) );
  buffer buf_n4018( .i (n4017), .o (n4018) );
  buffer buf_n4019( .i (n4018), .o (n4019) );
  buffer buf_n4020( .i (n4019), .o (n4020) );
  buffer buf_n4021( .i (n4020), .o (n4021) );
  buffer buf_n4022( .i (n4021), .o (n4022) );
  buffer buf_n4023( .i (n4022), .o (n4023) );
  buffer buf_n4024( .i (n4023), .o (n4024) );
  buffer buf_n4025( .i (n4024), .o (n4025) );
  buffer buf_n4026( .i (n4025), .o (n4026) );
  buffer buf_n4027( .i (n4026), .o (n4027) );
  buffer buf_n4028( .i (n4027), .o (n4028) );
  buffer buf_n4029( .i (n4028), .o (n4029) );
  buffer buf_n4030( .i (n4029), .o (n4030) );
  buffer buf_n4031( .i (n4030), .o (n4031) );
  buffer buf_n4032( .i (n4031), .o (n4032) );
  buffer buf_n4033( .i (n4032), .o (n4033) );
  buffer buf_n450( .i (x10), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  assign n4789 = n3870 & n4353 ;
  buffer buf_n4790( .i (n4789), .o (n4790) );
  buffer buf_n4791( .i (n4790), .o (n4791) );
  assign n4792 = ~n3524 & n4791 ;
  assign n4793 = n3524 & ~n4791 ;
  assign n4794 = n4792 | n4793 ;
  buffer buf_n4795( .i (n4794), .o (n4795) );
  buffer buf_n4796( .i (n4795), .o (n4796) );
  buffer buf_n4797( .i (n4796), .o (n4797) );
  buffer buf_n4798( .i (n4797), .o (n4798) );
  buffer buf_n4799( .i (n4798), .o (n4799) );
  buffer buf_n1272( .i (x22), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n2919( .i (x49), .o (n2919) );
  buffer buf_n2920( .i (n2919), .o (n2920) );
  buffer buf_n2921( .i (n2920), .o (n2921) );
  buffer buf_n2922( .i (n2921), .o (n2922) );
  buffer buf_n2923( .i (n2922), .o (n2923) );
  buffer buf_n2924( .i (n2923), .o (n2924) );
  buffer buf_n2156( .i (x36), .o (n2156) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n2158( .i (n2157), .o (n2158) );
  buffer buf_n2159( .i (n2158), .o (n2159) );
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n2532), .o (n2533) );
  buffer buf_n2534( .i (n2533), .o (n2534) );
  assign n4802 = n2159 & n2534 ;
  buffer buf_n4803( .i (n4802), .o (n4803) );
  assign n4834 = n2924 | n4803 ;
  buffer buf_n4835( .i (n4834), .o (n4835) );
  buffer buf_n4836( .i (n4835), .o (n4836) );
  assign n4837 = n2924 & n4803 ;
  buffer buf_n4838( .i (n4837), .o (n4838) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  assign n4839 = n6 & ~n3872 ;
  assign n4840 = n5 & n2534 ;
  assign n4841 = n4790 & ~n4840 ;
  assign n4842 = n4839 | n4841 ;
  buffer buf_n4843( .i (n4842), .o (n4843) );
  assign n4846 = n4838 | n4843 ;
  assign n4847 = n4836 & n4846 ;
  buffer buf_n4848( .i (n4847), .o (n4848) );
  assign n4849 = n1282 & n4848 ;
  buffer buf_n4850( .i (n4849), .o (n4850) );
  assign n4851 = n4799 | n4850 ;
  assign n4852 = n1282 | n4848 ;
  buffer buf_n4853( .i (n4852), .o (n4853) );
  buffer buf_n4854( .i (n4853), .o (n4854) );
  assign n4855 = n4851 & n4854 ;
  buffer buf_n4856( .i (n4855), .o (n4856) );
  assign n4857 = n465 | n4856 ;
  buffer buf_n4858( .i (n4857), .o (n4858) );
  buffer buf_n4859( .i (n4858), .o (n4859) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n4395( .i (n4394), .o (n4395) );
  buffer buf_n4396( .i (n4395), .o (n4396) );
  buffer buf_n4397( .i (n4396), .o (n4397) );
  buffer buf_n4398( .i (n4397), .o (n4398) );
  assign n4860 = n3880 & n4398 ;
  buffer buf_n4861( .i (n4860), .o (n4861) );
  assign n4862 = n1832 | n4861 ;
  assign n4863 = n1832 & n4861 ;
  assign n4864 = n4862 & ~n4863 ;
  buffer buf_n4865( .i (n4864), .o (n4865) );
  assign n4868 = n465 & n4856 ;
  buffer buf_n4869( .i (n4868), .o (n4869) );
  assign n4870 = n4865 | n4869 ;
  assign n4871 = n4859 & n4870 ;
  buffer buf_n4872( .i (n4871), .o (n4872) );
  assign n4873 = n4033 | n4872 ;
  buffer buf_n4874( .i (n4873), .o (n4874) );
  buffer buf_n4875( .i (n4874), .o (n4875) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n4423( .i (n4422), .o (n4423) );
  buffer buf_n4424( .i (n4423), .o (n4424) );
  buffer buf_n4425( .i (n4424), .o (n4425) );
  buffer buf_n4426( .i (n4425), .o (n4426) );
  buffer buf_n4427( .i (n4426), .o (n4427) );
  buffer buf_n4428( .i (n4427), .o (n4428) );
  buffer buf_n4429( .i (n4428), .o (n4429) );
  assign n4876 = n3885 & n4429 ;
  buffer buf_n4877( .i (n4876), .o (n4877) );
  assign n4878 = ~n104 & n4877 ;
  assign n4879 = n104 & ~n4877 ;
  assign n4880 = n4878 | n4879 ;
  buffer buf_n4881( .i (n4880), .o (n4881) );
  assign n4884 = n4033 & n4872 ;
  buffer buf_n4885( .i (n4884), .o (n4885) );
  assign n4886 = n4881 | n4885 ;
  assign n4887 = n4875 & n4886 ;
  buffer buf_n4888( .i (n4887), .o (n4888) );
  assign n4889 = n745 & n4888 ;
  buffer buf_n4890( .i (n4889), .o (n4890) );
  buffer buf_n2632( .i (n2631), .o (n2632) );
  buffer buf_n2633( .i (n2632), .o (n2633) );
  buffer buf_n2634( .i (n2633), .o (n2634) );
  buffer buf_n2635( .i (n2634), .o (n2635) );
  buffer buf_n2636( .i (n2635), .o (n2636) );
  buffer buf_n2637( .i (n2636), .o (n2637) );
  buffer buf_n2638( .i (n2637), .o (n2638) );
  buffer buf_n2639( .i (n2638), .o (n2639) );
  buffer buf_n2640( .i (n2639), .o (n2640) );
  buffer buf_n2641( .i (n2640), .o (n2641) );
  buffer buf_n2642( .i (n2641), .o (n2642) );
  buffer buf_n2643( .i (n2642), .o (n2643) );
  buffer buf_n4450( .i (n4449), .o (n4450) );
  buffer buf_n4451( .i (n4450), .o (n4451) );
  buffer buf_n4452( .i (n4451), .o (n4452) );
  buffer buf_n4453( .i (n4452), .o (n4453) );
  buffer buf_n4454( .i (n4453), .o (n4454) );
  buffer buf_n4455( .i (n4454), .o (n4455) );
  buffer buf_n4456( .i (n4455), .o (n4456) );
  buffer buf_n4457( .i (n4456), .o (n4457) );
  buffer buf_n4458( .i (n4457), .o (n4458) );
  buffer buf_n4459( .i (n4458), .o (n4459) );
  assign n4891 = n3890 & n4459 ;
  buffer buf_n4892( .i (n4891), .o (n4892) );
  assign n4893 = n2643 & n4892 ;
  assign n4894 = n2643 | n4892 ;
  assign n4895 = ~n4893 & n4894 ;
  buffer buf_n4896( .i (n4895), .o (n4896) );
  assign n4899 = n4890 | n4896 ;
  assign n4900 = n745 | n4888 ;
  buffer buf_n4901( .i (n4900), .o (n4901) );
  buffer buf_n4902( .i (n4901), .o (n4902) );
  assign n4903 = n4899 & n4902 ;
  buffer buf_n4904( .i (n4903), .o (n4904) );
  assign n4905 = n712 & n4904 ;
  buffer buf_n4906( .i (n4905), .o (n4906) );
  buffer buf_n4907( .i (n4906), .o (n4907) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n4475( .i (n4474), .o (n4475) );
  assign n4908 = n3883 & n4475 ;
  buffer buf_n4909( .i (n4908), .o (n4909) );
  assign n4910 = ~n1760 & n4909 ;
  assign n4911 = n1760 & ~n4909 ;
  assign n4912 = n4910 | n4911 ;
  buffer buf_n4913( .i (n4912), .o (n4913) );
  buffer buf_n4914( .i (n4913), .o (n4914) );
  buffer buf_n4915( .i (n4914), .o (n4915) );
  buffer buf_n4916( .i (n4915), .o (n4916) );
  buffer buf_n4917( .i (n4916), .o (n4917) );
  buffer buf_n4918( .i (n4917), .o (n4918) );
  buffer buf_n4919( .i (n4918), .o (n4919) );
  buffer buf_n4920( .i (n4919), .o (n4920) );
  buffer buf_n4921( .i (n4920), .o (n4921) );
  buffer buf_n4922( .i (n4921), .o (n4922) );
  buffer buf_n4923( .i (n4922), .o (n4923) );
  buffer buf_n4924( .i (n4923), .o (n4924) );
  buffer buf_n4925( .i (n4924), .o (n4925) );
  assign n4928 = n712 | n4904 ;
  buffer buf_n4929( .i (n4928), .o (n4929) );
  assign n4930 = n4925 & n4929 ;
  assign n4931 = n4907 | n4930 ;
  buffer buf_n4932( .i (n4931), .o (n4932) );
  assign n4933 = n82 & n4932 ;
  buffer buf_n4934( .i (n4933), .o (n4934) );
  buffer buf_n3497( .i (n3496), .o (n3497) );
  buffer buf_n3498( .i (n3497), .o (n3498) );
  buffer buf_n3499( .i (n3498), .o (n3499) );
  buffer buf_n4478( .i (n4477), .o (n4478) );
  assign n4935 = n3885 & n4478 ;
  buffer buf_n4936( .i (n4935), .o (n4936) );
  assign n4937 = n3499 | n4936 ;
  assign n4938 = n3499 & n4936 ;
  assign n4939 = n4937 & ~n4938 ;
  buffer buf_n4940( .i (n4939), .o (n4940) );
  buffer buf_n4941( .i (n4940), .o (n4941) );
  buffer buf_n4942( .i (n4941), .o (n4942) );
  buffer buf_n4943( .i (n4942), .o (n4943) );
  buffer buf_n4944( .i (n4943), .o (n4944) );
  buffer buf_n4945( .i (n4944), .o (n4945) );
  buffer buf_n4946( .i (n4945), .o (n4946) );
  buffer buf_n4947( .i (n4946), .o (n4947) );
  buffer buf_n4948( .i (n4947), .o (n4948) );
  buffer buf_n4949( .i (n4948), .o (n4949) );
  buffer buf_n4950( .i (n4949), .o (n4950) );
  buffer buf_n4951( .i (n4950), .o (n4951) );
  buffer buf_n4952( .i (n4951), .o (n4952) );
  buffer buf_n4953( .i (n4952), .o (n4953) );
  buffer buf_n4954( .i (n4953), .o (n4954) );
  buffer buf_n4955( .i (n4954), .o (n4955) );
  assign n4958 = n4934 | n4955 ;
  assign n4959 = n82 | n4932 ;
  buffer buf_n4960( .i (n4959), .o (n4960) );
  buffer buf_n4961( .i (n4960), .o (n4961) );
  assign n4962 = n4958 & n4961 ;
  buffer buf_n4963( .i (n4962), .o (n4963) );
  assign n4964 = n1481 & n4963 ;
  buffer buf_n4965( .i (n4964), .o (n4965) );
  buffer buf_n2437( .i (n2436), .o (n2437) );
  buffer buf_n2438( .i (n2437), .o (n2438) );
  buffer buf_n2439( .i (n2438), .o (n2439) );
  buffer buf_n4481( .i (n4480), .o (n4481) );
  assign n4966 = n3887 & n4481 ;
  buffer buf_n4967( .i (n4966), .o (n4967) );
  assign n4968 = ~n2439 & n4967 ;
  assign n4969 = n2439 & ~n4967 ;
  assign n4970 = n4968 | n4969 ;
  buffer buf_n4971( .i (n4970), .o (n4971) );
  buffer buf_n4972( .i (n4971), .o (n4972) );
  buffer buf_n4973( .i (n4972), .o (n4973) );
  buffer buf_n4974( .i (n4973), .o (n4974) );
  buffer buf_n4975( .i (n4974), .o (n4975) );
  buffer buf_n4976( .i (n4975), .o (n4976) );
  buffer buf_n4977( .i (n4976), .o (n4977) );
  buffer buf_n4978( .i (n4977), .o (n4978) );
  buffer buf_n4979( .i (n4978), .o (n4979) );
  buffer buf_n4980( .i (n4979), .o (n4980) );
  buffer buf_n4981( .i (n4980), .o (n4981) );
  buffer buf_n4982( .i (n4981), .o (n4982) );
  buffer buf_n4983( .i (n4982), .o (n4983) );
  buffer buf_n4984( .i (n4983), .o (n4984) );
  buffer buf_n4985( .i (n4984), .o (n4985) );
  buffer buf_n4986( .i (n4985), .o (n4986) );
  buffer buf_n4987( .i (n4986), .o (n4987) );
  buffer buf_n4988( .i (n4987), .o (n4988) );
  buffer buf_n4989( .i (n4988), .o (n4989) );
  assign n4992 = n4965 | n4989 ;
  assign n4993 = n1481 | n4963 ;
  buffer buf_n4994( .i (n4993), .o (n4994) );
  buffer buf_n4995( .i (n4994), .o (n4995) );
  assign n4996 = n4992 & n4995 ;
  buffer buf_n4997( .i (n4996), .o (n4997) );
  assign n4998 = n3278 | n4997 ;
  buffer buf_n4999( .i (n4998), .o (n4999) );
  buffer buf_n5000( .i (n4999), .o (n5000) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n4484( .i (n4483), .o (n4484) );
  assign n5001 = n3889 & n4484 ;
  buffer buf_n5002( .i (n5001), .o (n5002) );
  assign n5003 = n1803 | n5002 ;
  assign n5004 = n1803 & n5002 ;
  assign n5005 = n5003 & ~n5004 ;
  buffer buf_n5006( .i (n5005), .o (n5006) );
  buffer buf_n5007( .i (n5006), .o (n5007) );
  buffer buf_n5008( .i (n5007), .o (n5008) );
  buffer buf_n5009( .i (n5008), .o (n5009) );
  buffer buf_n5010( .i (n5009), .o (n5010) );
  buffer buf_n5011( .i (n5010), .o (n5011) );
  buffer buf_n5012( .i (n5011), .o (n5012) );
  buffer buf_n5013( .i (n5012), .o (n5013) );
  buffer buf_n5014( .i (n5013), .o (n5014) );
  buffer buf_n5015( .i (n5014), .o (n5015) );
  buffer buf_n5016( .i (n5015), .o (n5016) );
  buffer buf_n5017( .i (n5016), .o (n5017) );
  buffer buf_n5018( .i (n5017), .o (n5018) );
  buffer buf_n5019( .i (n5018), .o (n5019) );
  buffer buf_n5020( .i (n5019), .o (n5020) );
  buffer buf_n5021( .i (n5020), .o (n5021) );
  buffer buf_n5022( .i (n5021), .o (n5022) );
  buffer buf_n5023( .i (n5022), .o (n5023) );
  buffer buf_n5024( .i (n5023), .o (n5024) );
  buffer buf_n5025( .i (n5024), .o (n5025) );
  buffer buf_n5026( .i (n5025), .o (n5026) );
  buffer buf_n5027( .i (n5026), .o (n5027) );
  assign n5030 = n3278 & n4997 ;
  buffer buf_n5031( .i (n5030), .o (n5031) );
  assign n5032 = n5027 | n5031 ;
  assign n5033 = n5000 & n5032 ;
  buffer buf_n5034( .i (n5033), .o (n5034) );
  assign n5035 = n4237 & n5034 ;
  buffer buf_n5036( .i (n5035), .o (n5036) );
  assign n5037 = n4786 | n5036 ;
  assign n5038 = n4237 | n5034 ;
  buffer buf_n5039( .i (n5038), .o (n5039) );
  buffer buf_n5040( .i (n5039), .o (n5040) );
  assign n5041 = n5037 & n5040 ;
  buffer buf_n5042( .i (n5041), .o (n5042) );
  assign n5043 = n231 & n5042 ;
  buffer buf_n5044( .i (n5043), .o (n5044) );
  buffer buf_n3730( .i (n3729), .o (n3730) );
  buffer buf_n3731( .i (n3730), .o (n3731) );
  buffer buf_n3732( .i (n3731), .o (n3732) );
  buffer buf_n4490( .i (n4489), .o (n4490) );
  assign n5046 = n3893 & n4490 ;
  buffer buf_n5047( .i (n5046), .o (n5047) );
  assign n5048 = n3732 & n5047 ;
  assign n5049 = n3732 | n5047 ;
  assign n5050 = ~n5048 & n5049 ;
  buffer buf_n5051( .i (n5050), .o (n5051) );
  buffer buf_n5052( .i (n5051), .o (n5052) );
  buffer buf_n5053( .i (n5052), .o (n5053) );
  buffer buf_n5054( .i (n5053), .o (n5054) );
  buffer buf_n5055( .i (n5054), .o (n5055) );
  buffer buf_n5056( .i (n5055), .o (n5056) );
  buffer buf_n5057( .i (n5056), .o (n5057) );
  buffer buf_n5058( .i (n5057), .o (n5058) );
  buffer buf_n5059( .i (n5058), .o (n5059) );
  buffer buf_n5060( .i (n5059), .o (n5060) );
  buffer buf_n5061( .i (n5060), .o (n5061) );
  buffer buf_n5062( .i (n5061), .o (n5062) );
  buffer buf_n5063( .i (n5062), .o (n5063) );
  buffer buf_n5064( .i (n5063), .o (n5064) );
  buffer buf_n5065( .i (n5064), .o (n5065) );
  buffer buf_n5066( .i (n5065), .o (n5066) );
  buffer buf_n5067( .i (n5066), .o (n5067) );
  buffer buf_n5068( .i (n5067), .o (n5068) );
  buffer buf_n5069( .i (n5068), .o (n5069) );
  buffer buf_n5070( .i (n5069), .o (n5070) );
  buffer buf_n5071( .i (n5070), .o (n5071) );
  buffer buf_n5072( .i (n5071), .o (n5072) );
  buffer buf_n5073( .i (n5072), .o (n5073) );
  buffer buf_n5074( .i (n5073), .o (n5074) );
  buffer buf_n5075( .i (n5074), .o (n5075) );
  buffer buf_n5076( .i (n5075), .o (n5076) );
  buffer buf_n5077( .i (n5076), .o (n5077) );
  buffer buf_n5078( .i (n5077), .o (n5078) );
  assign n5081 = n5044 | n5078 ;
  buffer buf_n5082( .i (n5081), .o (n5082) );
  assign n5083 = n231 | n5042 ;
  buffer buf_n5084( .i (n5083), .o (n5084) );
  buffer buf_n5085( .i (n5084), .o (n5085) );
  buffer buf_n5086( .i (n5085), .o (n5086) );
  assign n5087 = n5082 & n5086 ;
  buffer buf_n5088( .i (n5087), .o (n5088) );
  assign n5089 = n2154 & n5088 ;
  buffer buf_n5090( .i (n5089), .o (n5090) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n4493( .i (n4492), .o (n4493) );
  assign n5091 = n3895 & n4493 ;
  buffer buf_n5092( .i (n5091), .o (n5092) );
  assign n5093 = n355 & ~n5092 ;
  assign n5094 = ~n355 & n5092 ;
  assign n5095 = n5093 | n5094 ;
  buffer buf_n5096( .i (n5095), .o (n5096) );
  buffer buf_n5097( .i (n5096), .o (n5097) );
  buffer buf_n5098( .i (n5097), .o (n5098) );
  buffer buf_n5099( .i (n5098), .o (n5099) );
  buffer buf_n5100( .i (n5099), .o (n5100) );
  buffer buf_n5101( .i (n5100), .o (n5101) );
  buffer buf_n5102( .i (n5101), .o (n5102) );
  buffer buf_n5103( .i (n5102), .o (n5103) );
  buffer buf_n5104( .i (n5103), .o (n5104) );
  buffer buf_n5105( .i (n5104), .o (n5105) );
  buffer buf_n5106( .i (n5105), .o (n5106) );
  buffer buf_n5107( .i (n5106), .o (n5107) );
  buffer buf_n5108( .i (n5107), .o (n5108) );
  buffer buf_n5109( .i (n5108), .o (n5109) );
  buffer buf_n5110( .i (n5109), .o (n5110) );
  buffer buf_n5111( .i (n5110), .o (n5111) );
  buffer buf_n5112( .i (n5111), .o (n5112) );
  buffer buf_n5113( .i (n5112), .o (n5113) );
  buffer buf_n5114( .i (n5113), .o (n5114) );
  buffer buf_n5115( .i (n5114), .o (n5115) );
  buffer buf_n5116( .i (n5115), .o (n5116) );
  buffer buf_n5117( .i (n5116), .o (n5117) );
  buffer buf_n5118( .i (n5117), .o (n5118) );
  buffer buf_n5119( .i (n5118), .o (n5119) );
  buffer buf_n5120( .i (n5119), .o (n5120) );
  buffer buf_n5121( .i (n5120), .o (n5121) );
  buffer buf_n5122( .i (n5121), .o (n5122) );
  buffer buf_n5123( .i (n5122), .o (n5123) );
  buffer buf_n5124( .i (n5123), .o (n5124) );
  buffer buf_n5125( .i (n5124), .o (n5125) );
  buffer buf_n5126( .i (n5125), .o (n5126) );
  buffer buf_n5127( .i (n5126), .o (n5127) );
  assign n5130 = n5090 | n5127 ;
  assign n5131 = n2154 | n5088 ;
  buffer buf_n5132( .i (n5131), .o (n5132) );
  buffer buf_n5133( .i (n5132), .o (n5133) );
  assign n5134 = n5130 & n5133 ;
  buffer buf_n5135( .i (n5134), .o (n5135) );
  assign n5136 = n1933 | n5135 ;
  buffer buf_n5137( .i (n5136), .o (n5137) );
  buffer buf_n5138( .i (n5137), .o (n5138) );
  buffer buf_n5139( .i (n5138), .o (n5139) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n4496( .i (n4495), .o (n4496) );
  assign n5140 = n3897 & n4496 ;
  buffer buf_n5141( .i (n5140), .o (n5141) );
  assign n5142 = n2085 & n5141 ;
  assign n5143 = n2085 | n5141 ;
  assign n5144 = ~n5142 & n5143 ;
  buffer buf_n5145( .i (n5144), .o (n5145) );
  buffer buf_n5146( .i (n5145), .o (n5146) );
  buffer buf_n5147( .i (n5146), .o (n5147) );
  buffer buf_n5148( .i (n5147), .o (n5148) );
  buffer buf_n5149( .i (n5148), .o (n5149) );
  buffer buf_n5150( .i (n5149), .o (n5150) );
  buffer buf_n5151( .i (n5150), .o (n5151) );
  buffer buf_n5152( .i (n5151), .o (n5152) );
  buffer buf_n5153( .i (n5152), .o (n5153) );
  buffer buf_n5154( .i (n5153), .o (n5154) );
  buffer buf_n5155( .i (n5154), .o (n5155) );
  buffer buf_n5156( .i (n5155), .o (n5156) );
  buffer buf_n5157( .i (n5156), .o (n5157) );
  buffer buf_n5158( .i (n5157), .o (n5158) );
  buffer buf_n5159( .i (n5158), .o (n5159) );
  buffer buf_n5160( .i (n5159), .o (n5160) );
  buffer buf_n5161( .i (n5160), .o (n5161) );
  buffer buf_n5162( .i (n5161), .o (n5162) );
  buffer buf_n5163( .i (n5162), .o (n5163) );
  buffer buf_n5164( .i (n5163), .o (n5164) );
  buffer buf_n5165( .i (n5164), .o (n5165) );
  buffer buf_n5166( .i (n5165), .o (n5166) );
  buffer buf_n5167( .i (n5166), .o (n5167) );
  buffer buf_n5168( .i (n5167), .o (n5168) );
  buffer buf_n5169( .i (n5168), .o (n5169) );
  buffer buf_n5170( .i (n5169), .o (n5170) );
  buffer buf_n5171( .i (n5170), .o (n5171) );
  buffer buf_n5172( .i (n5171), .o (n5172) );
  buffer buf_n5173( .i (n5172), .o (n5173) );
  buffer buf_n5174( .i (n5173), .o (n5174) );
  buffer buf_n5175( .i (n5174), .o (n5175) );
  buffer buf_n5176( .i (n5175), .o (n5176) );
  buffer buf_n5177( .i (n5176), .o (n5177) );
  buffer buf_n5178( .i (n5177), .o (n5178) );
  buffer buf_n5179( .i (n5178), .o (n5179) );
  assign n5182 = n1933 & n5135 ;
  buffer buf_n5183( .i (n5182), .o (n5183) );
  assign n5185 = n5179 | n5183 ;
  buffer buf_n5186( .i (n5185), .o (n5186) );
  assign n5187 = n5139 & n5186 ;
  buffer buf_n5188( .i (n5187), .o (n5188) );
  assign n5189 = n1101 & n5188 ;
  buffer buf_n5190( .i (n5189), .o (n5190) );
  assign n5191 = n4754 | n5190 ;
  assign n5192 = n1101 | n5188 ;
  buffer buf_n5193( .i (n5192), .o (n5193) );
  buffer buf_n5194( .i (n5193), .o (n5194) );
  assign n5195 = n5191 & n5194 ;
  buffer buf_n5196( .i (n5195), .o (n5196) );
  assign n5197 = n1389 & n5196 ;
  buffer buf_n5198( .i (n5197), .o (n5198) );
  buffer buf_n2231( .i (n2230), .o (n2231) );
  buffer buf_n2232( .i (n2231), .o (n2232) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n4502( .i (n4501), .o (n4502) );
  assign n5199 = n3901 & n4502 ;
  buffer buf_n5200( .i (n5199), .o (n5200) );
  assign n5201 = n2233 & n5200 ;
  assign n5202 = n2233 | n5200 ;
  assign n5203 = ~n5201 & n5202 ;
  buffer buf_n5204( .i (n5203), .o (n5204) );
  buffer buf_n5205( .i (n5204), .o (n5205) );
  buffer buf_n5206( .i (n5205), .o (n5206) );
  buffer buf_n5207( .i (n5206), .o (n5207) );
  buffer buf_n5208( .i (n5207), .o (n5208) );
  buffer buf_n5209( .i (n5208), .o (n5209) );
  buffer buf_n5210( .i (n5209), .o (n5210) );
  buffer buf_n5211( .i (n5210), .o (n5211) );
  buffer buf_n5212( .i (n5211), .o (n5212) );
  buffer buf_n5213( .i (n5212), .o (n5213) );
  buffer buf_n5214( .i (n5213), .o (n5214) );
  buffer buf_n5215( .i (n5214), .o (n5215) );
  buffer buf_n5216( .i (n5215), .o (n5216) );
  buffer buf_n5217( .i (n5216), .o (n5217) );
  buffer buf_n5218( .i (n5217), .o (n5218) );
  buffer buf_n5219( .i (n5218), .o (n5219) );
  buffer buf_n5220( .i (n5219), .o (n5220) );
  buffer buf_n5221( .i (n5220), .o (n5221) );
  buffer buf_n5222( .i (n5221), .o (n5222) );
  buffer buf_n5223( .i (n5222), .o (n5223) );
  buffer buf_n5224( .i (n5223), .o (n5224) );
  buffer buf_n5225( .i (n5224), .o (n5225) );
  buffer buf_n5226( .i (n5225), .o (n5226) );
  buffer buf_n5227( .i (n5226), .o (n5227) );
  buffer buf_n5228( .i (n5227), .o (n5228) );
  buffer buf_n5229( .i (n5228), .o (n5229) );
  buffer buf_n5230( .i (n5229), .o (n5230) );
  buffer buf_n5231( .i (n5230), .o (n5231) );
  buffer buf_n5232( .i (n5231), .o (n5232) );
  buffer buf_n5233( .i (n5232), .o (n5233) );
  buffer buf_n5234( .i (n5233), .o (n5234) );
  buffer buf_n5235( .i (n5234), .o (n5235) );
  buffer buf_n5236( .i (n5235), .o (n5236) );
  buffer buf_n5237( .i (n5236), .o (n5237) );
  buffer buf_n5238( .i (n5237), .o (n5238) );
  buffer buf_n5239( .i (n5238), .o (n5239) );
  buffer buf_n5240( .i (n5239), .o (n5240) );
  buffer buf_n5241( .i (n5240), .o (n5241) );
  buffer buf_n5242( .i (n5241), .o (n5242) );
  buffer buf_n5243( .i (n5242), .o (n5243) );
  buffer buf_n5244( .i (n5243), .o (n5244) );
  buffer buf_n5245( .i (n5244), .o (n5245) );
  assign n5248 = n5198 | n5245 ;
  assign n5249 = n1389 | n5196 ;
  buffer buf_n5250( .i (n5249), .o (n5250) );
  buffer buf_n5251( .i (n5250), .o (n5251) );
  assign n5252 = n5248 & n5251 ;
  buffer buf_n5253( .i (n5252), .o (n5253) );
  assign n5254 = n2917 | n5253 ;
  buffer buf_n5255( .i (n5254), .o (n5255) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n4505( .i (n4504), .o (n4505) );
  assign n5256 = n3903 & n4505 ;
  buffer buf_n5257( .i (n5256), .o (n5257) );
  assign n5258 = n174 & ~n5257 ;
  assign n5259 = ~n174 & n5257 ;
  assign n5260 = n5258 | n5259 ;
  buffer buf_n5261( .i (n5260), .o (n5261) );
  buffer buf_n5262( .i (n5261), .o (n5262) );
  buffer buf_n5263( .i (n5262), .o (n5263) );
  buffer buf_n5264( .i (n5263), .o (n5264) );
  buffer buf_n5265( .i (n5264), .o (n5265) );
  buffer buf_n5266( .i (n5265), .o (n5266) );
  buffer buf_n5267( .i (n5266), .o (n5267) );
  buffer buf_n5268( .i (n5267), .o (n5268) );
  buffer buf_n5269( .i (n5268), .o (n5269) );
  buffer buf_n5270( .i (n5269), .o (n5270) );
  buffer buf_n5271( .i (n5270), .o (n5271) );
  buffer buf_n5272( .i (n5271), .o (n5272) );
  buffer buf_n5273( .i (n5272), .o (n5273) );
  buffer buf_n5274( .i (n5273), .o (n5274) );
  buffer buf_n5275( .i (n5274), .o (n5275) );
  buffer buf_n5276( .i (n5275), .o (n5276) );
  buffer buf_n5277( .i (n5276), .o (n5277) );
  buffer buf_n5278( .i (n5277), .o (n5278) );
  buffer buf_n5279( .i (n5278), .o (n5279) );
  buffer buf_n5280( .i (n5279), .o (n5280) );
  buffer buf_n5281( .i (n5280), .o (n5281) );
  buffer buf_n5282( .i (n5281), .o (n5282) );
  buffer buf_n5283( .i (n5282), .o (n5283) );
  buffer buf_n5284( .i (n5283), .o (n5284) );
  buffer buf_n5285( .i (n5284), .o (n5285) );
  buffer buf_n5286( .i (n5285), .o (n5286) );
  buffer buf_n5287( .i (n5286), .o (n5287) );
  buffer buf_n5288( .i (n5287), .o (n5288) );
  buffer buf_n5289( .i (n5288), .o (n5289) );
  buffer buf_n5290( .i (n5289), .o (n5290) );
  buffer buf_n5291( .i (n5290), .o (n5291) );
  buffer buf_n5292( .i (n5291), .o (n5292) );
  buffer buf_n5293( .i (n5292), .o (n5293) );
  buffer buf_n5294( .i (n5293), .o (n5294) );
  buffer buf_n5295( .i (n5294), .o (n5295) );
  buffer buf_n5296( .i (n5295), .o (n5296) );
  buffer buf_n5297( .i (n5296), .o (n5297) );
  buffer buf_n5298( .i (n5297), .o (n5298) );
  buffer buf_n5299( .i (n5298), .o (n5299) );
  buffer buf_n5300( .i (n5299), .o (n5300) );
  buffer buf_n5301( .i (n5300), .o (n5301) );
  buffer buf_n5302( .i (n5301), .o (n5302) );
  buffer buf_n5303( .i (n5302), .o (n5303) );
  buffer buf_n5304( .i (n5303), .o (n5304) );
  buffer buf_n5305( .i (n5304), .o (n5305) );
  assign n5308 = n5255 & n5305 ;
  assign n5309 = n2917 & n5253 ;
  buffer buf_n5310( .i (n5309), .o (n5310) );
  buffer buf_n5311( .i (n5310), .o (n5311) );
  assign n5312 = n5308 | n5311 ;
  buffer buf_n5313( .i (n5312), .o (n5313) );
  assign n5314 = n576 & n5313 ;
  buffer buf_n5315( .i (n5314), .o (n5315) );
  buffer buf_n5316( .i (n5315), .o (n5316) );
  assign n5317 = n576 | n5313 ;
  buffer buf_n5318( .i (n5317), .o (n5318) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  assign n5319 = n3904 & n4507 ;
  buffer buf_n5320( .i (n5319), .o (n5320) );
  assign n5321 = n1141 | n5320 ;
  assign n5322 = n1141 & n5320 ;
  assign n5323 = n5321 & ~n5322 ;
  buffer buf_n5324( .i (n5323), .o (n5324) );
  buffer buf_n5325( .i (n5324), .o (n5325) );
  buffer buf_n5326( .i (n5325), .o (n5326) );
  buffer buf_n5327( .i (n5326), .o (n5327) );
  buffer buf_n5328( .i (n5327), .o (n5328) );
  buffer buf_n5329( .i (n5328), .o (n5329) );
  buffer buf_n5330( .i (n5329), .o (n5330) );
  buffer buf_n5331( .i (n5330), .o (n5331) );
  buffer buf_n5332( .i (n5331), .o (n5332) );
  buffer buf_n5333( .i (n5332), .o (n5333) );
  buffer buf_n5334( .i (n5333), .o (n5334) );
  buffer buf_n5335( .i (n5334), .o (n5335) );
  buffer buf_n5336( .i (n5335), .o (n5336) );
  buffer buf_n5337( .i (n5336), .o (n5337) );
  buffer buf_n5338( .i (n5337), .o (n5338) );
  buffer buf_n5339( .i (n5338), .o (n5339) );
  buffer buf_n5340( .i (n5339), .o (n5340) );
  buffer buf_n5341( .i (n5340), .o (n5341) );
  buffer buf_n5342( .i (n5341), .o (n5342) );
  buffer buf_n5343( .i (n5342), .o (n5343) );
  buffer buf_n5344( .i (n5343), .o (n5344) );
  buffer buf_n5345( .i (n5344), .o (n5345) );
  buffer buf_n5346( .i (n5345), .o (n5346) );
  buffer buf_n5347( .i (n5346), .o (n5347) );
  buffer buf_n5348( .i (n5347), .o (n5348) );
  buffer buf_n5349( .i (n5348), .o (n5349) );
  buffer buf_n5350( .i (n5349), .o (n5350) );
  buffer buf_n5351( .i (n5350), .o (n5351) );
  buffer buf_n5352( .i (n5351), .o (n5352) );
  buffer buf_n5353( .i (n5352), .o (n5353) );
  buffer buf_n5354( .i (n5353), .o (n5354) );
  buffer buf_n5355( .i (n5354), .o (n5355) );
  buffer buf_n5356( .i (n5355), .o (n5356) );
  buffer buf_n5357( .i (n5356), .o (n5357) );
  buffer buf_n5358( .i (n5357), .o (n5358) );
  buffer buf_n5359( .i (n5358), .o (n5359) );
  buffer buf_n5360( .i (n5359), .o (n5360) );
  buffer buf_n5361( .i (n5360), .o (n5361) );
  buffer buf_n5362( .i (n5361), .o (n5362) );
  buffer buf_n5363( .i (n5362), .o (n5363) );
  buffer buf_n5364( .i (n5363), .o (n5364) );
  buffer buf_n5365( .i (n5364), .o (n5365) );
  buffer buf_n5366( .i (n5365), .o (n5366) );
  buffer buf_n5367( .i (n5366), .o (n5367) );
  buffer buf_n5368( .i (n5367), .o (n5368) );
  buffer buf_n5369( .i (n5368), .o (n5369) );
  buffer buf_n5370( .i (n5369), .o (n5370) );
  buffer buf_n5371( .i (n5370), .o (n5371) );
  buffer buf_n5372( .i (n5371), .o (n5372) );
  assign n5375 = n5318 & n5372 ;
  assign n5376 = n5316 | n5375 ;
  buffer buf_n5377( .i (n5376), .o (n5377) );
  assign n5378 = n850 & n5377 ;
  buffer buf_n5379( .i (n5378), .o (n5379) );
  buffer buf_n5380( .i (n5379), .o (n5380) );
  assign n5381 = n850 | n5377 ;
  buffer buf_n5382( .i (n5381), .o (n5382) );
  buffer buf_n2832( .i (n2831), .o (n2832) );
  buffer buf_n2833( .i (n2832), .o (n2833) );
  assign n5383 = n3906 & n4509 ;
  buffer buf_n5384( .i (n5383), .o (n5384) );
  assign n5385 = n2833 & ~n5384 ;
  assign n5386 = ~n2833 & n5384 ;
  assign n5387 = n5385 | n5386 ;
  buffer buf_n5388( .i (n5387), .o (n5388) );
  buffer buf_n5389( .i (n5388), .o (n5389) );
  buffer buf_n5390( .i (n5389), .o (n5390) );
  buffer buf_n5391( .i (n5390), .o (n5391) );
  buffer buf_n5392( .i (n5391), .o (n5392) );
  buffer buf_n5393( .i (n5392), .o (n5393) );
  buffer buf_n5394( .i (n5393), .o (n5394) );
  buffer buf_n5395( .i (n5394), .o (n5395) );
  buffer buf_n5396( .i (n5395), .o (n5396) );
  buffer buf_n5397( .i (n5396), .o (n5397) );
  buffer buf_n5398( .i (n5397), .o (n5398) );
  buffer buf_n5399( .i (n5398), .o (n5399) );
  buffer buf_n5400( .i (n5399), .o (n5400) );
  buffer buf_n5401( .i (n5400), .o (n5401) );
  buffer buf_n5402( .i (n5401), .o (n5402) );
  buffer buf_n5403( .i (n5402), .o (n5403) );
  buffer buf_n5404( .i (n5403), .o (n5404) );
  buffer buf_n5405( .i (n5404), .o (n5405) );
  buffer buf_n5406( .i (n5405), .o (n5406) );
  buffer buf_n5407( .i (n5406), .o (n5407) );
  buffer buf_n5408( .i (n5407), .o (n5408) );
  buffer buf_n5409( .i (n5408), .o (n5409) );
  buffer buf_n5410( .i (n5409), .o (n5410) );
  buffer buf_n5411( .i (n5410), .o (n5411) );
  buffer buf_n5412( .i (n5411), .o (n5412) );
  buffer buf_n5413( .i (n5412), .o (n5413) );
  buffer buf_n5414( .i (n5413), .o (n5414) );
  buffer buf_n5415( .i (n5414), .o (n5415) );
  buffer buf_n5416( .i (n5415), .o (n5416) );
  buffer buf_n5417( .i (n5416), .o (n5417) );
  buffer buf_n5418( .i (n5417), .o (n5418) );
  buffer buf_n5419( .i (n5418), .o (n5419) );
  buffer buf_n5420( .i (n5419), .o (n5420) );
  buffer buf_n5421( .i (n5420), .o (n5421) );
  buffer buf_n5422( .i (n5421), .o (n5422) );
  buffer buf_n5423( .i (n5422), .o (n5423) );
  buffer buf_n5424( .i (n5423), .o (n5424) );
  buffer buf_n5425( .i (n5424), .o (n5425) );
  buffer buf_n5426( .i (n5425), .o (n5426) );
  buffer buf_n5427( .i (n5426), .o (n5427) );
  buffer buf_n5428( .i (n5427), .o (n5428) );
  buffer buf_n5429( .i (n5428), .o (n5429) );
  buffer buf_n5430( .i (n5429), .o (n5430) );
  buffer buf_n5431( .i (n5430), .o (n5431) );
  buffer buf_n5432( .i (n5431), .o (n5432) );
  buffer buf_n5433( .i (n5432), .o (n5433) );
  buffer buf_n5434( .i (n5433), .o (n5434) );
  buffer buf_n5435( .i (n5434), .o (n5435) );
  buffer buf_n5436( .i (n5435), .o (n5436) );
  buffer buf_n5437( .i (n5436), .o (n5437) );
  buffer buf_n5438( .i (n5437), .o (n5438) );
  buffer buf_n5439( .i (n5438), .o (n5439) );
  assign n5442 = n5382 & n5439 ;
  assign n5443 = n5380 | n5442 ;
  buffer buf_n5444( .i (n5443), .o (n5444) );
  assign n5445 = n1741 & n5444 ;
  buffer buf_n5446( .i (n5445), .o (n5446) );
  assign n5447 = n4708 | n5446 ;
  assign n5448 = n1741 | n5444 ;
  buffer buf_n5449( .i (n5448), .o (n5449) );
  buffer buf_n5450( .i (n5449), .o (n5450) );
  assign n5451 = n5447 & n5450 ;
  buffer buf_n5452( .i (n5451), .o (n5452) );
  assign n5453 = n680 & n5452 ;
  buffer buf_n5454( .i (n5453), .o (n5454) );
  assign n5455 = n4646 | n5454 ;
  assign n5456 = n680 | n5452 ;
  buffer buf_n5457( .i (n5456), .o (n5457) );
  buffer buf_n5458( .i (n5457), .o (n5458) );
  assign n5459 = n5455 & n5458 ;
  buffer buf_n5460( .i (n5459), .o (n5460) );
  assign n5461 = n1590 & n5460 ;
  buffer buf_n5462( .i (n5461), .o (n5462) );
  assign n5463 = n4581 | n5462 ;
  assign n5464 = n1590 | n5460 ;
  buffer buf_n5465( .i (n5464), .o (n5465) );
  buffer buf_n5466( .i (n5465), .o (n5466) );
  assign n5467 = n5463 & n5466 ;
  buffer buf_n5468( .i (n5467), .o (n5468) );
  assign n5469 = n4351 & n5468 ;
  buffer buf_n5470( .i (n5469), .o (n5470) );
  assign n5472 = n4351 | n5468 ;
  buffer buf_n5473( .i (n5472), .o (n5473) );
  assign n5474 = ~n5470 & n5473 ;
  buffer buf_n5475( .i (n5474), .o (n5475) );
  buffer buf_n1391( .i (x24), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n3913( .i (n3912), .o (n3913) );
  buffer buf_n3914( .i (n3913), .o (n3914) );
  assign n5476 = n409 | n4515 ;
  buffer buf_n5477( .i (n5476), .o (n5477) );
  assign n5478 = n3914 & n5477 ;
  buffer buf_n5479( .i (n5478), .o (n5479) );
  assign n5480 = n1439 & ~n5479 ;
  assign n5481 = ~n1439 & n5479 ;
  assign n5482 = n5480 | n5481 ;
  buffer buf_n5483( .i (n5482), .o (n5483) );
  buffer buf_n5484( .i (n5483), .o (n5484) );
  buffer buf_n5485( .i (n5484), .o (n5485) );
  buffer buf_n5486( .i (n5485), .o (n5486) );
  buffer buf_n5487( .i (n5486), .o (n5487) );
  buffer buf_n5488( .i (n5487), .o (n5488) );
  buffer buf_n5489( .i (n5488), .o (n5489) );
  buffer buf_n5490( .i (n5489), .o (n5490) );
  buffer buf_n5491( .i (n5490), .o (n5491) );
  buffer buf_n5492( .i (n5491), .o (n5492) );
  buffer buf_n5493( .i (n5492), .o (n5493) );
  buffer buf_n5494( .i (n5493), .o (n5494) );
  buffer buf_n5495( .i (n5494), .o (n5495) );
  buffer buf_n5496( .i (n5495), .o (n5496) );
  buffer buf_n5497( .i (n5496), .o (n5497) );
  buffer buf_n5498( .i (n5497), .o (n5498) );
  buffer buf_n5499( .i (n5498), .o (n5499) );
  buffer buf_n5500( .i (n5499), .o (n5500) );
  buffer buf_n5501( .i (n5500), .o (n5501) );
  buffer buf_n5502( .i (n5501), .o (n5502) );
  buffer buf_n5503( .i (n5502), .o (n5503) );
  buffer buf_n5504( .i (n5503), .o (n5504) );
  buffer buf_n5505( .i (n5504), .o (n5505) );
  buffer buf_n5506( .i (n5505), .o (n5506) );
  buffer buf_n5507( .i (n5506), .o (n5507) );
  buffer buf_n5508( .i (n5507), .o (n5508) );
  buffer buf_n5509( .i (n5508), .o (n5509) );
  buffer buf_n5510( .i (n5509), .o (n5510) );
  buffer buf_n5511( .i (n5510), .o (n5511) );
  buffer buf_n5512( .i (n5511), .o (n5512) );
  buffer buf_n5513( .i (n5512), .o (n5513) );
  buffer buf_n5514( .i (n5513), .o (n5514) );
  buffer buf_n5515( .i (n5514), .o (n5515) );
  buffer buf_n5516( .i (n5515), .o (n5516) );
  buffer buf_n5517( .i (n5516), .o (n5517) );
  buffer buf_n5518( .i (n5517), .o (n5518) );
  buffer buf_n5519( .i (n5518), .o (n5519) );
  buffer buf_n5520( .i (n5519), .o (n5520) );
  buffer buf_n5521( .i (n5520), .o (n5521) );
  buffer buf_n5522( .i (n5521), .o (n5522) );
  buffer buf_n5523( .i (n5522), .o (n5523) );
  buffer buf_n5524( .i (n5523), .o (n5524) );
  buffer buf_n5525( .i (n5524), .o (n5525) );
  buffer buf_n5526( .i (n5525), .o (n5526) );
  buffer buf_n5527( .i (n5526), .o (n5527) );
  buffer buf_n5528( .i (n5527), .o (n5528) );
  buffer buf_n5529( .i (n5528), .o (n5529) );
  buffer buf_n5530( .i (n5529), .o (n5530) );
  buffer buf_n5531( .i (n5530), .o (n5531) );
  buffer buf_n5532( .i (n5531), .o (n5532) );
  buffer buf_n5533( .i (n5532), .o (n5533) );
  buffer buf_n5534( .i (n5533), .o (n5534) );
  buffer buf_n5535( .i (n5534), .o (n5535) );
  buffer buf_n5536( .i (n5535), .o (n5536) );
  buffer buf_n5537( .i (n5536), .o (n5537) );
  buffer buf_n5538( .i (n5537), .o (n5538) );
  buffer buf_n5539( .i (n5538), .o (n5539) );
  buffer buf_n5540( .i (n5539), .o (n5540) );
  buffer buf_n5541( .i (n5540), .o (n5541) );
  buffer buf_n5542( .i (n5541), .o (n5542) );
  buffer buf_n5543( .i (n5542), .o (n5543) );
  buffer buf_n5544( .i (n5543), .o (n5544) );
  buffer buf_n5545( .i (n5544), .o (n5545) );
  buffer buf_n5546( .i (n5545), .o (n5546) );
  buffer buf_n5547( .i (n5546), .o (n5547) );
  buffer buf_n5548( .i (n5547), .o (n5548) );
  assign n5549 = n5475 & n5548 ;
  assign n5550 = n5475 | n5548 ;
  assign n5551 = ~n5549 & n5550 ;
  buffer buf_n5552( .i (n5551), .o (n5552) );
  buffer buf_n2236( .i (x38), .o (n2236) );
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  buffer buf_n2250( .i (n2249), .o (n2250) );
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  buffer buf_n2265( .i (n2264), .o (n2265) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  buffer buf_n2269( .i (n2268), .o (n2269) );
  buffer buf_n2270( .i (n2269), .o (n2270) );
  buffer buf_n3974( .i (x63), .o (n3974) );
  buffer buf_n3975( .i (n3974), .o (n3975) );
  buffer buf_n3976( .i (n3975), .o (n3976) );
  buffer buf_n3977( .i (n3976), .o (n3977) );
  buffer buf_n3978( .i (n3977), .o (n3978) );
  buffer buf_n3979( .i (n3978), .o (n3979) );
  buffer buf_n3980( .i (n3979), .o (n3980) );
  buffer buf_n3981( .i (n3980), .o (n3981) );
  buffer buf_n3982( .i (n3981), .o (n3982) );
  buffer buf_n3983( .i (n3982), .o (n3983) );
  buffer buf_n3984( .i (n3983), .o (n3984) );
  buffer buf_n3985( .i (n3984), .o (n3985) );
  buffer buf_n3986( .i (n3985), .o (n3986) );
  buffer buf_n3987( .i (n3986), .o (n3987) );
  buffer buf_n3988( .i (n3987), .o (n3988) );
  buffer buf_n3989( .i (n3988), .o (n3989) );
  buffer buf_n3990( .i (n3989), .o (n3990) );
  buffer buf_n3991( .i (n3990), .o (n3991) );
  buffer buf_n3992( .i (n3991), .o (n3992) );
  buffer buf_n3993( .i (n3992), .o (n3993) );
  buffer buf_n3994( .i (n3993), .o (n3994) );
  buffer buf_n3995( .i (n3994), .o (n3995) );
  buffer buf_n3996( .i (n3995), .o (n3996) );
  buffer buf_n3997( .i (n3996), .o (n3997) );
  buffer buf_n3998( .i (n3997), .o (n3998) );
  buffer buf_n3999( .i (n3998), .o (n3999) );
  buffer buf_n4000( .i (n3999), .o (n4000) );
  buffer buf_n4001( .i (n4000), .o (n4001) );
  buffer buf_n4002( .i (n4001), .o (n4002) );
  buffer buf_n4003( .i (n4002), .o (n4003) );
  buffer buf_n4004( .i (n4003), .o (n4004) );
  buffer buf_n4005( .i (n4004), .o (n4005) );
  buffer buf_n4006( .i (n4005), .o (n4006) );
  buffer buf_n4007( .i (n4006), .o (n4007) );
  buffer buf_n4008( .i (n4007), .o (n4008) );
  assign n5602 = ~n2270 & n4008 ;
  buffer buf_n291( .i (x6), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  assign n5603 = ~n324 & n3901 ;
  buffer buf_n5604( .i (n5603), .o (n5604) );
  assign n5605 = n5602 & n5604 ;
  assign n5606 = n321 | n4004 ;
  buffer buf_n5607( .i (n5606), .o (n5607) );
  buffer buf_n5608( .i (n5607), .o (n5608) );
  buffer buf_n5609( .i (n5608), .o (n5609) );
  buffer buf_n5610( .i (n5609), .o (n5610) );
  assign n5611 = n2269 | n3901 ;
  buffer buf_n5612( .i (n5611), .o (n5612) );
  assign n5613 = n5610 | n5612 ;
  assign n5614 = ~n5605 & n5613 ;
  buffer buf_n5615( .i (n5614), .o (n5615) );
  buffer buf_n5616( .i (n5615), .o (n5616) );
  buffer buf_n5617( .i (n5616), .o (n5617) );
  buffer buf_n5618( .i (n5617), .o (n5618) );
  buffer buf_n5619( .i (n5618), .o (n5619) );
  buffer buf_n5620( .i (n5619), .o (n5620) );
  buffer buf_n5621( .i (n5620), .o (n5621) );
  buffer buf_n5622( .i (n5621), .o (n5622) );
  buffer buf_n5623( .i (n5622), .o (n5623) );
  buffer buf_n5624( .i (n5623), .o (n5624) );
  buffer buf_n5625( .i (n5624), .o (n5625) );
  buffer buf_n5626( .i (n5625), .o (n5626) );
  buffer buf_n5627( .i (n5626), .o (n5627) );
  buffer buf_n5628( .i (n5627), .o (n5628) );
  buffer buf_n5629( .i (n5628), .o (n5629) );
  buffer buf_n5630( .i (n5629), .o (n5630) );
  buffer buf_n5631( .i (n5630), .o (n5631) );
  buffer buf_n5632( .i (n5631), .o (n5632) );
  buffer buf_n5633( .i (n5632), .o (n5633) );
  buffer buf_n5634( .i (n5633), .o (n5634) );
  buffer buf_n5635( .i (n5634), .o (n5635) );
  buffer buf_n5636( .i (n5635), .o (n5636) );
  buffer buf_n5637( .i (n5636), .o (n5637) );
  buffer buf_n5638( .i (n5637), .o (n5638) );
  buffer buf_n5639( .i (n5638), .o (n5639) );
  buffer buf_n5640( .i (n5639), .o (n5640) );
  buffer buf_n5641( .i (n5640), .o (n5641) );
  buffer buf_n5642( .i (n5641), .o (n5642) );
  buffer buf_n5643( .i (n5642), .o (n5643) );
  buffer buf_n5644( .i (n5643), .o (n5644) );
  buffer buf_n5645( .i (n5644), .o (n5645) );
  buffer buf_n5646( .i (n5645), .o (n5646) );
  buffer buf_n5647( .i (n5646), .o (n5647) );
  buffer buf_n5648( .i (n5647), .o (n5648) );
  buffer buf_n5649( .i (n5648), .o (n5649) );
  buffer buf_n5650( .i (n5649), .o (n5650) );
  buffer buf_n5651( .i (n5650), .o (n5651) );
  buffer buf_n5652( .i (n5651), .o (n5652) );
  buffer buf_n5653( .i (n5652), .o (n5653) );
  buffer buf_n5654( .i (n5653), .o (n5654) );
  buffer buf_n5655( .i (n5654), .o (n5655) );
  buffer buf_n5656( .i (n5655), .o (n5656) );
  buffer buf_n5657( .i (n5656), .o (n5657) );
  buffer buf_n5658( .i (n5657), .o (n5658) );
  buffer buf_n5659( .i (n5658), .o (n5659) );
  buffer buf_n5660( .i (n5659), .o (n5660) );
  buffer buf_n5661( .i (n5660), .o (n5661) );
  buffer buf_n5662( .i (n5661), .o (n5662) );
  buffer buf_n5663( .i (n5662), .o (n5663) );
  buffer buf_n5664( .i (n5663), .o (n5664) );
  buffer buf_n5665( .i (n5664), .o (n5665) );
  buffer buf_n5666( .i (n5665), .o (n5666) );
  buffer buf_n5667( .i (n5666), .o (n5667) );
  buffer buf_n5668( .i (n5667), .o (n5668) );
  buffer buf_n5669( .i (n5668), .o (n5669) );
  buffer buf_n5670( .i (n5669), .o (n5670) );
  buffer buf_n5671( .i (n5670), .o (n5671) );
  buffer buf_n5672( .i (n5671), .o (n5672) );
  buffer buf_n5673( .i (n5672), .o (n5673) );
  buffer buf_n5674( .i (n5673), .o (n5674) );
  buffer buf_n5675( .i (n5674), .o (n5675) );
  buffer buf_n5676( .i (n5675), .o (n5676) );
  buffer buf_n5677( .i (n5676), .o (n5677) );
  buffer buf_n5678( .i (n5677), .o (n5678) );
  buffer buf_n5679( .i (n5678), .o (n5679) );
  buffer buf_n5680( .i (n5679), .o (n5680) );
  buffer buf_n5681( .i (n5680), .o (n5681) );
  buffer buf_n5682( .i (n5681), .o (n5682) );
  buffer buf_n5683( .i (n5682), .o (n5683) );
  buffer buf_n5684( .i (n5683), .o (n5684) );
  buffer buf_n5685( .i (n5684), .o (n5685) );
  buffer buf_n5686( .i (n5685), .o (n5686) );
  buffer buf_n5687( .i (n5686), .o (n5687) );
  buffer buf_n5688( .i (n5687), .o (n5688) );
  buffer buf_n5689( .i (n5688), .o (n5689) );
  buffer buf_n5690( .i (n5689), .o (n5690) );
  buffer buf_n5691( .i (n5690), .o (n5691) );
  buffer buf_n5692( .i (n5691), .o (n5692) );
  buffer buf_n5693( .i (n5692), .o (n5693) );
  buffer buf_n5694( .i (n5693), .o (n5694) );
  buffer buf_n5695( .i (n5694), .o (n5695) );
  buffer buf_n5696( .i (n5695), .o (n5696) );
  assign n5744 = n5552 & ~n5696 ;
  buffer buf_n2271( .i (n2270), .o (n2271) );
  assign n5745 = n2271 & n5604 ;
  buffer buf_n5746( .i (n5745), .o (n5746) );
  buffer buf_n5747( .i (n5746), .o (n5747) );
  buffer buf_n5748( .i (n5747), .o (n5748) );
  buffer buf_n5749( .i (n5748), .o (n5749) );
  buffer buf_n5750( .i (n5749), .o (n5750) );
  buffer buf_n5751( .i (n5750), .o (n5751) );
  buffer buf_n5752( .i (n5751), .o (n5752) );
  assign n5875 = n5620 & ~n5752 ;
  buffer buf_n5876( .i (n5875), .o (n5876) );
  buffer buf_n5877( .i (n5876), .o (n5877) );
  buffer buf_n5878( .i (n5877), .o (n5878) );
  buffer buf_n5879( .i (n5878), .o (n5879) );
  buffer buf_n5880( .i (n5879), .o (n5880) );
  buffer buf_n5881( .i (n5880), .o (n5881) );
  buffer buf_n5882( .i (n5881), .o (n5882) );
  buffer buf_n5883( .i (n5882), .o (n5883) );
  buffer buf_n5884( .i (n5883), .o (n5884) );
  buffer buf_n5885( .i (n5884), .o (n5885) );
  assign n5886 = n318 & ~n4001 ;
  buffer buf_n5887( .i (n5886), .o (n5887) );
  assign n5894 = n2263 & ~n3895 ;
  buffer buf_n5895( .i (n5894), .o (n5895) );
  assign n5899 = n5887 & n5895 ;
  assign n5900 = ~n2264 & n3896 ;
  assign n5901 = n318 & n4001 ;
  buffer buf_n5902( .i (n5901), .o (n5902) );
  assign n5905 = n5900 & n5902 ;
  assign n5906 = n5899 | n5905 ;
  buffer buf_n5907( .i (n5906), .o (n5907) );
  buffer buf_n5908( .i (n5907), .o (n5908) );
  buffer buf_n5909( .i (n5908), .o (n5909) );
  buffer buf_n5910( .i (n5909), .o (n5910) );
  buffer buf_n5911( .i (n5910), .o (n5911) );
  buffer buf_n5912( .i (n5911), .o (n5912) );
  buffer buf_n5913( .i (n5912), .o (n5913) );
  buffer buf_n5914( .i (n5913), .o (n5914) );
  buffer buf_n5915( .i (n5914), .o (n5915) );
  buffer buf_n5916( .i (n5915), .o (n5916) );
  buffer buf_n5917( .i (n5916), .o (n5917) );
  buffer buf_n5918( .i (n5917), .o (n5918) );
  buffer buf_n5919( .i (n5918), .o (n5919) );
  buffer buf_n5920( .i (n5919), .o (n5920) );
  buffer buf_n5921( .i (n5920), .o (n5921) );
  buffer buf_n5922( .i (n5921), .o (n5922) );
  buffer buf_n5923( .i (n5922), .o (n5923) );
  buffer buf_n5924( .i (n5923), .o (n5924) );
  buffer buf_n5925( .i (n5924), .o (n5925) );
  buffer buf_n5926( .i (n5925), .o (n5926) );
  buffer buf_n5927( .i (n5926), .o (n5927) );
  buffer buf_n5928( .i (n5927), .o (n5928) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n2457( .i (x41), .o (n2457) );
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n2460( .i (n2459), .o (n2460) );
  buffer buf_n2461( .i (n2460), .o (n2461) );
  buffer buf_n2462( .i (n2461), .o (n2462) );
  buffer buf_n2463( .i (n2462), .o (n2463) );
  buffer buf_n2464( .i (n2463), .o (n2464) );
  buffer buf_n2465( .i (n2464), .o (n2465) );
  buffer buf_n2466( .i (n2465), .o (n2466) );
  buffer buf_n2467( .i (n2466), .o (n2467) );
  buffer buf_n2468( .i (n2467), .o (n2468) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  buffer buf_n2470( .i (n2469), .o (n2470) );
  buffer buf_n2471( .i (n2470), .o (n2471) );
  buffer buf_n2472( .i (n2471), .o (n2472) );
  buffer buf_n2473( .i (n2472), .o (n2473) );
  buffer buf_n2474( .i (n2473), .o (n2474) );
  buffer buf_n2475( .i (n2474), .o (n2475) );
  buffer buf_n2476( .i (n2475), .o (n2476) );
  buffer buf_n2477( .i (n2476), .o (n2477) );
  buffer buf_n2478( .i (n2477), .o (n2478) );
  buffer buf_n2479( .i (n2478), .o (n2479) );
  buffer buf_n2480( .i (n2479), .o (n2480) );
  buffer buf_n2481( .i (n2480), .o (n2481) );
  buffer buf_n2482( .i (n2481), .o (n2482) );
  buffer buf_n2483( .i (n2482), .o (n2483) );
  buffer buf_n2484( .i (n2483), .o (n2484) );
  buffer buf_n2485( .i (n2484), .o (n2485) );
  buffer buf_n2486( .i (n2485), .o (n2486) );
  buffer buf_n2487( .i (n2486), .o (n2487) );
  buffer buf_n2488( .i (n2487), .o (n2488) );
  buffer buf_n2489( .i (n2488), .o (n2489) );
  buffer buf_n2490( .i (n2489), .o (n2490) );
  buffer buf_n2491( .i (n2490), .o (n2491) );
  assign n5929 = n2491 & n5909 ;
  buffer buf_n2160( .i (n2159), .o (n2160) );
  buffer buf_n2161( .i (n2160), .o (n2161) );
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n2163( .i (n2162), .o (n2163) );
  buffer buf_n2164( .i (n2163), .o (n2164) );
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n2166( .i (n2165), .o (n2166) );
  buffer buf_n2167( .i (n2166), .o (n2167) );
  buffer buf_n2168( .i (n2167), .o (n2168) );
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  buffer buf_n2171( .i (n2170), .o (n2171) );
  buffer buf_n2172( .i (n2171), .o (n2172) );
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n2175( .i (n2174), .o (n2175) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n2177), .o (n2178) );
  buffer buf_n2179( .i (n2178), .o (n2179) );
  buffer buf_n2180( .i (n2179), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  buffer buf_n2182( .i (n2181), .o (n2182) );
  buffer buf_n2183( .i (n2182), .o (n2183) );
  buffer buf_n2184( .i (n2183), .o (n2184) );
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  buffer buf_n2187( .i (n2186), .o (n2187) );
  buffer buf_n2188( .i (n2187), .o (n2188) );
  buffer buf_n2189( .i (n2188), .o (n2189) );
  buffer buf_n2190( .i (n2189), .o (n2190) );
  assign n5930 = n2190 & ~n5909 ;
  assign n5931 = n5929 | n5930 ;
  buffer buf_n5932( .i (n5931), .o (n5932) );
  assign n5938 = n3905 & n5932 ;
  buffer buf_n5939( .i (n5938), .o (n5939) );
  buffer buf_n5940( .i (n5939), .o (n5940) );
  buffer buf_n5941( .i (n5940), .o (n5941) );
  buffer buf_n5942( .i (n5941), .o (n5942) );
  buffer buf_n5943( .i (n5942), .o (n5943) );
  buffer buf_n5944( .i (n5943), .o (n5944) );
  buffer buf_n5945( .i (n5944), .o (n5945) );
  assign n5946 = n130 & n5945 ;
  buffer buf_n5947( .i (n5946), .o (n5947) );
  buffer buf_n5948( .i (n5947), .o (n5948) );
  buffer buf_n5949( .i (n5948), .o (n5949) );
  buffer buf_n5950( .i (n5949), .o (n5950) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  buffer buf_n1846( .i (n1845), .o (n1846) );
  buffer buf_n1847( .i (n1846), .o (n1847) );
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n3526( .i (n3525), .o (n3526) );
  buffer buf_n3527( .i (n3526), .o (n3527) );
  buffer buf_n3528( .i (n3527), .o (n3528) );
  buffer buf_n3529( .i (n3528), .o (n3529) );
  buffer buf_n3530( .i (n3529), .o (n3530) );
  buffer buf_n3531( .i (n3530), .o (n3531) );
  buffer buf_n3532( .i (n3531), .o (n3532) );
  buffer buf_n3533( .i (n3532), .o (n3533) );
  buffer buf_n3534( .i (n3533), .o (n3534) );
  buffer buf_n3535( .i (n3534), .o (n3535) );
  buffer buf_n3536( .i (n3535), .o (n3536) );
  buffer buf_n3537( .i (n3536), .o (n3537) );
  buffer buf_n3538( .i (n3537), .o (n3538) );
  buffer buf_n3539( .i (n3538), .o (n3539) );
  buffer buf_n3540( .i (n3539), .o (n3540) );
  buffer buf_n3541( .i (n3540), .o (n3541) );
  buffer buf_n3542( .i (n3541), .o (n3542) );
  buffer buf_n3543( .i (n3542), .o (n3543) );
  buffer buf_n3544( .i (n3543), .o (n3544) );
  buffer buf_n3545( .i (n3544), .o (n3545) );
  buffer buf_n3546( .i (n3545), .o (n3546) );
  buffer buf_n3547( .i (n3546), .o (n3547) );
  buffer buf_n3548( .i (n3547), .o (n3548) );
  buffer buf_n3549( .i (n3548), .o (n3549) );
  buffer buf_n3550( .i (n3549), .o (n3550) );
  buffer buf_n3551( .i (n3550), .o (n3551) );
  buffer buf_n3552( .i (n3551), .o (n3552) );
  buffer buf_n3553( .i (n3552), .o (n3553) );
  buffer buf_n3554( .i (n3553), .o (n3554) );
  buffer buf_n3555( .i (n3554), .o (n3555) );
  buffer buf_n3556( .i (n3555), .o (n3556) );
  buffer buf_n3557( .i (n3556), .o (n3557) );
  buffer buf_n3558( .i (n3557), .o (n3558) );
  buffer buf_n3559( .i (n3558), .o (n3559) );
  buffer buf_n3560( .i (n3559), .o (n3560) );
  buffer buf_n3561( .i (n3560), .o (n3561) );
  buffer buf_n3562( .i (n3561), .o (n3562) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  assign n5952 = n41 & ~n5939 ;
  buffer buf_n5953( .i (n5952), .o (n5953) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  buffer buf_n2536( .i (n2535), .o (n2536) );
  buffer buf_n2537( .i (n2536), .o (n2537) );
  buffer buf_n2538( .i (n2537), .o (n2538) );
  buffer buf_n2539( .i (n2538), .o (n2539) );
  buffer buf_n2540( .i (n2539), .o (n2540) );
  buffer buf_n2541( .i (n2540), .o (n2541) );
  buffer buf_n2542( .i (n2541), .o (n2542) );
  buffer buf_n2543( .i (n2542), .o (n2543) );
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  buffer buf_n2551( .i (n2550), .o (n2551) );
  buffer buf_n2552( .i (n2551), .o (n2552) );
  buffer buf_n2553( .i (n2552), .o (n2553) );
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2555( .i (n2554), .o (n2555) );
  buffer buf_n2556( .i (n2555), .o (n2556) );
  buffer buf_n2557( .i (n2556), .o (n2557) );
  buffer buf_n2558( .i (n2557), .o (n2558) );
  buffer buf_n2559( .i (n2558), .o (n2559) );
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  buffer buf_n2563( .i (n2562), .o (n2563) );
  buffer buf_n2564( .i (n2563), .o (n2564) );
  buffer buf_n2565( .i (n2564), .o (n2565) );
  buffer buf_n2566( .i (n2565), .o (n2566) );
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n2568( .i (n2567), .o (n2568) );
  buffer buf_n2925( .i (n2924), .o (n2925) );
  buffer buf_n2926( .i (n2925), .o (n2926) );
  buffer buf_n2927( .i (n2926), .o (n2927) );
  buffer buf_n2928( .i (n2927), .o (n2928) );
  buffer buf_n2929( .i (n2928), .o (n2929) );
  buffer buf_n2930( .i (n2929), .o (n2930) );
  buffer buf_n2931( .i (n2930), .o (n2931) );
  buffer buf_n2932( .i (n2931), .o (n2932) );
  buffer buf_n2933( .i (n2932), .o (n2933) );
  buffer buf_n2934( .i (n2933), .o (n2934) );
  buffer buf_n2935( .i (n2934), .o (n2935) );
  buffer buf_n2936( .i (n2935), .o (n2936) );
  buffer buf_n2937( .i (n2936), .o (n2937) );
  buffer buf_n2938( .i (n2937), .o (n2938) );
  buffer buf_n2939( .i (n2938), .o (n2939) );
  buffer buf_n2940( .i (n2939), .o (n2940) );
  buffer buf_n2941( .i (n2940), .o (n2941) );
  buffer buf_n2942( .i (n2941), .o (n2942) );
  buffer buf_n2943( .i (n2942), .o (n2943) );
  buffer buf_n2944( .i (n2943), .o (n2944) );
  buffer buf_n2945( .i (n2944), .o (n2945) );
  buffer buf_n2946( .i (n2945), .o (n2946) );
  buffer buf_n2947( .i (n2946), .o (n2947) );
  buffer buf_n2948( .i (n2947), .o (n2948) );
  buffer buf_n2949( .i (n2948), .o (n2949) );
  buffer buf_n2950( .i (n2949), .o (n2950) );
  buffer buf_n2951( .i (n2950), .o (n2951) );
  buffer buf_n2952( .i (n2951), .o (n2952) );
  buffer buf_n2953( .i (n2952), .o (n2953) );
  assign n5954 = n2953 & ~n5909 ;
  buffer buf_n3280( .i (x54), .o (n3280) );
  buffer buf_n3281( .i (n3280), .o (n3281) );
  buffer buf_n3282( .i (n3281), .o (n3282) );
  buffer buf_n3283( .i (n3282), .o (n3283) );
  buffer buf_n3284( .i (n3283), .o (n3284) );
  buffer buf_n3285( .i (n3284), .o (n3285) );
  buffer buf_n3286( .i (n3285), .o (n3286) );
  buffer buf_n3287( .i (n3286), .o (n3287) );
  buffer buf_n3288( .i (n3287), .o (n3288) );
  buffer buf_n3289( .i (n3288), .o (n3289) );
  buffer buf_n3290( .i (n3289), .o (n3290) );
  buffer buf_n3291( .i (n3290), .o (n3291) );
  buffer buf_n3292( .i (n3291), .o (n3292) );
  buffer buf_n3293( .i (n3292), .o (n3293) );
  buffer buf_n3294( .i (n3293), .o (n3294) );
  buffer buf_n3295( .i (n3294), .o (n3295) );
  buffer buf_n3296( .i (n3295), .o (n3296) );
  buffer buf_n3297( .i (n3296), .o (n3297) );
  buffer buf_n3298( .i (n3297), .o (n3298) );
  buffer buf_n3299( .i (n3298), .o (n3299) );
  buffer buf_n3300( .i (n3299), .o (n3300) );
  buffer buf_n3301( .i (n3300), .o (n3301) );
  buffer buf_n3302( .i (n3301), .o (n3302) );
  buffer buf_n3303( .i (n3302), .o (n3303) );
  buffer buf_n3304( .i (n3303), .o (n3304) );
  buffer buf_n3305( .i (n3304), .o (n3305) );
  buffer buf_n3306( .i (n3305), .o (n3306) );
  buffer buf_n3307( .i (n3306), .o (n3307) );
  buffer buf_n3308( .i (n3307), .o (n3308) );
  buffer buf_n3309( .i (n3308), .o (n3309) );
  buffer buf_n3310( .i (n3309), .o (n3310) );
  buffer buf_n3311( .i (n3310), .o (n3311) );
  buffer buf_n3312( .i (n3311), .o (n3312) );
  buffer buf_n3313( .i (n3312), .o (n3313) );
  buffer buf_n3314( .i (n3313), .o (n3314) );
  buffer buf_n5955( .i (n5908), .o (n5955) );
  assign n5956 = n3314 & n5955 ;
  assign n5957 = n5954 | n5956 ;
  buffer buf_n5958( .i (n5957), .o (n5958) );
  assign n5959 = ~n2568 & n5958 ;
  assign n5960 = n2568 & n5932 ;
  assign n5961 = n5959 | n5960 ;
  buffer buf_n5962( .i (n5961), .o (n5962) );
  assign n5963 = n42 | n5962 ;
  assign n5964 = ~n5953 & n5963 ;
  buffer buf_n5965( .i (n5964), .o (n5965) );
  assign n5966 = ~n3562 & n5965 ;
  assign n5967 = n3561 & n5942 ;
  buffer buf_n5968( .i (n5967), .o (n5968) );
  assign n5970 = n5966 | n5968 ;
  buffer buf_n5971( .i (n5970), .o (n5971) );
  assign n5972 = n1864 & ~n5971 ;
  assign n5973 = n3267 & ~n5955 ;
  assign n5974 = n4273 & n5955 ;
  assign n5975 = n5973 | n5974 ;
  buffer buf_n5976( .i (n5975), .o (n5976) );
  assign n5977 = ~n2568 & n5976 ;
  assign n5978 = n1475 & ~n5955 ;
  buffer buf_n1935( .i (x33), .o (n1935) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  buffer buf_n1954( .i (n1953), .o (n1954) );
  buffer buf_n1955( .i (n1954), .o (n1955) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  buffer buf_n1960( .i (n1959), .o (n1960) );
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n1967( .i (n1966), .o (n1967) );
  buffer buf_n1968( .i (n1967), .o (n1968) );
  buffer buf_n1969( .i (n1968), .o (n1969) );
  buffer buf_n5979( .i (n5908), .o (n5979) );
  assign n5980 = n1969 & n5979 ;
  assign n5981 = n5978 | n5980 ;
  buffer buf_n5982( .i (n5981), .o (n5982) );
  buffer buf_n5983( .i (n2567), .o (n5983) );
  assign n5984 = n5982 & n5983 ;
  assign n5985 = n5977 | n5984 ;
  buffer buf_n5986( .i (n5985), .o (n5986) );
  assign n5987 = ~n42 & n5986 ;
  buffer buf_n3744( .i (x60), .o (n3744) );
  buffer buf_n3745( .i (n3744), .o (n3745) );
  buffer buf_n3746( .i (n3745), .o (n3746) );
  buffer buf_n3747( .i (n3746), .o (n3747) );
  buffer buf_n3748( .i (n3747), .o (n3748) );
  buffer buf_n3749( .i (n3748), .o (n3749) );
  buffer buf_n3750( .i (n3749), .o (n3750) );
  buffer buf_n3751( .i (n3750), .o (n3751) );
  buffer buf_n3752( .i (n3751), .o (n3752) );
  buffer buf_n3753( .i (n3752), .o (n3753) );
  buffer buf_n3754( .i (n3753), .o (n3754) );
  buffer buf_n3755( .i (n3754), .o (n3755) );
  buffer buf_n3756( .i (n3755), .o (n3756) );
  buffer buf_n3757( .i (n3756), .o (n3757) );
  buffer buf_n3758( .i (n3757), .o (n3758) );
  buffer buf_n3759( .i (n3758), .o (n3759) );
  buffer buf_n3760( .i (n3759), .o (n3760) );
  buffer buf_n3761( .i (n3760), .o (n3761) );
  buffer buf_n3762( .i (n3761), .o (n3762) );
  buffer buf_n3763( .i (n3762), .o (n3763) );
  buffer buf_n3764( .i (n3763), .o (n3764) );
  buffer buf_n3765( .i (n3764), .o (n3765) );
  buffer buf_n3766( .i (n3765), .o (n3766) );
  buffer buf_n3767( .i (n3766), .o (n3767) );
  buffer buf_n3768( .i (n3767), .o (n3768) );
  buffer buf_n3769( .i (n3768), .o (n3769) );
  buffer buf_n3770( .i (n3769), .o (n3770) );
  buffer buf_n3771( .i (n3770), .o (n3771) );
  buffer buf_n3772( .i (n3771), .o (n3772) );
  buffer buf_n3773( .i (n3772), .o (n3773) );
  buffer buf_n3774( .i (n3773), .o (n3774) );
  buffer buf_n3775( .i (n3774), .o (n3775) );
  buffer buf_n3776( .i (n3775), .o (n3776) );
  buffer buf_n3777( .i (n3776), .o (n3777) );
  buffer buf_n3778( .i (n3777), .o (n3778) );
  assign n5988 = n3778 & n5979 ;
  assign n5989 = n81 & ~n5979 ;
  assign n5990 = n5988 | n5989 ;
  buffer buf_n5991( .i (n5990), .o (n5991) );
  assign n5992 = ~n5983 & n5991 ;
  buffer buf_n1143( .i (x21), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  assign n5993 = n1177 & n5979 ;
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n5994( .i (n5908), .o (n5994) );
  assign n5995 = n716 & ~n5994 ;
  assign n5996 = n5993 | n5995 ;
  buffer buf_n5997( .i (n5996), .o (n5997) );
  assign n5998 = n5983 & n5997 ;
  assign n5999 = n5992 | n5998 ;
  buffer buf_n6000( .i (n5999), .o (n6000) );
  assign n6001 = n42 & n6000 ;
  assign n6002 = n5987 | n6001 ;
  buffer buf_n6003( .i (n6002), .o (n6003) );
  assign n6004 = ~n3562 & n6003 ;
  buffer buf_n2273( .i (x39), .o (n2273) );
  buffer buf_n2274( .i (n2273), .o (n2274) );
  buffer buf_n2275( .i (n2274), .o (n2275) );
  buffer buf_n2276( .i (n2275), .o (n2276) );
  buffer buf_n2277( .i (n2276), .o (n2277) );
  buffer buf_n2278( .i (n2277), .o (n2278) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  buffer buf_n2280( .i (n2279), .o (n2280) );
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n2289( .i (n2288), .o (n2289) );
  buffer buf_n2290( .i (n2289), .o (n2290) );
  buffer buf_n2291( .i (n2290), .o (n2291) );
  buffer buf_n2292( .i (n2291), .o (n2292) );
  buffer buf_n2293( .i (n2292), .o (n2293) );
  buffer buf_n2294( .i (n2293), .o (n2294) );
  buffer buf_n2295( .i (n2294), .o (n2295) );
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n2297( .i (n2296), .o (n2297) );
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  buffer buf_n2307( .i (n2306), .o (n2307) );
  assign n6005 = n2307 & n5994 ;
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  assign n6006 = n484 & ~n5994 ;
  assign n6007 = n6005 | n6006 ;
  buffer buf_n6008( .i (n6007), .o (n6008) );
  assign n6009 = ~n5983 & n6008 ;
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  assign n6010 = n1306 & ~n5994 ;
  buffer buf_n2959( .i (x50), .o (n2959) );
  buffer buf_n2960( .i (n2959), .o (n2960) );
  buffer buf_n2961( .i (n2960), .o (n2961) );
  buffer buf_n2962( .i (n2961), .o (n2962) );
  buffer buf_n2963( .i (n2962), .o (n2963) );
  buffer buf_n2964( .i (n2963), .o (n2964) );
  buffer buf_n2965( .i (n2964), .o (n2965) );
  buffer buf_n2966( .i (n2965), .o (n2966) );
  buffer buf_n2967( .i (n2966), .o (n2967) );
  buffer buf_n2968( .i (n2967), .o (n2968) );
  buffer buf_n2969( .i (n2968), .o (n2969) );
  buffer buf_n2970( .i (n2969), .o (n2970) );
  buffer buf_n2971( .i (n2970), .o (n2971) );
  buffer buf_n2972( .i (n2971), .o (n2972) );
  buffer buf_n2973( .i (n2972), .o (n2973) );
  buffer buf_n2974( .i (n2973), .o (n2974) );
  buffer buf_n2975( .i (n2974), .o (n2975) );
  buffer buf_n2976( .i (n2975), .o (n2976) );
  buffer buf_n2977( .i (n2976), .o (n2977) );
  buffer buf_n2978( .i (n2977), .o (n2978) );
  buffer buf_n2979( .i (n2978), .o (n2979) );
  buffer buf_n2980( .i (n2979), .o (n2980) );
  buffer buf_n2981( .i (n2980), .o (n2981) );
  buffer buf_n2982( .i (n2981), .o (n2982) );
  buffer buf_n2983( .i (n2982), .o (n2983) );
  buffer buf_n2984( .i (n2983), .o (n2984) );
  buffer buf_n2985( .i (n2984), .o (n2985) );
  buffer buf_n2986( .i (n2985), .o (n2986) );
  buffer buf_n2987( .i (n2986), .o (n2987) );
  buffer buf_n2988( .i (n2987), .o (n2988) );
  buffer buf_n2989( .i (n2988), .o (n2989) );
  buffer buf_n2990( .i (n2989), .o (n2990) );
  buffer buf_n2991( .i (n2990), .o (n2991) );
  buffer buf_n2992( .i (n2991), .o (n2992) );
  buffer buf_n2993( .i (n2992), .o (n2993) );
  buffer buf_n6011( .i (n5907), .o (n6011) );
  buffer buf_n6012( .i (n6011), .o (n6012) );
  assign n6013 = n2993 & n6012 ;
  assign n6014 = n6010 | n6013 ;
  buffer buf_n6015( .i (n6014), .o (n6015) );
  buffer buf_n6016( .i (n2567), .o (n6016) );
  assign n6017 = n6015 & n6016 ;
  assign n6018 = n6009 | n6017 ;
  buffer buf_n6019( .i (n6018), .o (n6019) );
  buffer buf_n6020( .i (n41), .o (n6020) );
  assign n6021 = n6019 & n6020 ;
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  assign n6022 = n754 & ~n6012 ;
  buffer buf_n4053( .i (x65), .o (n4053) );
  buffer buf_n4054( .i (n4053), .o (n4054) );
  buffer buf_n4055( .i (n4054), .o (n4055) );
  buffer buf_n4056( .i (n4055), .o (n4056) );
  buffer buf_n4057( .i (n4056), .o (n4057) );
  buffer buf_n4058( .i (n4057), .o (n4058) );
  buffer buf_n4059( .i (n4058), .o (n4059) );
  buffer buf_n4060( .i (n4059), .o (n4060) );
  buffer buf_n4061( .i (n4060), .o (n4061) );
  buffer buf_n4062( .i (n4061), .o (n4062) );
  buffer buf_n4063( .i (n4062), .o (n4063) );
  buffer buf_n4064( .i (n4063), .o (n4064) );
  buffer buf_n4065( .i (n4064), .o (n4065) );
  buffer buf_n4066( .i (n4065), .o (n4066) );
  buffer buf_n4067( .i (n4066), .o (n4067) );
  buffer buf_n4068( .i (n4067), .o (n4068) );
  buffer buf_n4069( .i (n4068), .o (n4069) );
  buffer buf_n4070( .i (n4069), .o (n4070) );
  buffer buf_n4071( .i (n4070), .o (n4071) );
  buffer buf_n4072( .i (n4071), .o (n4072) );
  buffer buf_n4073( .i (n4072), .o (n4073) );
  buffer buf_n4074( .i (n4073), .o (n4074) );
  buffer buf_n4075( .i (n4074), .o (n4075) );
  buffer buf_n4076( .i (n4075), .o (n4076) );
  buffer buf_n4077( .i (n4076), .o (n4077) );
  buffer buf_n4078( .i (n4077), .o (n4078) );
  buffer buf_n4079( .i (n4078), .o (n4079) );
  buffer buf_n4080( .i (n4079), .o (n4080) );
  buffer buf_n4081( .i (n4080), .o (n4081) );
  buffer buf_n4082( .i (n4081), .o (n4082) );
  buffer buf_n4083( .i (n4082), .o (n4083) );
  buffer buf_n4084( .i (n4083), .o (n4084) );
  buffer buf_n4085( .i (n4084), .o (n4085) );
  buffer buf_n4086( .i (n4085), .o (n4086) );
  buffer buf_n4087( .i (n4086), .o (n4087) );
  assign n6023 = n4087 & n6012 ;
  assign n6024 = n6022 | n6023 ;
  buffer buf_n6025( .i (n6024), .o (n6025) );
  assign n6026 = ~n6016 & n6025 ;
  buffer buf_n4034( .i (n4033), .o (n4034) );
  buffer buf_n4035( .i (n4034), .o (n4035) );
  buffer buf_n4036( .i (n4035), .o (n4036) );
  buffer buf_n4037( .i (n4036), .o (n4037) );
  buffer buf_n4038( .i (n4037), .o (n4038) );
  buffer buf_n4039( .i (n4038), .o (n4039) );
  buffer buf_n4040( .i (n4039), .o (n4040) );
  buffer buf_n4041( .i (n4040), .o (n4041) );
  buffer buf_n4042( .i (n4041), .o (n4042) );
  buffer buf_n4043( .i (n4042), .o (n4043) );
  buffer buf_n4044( .i (n4043), .o (n4044) );
  buffer buf_n4045( .i (n4044), .o (n4045) );
  buffer buf_n4046( .i (n4045), .o (n4046) );
  buffer buf_n4047( .i (n4046), .o (n4047) );
  assign n6027 = n4047 & ~n6012 ;
  buffer buf_n3566( .i (x58), .o (n3566) );
  buffer buf_n3567( .i (n3566), .o (n3567) );
  buffer buf_n3568( .i (n3567), .o (n3568) );
  buffer buf_n3569( .i (n3568), .o (n3569) );
  buffer buf_n3570( .i (n3569), .o (n3570) );
  buffer buf_n3571( .i (n3570), .o (n3571) );
  buffer buf_n3572( .i (n3571), .o (n3572) );
  buffer buf_n3573( .i (n3572), .o (n3573) );
  buffer buf_n3574( .i (n3573), .o (n3574) );
  buffer buf_n3575( .i (n3574), .o (n3575) );
  buffer buf_n3576( .i (n3575), .o (n3576) );
  buffer buf_n3577( .i (n3576), .o (n3577) );
  buffer buf_n3578( .i (n3577), .o (n3578) );
  buffer buf_n3579( .i (n3578), .o (n3579) );
  buffer buf_n3580( .i (n3579), .o (n3580) );
  buffer buf_n3581( .i (n3580), .o (n3581) );
  buffer buf_n3582( .i (n3581), .o (n3582) );
  buffer buf_n3583( .i (n3582), .o (n3583) );
  buffer buf_n3584( .i (n3583), .o (n3584) );
  buffer buf_n3585( .i (n3584), .o (n3585) );
  buffer buf_n3586( .i (n3585), .o (n3586) );
  buffer buf_n3587( .i (n3586), .o (n3587) );
  buffer buf_n3588( .i (n3587), .o (n3588) );
  buffer buf_n3589( .i (n3588), .o (n3589) );
  buffer buf_n3590( .i (n3589), .o (n3590) );
  buffer buf_n3591( .i (n3590), .o (n3591) );
  buffer buf_n3592( .i (n3591), .o (n3592) );
  buffer buf_n3593( .i (n3592), .o (n3593) );
  buffer buf_n3594( .i (n3593), .o (n3594) );
  buffer buf_n3595( .i (n3594), .o (n3595) );
  buffer buf_n3596( .i (n3595), .o (n3596) );
  buffer buf_n3597( .i (n3596), .o (n3597) );
  buffer buf_n3598( .i (n3597), .o (n3598) );
  buffer buf_n3599( .i (n3598), .o (n3599) );
  buffer buf_n3600( .i (n3599), .o (n3600) );
  buffer buf_n6028( .i (n6011), .o (n6028) );
  assign n6029 = n3600 & n6028 ;
  assign n6030 = n6027 | n6029 ;
  buffer buf_n6031( .i (n6030), .o (n6031) );
  assign n6032 = n6016 & n6031 ;
  assign n6033 = n6026 | n6032 ;
  buffer buf_n6034( .i (n6033), .o (n6034) );
  assign n6035 = ~n6020 & n6034 ;
  assign n6036 = n6021 | n6035 ;
  buffer buf_n6037( .i (n6036), .o (n6037) );
  assign n6038 = n3562 & n6037 ;
  assign n6039 = n6004 | n6038 ;
  buffer buf_n6040( .i (n6039), .o (n6040) );
  assign n6042 = n1864 | n6040 ;
  assign n6043 = ~n5972 & n6042 ;
  buffer buf_n6044( .i (n6043), .o (n6044) );
  assign n6045 = ~n134 & n6044 ;
  assign n6046 = n5950 | n6045 ;
  buffer buf_n6047( .i (n6046), .o (n6047) );
  buffer buf_n6048( .i (n6047), .o (n6048) );
  assign n6049 = n5928 & ~n6048 ;
  assign n6050 = n5885 & ~n6049 ;
  buffer buf_n5896( .i (n5895), .o (n5896) );
  buffer buf_n5897( .i (n5896), .o (n5897) );
  buffer buf_n5903( .i (n5902), .o (n5903) );
  buffer buf_n5904( .i (n5903), .o (n5904) );
  assign n6051 = n5897 & n5904 ;
  buffer buf_n6052( .i (n6051), .o (n6052) );
  buffer buf_n6053( .i (n6052), .o (n6053) );
  buffer buf_n6054( .i (n6053), .o (n6054) );
  buffer buf_n6055( .i (n6054), .o (n6055) );
  buffer buf_n6056( .i (n6055), .o (n6056) );
  buffer buf_n6057( .i (n6056), .o (n6057) );
  buffer buf_n6058( .i (n6057), .o (n6058) );
  assign n6060 = n4278 & ~n6058 ;
  buffer buf_n6061( .i (n6060), .o (n6061) );
  assign n6062 = ~n322 & n5897 ;
  buffer buf_n6063( .i (n6062), .o (n6063) );
  buffer buf_n6064( .i (n6063), .o (n6064) );
  buffer buf_n6065( .i (n6064), .o (n6065) );
  buffer buf_n6066( .i (n6065), .o (n6066) );
  buffer buf_n6067( .i (n6066), .o (n6067) );
  buffer buf_n6068( .i (n6067), .o (n6068) );
  buffer buf_n6069( .i (n6068), .o (n6069) );
  assign n6071 = n4278 | n6069 ;
  assign n6072 = n1431 & n6071 ;
  assign n6073 = n6061 | n6072 ;
  buffer buf_n6074( .i (n6073), .o (n6074) );
  buffer buf_n5898( .i (n5897), .o (n5898) );
  assign n6075 = ~n5607 & n5898 ;
  buffer buf_n6076( .i (n6075), .o (n6076) );
  buffer buf_n6077( .i (n6076), .o (n6077) );
  buffer buf_n6078( .i (n6077), .o (n6078) );
  buffer buf_n6079( .i (n6078), .o (n6079) );
  buffer buf_n6080( .i (n6079), .o (n6080) );
  buffer buf_n6081( .i (n6080), .o (n6081) );
  buffer buf_n6082( .i (n6081), .o (n6082) );
  assign n6083 = n1431 & n6082 ;
  assign n6084 = n6061 & n6083 ;
  buffer buf_n5888( .i (n5887), .o (n5888) );
  buffer buf_n5889( .i (n5888), .o (n5889) );
  buffer buf_n5890( .i (n5889), .o (n5890) );
  buffer buf_n5891( .i (n5890), .o (n5891) );
  buffer buf_n5892( .i (n5891), .o (n5892) );
  buffer buf_n5893( .i (n5892), .o (n5893) );
  assign n6085 = ~n5612 & n5893 ;
  buffer buf_n6086( .i (n6085), .o (n6086) );
  buffer buf_n6087( .i (n6086), .o (n6087) );
  buffer buf_n6088( .i (n6087), .o (n6088) );
  buffer buf_n6089( .i (n6088), .o (n6089) );
  buffer buf_n6090( .i (n6089), .o (n6090) );
  buffer buf_n6091( .i (n6090), .o (n6091) );
  assign n6103 = n6084 | n6091 ;
  assign n6104 = n6074 & ~n6103 ;
  assign n6105 = n5919 | n6104 ;
  buffer buf_n6106( .i (n6105), .o (n6106) );
  buffer buf_n6107( .i (n6106), .o (n6107) );
  buffer buf_n6108( .i (n6107), .o (n6108) );
  buffer buf_n6109( .i (n6108), .o (n6109) );
  buffer buf_n6110( .i (n6109), .o (n6110) );
  buffer buf_n6111( .i (n6110), .o (n6111) );
  buffer buf_n6112( .i (n6111), .o (n6112) );
  buffer buf_n6113( .i (n6112), .o (n6113) );
  buffer buf_n6114( .i (n6113), .o (n6114) );
  buffer buf_n6092( .i (n6091), .o (n6092) );
  buffer buf_n6093( .i (n6092), .o (n6093) );
  buffer buf_n6094( .i (n6093), .o (n6094) );
  buffer buf_n6095( .i (n6094), .o (n6095) );
  buffer buf_n6096( .i (n6095), .o (n6096) );
  buffer buf_n6097( .i (n6096), .o (n6097) );
  buffer buf_n6098( .i (n6097), .o (n6098) );
  buffer buf_n6099( .i (n6098), .o (n6099) );
  buffer buf_n6100( .i (n6099), .o (n6100) );
  buffer buf_n6101( .i (n6100), .o (n6101) );
  buffer buf_n6102( .i (n6101), .o (n6102) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n3563( .i (n3562), .o (n3563) );
  buffer buf_n43( .i (n42), .o (n43) );
  assign n6115 = n6016 & n6025 ;
  buffer buf_n6116( .i (n2567), .o (n6116) );
  assign n6117 = n5997 & ~n6116 ;
  assign n6118 = n6115 | n6117 ;
  buffer buf_n6119( .i (n6118), .o (n6119) );
  buffer buf_n6120( .i (n6119), .o (n6120) );
  assign n6121 = ~n43 & n6120 ;
  assign n6122 = n6008 & n6116 ;
  assign n6123 = n6031 & ~n6116 ;
  assign n6124 = n6122 | n6123 ;
  buffer buf_n6125( .i (n6124), .o (n6125) );
  buffer buf_n6126( .i (n6125), .o (n6126) );
  assign n6127 = n43 & n6126 ;
  assign n6128 = n6121 | n6127 ;
  buffer buf_n6129( .i (n6128), .o (n6129) );
  assign n6130 = ~n3563 & n6129 ;
  buffer buf_n2569( .i (n2568), .o (n2569) );
  buffer buf_n2570( .i (n2569), .o (n2570) );
  buffer buf_n5933( .i (n5932), .o (n5933) );
  buffer buf_n5934( .i (n5933), .o (n5934) );
  assign n6131 = ~n2570 & n5934 ;
  buffer buf_n6132( .i (n6131), .o (n6132) );
  assign n6133 = n5953 & ~n6132 ;
  assign n6134 = n6015 & ~n6116 ;
  buffer buf_n6135( .i (n2566), .o (n6135) );
  buffer buf_n6136( .i (n6135), .o (n6136) );
  assign n6137 = n5958 & n6136 ;
  assign n6138 = n6134 | n6137 ;
  buffer buf_n6139( .i (n6138), .o (n6139) );
  buffer buf_n6140( .i (n6139), .o (n6140) );
  assign n6141 = n43 | n6140 ;
  assign n6142 = ~n6133 & n6141 ;
  buffer buf_n6143( .i (n6142), .o (n6143) );
  assign n6144 = n3563 & n6143 ;
  assign n6145 = n6130 | n6144 ;
  buffer buf_n6146( .i (n6145), .o (n6146) );
  assign n6147 = ~n1865 & n6146 ;
  assign n6148 = n1862 & n5944 ;
  buffer buf_n6149( .i (n6148), .o (n6149) );
  buffer buf_n6150( .i (n6149), .o (n6150) );
  buffer buf_n6151( .i (n6150), .o (n6151) );
  assign n6152 = n6147 | n6151 ;
  buffer buf_n6153( .i (n6152), .o (n6153) );
  assign n6154 = n135 & ~n6153 ;
  assign n6155 = n4222 & n5910 ;
  assign n6156 = n1518 & ~n5910 ;
  assign n6157 = n6155 | n6156 ;
  buffer buf_n6158( .i (n6157), .o (n6158) );
  assign n6159 = n2569 & n6158 ;
  assign n6160 = n4274 & ~n5910 ;
  buffer buf_n6161( .i (n6028), .o (n6161) );
  assign n6162 = n3268 & n6161 ;
  assign n6163 = n6160 | n6162 ;
  buffer buf_n6164( .i (n6163), .o (n6164) );
  assign n6165 = ~n2569 & n6164 ;
  assign n6166 = n6159 | n6165 ;
  buffer buf_n6167( .i (n6166), .o (n6167) );
  buffer buf_n6169( .i (n6020), .o (n6169) );
  assign n6170 = n6167 & ~n6169 ;
  assign n6171 = n1679 & ~n6161 ;
  assign n6172 = n2128 & n6161 ;
  assign n6173 = n6171 | n6172 ;
  buffer buf_n6174( .i (n6173), .o (n6174) );
  assign n6175 = n2569 & n6174 ;
  assign n6176 = n613 & ~n6161 ;
  buffer buf_n6177( .i (n6028), .o (n6177) );
  assign n6178 = n211 & n6177 ;
  assign n6179 = n6176 | n6178 ;
  buffer buf_n6180( .i (n6179), .o (n6180) );
  buffer buf_n6181( .i (n6136), .o (n6181) );
  assign n6182 = n6180 & ~n6181 ;
  assign n6183 = n6175 | n6182 ;
  buffer buf_n6184( .i (n6183), .o (n6184) );
  assign n6185 = n6169 & n6184 ;
  assign n6186 = n6170 | n6185 ;
  buffer buf_n6187( .i (n6186), .o (n6187) );
  assign n6189 = ~n3563 & n6187 ;
  assign n6190 = n1346 & ~n6028 ;
  buffer buf_n6191( .i (n6011), .o (n6191) );
  assign n6192 = n2869 & n6191 ;
  assign n6193 = n6190 | n6192 ;
  buffer buf_n6194( .i (n6193), .o (n6194) );
  buffer buf_n6195( .i (n6194), .o (n6195) );
  assign n6196 = n6181 & ~n6195 ;
  assign n6197 = n1347 & n6177 ;
  assign n6198 = n2870 & ~n6177 ;
  assign n6199 = n6197 | n6198 ;
  buffer buf_n6200( .i (n6199), .o (n6200) );
  assign n6201 = n6181 | n6200 ;
  assign n6202 = ~n6196 & n6201 ;
  buffer buf_n6203( .i (n6202), .o (n6203) );
  assign n6204 = n6169 & n6203 ;
  assign n6205 = n1902 & n6177 ;
  buffer buf_n6206( .i (n6191), .o (n6206) );
  assign n6207 = n793 & ~n6206 ;
  assign n6208 = n6205 | n6207 ;
  buffer buf_n6209( .i (n6208), .o (n6209) );
  assign n6210 = ~n6181 & n6209 ;
  assign n6211 = n524 & ~n6206 ;
  assign n6212 = n1064 & n6206 ;
  assign n6213 = n6211 | n6212 ;
  buffer buf_n6214( .i (n6213), .o (n6214) );
  buffer buf_n6215( .i (n6136), .o (n6215) );
  assign n6216 = n6214 & n6215 ;
  assign n6217 = n6210 | n6216 ;
  buffer buf_n6218( .i (n6217), .o (n6218) );
  assign n6219 = ~n6169 & n6218 ;
  assign n6220 = n6204 | n6219 ;
  buffer buf_n6221( .i (n6220), .o (n6221) );
  buffer buf_n6222( .i (n3561), .o (n6222) );
  buffer buf_n6223( .i (n6222), .o (n6223) );
  assign n6224 = n6221 & n6223 ;
  assign n6225 = n6189 | n6224 ;
  buffer buf_n6226( .i (n6225), .o (n6226) );
  assign n6227 = ~n1865 & n6226 ;
  assign n6228 = n1901 & ~n6191 ;
  assign n6229 = n792 & n6191 ;
  assign n6230 = n6228 | n6229 ;
  buffer buf_n6231( .i (n6230), .o (n6231) );
  assign n6232 = n6136 & n6231 ;
  buffer buf_n6233( .i (n6011), .o (n6233) );
  assign n6234 = n523 & n6233 ;
  assign n6235 = n1063 & ~n6233 ;
  assign n6236 = n6234 | n6235 ;
  buffer buf_n6237( .i (n6236), .o (n6237) );
  buffer buf_n6238( .i (n6135), .o (n6238) );
  assign n6239 = n6237 & ~n6238 ;
  assign n6240 = n6232 | n6239 ;
  buffer buf_n6241( .i (n6240), .o (n6241) );
  assign n6243 = ~n6020 & n6241 ;
  assign n6244 = n210 & ~n6233 ;
  assign n6245 = n612 & n6233 ;
  assign n6246 = n6244 | n6245 ;
  buffer buf_n6247( .i (n6246), .o (n6247) );
  assign n6248 = n6238 & n6247 ;
  buffer buf_n6249( .i (n5907), .o (n6249) );
  buffer buf_n6250( .i (n6249), .o (n6250) );
  assign n6251 = n1678 & n6250 ;
  assign n6252 = n2127 & ~n6250 ;
  assign n6253 = n6251 | n6252 ;
  buffer buf_n6254( .i (n6253), .o (n6254) );
  assign n6255 = ~n6238 & n6254 ;
  assign n6256 = n6248 | n6255 ;
  buffer buf_n6257( .i (n6256), .o (n6257) );
  buffer buf_n6258( .i (n41), .o (n6258) );
  assign n6259 = n6257 & n6258 ;
  assign n6260 = n6243 | n6259 ;
  buffer buf_n6261( .i (n6260), .o (n6261) );
  assign n6263 = ~n6222 & n6261 ;
  assign n6264 = n5976 & n6238 ;
  assign n6265 = n1517 & n6250 ;
  assign n6266 = n4221 & ~n6250 ;
  assign n6267 = n6265 | n6266 ;
  buffer buf_n6268( .i (n6267), .o (n6268) );
  buffer buf_n6269( .i (n6135), .o (n6269) );
  assign n6270 = n6268 & ~n6269 ;
  assign n6271 = n6264 | n6270 ;
  buffer buf_n6272( .i (n6271), .o (n6272) );
  assign n6273 = ~n6258 & n6272 ;
  assign n6274 = n5991 & n6269 ;
  assign n6275 = n5982 & ~n6269 ;
  assign n6276 = n6274 | n6275 ;
  buffer buf_n6277( .i (n6276), .o (n6277) );
  assign n6278 = n6258 & n6277 ;
  assign n6279 = n6273 | n6278 ;
  buffer buf_n6280( .i (n6279), .o (n6280) );
  assign n6282 = n6222 & n6280 ;
  assign n6283 = n6263 | n6282 ;
  buffer buf_n6284( .i (n6283), .o (n6284) );
  assign n6286 = n1864 & n6284 ;
  assign n6287 = n132 | n6286 ;
  assign n6288 = n6227 | n6287 ;
  buffer buf_n6289( .i (n6288), .o (n6289) );
  buffer buf_n6290( .i (n6289), .o (n6290) );
  assign n6291 = ~n6154 & n6290 ;
  buffer buf_n6292( .i (n6291), .o (n6292) );
  assign n6293 = n6102 & n6292 ;
  assign n6294 = n6114 | n6293 ;
  assign n6295 = n6050 & n6294 ;
  buffer buf_n6296( .i (n6295), .o (n6296) );
  buffer buf_n6297( .i (n6296), .o (n6297) );
  buffer buf_n6298( .i (n6297), .o (n6298) );
  buffer buf_n6299( .i (n6298), .o (n6299) );
  buffer buf_n6300( .i (n6299), .o (n6300) );
  buffer buf_n6301( .i (n6300), .o (n6301) );
  buffer buf_n6302( .i (n6301), .o (n6302) );
  buffer buf_n6303( .i (n6302), .o (n6303) );
  buffer buf_n6304( .i (n6303), .o (n6304) );
  buffer buf_n6305( .i (n6304), .o (n6305) );
  buffer buf_n6306( .i (n6305), .o (n6306) );
  buffer buf_n6307( .i (n6306), .o (n6307) );
  buffer buf_n6308( .i (n6307), .o (n6308) );
  buffer buf_n6309( .i (n6308), .o (n6309) );
  buffer buf_n6310( .i (n6309), .o (n6310) );
  buffer buf_n6311( .i (n6310), .o (n6311) );
  buffer buf_n6312( .i (n6311), .o (n6312) );
  buffer buf_n6313( .i (n6312), .o (n6313) );
  buffer buf_n6314( .i (n6313), .o (n6314) );
  buffer buf_n6315( .i (n6314), .o (n6315) );
  buffer buf_n6316( .i (n6315), .o (n6316) );
  buffer buf_n6317( .i (n6316), .o (n6317) );
  buffer buf_n6318( .i (n6317), .o (n6318) );
  buffer buf_n6319( .i (n6318), .o (n6319) );
  buffer buf_n6320( .i (n6319), .o (n6320) );
  buffer buf_n6321( .i (n6320), .o (n6321) );
  buffer buf_n6322( .i (n6321), .o (n6322) );
  buffer buf_n6323( .i (n6322), .o (n6323) );
  buffer buf_n6324( .i (n6323), .o (n6324) );
  buffer buf_n6325( .i (n6324), .o (n6325) );
  buffer buf_n6326( .i (n6325), .o (n6326) );
  buffer buf_n6327( .i (n6326), .o (n6327) );
  buffer buf_n6328( .i (n6327), .o (n6328) );
  buffer buf_n6329( .i (n6328), .o (n6329) );
  buffer buf_n6330( .i (n6329), .o (n6330) );
  buffer buf_n6331( .i (n6330), .o (n6331) );
  buffer buf_n6332( .i (n6331), .o (n6332) );
  buffer buf_n6333( .i (n6332), .o (n6333) );
  buffer buf_n6334( .i (n6333), .o (n6334) );
  buffer buf_n6335( .i (n6334), .o (n6335) );
  buffer buf_n6336( .i (n6335), .o (n6336) );
  buffer buf_n6337( .i (n6336), .o (n6337) );
  buffer buf_n6338( .i (n6337), .o (n6338) );
  buffer buf_n6339( .i (n6338), .o (n6339) );
  buffer buf_n6340( .i (n6339), .o (n6340) );
  buffer buf_n6341( .i (n6340), .o (n6341) );
  buffer buf_n6342( .i (n6341), .o (n6342) );
  buffer buf_n6343( .i (n6342), .o (n6343) );
  buffer buf_n6344( .i (n6343), .o (n6344) );
  buffer buf_n6345( .i (n6344), .o (n6345) );
  buffer buf_n6346( .i (n6345), .o (n6346) );
  buffer buf_n6347( .i (n6346), .o (n6347) );
  buffer buf_n6348( .i (n6347), .o (n6348) );
  buffer buf_n6349( .i (n6348), .o (n6349) );
  buffer buf_n6350( .i (n6349), .o (n6350) );
  buffer buf_n6351( .i (n6350), .o (n6351) );
  buffer buf_n6352( .i (n6351), .o (n6352) );
  buffer buf_n6353( .i (n6352), .o (n6353) );
  buffer buf_n6354( .i (n6353), .o (n6354) );
  buffer buf_n6355( .i (n6354), .o (n6355) );
  buffer buf_n6356( .i (n6355), .o (n6356) );
  buffer buf_n6357( .i (n6356), .o (n6357) );
  buffer buf_n6358( .i (n6357), .o (n6358) );
  buffer buf_n6359( .i (n6358), .o (n6359) );
  assign n6360 = n5744 | n6359 ;
  buffer buf_n6361( .i (n6360), .o (n6361) );
  buffer buf_n6362( .i (n6361), .o (n6362) );
  buffer buf_n6363( .i (n6362), .o (n6363) );
  buffer buf_n6364( .i (n6363), .o (n6364) );
  buffer buf_n6365( .i (n6364), .o (n6365) );
  buffer buf_n6366( .i (n6365), .o (n6366) );
  buffer buf_n6367( .i (n6366), .o (n6367) );
  buffer buf_n6368( .i (n6367), .o (n6368) );
  buffer buf_n6369( .i (n6368), .o (n6369) );
  buffer buf_n6370( .i (n6369), .o (n6370) );
  buffer buf_n6371( .i (n6370), .o (n6371) );
  buffer buf_n6372( .i (n6371), .o (n6372) );
  buffer buf_n6373( .i (n6372), .o (n6373) );
  buffer buf_n6374( .i (n6373), .o (n6374) );
  buffer buf_n6375( .i (n6374), .o (n6375) );
  buffer buf_n6376( .i (n6375), .o (n6376) );
  buffer buf_n6377( .i (n6376), .o (n6377) );
  buffer buf_n6378( .i (n6377), .o (n6378) );
  buffer buf_n6379( .i (n6378), .o (n6379) );
  buffer buf_n6380( .i (n6379), .o (n6380) );
  buffer buf_n6381( .i (n6380), .o (n6381) );
  buffer buf_n6382( .i (n6381), .o (n6382) );
  buffer buf_n6383( .i (n6382), .o (n6383) );
  buffer buf_n6384( .i (n6383), .o (n6384) );
  buffer buf_n6385( .i (n6384), .o (n6385) );
  buffer buf_n6386( .i (n6385), .o (n6386) );
  buffer buf_n6387( .i (n6386), .o (n6387) );
  buffer buf_n6388( .i (n6387), .o (n6388) );
  buffer buf_n6389( .i (n6388), .o (n6389) );
  buffer buf_n6390( .i (n6389), .o (n6390) );
  buffer buf_n6391( .i (n6390), .o (n6391) );
  buffer buf_n6392( .i (n6391), .o (n6392) );
  buffer buf_n6393( .i (n6392), .o (n6393) );
  buffer buf_n6394( .i (n6393), .o (n6394) );
  buffer buf_n6395( .i (n6394), .o (n6395) );
  buffer buf_n6396( .i (n6395), .o (n6396) );
  buffer buf_n6397( .i (n6396), .o (n6397) );
  buffer buf_n6398( .i (n6397), .o (n6398) );
  buffer buf_n6399( .i (n6398), .o (n6399) );
  buffer buf_n6400( .i (n6399), .o (n6400) );
  buffer buf_n6401( .i (n6400), .o (n6401) );
  buffer buf_n6402( .i (n6401), .o (n6402) );
  buffer buf_n6403( .i (n6402), .o (n6403) );
  buffer buf_n6404( .i (n6403), .o (n6404) );
  buffer buf_n6405( .i (n6404), .o (n6405) );
  buffer buf_n6406( .i (n6405), .o (n6406) );
  buffer buf_n6407( .i (n6406), .o (n6407) );
  buffer buf_n5553( .i (n5552), .o (n5553) );
  buffer buf_n5554( .i (n5553), .o (n5554) );
  buffer buf_n5555( .i (n5554), .o (n5555) );
  buffer buf_n5556( .i (n5555), .o (n5556) );
  buffer buf_n5557( .i (n5556), .o (n5557) );
  buffer buf_n5558( .i (n5557), .o (n5558) );
  buffer buf_n5559( .i (n5558), .o (n5559) );
  buffer buf_n5560( .i (n5559), .o (n5560) );
  buffer buf_n5561( .i (n5560), .o (n5561) );
  buffer buf_n5562( .i (n5561), .o (n5562) );
  buffer buf_n5563( .i (n5562), .o (n5563) );
  buffer buf_n5564( .i (n5563), .o (n5564) );
  buffer buf_n5565( .i (n5564), .o (n5565) );
  buffer buf_n5566( .i (n5565), .o (n5566) );
  buffer buf_n5567( .i (n5566), .o (n5567) );
  buffer buf_n5568( .i (n5567), .o (n5568) );
  buffer buf_n5569( .i (n5568), .o (n5569) );
  buffer buf_n5570( .i (n5569), .o (n5570) );
  buffer buf_n5571( .i (n5570), .o (n5571) );
  buffer buf_n5572( .i (n5571), .o (n5572) );
  buffer buf_n5573( .i (n5572), .o (n5573) );
  buffer buf_n5574( .i (n5573), .o (n5574) );
  buffer buf_n5575( .i (n5574), .o (n5575) );
  buffer buf_n5576( .i (n5575), .o (n5576) );
  buffer buf_n5577( .i (n5576), .o (n5577) );
  buffer buf_n5578( .i (n5577), .o (n5578) );
  buffer buf_n5579( .i (n5578), .o (n5579) );
  buffer buf_n5580( .i (n5579), .o (n5580) );
  buffer buf_n5581( .i (n5580), .o (n5581) );
  buffer buf_n5582( .i (n5581), .o (n5582) );
  buffer buf_n5583( .i (n5582), .o (n5583) );
  buffer buf_n5584( .i (n5583), .o (n5584) );
  buffer buf_n5585( .i (n5584), .o (n5585) );
  buffer buf_n5586( .i (n5585), .o (n5586) );
  buffer buf_n5587( .i (n5586), .o (n5587) );
  buffer buf_n5588( .i (n5587), .o (n5588) );
  buffer buf_n5589( .i (n5588), .o (n5589) );
  buffer buf_n5590( .i (n5589), .o (n5590) );
  buffer buf_n5591( .i (n5590), .o (n5591) );
  buffer buf_n5592( .i (n5591), .o (n5592) );
  buffer buf_n5593( .i (n5592), .o (n5593) );
  buffer buf_n5594( .i (n5593), .o (n5594) );
  buffer buf_n5595( .i (n5594), .o (n5595) );
  buffer buf_n5596( .i (n5595), .o (n5596) );
  buffer buf_n5597( .i (n5596), .o (n5597) );
  buffer buf_n5598( .i (n5597), .o (n5598) );
  buffer buf_n5599( .i (n5598), .o (n5599) );
  buffer buf_n5600( .i (n5599), .o (n5600) );
  buffer buf_n5601( .i (n5600), .o (n5601) );
  buffer buf_n4956( .i (n4955), .o (n4956) );
  buffer buf_n4957( .i (n4956), .o (n4957) );
  assign n6408 = ~n4934 & n4960 ;
  buffer buf_n6409( .i (n6408), .o (n6409) );
  assign n6410 = n4957 & ~n6409 ;
  assign n6411 = ~n4957 & n6409 ;
  assign n6412 = n6410 | n6411 ;
  buffer buf_n6413( .i (n6412), .o (n6413) );
  buffer buf_n6414( .i (n6413), .o (n6414) );
  buffer buf_n6415( .i (n6414), .o (n6415) );
  buffer buf_n6416( .i (n6415), .o (n6416) );
  buffer buf_n6417( .i (n6416), .o (n6417) );
  buffer buf_n6418( .i (n6417), .o (n6418) );
  buffer buf_n6419( .i (n6418), .o (n6419) );
  buffer buf_n6420( .i (n6419), .o (n6420) );
  buffer buf_n6421( .i (n6420), .o (n6421) );
  buffer buf_n6422( .i (n6421), .o (n6422) );
  buffer buf_n6423( .i (n6422), .o (n6423) );
  buffer buf_n6424( .i (n6423), .o (n6424) );
  buffer buf_n6425( .i (n6424), .o (n6425) );
  assign n6540 = ~n5631 & n6425 ;
  assign n6541 = n6125 & ~n6258 ;
  buffer buf_n6542( .i (n40), .o (n6542) );
  buffer buf_n6543( .i (n6542), .o (n6543) );
  assign n6544 = n6139 & n6543 ;
  assign n6545 = n6541 | n6544 ;
  buffer buf_n6546( .i (n6545), .o (n6546) );
  assign n6547 = n6222 & n6546 ;
  assign n6548 = n6277 & ~n6543 ;
  assign n6549 = n6119 & n6543 ;
  assign n6550 = n6548 | n6549 ;
  buffer buf_n6551( .i (n6550), .o (n6551) );
  buffer buf_n6552( .i (n3561), .o (n6552) );
  assign n6553 = n6551 & ~n6552 ;
  assign n6554 = n6547 | n6553 ;
  buffer buf_n6555( .i (n6554), .o (n6555) );
  buffer buf_n6557( .i (n1863), .o (n6557) );
  assign n6558 = n6555 & ~n6557 ;
  buffer buf_n5935( .i (n5934), .o (n5935) );
  buffer buf_n4399( .i (n4398), .o (n4399) );
  buffer buf_n4400( .i (n4399), .o (n4400) );
  buffer buf_n4401( .i (n4400), .o (n4401) );
  buffer buf_n4402( .i (n4401), .o (n4402) );
  buffer buf_n4403( .i (n4402), .o (n4403) );
  buffer buf_n4404( .i (n4403), .o (n4404) );
  buffer buf_n4405( .i (n4404), .o (n4405) );
  buffer buf_n4406( .i (n4405), .o (n4406) );
  buffer buf_n4407( .i (n4406), .o (n4407) );
  buffer buf_n4408( .i (n4407), .o (n4408) );
  buffer buf_n4409( .i (n4408), .o (n4409) );
  buffer buf_n4410( .i (n4409), .o (n4410) );
  buffer buf_n4411( .i (n4410), .o (n4411) );
  buffer buf_n4412( .i (n4411), .o (n4412) );
  buffer buf_n4413( .i (n4412), .o (n4413) );
  buffer buf_n4414( .i (n4413), .o (n4414) );
  buffer buf_n4415( .i (n4414), .o (n4415) );
  buffer buf_n4416( .i (n4415), .o (n4416) );
  buffer buf_n4417( .i (n4416), .o (n4417) );
  buffer buf_n4418( .i (n4417), .o (n4418) );
  buffer buf_n4419( .i (n4418), .o (n4419) );
  buffer buf_n4420( .i (n4419), .o (n4420) );
  assign n6559 = ~n3902 & n4420 ;
  assign n6560 = n1853 & ~n6559 ;
  buffer buf_n6561( .i (n6560), .o (n6561) );
  buffer buf_n6562( .i (n6561), .o (n6562) );
  buffer buf_n6563( .i (n6562), .o (n6563) );
  buffer buf_n6564( .i (n6563), .o (n6564) );
  assign n6565 = n5935 & n6564 ;
  buffer buf_n6566( .i (n6565), .o (n6566) );
  buffer buf_n6567( .i (n6566), .o (n6567) );
  buffer buf_n6568( .i (n6567), .o (n6568) );
  buffer buf_n6569( .i (n6568), .o (n6569) );
  buffer buf_n6570( .i (n6569), .o (n6570) );
  buffer buf_n6571( .i (n6570), .o (n6571) );
  assign n6572 = n6558 | n6571 ;
  buffer buf_n6573( .i (n6572), .o (n6573) );
  assign n6574 = n134 & ~n6573 ;
  buffer buf_n3564( .i (n3563), .o (n3564) );
  buffer buf_n44( .i (n43), .o (n44) );
  assign n6575 = n1476 & n6206 ;
  buffer buf_n1970( .i (n1969), .o (n1970) );
  buffer buf_n6576( .i (n6249), .o (n6576) );
  buffer buf_n6577( .i (n6576), .o (n6577) );
  assign n6578 = n1970 & ~n6577 ;
  assign n6579 = n6575 | n6578 ;
  buffer buf_n6580( .i (n6579), .o (n6580) );
  buffer buf_n6581( .i (n6580), .o (n6581) );
  assign n6582 = n2570 & n6581 ;
  buffer buf_n3779( .i (n3778), .o (n3779) );
  buffer buf_n3780( .i (n3779), .o (n3780) );
  assign n6583 = n3780 & ~n5911 ;
  buffer buf_n83( .i (n82), .o (n83) );
  assign n6584 = n83 & n5911 ;
  assign n6585 = n6583 | n6584 ;
  buffer buf_n6586( .i (n6585), .o (n6586) );
  assign n6587 = ~n2570 & n6586 ;
  assign n6588 = n6582 | n6587 ;
  buffer buf_n6589( .i (n6588), .o (n6589) );
  assign n6590 = ~n44 & n6589 ;
  buffer buf_n6168( .i (n6167), .o (n6168) );
  assign n6591 = n44 & n6168 ;
  assign n6592 = n6590 | n6591 ;
  buffer buf_n6593( .i (n6592), .o (n6593) );
  assign n6594 = ~n3564 & n6593 ;
  buffer buf_n6595( .i (n6543), .o (n6595) );
  assign n6596 = n6218 & n6595 ;
  assign n6597 = n6184 & ~n6595 ;
  assign n6598 = n6596 | n6597 ;
  buffer buf_n6599( .i (n6598), .o (n6599) );
  buffer buf_n6600( .i (n6599), .o (n6600) );
  assign n6601 = n3564 & n6600 ;
  assign n6602 = n6594 | n6601 ;
  assign n6603 = ~n1865 & n6602 ;
  buffer buf_n6242( .i (n6241), .o (n6242) );
  assign n6604 = n6242 & n6595 ;
  assign n6605 = n6203 & ~n6595 ;
  assign n6606 = n6604 | n6605 ;
  buffer buf_n6607( .i (n6606), .o (n6607) );
  assign n6608 = ~n6223 & n6607 ;
  buffer buf_n6609( .i (n6542), .o (n6609) );
  assign n6610 = n6257 & ~n6609 ;
  assign n6611 = n6272 & n6609 ;
  assign n6612 = n6610 | n6611 ;
  buffer buf_n6613( .i (n6612), .o (n6613) );
  buffer buf_n6614( .i (n6613), .o (n6614) );
  assign n6615 = n6223 & n6614 ;
  assign n6616 = n6608 | n6615 ;
  buffer buf_n6617( .i (n6616), .o (n6617) );
  assign n6618 = n1865 & n6617 ;
  assign n6619 = n6603 | n6618 ;
  assign n6620 = n134 | n6619 ;
  assign n6621 = ~n6574 & n6620 ;
  buffer buf_n6622( .i (n6621), .o (n6622) );
  assign n6623 = n5927 & ~n6622 ;
  assign n6624 = n5884 & ~n6623 ;
  assign n6625 = n6019 & ~n6609 ;
  assign n6626 = n5962 & n6609 ;
  assign n6627 = n6625 | n6626 ;
  buffer buf_n6628( .i (n6627), .o (n6628) );
  assign n6629 = n6552 & n6628 ;
  buffer buf_n6630( .i (n6542), .o (n6630) );
  assign n6631 = n6034 & n6630 ;
  assign n6632 = n6000 & ~n6630 ;
  assign n6633 = n6631 | n6632 ;
  buffer buf_n6634( .i (n6633), .o (n6634) );
  assign n6635 = ~n6552 & n6634 ;
  assign n6636 = n6629 | n6635 ;
  buffer buf_n6637( .i (n6636), .o (n6637) );
  assign n6638 = ~n6557 & n6637 ;
  assign n6639 = n6150 | n6638 ;
  buffer buf_n6640( .i (n6639), .o (n6640) );
  buffer buf_n6641( .i (n133), .o (n6641) );
  assign n6642 = n6640 & ~n6641 ;
  assign n6643 = n5950 | n6642 ;
  buffer buf_n6644( .i (n6643), .o (n6644) );
  assign n6645 = n6101 & n6644 ;
  assign n6646 = n83 & ~n6055 ;
  buffer buf_n6647( .i (n6646), .o (n6647) );
  buffer buf_n3500( .i (n3499), .o (n3500) );
  buffer buf_n3501( .i (n3500), .o (n3501) );
  buffer buf_n3502( .i (n3501), .o (n3502) );
  buffer buf_n3503( .i (n3502), .o (n3503) );
  buffer buf_n3504( .i (n3503), .o (n3504) );
  buffer buf_n3505( .i (n3504), .o (n3505) );
  buffer buf_n3506( .i (n3505), .o (n3506) );
  buffer buf_n3507( .i (n3506), .o (n3507) );
  buffer buf_n3508( .i (n3507), .o (n3508) );
  buffer buf_n3509( .i (n3508), .o (n3509) );
  buffer buf_n3510( .i (n3509), .o (n3510) );
  buffer buf_n3511( .i (n3510), .o (n3511) );
  buffer buf_n3512( .i (n3511), .o (n3512) );
  buffer buf_n3513( .i (n3512), .o (n3513) );
  buffer buf_n3514( .i (n3513), .o (n3514) );
  buffer buf_n3515( .i (n3514), .o (n3515) );
  buffer buf_n3516( .i (n3515), .o (n3516) );
  buffer buf_n3517( .i (n3516), .o (n3517) );
  assign n6648 = n83 | n6066 ;
  assign n6649 = n3517 & n6648 ;
  assign n6650 = n6647 | n6649 ;
  buffer buf_n6651( .i (n6650), .o (n6651) );
  assign n6652 = n3517 & n6079 ;
  assign n6653 = n6647 & n6652 ;
  assign n6654 = n6088 | n6653 ;
  assign n6655 = n6651 & ~n6654 ;
  buffer buf_n6656( .i (n6655), .o (n6656) );
  buffer buf_n6657( .i (n6656), .o (n6657) );
  buffer buf_n6658( .i (n6657), .o (n6658) );
  assign n6659 = n5919 | n6658 ;
  buffer buf_n6660( .i (n6659), .o (n6660) );
  buffer buf_n6661( .i (n6660), .o (n6661) );
  buffer buf_n6662( .i (n6661), .o (n6662) );
  buffer buf_n6663( .i (n6662), .o (n6663) );
  buffer buf_n6664( .i (n6663), .o (n6664) );
  buffer buf_n6665( .i (n6664), .o (n6665) );
  buffer buf_n6666( .i (n6665), .o (n6666) );
  buffer buf_n6667( .i (n6666), .o (n6667) );
  assign n6668 = n6645 | n6667 ;
  assign n6669 = n6624 & n6668 ;
  assign n6670 = n6540 | n6669 ;
  buffer buf_n6671( .i (n6670), .o (n6671) );
  buffer buf_n6672( .i (n6671), .o (n6672) );
  buffer buf_n6673( .i (n6672), .o (n6673) );
  buffer buf_n6674( .i (n6673), .o (n6674) );
  buffer buf_n6675( .i (n6674), .o (n6675) );
  buffer buf_n6676( .i (n6675), .o (n6676) );
  buffer buf_n6677( .i (n6676), .o (n6677) );
  buffer buf_n6678( .i (n6677), .o (n6678) );
  buffer buf_n6679( .i (n6678), .o (n6679) );
  buffer buf_n6680( .i (n6679), .o (n6680) );
  buffer buf_n6681( .i (n6680), .o (n6681) );
  buffer buf_n6682( .i (n6681), .o (n6682) );
  buffer buf_n6683( .i (n6682), .o (n6683) );
  buffer buf_n6684( .i (n6683), .o (n6684) );
  buffer buf_n6685( .i (n6684), .o (n6685) );
  buffer buf_n6686( .i (n6685), .o (n6686) );
  buffer buf_n6687( .i (n6686), .o (n6687) );
  buffer buf_n6688( .i (n6687), .o (n6688) );
  buffer buf_n6689( .i (n6688), .o (n6689) );
  buffer buf_n6690( .i (n6689), .o (n6690) );
  buffer buf_n6691( .i (n6690), .o (n6691) );
  buffer buf_n6692( .i (n6691), .o (n6692) );
  buffer buf_n6693( .i (n6692), .o (n6693) );
  buffer buf_n6694( .i (n6693), .o (n6694) );
  buffer buf_n6695( .i (n6694), .o (n6695) );
  buffer buf_n6696( .i (n6695), .o (n6696) );
  buffer buf_n6697( .i (n6696), .o (n6697) );
  buffer buf_n6698( .i (n6697), .o (n6698) );
  buffer buf_n6699( .i (n6698), .o (n6699) );
  buffer buf_n6700( .i (n6699), .o (n6700) );
  buffer buf_n6701( .i (n6700), .o (n6701) );
  buffer buf_n6702( .i (n6701), .o (n6702) );
  buffer buf_n6703( .i (n6702), .o (n6703) );
  buffer buf_n6704( .i (n6703), .o (n6704) );
  buffer buf_n6705( .i (n6704), .o (n6705) );
  buffer buf_n6706( .i (n6705), .o (n6706) );
  buffer buf_n6707( .i (n6706), .o (n6707) );
  buffer buf_n6708( .i (n6707), .o (n6708) );
  buffer buf_n6709( .i (n6708), .o (n6709) );
  buffer buf_n6710( .i (n6709), .o (n6710) );
  buffer buf_n6711( .i (n6710), .o (n6711) );
  buffer buf_n6712( .i (n6711), .o (n6712) );
  buffer buf_n6713( .i (n6712), .o (n6713) );
  buffer buf_n6714( .i (n6713), .o (n6714) );
  buffer buf_n6715( .i (n6714), .o (n6715) );
  buffer buf_n6716( .i (n6715), .o (n6716) );
  buffer buf_n6717( .i (n6716), .o (n6717) );
  buffer buf_n6718( .i (n6717), .o (n6718) );
  buffer buf_n6719( .i (n6718), .o (n6719) );
  buffer buf_n6720( .i (n6719), .o (n6720) );
  buffer buf_n6721( .i (n6720), .o (n6721) );
  buffer buf_n6722( .i (n6721), .o (n6722) );
  buffer buf_n6723( .i (n6722), .o (n6723) );
  buffer buf_n6724( .i (n6723), .o (n6724) );
  buffer buf_n6725( .i (n6724), .o (n6725) );
  buffer buf_n6726( .i (n6725), .o (n6726) );
  buffer buf_n6727( .i (n6726), .o (n6727) );
  buffer buf_n6728( .i (n6727), .o (n6728) );
  buffer buf_n6729( .i (n6728), .o (n6729) );
  buffer buf_n6730( .i (n6729), .o (n6730) );
  buffer buf_n6731( .i (n6730), .o (n6731) );
  buffer buf_n6732( .i (n6731), .o (n6732) );
  buffer buf_n6733( .i (n6732), .o (n6733) );
  buffer buf_n6734( .i (n6733), .o (n6734) );
  buffer buf_n6735( .i (n6734), .o (n6735) );
  buffer buf_n6736( .i (n6735), .o (n6736) );
  buffer buf_n6737( .i (n6736), .o (n6737) );
  buffer buf_n6738( .i (n6737), .o (n6738) );
  buffer buf_n6739( .i (n6738), .o (n6739) );
  buffer buf_n6740( .i (n6739), .o (n6740) );
  buffer buf_n6741( .i (n6740), .o (n6741) );
  buffer buf_n6742( .i (n6741), .o (n6742) );
  buffer buf_n6743( .i (n6742), .o (n6743) );
  buffer buf_n6744( .i (n6743), .o (n6744) );
  buffer buf_n6745( .i (n6744), .o (n6745) );
  buffer buf_n6746( .i (n6745), .o (n6746) );
  buffer buf_n6747( .i (n6746), .o (n6747) );
  buffer buf_n6748( .i (n6747), .o (n6748) );
  buffer buf_n6749( .i (n6748), .o (n6749) );
  buffer buf_n6750( .i (n6749), .o (n6750) );
  buffer buf_n6751( .i (n6750), .o (n6751) );
  buffer buf_n6752( .i (n6751), .o (n6752) );
  buffer buf_n6753( .i (n6752), .o (n6753) );
  buffer buf_n6754( .i (n6753), .o (n6754) );
  buffer buf_n6755( .i (n6754), .o (n6755) );
  buffer buf_n6756( .i (n6755), .o (n6756) );
  buffer buf_n6757( .i (n6756), .o (n6757) );
  buffer buf_n6758( .i (n6757), .o (n6758) );
  buffer buf_n6759( .i (n6758), .o (n6759) );
  buffer buf_n6760( .i (n6759), .o (n6760) );
  buffer buf_n6761( .i (n6760), .o (n6761) );
  buffer buf_n6762( .i (n6761), .o (n6762) );
  buffer buf_n6763( .i (n6762), .o (n6763) );
  buffer buf_n6764( .i (n6763), .o (n6764) );
  buffer buf_n6765( .i (n6764), .o (n6765) );
  buffer buf_n6766( .i (n6765), .o (n6766) );
  buffer buf_n6767( .i (n6766), .o (n6767) );
  buffer buf_n6768( .i (n6767), .o (n6768) );
  buffer buf_n6769( .i (n6768), .o (n6769) );
  buffer buf_n6770( .i (n6769), .o (n6770) );
  buffer buf_n6771( .i (n6770), .o (n6771) );
  buffer buf_n6772( .i (n6771), .o (n6772) );
  buffer buf_n6773( .i (n6772), .o (n6773) );
  buffer buf_n6774( .i (n6773), .o (n6774) );
  buffer buf_n6775( .i (n6774), .o (n6775) );
  buffer buf_n6776( .i (n6775), .o (n6776) );
  buffer buf_n6777( .i (n6776), .o (n6777) );
  buffer buf_n6778( .i (n6777), .o (n6778) );
  buffer buf_n6779( .i (n6778), .o (n6779) );
  buffer buf_n6780( .i (n6779), .o (n6780) );
  buffer buf_n6781( .i (n6780), .o (n6781) );
  buffer buf_n6782( .i (n6781), .o (n6782) );
  buffer buf_n2492( .i (n2491), .o (n2492) );
  buffer buf_n2493( .i (n2492), .o (n2493) );
  buffer buf_n2494( .i (n2493), .o (n2494) );
  buffer buf_n2495( .i (n2494), .o (n2495) );
  buffer buf_n2496( .i (n2495), .o (n2496) );
  buffer buf_n2497( .i (n2496), .o (n2497) );
  buffer buf_n2498( .i (n2497), .o (n2498) );
  buffer buf_n2499( .i (n2498), .o (n2499) );
  buffer buf_n2500( .i (n2499), .o (n2500) );
  buffer buf_n2501( .i (n2500), .o (n2501) );
  buffer buf_n2502( .i (n2501), .o (n2502) );
  buffer buf_n2503( .i (n2502), .o (n2503) );
  buffer buf_n2504( .i (n2503), .o (n2504) );
  buffer buf_n2505( .i (n2504), .o (n2505) );
  buffer buf_n2506( .i (n2505), .o (n2506) );
  buffer buf_n2507( .i (n2506), .o (n2507) );
  buffer buf_n2508( .i (n2507), .o (n2508) );
  buffer buf_n2509( .i (n2508), .o (n2509) );
  buffer buf_n2510( .i (n2509), .o (n2510) );
  buffer buf_n2511( .i (n2510), .o (n2511) );
  buffer buf_n2512( .i (n2511), .o (n2512) );
  buffer buf_n2513( .i (n2512), .o (n2513) );
  buffer buf_n2514( .i (n2513), .o (n2514) );
  buffer buf_n2515( .i (n2514), .o (n2515) );
  buffer buf_n2516( .i (n2515), .o (n2516) );
  buffer buf_n2517( .i (n2516), .o (n2517) );
  buffer buf_n2518( .i (n2517), .o (n2518) );
  buffer buf_n2519( .i (n2518), .o (n2519) );
  buffer buf_n2520( .i (n2519), .o (n2520) );
  buffer buf_n2521( .i (n2520), .o (n2521) );
  buffer buf_n2522( .i (n2521), .o (n2522) );
  buffer buf_n2523( .i (n2522), .o (n2523) );
  buffer buf_n2524( .i (n2523), .o (n2524) );
  buffer buf_n2525( .i (n2524), .o (n2525) );
  buffer buf_n2526( .i (n2525), .o (n2526) );
  buffer buf_n2527( .i (n2526), .o (n2527) );
  buffer buf_n2528( .i (n2527), .o (n2528) );
  buffer buf_n2529( .i (n2528), .o (n2529) );
  buffer buf_n2722( .i (x46), .o (n2722) );
  buffer buf_n2723( .i (n2722), .o (n2723) );
  buffer buf_n2724( .i (n2723), .o (n2724) );
  buffer buf_n2725( .i (n2724), .o (n2725) );
  buffer buf_n2726( .i (n2725), .o (n2726) );
  buffer buf_n2727( .i (n2726), .o (n2727) );
  buffer buf_n2728( .i (n2727), .o (n2728) );
  buffer buf_n2729( .i (n2728), .o (n2729) );
  buffer buf_n2730( .i (n2729), .o (n2730) );
  buffer buf_n2731( .i (n2730), .o (n2731) );
  buffer buf_n2732( .i (n2731), .o (n2732) );
  buffer buf_n2733( .i (n2732), .o (n2733) );
  buffer buf_n2734( .i (n2733), .o (n2734) );
  buffer buf_n2735( .i (n2734), .o (n2735) );
  buffer buf_n2736( .i (n2735), .o (n2736) );
  buffer buf_n2737( .i (n2736), .o (n2737) );
  buffer buf_n2738( .i (n2737), .o (n2738) );
  buffer buf_n2739( .i (n2738), .o (n2739) );
  buffer buf_n2740( .i (n2739), .o (n2740) );
  buffer buf_n2741( .i (n2740), .o (n2741) );
  buffer buf_n2742( .i (n2741), .o (n2742) );
  buffer buf_n2743( .i (n2742), .o (n2743) );
  buffer buf_n2744( .i (n2743), .o (n2744) );
  buffer buf_n2745( .i (n2744), .o (n2745) );
  buffer buf_n2746( .i (n2745), .o (n2746) );
  buffer buf_n2747( .i (n2746), .o (n2747) );
  buffer buf_n2748( .i (n2747), .o (n2748) );
  buffer buf_n2749( .i (n2748), .o (n2749) );
  buffer buf_n2750( .i (n2749), .o (n2750) );
  buffer buf_n2751( .i (n2750), .o (n2751) );
  buffer buf_n2752( .i (n2751), .o (n2752) );
  buffer buf_n2753( .i (n2752), .o (n2753) );
  buffer buf_n2754( .i (n2753), .o (n2754) );
  buffer buf_n2755( .i (n2754), .o (n2755) );
  buffer buf_n2756( .i (n2755), .o (n2756) );
  buffer buf_n2757( .i (n2756), .o (n2757) );
  buffer buf_n2758( .i (n2757), .o (n2758) );
  buffer buf_n2759( .i (n2758), .o (n2759) );
  buffer buf_n2760( .i (n2759), .o (n2760) );
  buffer buf_n2761( .i (n2760), .o (n2761) );
  buffer buf_n2762( .i (n2761), .o (n2762) );
  buffer buf_n2763( .i (n2762), .o (n2763) );
  buffer buf_n2764( .i (n2763), .o (n2764) );
  buffer buf_n2765( .i (n2764), .o (n2765) );
  buffer buf_n2766( .i (n2765), .o (n2766) );
  buffer buf_n2767( .i (n2766), .o (n2767) );
  buffer buf_n2768( .i (n2767), .o (n2768) );
  buffer buf_n2769( .i (n2768), .o (n2769) );
  buffer buf_n2770( .i (n2769), .o (n2770) );
  buffer buf_n2771( .i (n2770), .o (n2771) );
  buffer buf_n2772( .i (n2771), .o (n2772) );
  buffer buf_n2773( .i (n2772), .o (n2773) );
  buffer buf_n2774( .i (n2773), .o (n2774) );
  buffer buf_n2775( .i (n2774), .o (n2775) );
  buffer buf_n2776( .i (n2775), .o (n2776) );
  buffer buf_n2777( .i (n2776), .o (n2777) );
  buffer buf_n2778( .i (n2777), .o (n2778) );
  buffer buf_n2779( .i (n2778), .o (n2779) );
  buffer buf_n2780( .i (n2779), .o (n2780) );
  buffer buf_n2781( .i (n2780), .o (n2781) );
  buffer buf_n2782( .i (n2781), .o (n2782) );
  buffer buf_n2783( .i (n2782), .o (n2783) );
  buffer buf_n2784( .i (n2783), .o (n2784) );
  buffer buf_n2785( .i (n2784), .o (n2785) );
  buffer buf_n2786( .i (n2785), .o (n2786) );
  buffer buf_n2787( .i (n2786), .o (n2787) );
  buffer buf_n2788( .i (n2787), .o (n2788) );
  buffer buf_n2789( .i (n2788), .o (n2789) );
  buffer buf_n2790( .i (n2789), .o (n2790) );
  buffer buf_n2791( .i (n2790), .o (n2791) );
  buffer buf_n3164( .i (x52), .o (n3164) );
  buffer buf_n3165( .i (n3164), .o (n3165) );
  buffer buf_n3166( .i (n3165), .o (n3166) );
  buffer buf_n3167( .i (n3166), .o (n3167) );
  buffer buf_n3168( .i (n3167), .o (n3168) );
  buffer buf_n3169( .i (n3168), .o (n3169) );
  buffer buf_n3170( .i (n3169), .o (n3170) );
  buffer buf_n3171( .i (n3170), .o (n3171) );
  buffer buf_n3172( .i (n3171), .o (n3172) );
  buffer buf_n3173( .i (n3172), .o (n3173) );
  buffer buf_n3174( .i (n3173), .o (n3174) );
  buffer buf_n3175( .i (n3174), .o (n3175) );
  buffer buf_n3176( .i (n3175), .o (n3176) );
  buffer buf_n3177( .i (n3176), .o (n3177) );
  buffer buf_n3178( .i (n3177), .o (n3178) );
  buffer buf_n3179( .i (n3178), .o (n3179) );
  buffer buf_n3180( .i (n3179), .o (n3180) );
  buffer buf_n3181( .i (n3180), .o (n3181) );
  buffer buf_n3182( .i (n3181), .o (n3182) );
  buffer buf_n3183( .i (n3182), .o (n3183) );
  buffer buf_n3184( .i (n3183), .o (n3184) );
  buffer buf_n3185( .i (n3184), .o (n3185) );
  buffer buf_n3186( .i (n3185), .o (n3186) );
  buffer buf_n3187( .i (n3186), .o (n3187) );
  buffer buf_n3188( .i (n3187), .o (n3188) );
  buffer buf_n3189( .i (n3188), .o (n3189) );
  buffer buf_n3190( .i (n3189), .o (n3190) );
  buffer buf_n3191( .i (n3190), .o (n3191) );
  buffer buf_n3192( .i (n3191), .o (n3192) );
  buffer buf_n3193( .i (n3192), .o (n3193) );
  buffer buf_n3194( .i (n3193), .o (n3194) );
  buffer buf_n3195( .i (n3194), .o (n3195) );
  buffer buf_n3196( .i (n3195), .o (n3196) );
  buffer buf_n3197( .i (n3196), .o (n3197) );
  buffer buf_n3198( .i (n3197), .o (n3198) );
  buffer buf_n3199( .i (n3198), .o (n3199) );
  buffer buf_n3200( .i (n3199), .o (n3200) );
  buffer buf_n3201( .i (n3200), .o (n3201) );
  buffer buf_n3202( .i (n3201), .o (n3202) );
  buffer buf_n3203( .i (n3202), .o (n3203) );
  buffer buf_n3204( .i (n3203), .o (n3204) );
  buffer buf_n3205( .i (n3204), .o (n3205) );
  buffer buf_n3206( .i (n3205), .o (n3206) );
  buffer buf_n3207( .i (n3206), .o (n3207) );
  buffer buf_n3208( .i (n3207), .o (n3208) );
  buffer buf_n3209( .i (n3208), .o (n3209) );
  buffer buf_n3210( .i (n3209), .o (n3210) );
  buffer buf_n3211( .i (n3210), .o (n3211) );
  buffer buf_n3212( .i (n3211), .o (n3212) );
  buffer buf_n3213( .i (n3212), .o (n3213) );
  buffer buf_n3214( .i (n3213), .o (n3214) );
  buffer buf_n3215( .i (n3214), .o (n3215) );
  buffer buf_n3216( .i (n3215), .o (n3216) );
  buffer buf_n3217( .i (n3216), .o (n3217) );
  buffer buf_n3218( .i (n3217), .o (n3218) );
  buffer buf_n3219( .i (n3218), .o (n3219) );
  buffer buf_n3220( .i (n3219), .o (n3220) );
  buffer buf_n3221( .i (n3220), .o (n3221) );
  buffer buf_n3222( .i (n3221), .o (n3222) );
  buffer buf_n3223( .i (n3222), .o (n3223) );
  buffer buf_n3224( .i (n3223), .o (n3224) );
  buffer buf_n3225( .i (n3224), .o (n3225) );
  buffer buf_n3226( .i (n3225), .o (n3226) );
  buffer buf_n3227( .i (n3226), .o (n3227) );
  buffer buf_n3228( .i (n3227), .o (n3228) );
  buffer buf_n3229( .i (n3228), .o (n3229) );
  buffer buf_n3230( .i (n3229), .o (n3230) );
  buffer buf_n3915( .i (n3914), .o (n3915) );
  buffer buf_n3916( .i (n3915), .o (n3916) );
  buffer buf_n3917( .i (n3916), .o (n3917) );
  buffer buf_n3918( .i (n3917), .o (n3918) );
  buffer buf_n3919( .i (n3918), .o (n3919) );
  buffer buf_n3920( .i (n3919), .o (n3920) );
  buffer buf_n3921( .i (n3920), .o (n3921) );
  buffer buf_n3922( .i (n3921), .o (n3922) );
  buffer buf_n3923( .i (n3922), .o (n3923) );
  buffer buf_n3924( .i (n3923), .o (n3924) );
  buffer buf_n3925( .i (n3924), .o (n3925) );
  buffer buf_n3926( .i (n3925), .o (n3926) );
  buffer buf_n3927( .i (n3926), .o (n3927) );
  buffer buf_n3928( .i (n3927), .o (n3928) );
  buffer buf_n3929( .i (n3928), .o (n3929) );
  buffer buf_n3930( .i (n3929), .o (n3930) );
  buffer buf_n3931( .i (n3930), .o (n3931) );
  buffer buf_n3932( .i (n3931), .o (n3932) );
  buffer buf_n3933( .i (n3932), .o (n3933) );
  buffer buf_n3934( .i (n3933), .o (n3934) );
  assign n6783 = n3230 & n3934 ;
  buffer buf_n2657( .i (x45), .o (n2657) );
  buffer buf_n2658( .i (n2657), .o (n2658) );
  buffer buf_n2659( .i (n2658), .o (n2659) );
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2660), .o (n2661) );
  buffer buf_n2662( .i (n2661), .o (n2662) );
  buffer buf_n2663( .i (n2662), .o (n2663) );
  buffer buf_n2664( .i (n2663), .o (n2664) );
  buffer buf_n2665( .i (n2664), .o (n2665) );
  buffer buf_n2666( .i (n2665), .o (n2666) );
  buffer buf_n2667( .i (n2666), .o (n2667) );
  buffer buf_n2668( .i (n2667), .o (n2668) );
  buffer buf_n2669( .i (n2668), .o (n2669) );
  buffer buf_n2670( .i (n2669), .o (n2670) );
  buffer buf_n2671( .i (n2670), .o (n2671) );
  buffer buf_n2672( .i (n2671), .o (n2672) );
  buffer buf_n2673( .i (n2672), .o (n2673) );
  buffer buf_n2674( .i (n2673), .o (n2674) );
  buffer buf_n2675( .i (n2674), .o (n2675) );
  buffer buf_n2676( .i (n2675), .o (n2676) );
  buffer buf_n2677( .i (n2676), .o (n2677) );
  buffer buf_n2678( .i (n2677), .o (n2678) );
  buffer buf_n2679( .i (n2678), .o (n2679) );
  buffer buf_n2680( .i (n2679), .o (n2680) );
  buffer buf_n2681( .i (n2680), .o (n2681) );
  buffer buf_n2682( .i (n2681), .o (n2682) );
  buffer buf_n2683( .i (n2682), .o (n2683) );
  buffer buf_n2684( .i (n2683), .o (n2684) );
  buffer buf_n2685( .i (n2684), .o (n2685) );
  buffer buf_n2686( .i (n2685), .o (n2686) );
  buffer buf_n2687( .i (n2686), .o (n2687) );
  buffer buf_n2688( .i (n2687), .o (n2688) );
  buffer buf_n2689( .i (n2688), .o (n2689) );
  buffer buf_n2690( .i (n2689), .o (n2690) );
  buffer buf_n2691( .i (n2690), .o (n2691) );
  buffer buf_n2692( .i (n2691), .o (n2692) );
  buffer buf_n2693( .i (n2692), .o (n2693) );
  buffer buf_n2694( .i (n2693), .o (n2694) );
  buffer buf_n2695( .i (n2694), .o (n2695) );
  buffer buf_n2696( .i (n2695), .o (n2696) );
  buffer buf_n2697( .i (n2696), .o (n2697) );
  buffer buf_n2698( .i (n2697), .o (n2698) );
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n2700( .i (n2699), .o (n2700) );
  buffer buf_n2701( .i (n2700), .o (n2701) );
  buffer buf_n2702( .i (n2701), .o (n2702) );
  buffer buf_n2703( .i (n2702), .o (n2703) );
  buffer buf_n2704( .i (n2703), .o (n2704) );
  buffer buf_n2705( .i (n2704), .o (n2705) );
  buffer buf_n2706( .i (n2705), .o (n2706) );
  buffer buf_n2707( .i (n2706), .o (n2707) );
  buffer buf_n2708( .i (n2707), .o (n2708) );
  buffer buf_n2709( .i (n2708), .o (n2709) );
  buffer buf_n2710( .i (n2709), .o (n2710) );
  buffer buf_n2711( .i (n2710), .o (n2711) );
  buffer buf_n2712( .i (n2711), .o (n2712) );
  buffer buf_n2713( .i (n2712), .o (n2713) );
  buffer buf_n2714( .i (n2713), .o (n2714) );
  buffer buf_n2715( .i (n2714), .o (n2715) );
  buffer buf_n2716( .i (n2715), .o (n2716) );
  buffer buf_n2717( .i (n2716), .o (n2717) );
  buffer buf_n2718( .i (n2717), .o (n2718) );
  buffer buf_n2719( .i (n2718), .o (n2719) );
  buffer buf_n2720( .i (n2719), .o (n2720) );
  buffer buf_n912( .i (x17), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n852( .i (x16), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n233( .i (x5), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n973( .i (x18), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n3110( .i (x51), .o (n3110) );
  buffer buf_n3111( .i (n3110), .o (n3111) );
  buffer buf_n3112( .i (n3111), .o (n3112) );
  buffer buf_n3113( .i (n3112), .o (n3113) );
  buffer buf_n3114( .i (n3113), .o (n3114) );
  buffer buf_n3115( .i (n3114), .o (n3115) );
  buffer buf_n3116( .i (n3115), .o (n3116) );
  buffer buf_n3117( .i (n3116), .o (n3117) );
  buffer buf_n3118( .i (n3117), .o (n3118) );
  buffer buf_n3119( .i (n3118), .o (n3119) );
  buffer buf_n3120( .i (n3119), .o (n3120) );
  buffer buf_n3121( .i (n3120), .o (n3121) );
  buffer buf_n3122( .i (n3121), .o (n3122) );
  buffer buf_n3123( .i (n3122), .o (n3123) );
  buffer buf_n3124( .i (n3123), .o (n3124) );
  buffer buf_n3125( .i (n3124), .o (n3125) );
  buffer buf_n3126( .i (n3125), .o (n3126) );
  buffer buf_n3127( .i (n3126), .o (n3127) );
  buffer buf_n3128( .i (n3127), .o (n3128) );
  buffer buf_n3129( .i (n3128), .o (n3129) );
  buffer buf_n3130( .i (n3129), .o (n3130) );
  buffer buf_n3131( .i (n3130), .o (n3131) );
  buffer buf_n3132( .i (n3131), .o (n3132) );
  buffer buf_n3133( .i (n3132), .o (n3133) );
  buffer buf_n3134( .i (n3133), .o (n3134) );
  buffer buf_n3135( .i (n3134), .o (n3135) );
  buffer buf_n3136( .i (n3135), .o (n3136) );
  buffer buf_n3137( .i (n3136), .o (n3137) );
  buffer buf_n3138( .i (n3137), .o (n3138) );
  buffer buf_n3139( .i (n3138), .o (n3139) );
  buffer buf_n3140( .i (n3139), .o (n3140) );
  buffer buf_n3141( .i (n3140), .o (n3141) );
  buffer buf_n3142( .i (n3141), .o (n3142) );
  buffer buf_n3143( .i (n3142), .o (n3143) );
  buffer buf_n3144( .i (n3143), .o (n3144) );
  buffer buf_n3145( .i (n3144), .o (n3145) );
  buffer buf_n3146( .i (n3145), .o (n3146) );
  buffer buf_n3147( .i (n3146), .o (n3147) );
  buffer buf_n3148( .i (n3147), .o (n3148) );
  buffer buf_n3149( .i (n3148), .o (n3149) );
  buffer buf_n3150( .i (n3149), .o (n3150) );
  buffer buf_n3151( .i (n3150), .o (n3151) );
  buffer buf_n3152( .i (n3151), .o (n3152) );
  buffer buf_n3153( .i (n3152), .o (n3153) );
  buffer buf_n3154( .i (n3153), .o (n3154) );
  buffer buf_n3155( .i (n3154), .o (n3155) );
  buffer buf_n3156( .i (n3155), .o (n3156) );
  buffer buf_n3157( .i (n3156), .o (n3157) );
  buffer buf_n3158( .i (n3157), .o (n3158) );
  buffer buf_n3159( .i (n3158), .o (n3159) );
  buffer buf_n3160( .i (n3159), .o (n3160) );
  buffer buf_n1592( .i (x27), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n1633( .i (n1632), .o (n1633) );
  buffer buf_n1634( .i (n1633), .o (n1634) );
  buffer buf_n1635( .i (n1634), .o (n1635) );
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n1637( .i (n1636), .o (n1637) );
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  assign n6784 = n1437 | n5477 ;
  buffer buf_n6785( .i (n6784), .o (n6785) );
  assign n6786 = n1640 | n6785 ;
  buffer buf_n6787( .i (n6786), .o (n6787) );
  assign n6788 = n3160 | n6787 ;
  buffer buf_n6789( .i (n6788), .o (n6789) );
  assign n6790 = n1025 | n6789 ;
  buffer buf_n6791( .i (n6790), .o (n6791) );
  assign n6792 = n287 | n6791 ;
  buffer buf_n6793( .i (n6792), .o (n6793) );
  assign n6794 = n908 | n6793 ;
  assign n6795 = n3925 & n6794 ;
  buffer buf_n6796( .i (n6795), .o (n6796) );
  assign n6797 = n971 | n6796 ;
  buffer buf_n6798( .i (n6797), .o (n6798) );
  assign n6799 = n3929 & n6798 ;
  buffer buf_n6800( .i (n6799), .o (n6800) );
  assign n6801 = n2720 | n6800 ;
  buffer buf_n6802( .i (n6801), .o (n6802) );
  assign n6803 = n3933 & n6802 ;
  buffer buf_n6804( .i (n6803), .o (n6804) );
  assign n6805 = n6783 | n6804 ;
  buffer buf_n6806( .i (n6805), .o (n6806) );
  assign n6807 = ~n2791 & n6806 ;
  assign n6808 = n2791 & ~n6806 ;
  assign n6809 = n6807 | n6808 ;
  buffer buf_n6810( .i (n6809), .o (n6810) );
  assign n6811 = n2529 & n6810 ;
  buffer buf_n6812( .i (n6811), .o (n6812) );
  buffer buf_n6813( .i (n6812), .o (n6813) );
  buffer buf_n6814( .i (n6813), .o (n6814) );
  buffer buf_n6815( .i (n6814), .o (n6815) );
  buffer buf_n6816( .i (n6815), .o (n6816) );
  buffer buf_n6817( .i (n6816), .o (n6817) );
  buffer buf_n6818( .i (n6817), .o (n6818) );
  buffer buf_n6819( .i (n6818), .o (n6819) );
  buffer buf_n6820( .i (n6819), .o (n6820) );
  buffer buf_n6821( .i (n6820), .o (n6821) );
  buffer buf_n6822( .i (n6821), .o (n6822) );
  buffer buf_n6823( .i (n6822), .o (n6823) );
  buffer buf_n6824( .i (n6823), .o (n6824) );
  buffer buf_n6825( .i (n6824), .o (n6825) );
  buffer buf_n6826( .i (n6825), .o (n6826) );
  buffer buf_n6827( .i (n6826), .o (n6827) );
  buffer buf_n6828( .i (n6827), .o (n6828) );
  buffer buf_n6829( .i (n6828), .o (n6829) );
  buffer buf_n6830( .i (n6829), .o (n6830) );
  buffer buf_n6831( .i (n6830), .o (n6831) );
  buffer buf_n6832( .i (n6831), .o (n6832) );
  buffer buf_n6833( .i (n6832), .o (n6833) );
  buffer buf_n6834( .i (n6833), .o (n6834) );
  buffer buf_n6835( .i (n6834), .o (n6835) );
  buffer buf_n6836( .i (n6835), .o (n6836) );
  buffer buf_n6837( .i (n6836), .o (n6837) );
  buffer buf_n6838( .i (n6837), .o (n6838) );
  buffer buf_n6839( .i (n6838), .o (n6839) );
  buffer buf_n6840( .i (n6839), .o (n6840) );
  buffer buf_n6841( .i (n6840), .o (n6841) );
  buffer buf_n6842( .i (n6841), .o (n6842) );
  buffer buf_n6843( .i (n6842), .o (n6843) );
  buffer buf_n6844( .i (n6843), .o (n6844) );
  buffer buf_n6845( .i (n6844), .o (n6845) );
  buffer buf_n6846( .i (n6845), .o (n6846) );
  buffer buf_n6847( .i (n6846), .o (n6847) );
  buffer buf_n6848( .i (n6847), .o (n6848) );
  buffer buf_n6849( .i (n6848), .o (n6849) );
  buffer buf_n6850( .i (n6849), .o (n6850) );
  buffer buf_n6851( .i (n6850), .o (n6851) );
  buffer buf_n6852( .i (n6851), .o (n6852) );
  buffer buf_n6853( .i (n6852), .o (n6853) );
  buffer buf_n6854( .i (n6853), .o (n6854) );
  buffer buf_n6855( .i (n6854), .o (n6855) );
  buffer buf_n6856( .i (n6855), .o (n6856) );
  buffer buf_n6857( .i (n6856), .o (n6857) );
  buffer buf_n6858( .i (n6857), .o (n6858) );
  buffer buf_n6859( .i (n6858), .o (n6859) );
  buffer buf_n6860( .i (n6859), .o (n6860) );
  buffer buf_n6861( .i (n6860), .o (n6861) );
  buffer buf_n6862( .i (n6861), .o (n6862) );
  buffer buf_n6863( .i (n6862), .o (n6863) );
  buffer buf_n6864( .i (n6863), .o (n6864) );
  buffer buf_n6865( .i (n6864), .o (n6865) );
  buffer buf_n6866( .i (n6865), .o (n6866) );
  buffer buf_n6867( .i (n6866), .o (n6867) );
  buffer buf_n6868( .i (n6867), .o (n6868) );
  buffer buf_n6869( .i (n6868), .o (n6869) );
  buffer buf_n6870( .i (n6869), .o (n6870) );
  buffer buf_n6871( .i (n6870), .o (n6871) );
  buffer buf_n6872( .i (n6871), .o (n6872) );
  buffer buf_n6873( .i (n6872), .o (n6873) );
  buffer buf_n6874( .i (n6873), .o (n6874) );
  buffer buf_n6875( .i (n6874), .o (n6875) );
  buffer buf_n6876( .i (n6875), .o (n6876) );
  buffer buf_n6877( .i (n6876), .o (n6877) );
  buffer buf_n6878( .i (n6877), .o (n6878) );
  buffer buf_n6879( .i (n6878), .o (n6879) );
  buffer buf_n6880( .i (n6879), .o (n6880) );
  buffer buf_n6881( .i (n6880), .o (n6881) );
  buffer buf_n6882( .i (n6881), .o (n6882) );
  buffer buf_n6883( .i (n6882), .o (n6883) );
  buffer buf_n6884( .i (n6883), .o (n6884) );
  buffer buf_n6885( .i (n6884), .o (n6885) );
  buffer buf_n6886( .i (n6885), .o (n6886) );
  buffer buf_n6887( .i (n6886), .o (n6887) );
  buffer buf_n6888( .i (n6887), .o (n6888) );
  buffer buf_n6889( .i (n6888), .o (n6889) );
  buffer buf_n6890( .i (n6889), .o (n6890) );
  buffer buf_n6891( .i (n6890), .o (n6891) );
  buffer buf_n6892( .i (n6891), .o (n6892) );
  buffer buf_n6893( .i (n6892), .o (n6893) );
  buffer buf_n6894( .i (n6893), .o (n6894) );
  buffer buf_n6895( .i (n6894), .o (n6895) );
  buffer buf_n6896( .i (n6895), .o (n6896) );
  buffer buf_n6897( .i (n6896), .o (n6897) );
  buffer buf_n6898( .i (n6897), .o (n6898) );
  buffer buf_n3315( .i (n3314), .o (n3315) );
  buffer buf_n3316( .i (n3315), .o (n3316) );
  buffer buf_n3317( .i (n3316), .o (n3317) );
  buffer buf_n3318( .i (n3317), .o (n3318) );
  buffer buf_n3319( .i (n3318), .o (n3319) );
  buffer buf_n3320( .i (n3319), .o (n3320) );
  buffer buf_n3321( .i (n3320), .o (n3321) );
  buffer buf_n3322( .i (n3321), .o (n3322) );
  buffer buf_n3323( .i (n3322), .o (n3323) );
  buffer buf_n3324( .i (n3323), .o (n3324) );
  buffer buf_n3325( .i (n3324), .o (n3325) );
  buffer buf_n3326( .i (n3325), .o (n3326) );
  buffer buf_n3327( .i (n3326), .o (n3327) );
  buffer buf_n3328( .i (n3327), .o (n3328) );
  buffer buf_n3329( .i (n3328), .o (n3329) );
  buffer buf_n3330( .i (n3329), .o (n3330) );
  buffer buf_n3331( .i (n3330), .o (n3331) );
  buffer buf_n3332( .i (n3331), .o (n3332) );
  buffer buf_n3333( .i (n3332), .o (n3333) );
  buffer buf_n3334( .i (n3333), .o (n3334) );
  buffer buf_n3335( .i (n3334), .o (n3335) );
  buffer buf_n3336( .i (n3335), .o (n3336) );
  buffer buf_n3337( .i (n3336), .o (n3337) );
  buffer buf_n3338( .i (n3337), .o (n3338) );
  buffer buf_n3339( .i (n3338), .o (n3339) );
  buffer buf_n3340( .i (n3339), .o (n3340) );
  buffer buf_n3341( .i (n3340), .o (n3341) );
  buffer buf_n3342( .i (n3341), .o (n3342) );
  buffer buf_n3343( .i (n3342), .o (n3343) );
  buffer buf_n3344( .i (n3343), .o (n3344) );
  buffer buf_n3345( .i (n3344), .o (n3345) );
  buffer buf_n3346( .i (n3345), .o (n3346) );
  buffer buf_n3347( .i (n3346), .o (n3347) );
  buffer buf_n3348( .i (n3347), .o (n3348) );
  buffer buf_n3349( .i (n3348), .o (n3349) );
  buffer buf_n3350( .i (n3349), .o (n3350) );
  buffer buf_n3351( .i (n3350), .o (n3351) );
  buffer buf_n3352( .i (n3351), .o (n3352) );
  buffer buf_n3353( .i (n3352), .o (n3353) );
  buffer buf_n3354( .i (n3353), .o (n3354) );
  buffer buf_n3355( .i (n3354), .o (n3355) );
  buffer buf_n3356( .i (n3355), .o (n3356) );
  buffer buf_n3357( .i (n3356), .o (n3357) );
  buffer buf_n3358( .i (n3357), .o (n3358) );
  buffer buf_n3359( .i (n3358), .o (n3359) );
  buffer buf_n3360( .i (n3359), .o (n3360) );
  buffer buf_n3361( .i (n3360), .o (n3361) );
  buffer buf_n3362( .i (n3361), .o (n3362) );
  buffer buf_n3363( .i (n3362), .o (n3363) );
  buffer buf_n3364( .i (n3363), .o (n3364) );
  buffer buf_n3365( .i (n3364), .o (n3365) );
  buffer buf_n3366( .i (n3365), .o (n3366) );
  buffer buf_n3367( .i (n3366), .o (n3367) );
  buffer buf_n3368( .i (n3367), .o (n3368) );
  buffer buf_n3369( .i (n3368), .o (n3369) );
  buffer buf_n3370( .i (n3369), .o (n3370) );
  buffer buf_n3371( .i (n3370), .o (n3371) );
  buffer buf_n3372( .i (n3371), .o (n3372) );
  buffer buf_n3373( .i (n3372), .o (n3373) );
  buffer buf_n3374( .i (n3373), .o (n3374) );
  buffer buf_n3375( .i (n3374), .o (n3375) );
  buffer buf_n3376( .i (n3375), .o (n3376) );
  buffer buf_n3377( .i (n3376), .o (n3377) );
  buffer buf_n3378( .i (n3377), .o (n3378) );
  buffer buf_n3379( .i (n3378), .o (n3379) );
  buffer buf_n3380( .i (n3379), .o (n3380) );
  buffer buf_n3381( .i (n3380), .o (n3381) );
  buffer buf_n3382( .i (n3381), .o (n3382) );
  buffer buf_n3383( .i (n3382), .o (n3383) );
  buffer buf_n3384( .i (n3383), .o (n3384) );
  buffer buf_n3385( .i (n3384), .o (n3385) );
  buffer buf_n3386( .i (n3385), .o (n3386) );
  buffer buf_n3387( .i (n3386), .o (n3387) );
  buffer buf_n3388( .i (n3387), .o (n3388) );
  buffer buf_n3389( .i (n3388), .o (n3389) );
  buffer buf_n3390( .i (n3389), .o (n3390) );
  buffer buf_n3391( .i (n3390), .o (n3391) );
  buffer buf_n3392( .i (n3391), .o (n3392) );
  buffer buf_n3393( .i (n3392), .o (n3393) );
  buffer buf_n3394( .i (n3393), .o (n3394) );
  buffer buf_n3395( .i (n3394), .o (n3395) );
  buffer buf_n3396( .i (n3395), .o (n3396) );
  buffer buf_n3397( .i (n3396), .o (n3397) );
  buffer buf_n3398( .i (n3397), .o (n3398) );
  buffer buf_n3399( .i (n3398), .o (n3399) );
  buffer buf_n3400( .i (n3399), .o (n3400) );
  buffer buf_n3401( .i (n3400), .o (n3401) );
  buffer buf_n3402( .i (n3401), .o (n3402) );
  buffer buf_n3403( .i (n3402), .o (n3403) );
  buffer buf_n3404( .i (n3403), .o (n3404) );
  buffer buf_n3405( .i (n3404), .o (n3405) );
  buffer buf_n3406( .i (n3405), .o (n3406) );
  buffer buf_n3407( .i (n3406), .o (n3407) );
  buffer buf_n3408( .i (n3407), .o (n3408) );
  buffer buf_n3409( .i (n3408), .o (n3409) );
  buffer buf_n3410( .i (n3409), .o (n3410) );
  buffer buf_n3411( .i (n3410), .o (n3411) );
  buffer buf_n3412( .i (n3411), .o (n3412) );
  buffer buf_n3413( .i (n3412), .o (n3413) );
  buffer buf_n3414( .i (n3413), .o (n3414) );
  buffer buf_n3415( .i (n3414), .o (n3415) );
  buffer buf_n3416( .i (n3415), .o (n3416) );
  buffer buf_n3417( .i (n3416), .o (n3417) );
  buffer buf_n3418( .i (n3417), .o (n3418) );
  buffer buf_n3419( .i (n3418), .o (n3419) );
  buffer buf_n3420( .i (n3419), .o (n3420) );
  buffer buf_n3421( .i (n3420), .o (n3421) );
  buffer buf_n3422( .i (n3421), .o (n3422) );
  buffer buf_n3423( .i (n3422), .o (n3423) );
  buffer buf_n3424( .i (n3423), .o (n3424) );
  buffer buf_n3425( .i (n3424), .o (n3425) );
  buffer buf_n3426( .i (n3425), .o (n3426) );
  buffer buf_n3427( .i (n3426), .o (n3427) );
  buffer buf_n3428( .i (n3427), .o (n3428) );
  buffer buf_n3429( .i (n3428), .o (n3429) );
  buffer buf_n3430( .i (n3429), .o (n3430) );
  buffer buf_n3431( .i (n3430), .o (n3431) );
  buffer buf_n3432( .i (n3431), .o (n3432) );
  buffer buf_n3433( .i (n3432), .o (n3433) );
  buffer buf_n3434( .i (n3433), .o (n3434) );
  buffer buf_n2994( .i (n2993), .o (n2994) );
  buffer buf_n2995( .i (n2994), .o (n2995) );
  buffer buf_n2996( .i (n2995), .o (n2996) );
  buffer buf_n2997( .i (n2996), .o (n2997) );
  buffer buf_n2998( .i (n2997), .o (n2998) );
  buffer buf_n2999( .i (n2998), .o (n2999) );
  buffer buf_n3000( .i (n2999), .o (n3000) );
  buffer buf_n3001( .i (n3000), .o (n3001) );
  buffer buf_n3002( .i (n3001), .o (n3002) );
  buffer buf_n3003( .i (n3002), .o (n3003) );
  buffer buf_n3004( .i (n3003), .o (n3004) );
  buffer buf_n3005( .i (n3004), .o (n3005) );
  buffer buf_n3006( .i (n3005), .o (n3006) );
  buffer buf_n3007( .i (n3006), .o (n3007) );
  buffer buf_n3008( .i (n3007), .o (n3008) );
  buffer buf_n3009( .i (n3008), .o (n3009) );
  buffer buf_n3010( .i (n3009), .o (n3010) );
  buffer buf_n3011( .i (n3010), .o (n3011) );
  buffer buf_n3012( .i (n3011), .o (n3012) );
  buffer buf_n3013( .i (n3012), .o (n3013) );
  buffer buf_n3014( .i (n3013), .o (n3014) );
  buffer buf_n3015( .i (n3014), .o (n3015) );
  buffer buf_n3016( .i (n3015), .o (n3016) );
  buffer buf_n3017( .i (n3016), .o (n3017) );
  buffer buf_n3018( .i (n3017), .o (n3018) );
  buffer buf_n3019( .i (n3018), .o (n3019) );
  buffer buf_n3020( .i (n3019), .o (n3020) );
  buffer buf_n3021( .i (n3020), .o (n3021) );
  buffer buf_n3022( .i (n3021), .o (n3022) );
  buffer buf_n3023( .i (n3022), .o (n3023) );
  buffer buf_n3024( .i (n3023), .o (n3024) );
  buffer buf_n3025( .i (n3024), .o (n3025) );
  buffer buf_n3026( .i (n3025), .o (n3026) );
  buffer buf_n3027( .i (n3026), .o (n3027) );
  buffer buf_n3028( .i (n3027), .o (n3028) );
  buffer buf_n3029( .i (n3028), .o (n3029) );
  buffer buf_n3030( .i (n3029), .o (n3030) );
  buffer buf_n3031( .i (n3030), .o (n3031) );
  buffer buf_n3032( .i (n3031), .o (n3032) );
  buffer buf_n3033( .i (n3032), .o (n3033) );
  buffer buf_n3034( .i (n3033), .o (n3034) );
  buffer buf_n3035( .i (n3034), .o (n3035) );
  buffer buf_n3036( .i (n3035), .o (n3036) );
  buffer buf_n3037( .i (n3036), .o (n3037) );
  buffer buf_n3038( .i (n3037), .o (n3038) );
  buffer buf_n3039( .i (n3038), .o (n3039) );
  buffer buf_n3040( .i (n3039), .o (n3040) );
  buffer buf_n3041( .i (n3040), .o (n3041) );
  buffer buf_n3042( .i (n3041), .o (n3042) );
  buffer buf_n3043( .i (n3042), .o (n3043) );
  buffer buf_n3044( .i (n3043), .o (n3044) );
  buffer buf_n3045( .i (n3044), .o (n3045) );
  buffer buf_n3046( .i (n3045), .o (n3046) );
  buffer buf_n3047( .i (n3046), .o (n3047) );
  buffer buf_n3048( .i (n3047), .o (n3048) );
  buffer buf_n3049( .i (n3048), .o (n3049) );
  buffer buf_n3050( .i (n3049), .o (n3050) );
  buffer buf_n3051( .i (n3050), .o (n3051) );
  buffer buf_n3052( .i (n3051), .o (n3052) );
  buffer buf_n3053( .i (n3052), .o (n3053) );
  buffer buf_n3054( .i (n3053), .o (n3054) );
  buffer buf_n3055( .i (n3054), .o (n3055) );
  buffer buf_n3056( .i (n3055), .o (n3056) );
  buffer buf_n3057( .i (n3056), .o (n3057) );
  buffer buf_n3058( .i (n3057), .o (n3058) );
  buffer buf_n3059( .i (n3058), .o (n3059) );
  buffer buf_n3060( .i (n3059), .o (n3060) );
  buffer buf_n3061( .i (n3060), .o (n3061) );
  buffer buf_n3062( .i (n3061), .o (n3062) );
  buffer buf_n3063( .i (n3062), .o (n3063) );
  buffer buf_n3064( .i (n3063), .o (n3064) );
  buffer buf_n3065( .i (n3064), .o (n3065) );
  buffer buf_n3066( .i (n3065), .o (n3066) );
  buffer buf_n3067( .i (n3066), .o (n3067) );
  buffer buf_n3068( .i (n3067), .o (n3068) );
  buffer buf_n3069( .i (n3068), .o (n3069) );
  buffer buf_n3070( .i (n3069), .o (n3070) );
  buffer buf_n3071( .i (n3070), .o (n3071) );
  buffer buf_n3072( .i (n3071), .o (n3072) );
  buffer buf_n3073( .i (n3072), .o (n3073) );
  buffer buf_n3074( .i (n3073), .o (n3074) );
  buffer buf_n3075( .i (n3074), .o (n3075) );
  buffer buf_n3076( .i (n3075), .o (n3076) );
  buffer buf_n3077( .i (n3076), .o (n3077) );
  buffer buf_n3078( .i (n3077), .o (n3078) );
  buffer buf_n3079( .i (n3078), .o (n3079) );
  buffer buf_n3080( .i (n3079), .o (n3080) );
  buffer buf_n3081( .i (n3080), .o (n3081) );
  buffer buf_n3082( .i (n3081), .o (n3082) );
  buffer buf_n3083( .i (n3082), .o (n3083) );
  buffer buf_n3084( .i (n3083), .o (n3084) );
  buffer buf_n3085( .i (n3084), .o (n3085) );
  buffer buf_n3086( .i (n3085), .o (n3086) );
  buffer buf_n3087( .i (n3086), .o (n3087) );
  buffer buf_n3088( .i (n3087), .o (n3088) );
  buffer buf_n3089( .i (n3088), .o (n3089) );
  buffer buf_n3090( .i (n3089), .o (n3090) );
  buffer buf_n3091( .i (n3090), .o (n3091) );
  buffer buf_n3092( .i (n3091), .o (n3092) );
  buffer buf_n3093( .i (n3092), .o (n3093) );
  buffer buf_n3094( .i (n3093), .o (n3094) );
  buffer buf_n3095( .i (n3094), .o (n3095) );
  buffer buf_n3096( .i (n3095), .o (n3096) );
  buffer buf_n3097( .i (n3096), .o (n3097) );
  buffer buf_n3098( .i (n3097), .o (n3098) );
  buffer buf_n3099( .i (n3098), .o (n3099) );
  buffer buf_n3100( .i (n3099), .o (n3100) );
  buffer buf_n3101( .i (n3100), .o (n3101) );
  buffer buf_n3102( .i (n3101), .o (n3102) );
  buffer buf_n3103( .i (n3102), .o (n3103) );
  buffer buf_n3104( .i (n3103), .o (n3104) );
  buffer buf_n3105( .i (n3104), .o (n3105) );
  buffer buf_n3106( .i (n3105), .o (n3106) );
  buffer buf_n3107( .i (n3106), .o (n3107) );
  buffer buf_n3108( .i (n3107), .o (n3108) );
  assign n6899 = n971 & n6796 ;
  buffer buf_n6900( .i (n6899), .o (n6900) );
  assign n6901 = n6798 & ~n6900 ;
  buffer buf_n6902( .i (n6901), .o (n6902) );
  buffer buf_n6903( .i (n6902), .o (n6903) );
  buffer buf_n6904( .i (n6903), .o (n6904) );
  buffer buf_n6905( .i (n6904), .o (n6905) );
  buffer buf_n6906( .i (n6905), .o (n6906) );
  buffer buf_n6907( .i (n6906), .o (n6907) );
  buffer buf_n6908( .i (n6907), .o (n6908) );
  buffer buf_n6909( .i (n6908), .o (n6909) );
  buffer buf_n6910( .i (n6909), .o (n6910) );
  buffer buf_n6911( .i (n6910), .o (n6911) );
  buffer buf_n6912( .i (n6911), .o (n6912) );
  buffer buf_n6913( .i (n6912), .o (n6913) );
  buffer buf_n6914( .i (n6913), .o (n6914) );
  buffer buf_n6915( .i (n6914), .o (n6915) );
  buffer buf_n6916( .i (n6915), .o (n6916) );
  buffer buf_n6917( .i (n6916), .o (n6917) );
  buffer buf_n6918( .i (n6917), .o (n6918) );
  buffer buf_n6919( .i (n6918), .o (n6919) );
  buffer buf_n6920( .i (n6919), .o (n6920) );
  buffer buf_n6921( .i (n6920), .o (n6921) );
  buffer buf_n6922( .i (n6921), .o (n6922) );
  buffer buf_n6923( .i (n6922), .o (n6923) );
  buffer buf_n6924( .i (n6923), .o (n6924) );
  buffer buf_n6925( .i (n6924), .o (n6925) );
  buffer buf_n6926( .i (n6925), .o (n6926) );
  buffer buf_n6927( .i (n6926), .o (n6927) );
  buffer buf_n6928( .i (n6927), .o (n6928) );
  buffer buf_n6929( .i (n6928), .o (n6929) );
  buffer buf_n6930( .i (n6929), .o (n6930) );
  buffer buf_n6931( .i (n6930), .o (n6931) );
  buffer buf_n6932( .i (n6931), .o (n6932) );
  buffer buf_n6933( .i (n6932), .o (n6933) );
  buffer buf_n6934( .i (n6933), .o (n6934) );
  buffer buf_n6935( .i (n6934), .o (n6935) );
  buffer buf_n6936( .i (n6935), .o (n6936) );
  buffer buf_n6937( .i (n6936), .o (n6937) );
  buffer buf_n6938( .i (n6937), .o (n6938) );
  buffer buf_n6939( .i (n6938), .o (n6939) );
  buffer buf_n6940( .i (n6939), .o (n6940) );
  buffer buf_n6941( .i (n6940), .o (n6941) );
  buffer buf_n6942( .i (n6941), .o (n6942) );
  buffer buf_n6943( .i (n6942), .o (n6943) );
  buffer buf_n6944( .i (n6943), .o (n6944) );
  buffer buf_n6945( .i (n6944), .o (n6945) );
  buffer buf_n6946( .i (n6945), .o (n6946) );
  buffer buf_n6947( .i (n6946), .o (n6947) );
  buffer buf_n6948( .i (n6947), .o (n6948) );
  buffer buf_n6949( .i (n6948), .o (n6949) );
  buffer buf_n6950( .i (n6949), .o (n6950) );
  buffer buf_n6951( .i (n6950), .o (n6951) );
  buffer buf_n6952( .i (n6951), .o (n6952) );
  buffer buf_n6953( .i (n6952), .o (n6953) );
  buffer buf_n6954( .i (n6953), .o (n6954) );
  buffer buf_n6955( .i (n6954), .o (n6955) );
  buffer buf_n6956( .i (n6955), .o (n6956) );
  buffer buf_n6957( .i (n6956), .o (n6957) );
  buffer buf_n6958( .i (n6957), .o (n6958) );
  buffer buf_n6959( .i (n6958), .o (n6959) );
  buffer buf_n6960( .i (n6959), .o (n6960) );
  buffer buf_n6961( .i (n6960), .o (n6961) );
  buffer buf_n6962( .i (n6961), .o (n6962) );
  buffer buf_n6963( .i (n6962), .o (n6963) );
  buffer buf_n6964( .i (n6963), .o (n6964) );
  buffer buf_n6965( .i (n6964), .o (n6965) );
  buffer buf_n6966( .i (n6965), .o (n6966) );
  buffer buf_n6967( .i (n6966), .o (n6967) );
  buffer buf_n6968( .i (n6967), .o (n6968) );
  buffer buf_n6969( .i (n6968), .o (n6969) );
  buffer buf_n6970( .i (n6969), .o (n6970) );
  buffer buf_n6971( .i (n6970), .o (n6971) );
  buffer buf_n6972( .i (n6971), .o (n6972) );
  buffer buf_n6973( .i (n6972), .o (n6973) );
  buffer buf_n6974( .i (n6973), .o (n6974) );
  buffer buf_n6975( .i (n6974), .o (n6975) );
  buffer buf_n6976( .i (n6975), .o (n6976) );
  buffer buf_n6977( .i (n6976), .o (n6977) );
  buffer buf_n6978( .i (n6977), .o (n6978) );
  buffer buf_n6979( .i (n6978), .o (n6979) );
  buffer buf_n6980( .i (n6979), .o (n6980) );
  buffer buf_n6981( .i (n6980), .o (n6981) );
  buffer buf_n6982( .i (n6981), .o (n6982) );
  buffer buf_n6983( .i (n6982), .o (n6983) );
  buffer buf_n6984( .i (n6983), .o (n6984) );
  buffer buf_n2308( .i (n2307), .o (n2308) );
  buffer buf_n2309( .i (n2308), .o (n2309) );
  buffer buf_n2310( .i (n2309), .o (n2310) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n2321( .i (n2320), .o (n2321) );
  buffer buf_n2322( .i (n2321), .o (n2322) );
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2325( .i (n2324), .o (n2325) );
  buffer buf_n2326( .i (n2325), .o (n2326) );
  buffer buf_n2327( .i (n2326), .o (n2327) );
  buffer buf_n2328( .i (n2327), .o (n2328) );
  buffer buf_n2329( .i (n2328), .o (n2329) );
  buffer buf_n2330( .i (n2329), .o (n2330) );
  buffer buf_n2331( .i (n2330), .o (n2331) );
  buffer buf_n2332( .i (n2331), .o (n2332) );
  buffer buf_n2333( .i (n2332), .o (n2333) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n2335( .i (n2334), .o (n2335) );
  buffer buf_n2336( .i (n2335), .o (n2336) );
  buffer buf_n2337( .i (n2336), .o (n2337) );
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  buffer buf_n2340( .i (n2339), .o (n2340) );
  buffer buf_n2341( .i (n2340), .o (n2341) );
  buffer buf_n2342( .i (n2341), .o (n2342) );
  buffer buf_n2343( .i (n2342), .o (n2343) );
  buffer buf_n2344( .i (n2343), .o (n2344) );
  buffer buf_n2345( .i (n2344), .o (n2345) );
  buffer buf_n2346( .i (n2345), .o (n2346) );
  buffer buf_n2347( .i (n2346), .o (n2347) );
  buffer buf_n2348( .i (n2347), .o (n2348) );
  buffer buf_n2349( .i (n2348), .o (n2349) );
  buffer buf_n2350( .i (n2349), .o (n2350) );
  buffer buf_n2351( .i (n2350), .o (n2351) );
  buffer buf_n2352( .i (n2351), .o (n2352) );
  buffer buf_n2353( .i (n2352), .o (n2353) );
  buffer buf_n2354( .i (n2353), .o (n2354) );
  buffer buf_n2355( .i (n2354), .o (n2355) );
  buffer buf_n2356( .i (n2355), .o (n2356) );
  buffer buf_n2357( .i (n2356), .o (n2357) );
  buffer buf_n2358( .i (n2357), .o (n2358) );
  buffer buf_n2359( .i (n2358), .o (n2359) );
  buffer buf_n2360( .i (n2359), .o (n2360) );
  buffer buf_n2361( .i (n2360), .o (n2361) );
  buffer buf_n2362( .i (n2361), .o (n2362) );
  buffer buf_n2363( .i (n2362), .o (n2363) );
  buffer buf_n2364( .i (n2363), .o (n2364) );
  buffer buf_n2365( .i (n2364), .o (n2365) );
  buffer buf_n2366( .i (n2365), .o (n2366) );
  buffer buf_n2367( .i (n2366), .o (n2367) );
  buffer buf_n2368( .i (n2367), .o (n2368) );
  buffer buf_n2369( .i (n2368), .o (n2369) );
  buffer buf_n2370( .i (n2369), .o (n2370) );
  buffer buf_n2371( .i (n2370), .o (n2371) );
  buffer buf_n2372( .i (n2371), .o (n2372) );
  buffer buf_n2373( .i (n2372), .o (n2373) );
  buffer buf_n2374( .i (n2373), .o (n2374) );
  buffer buf_n2375( .i (n2374), .o (n2375) );
  buffer buf_n2376( .i (n2375), .o (n2376) );
  buffer buf_n2377( .i (n2376), .o (n2377) );
  buffer buf_n2378( .i (n2377), .o (n2378) );
  buffer buf_n2379( .i (n2378), .o (n2379) );
  buffer buf_n2380( .i (n2379), .o (n2380) );
  buffer buf_n2381( .i (n2380), .o (n2381) );
  buffer buf_n2382( .i (n2381), .o (n2382) );
  buffer buf_n2383( .i (n2382), .o (n2383) );
  buffer buf_n2384( .i (n2383), .o (n2384) );
  buffer buf_n2385( .i (n2384), .o (n2385) );
  buffer buf_n2386( .i (n2385), .o (n2386) );
  buffer buf_n2387( .i (n2386), .o (n2387) );
  buffer buf_n2388( .i (n2387), .o (n2388) );
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2391( .i (n2390), .o (n2391) );
  buffer buf_n2392( .i (n2391), .o (n2392) );
  buffer buf_n2393( .i (n2392), .o (n2393) );
  buffer buf_n2394( .i (n2393), .o (n2394) );
  buffer buf_n2395( .i (n2394), .o (n2395) );
  buffer buf_n2396( .i (n2395), .o (n2396) );
  buffer buf_n2397( .i (n2396), .o (n2397) );
  buffer buf_n2398( .i (n2397), .o (n2398) );
  buffer buf_n2399( .i (n2398), .o (n2399) );
  buffer buf_n2400( .i (n2399), .o (n2400) );
  buffer buf_n2401( .i (n2400), .o (n2401) );
  buffer buf_n2402( .i (n2401), .o (n2402) );
  buffer buf_n2403( .i (n2402), .o (n2403) );
  buffer buf_n2404( .i (n2403), .o (n2404) );
  buffer buf_n2405( .i (n2404), .o (n2405) );
  buffer buf_n2406( .i (n2405), .o (n2406) );
  buffer buf_n2407( .i (n2406), .o (n2407) );
  buffer buf_n2408( .i (n2407), .o (n2408) );
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  buffer buf_n2411( .i (n2410), .o (n2411) );
  buffer buf_n2412( .i (n2411), .o (n2412) );
  buffer buf_n2413( .i (n2412), .o (n2413) );
  buffer buf_n2414( .i (n2413), .o (n2414) );
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n2416( .i (n2415), .o (n2416) );
  buffer buf_n3601( .i (n3600), .o (n3601) );
  buffer buf_n3602( .i (n3601), .o (n3602) );
  buffer buf_n3603( .i (n3602), .o (n3603) );
  buffer buf_n3604( .i (n3603), .o (n3604) );
  buffer buf_n3605( .i (n3604), .o (n3605) );
  buffer buf_n3606( .i (n3605), .o (n3606) );
  buffer buf_n3607( .i (n3606), .o (n3607) );
  buffer buf_n3608( .i (n3607), .o (n3608) );
  buffer buf_n3609( .i (n3608), .o (n3609) );
  buffer buf_n3610( .i (n3609), .o (n3610) );
  buffer buf_n3611( .i (n3610), .o (n3611) );
  buffer buf_n3612( .i (n3611), .o (n3612) );
  buffer buf_n3613( .i (n3612), .o (n3613) );
  buffer buf_n3614( .i (n3613), .o (n3614) );
  buffer buf_n3615( .i (n3614), .o (n3615) );
  buffer buf_n3616( .i (n3615), .o (n3616) );
  buffer buf_n3617( .i (n3616), .o (n3617) );
  buffer buf_n3618( .i (n3617), .o (n3618) );
  buffer buf_n3619( .i (n3618), .o (n3619) );
  buffer buf_n3620( .i (n3619), .o (n3620) );
  buffer buf_n3621( .i (n3620), .o (n3621) );
  buffer buf_n3622( .i (n3621), .o (n3622) );
  buffer buf_n3623( .i (n3622), .o (n3623) );
  buffer buf_n3624( .i (n3623), .o (n3624) );
  buffer buf_n3625( .i (n3624), .o (n3625) );
  buffer buf_n3626( .i (n3625), .o (n3626) );
  buffer buf_n3627( .i (n3626), .o (n3627) );
  buffer buf_n3628( .i (n3627), .o (n3628) );
  buffer buf_n3629( .i (n3628), .o (n3629) );
  buffer buf_n3630( .i (n3629), .o (n3630) );
  buffer buf_n3631( .i (n3630), .o (n3631) );
  buffer buf_n3632( .i (n3631), .o (n3632) );
  buffer buf_n3633( .i (n3632), .o (n3633) );
  buffer buf_n3634( .i (n3633), .o (n3634) );
  buffer buf_n3635( .i (n3634), .o (n3635) );
  buffer buf_n3636( .i (n3635), .o (n3636) );
  buffer buf_n3637( .i (n3636), .o (n3637) );
  buffer buf_n3638( .i (n3637), .o (n3638) );
  buffer buf_n3639( .i (n3638), .o (n3639) );
  buffer buf_n3640( .i (n3639), .o (n3640) );
  buffer buf_n3641( .i (n3640), .o (n3641) );
  buffer buf_n3642( .i (n3641), .o (n3642) );
  buffer buf_n3643( .i (n3642), .o (n3643) );
  buffer buf_n3644( .i (n3643), .o (n3644) );
  buffer buf_n3645( .i (n3644), .o (n3645) );
  buffer buf_n3646( .i (n3645), .o (n3646) );
  buffer buf_n3647( .i (n3646), .o (n3647) );
  buffer buf_n3648( .i (n3647), .o (n3648) );
  buffer buf_n3649( .i (n3648), .o (n3649) );
  buffer buf_n3650( .i (n3649), .o (n3650) );
  buffer buf_n3651( .i (n3650), .o (n3651) );
  buffer buf_n3652( .i (n3651), .o (n3652) );
  buffer buf_n3653( .i (n3652), .o (n3653) );
  buffer buf_n3654( .i (n3653), .o (n3654) );
  buffer buf_n3655( .i (n3654), .o (n3655) );
  buffer buf_n3656( .i (n3655), .o (n3656) );
  buffer buf_n3657( .i (n3656), .o (n3657) );
  buffer buf_n3658( .i (n3657), .o (n3658) );
  buffer buf_n3659( .i (n3658), .o (n3659) );
  buffer buf_n3660( .i (n3659), .o (n3660) );
  buffer buf_n3661( .i (n3660), .o (n3661) );
  buffer buf_n3662( .i (n3661), .o (n3662) );
  buffer buf_n3663( .i (n3662), .o (n3663) );
  buffer buf_n3664( .i (n3663), .o (n3664) );
  buffer buf_n3665( .i (n3664), .o (n3665) );
  buffer buf_n3666( .i (n3665), .o (n3666) );
  buffer buf_n3667( .i (n3666), .o (n3667) );
  buffer buf_n3668( .i (n3667), .o (n3668) );
  buffer buf_n3669( .i (n3668), .o (n3669) );
  buffer buf_n3670( .i (n3669), .o (n3670) );
  buffer buf_n3671( .i (n3670), .o (n3671) );
  buffer buf_n3672( .i (n3671), .o (n3672) );
  buffer buf_n3673( .i (n3672), .o (n3673) );
  buffer buf_n3674( .i (n3673), .o (n3674) );
  buffer buf_n3675( .i (n3674), .o (n3675) );
  buffer buf_n3676( .i (n3675), .o (n3676) );
  buffer buf_n3677( .i (n3676), .o (n3677) );
  buffer buf_n3678( .i (n3677), .o (n3678) );
  buffer buf_n3679( .i (n3678), .o (n3679) );
  buffer buf_n3680( .i (n3679), .o (n3680) );
  buffer buf_n3681( .i (n3680), .o (n3681) );
  buffer buf_n3682( .i (n3681), .o (n3682) );
  buffer buf_n3683( .i (n3682), .o (n3683) );
  buffer buf_n3684( .i (n3683), .o (n3684) );
  buffer buf_n3685( .i (n3684), .o (n3685) );
  buffer buf_n3686( .i (n3685), .o (n3686) );
  buffer buf_n3687( .i (n3686), .o (n3687) );
  buffer buf_n3688( .i (n3687), .o (n3688) );
  buffer buf_n3689( .i (n3688), .o (n3689) );
  buffer buf_n3690( .i (n3689), .o (n3690) );
  buffer buf_n3691( .i (n3690), .o (n3691) );
  buffer buf_n3692( .i (n3691), .o (n3692) );
  buffer buf_n3693( .i (n3692), .o (n3693) );
  buffer buf_n3694( .i (n3693), .o (n3694) );
  buffer buf_n3695( .i (n3694), .o (n3695) );
  buffer buf_n3696( .i (n3695), .o (n3696) );
  buffer buf_n3697( .i (n3696), .o (n3697) );
  buffer buf_n3698( .i (n3697), .o (n3698) );
  buffer buf_n3699( .i (n3698), .o (n3699) );
  buffer buf_n3700( .i (n3699), .o (n3700) );
  buffer buf_n3701( .i (n3700), .o (n3701) );
  buffer buf_n3702( .i (n3701), .o (n3702) );
  buffer buf_n3703( .i (n3702), .o (n3703) );
  buffer buf_n4088( .i (n4087), .o (n4088) );
  buffer buf_n4089( .i (n4088), .o (n4089) );
  buffer buf_n4090( .i (n4089), .o (n4090) );
  buffer buf_n4091( .i (n4090), .o (n4091) );
  buffer buf_n4092( .i (n4091), .o (n4092) );
  buffer buf_n4093( .i (n4092), .o (n4093) );
  buffer buf_n4094( .i (n4093), .o (n4094) );
  buffer buf_n4095( .i (n4094), .o (n4095) );
  buffer buf_n4096( .i (n4095), .o (n4096) );
  buffer buf_n4097( .i (n4096), .o (n4097) );
  buffer buf_n4098( .i (n4097), .o (n4098) );
  buffer buf_n4099( .i (n4098), .o (n4099) );
  buffer buf_n4100( .i (n4099), .o (n4100) );
  buffer buf_n4101( .i (n4100), .o (n4101) );
  buffer buf_n4102( .i (n4101), .o (n4102) );
  buffer buf_n4103( .i (n4102), .o (n4103) );
  buffer buf_n4104( .i (n4103), .o (n4104) );
  buffer buf_n4105( .i (n4104), .o (n4105) );
  buffer buf_n4106( .i (n4105), .o (n4106) );
  buffer buf_n4107( .i (n4106), .o (n4107) );
  buffer buf_n4108( .i (n4107), .o (n4108) );
  buffer buf_n4109( .i (n4108), .o (n4109) );
  buffer buf_n4110( .i (n4109), .o (n4110) );
  buffer buf_n4111( .i (n4110), .o (n4111) );
  buffer buf_n4112( .i (n4111), .o (n4112) );
  buffer buf_n4113( .i (n4112), .o (n4113) );
  buffer buf_n4114( .i (n4113), .o (n4114) );
  buffer buf_n4115( .i (n4114), .o (n4115) );
  buffer buf_n4116( .i (n4115), .o (n4116) );
  buffer buf_n4117( .i (n4116), .o (n4117) );
  buffer buf_n4118( .i (n4117), .o (n4118) );
  buffer buf_n4119( .i (n4118), .o (n4119) );
  buffer buf_n4120( .i (n4119), .o (n4120) );
  buffer buf_n4121( .i (n4120), .o (n4121) );
  buffer buf_n4122( .i (n4121), .o (n4122) );
  buffer buf_n4123( .i (n4122), .o (n4123) );
  buffer buf_n4124( .i (n4123), .o (n4124) );
  buffer buf_n4125( .i (n4124), .o (n4125) );
  buffer buf_n4126( .i (n4125), .o (n4126) );
  buffer buf_n4127( .i (n4126), .o (n4127) );
  buffer buf_n4128( .i (n4127), .o (n4128) );
  buffer buf_n4129( .i (n4128), .o (n4129) );
  buffer buf_n4130( .i (n4129), .o (n4130) );
  buffer buf_n4131( .i (n4130), .o (n4131) );
  buffer buf_n4132( .i (n4131), .o (n4132) );
  buffer buf_n4133( .i (n4132), .o (n4133) );
  buffer buf_n4134( .i (n4133), .o (n4134) );
  buffer buf_n4135( .i (n4134), .o (n4135) );
  buffer buf_n4136( .i (n4135), .o (n4136) );
  buffer buf_n4137( .i (n4136), .o (n4137) );
  buffer buf_n4138( .i (n4137), .o (n4138) );
  buffer buf_n4139( .i (n4138), .o (n4139) );
  buffer buf_n4140( .i (n4139), .o (n4140) );
  buffer buf_n4141( .i (n4140), .o (n4141) );
  buffer buf_n4142( .i (n4141), .o (n4142) );
  buffer buf_n4143( .i (n4142), .o (n4143) );
  buffer buf_n4144( .i (n4143), .o (n4144) );
  buffer buf_n4145( .i (n4144), .o (n4145) );
  buffer buf_n4146( .i (n4145), .o (n4146) );
  buffer buf_n4147( .i (n4146), .o (n4147) );
  buffer buf_n4148( .i (n4147), .o (n4148) );
  buffer buf_n4149( .i (n4148), .o (n4149) );
  buffer buf_n4150( .i (n4149), .o (n4150) );
  buffer buf_n4151( .i (n4150), .o (n4151) );
  buffer buf_n4152( .i (n4151), .o (n4152) );
  buffer buf_n4153( .i (n4152), .o (n4153) );
  buffer buf_n4154( .i (n4153), .o (n4154) );
  buffer buf_n4155( .i (n4154), .o (n4155) );
  buffer buf_n4156( .i (n4155), .o (n4156) );
  buffer buf_n4157( .i (n4156), .o (n4157) );
  buffer buf_n4158( .i (n4157), .o (n4158) );
  buffer buf_n4159( .i (n4158), .o (n4159) );
  buffer buf_n4160( .i (n4159), .o (n4160) );
  buffer buf_n4161( .i (n4160), .o (n4161) );
  buffer buf_n4162( .i (n4161), .o (n4162) );
  buffer buf_n4163( .i (n4162), .o (n4163) );
  buffer buf_n4164( .i (n4163), .o (n4164) );
  buffer buf_n4165( .i (n4164), .o (n4165) );
  buffer buf_n4166( .i (n4165), .o (n4166) );
  buffer buf_n4167( .i (n4166), .o (n4167) );
  buffer buf_n4168( .i (n4167), .o (n4168) );
  buffer buf_n4169( .i (n4168), .o (n4169) );
  buffer buf_n4170( .i (n4169), .o (n4170) );
  buffer buf_n4171( .i (n4170), .o (n4171) );
  buffer buf_n4172( .i (n4171), .o (n4172) );
  buffer buf_n4173( .i (n4172), .o (n4173) );
  buffer buf_n4174( .i (n4173), .o (n4174) );
  buffer buf_n4175( .i (n4174), .o (n4175) );
  buffer buf_n4176( .i (n4175), .o (n4176) );
  buffer buf_n4177( .i (n4176), .o (n4177) );
  buffer buf_n4178( .i (n4177), .o (n4178) );
  buffer buf_n4179( .i (n4178), .o (n4179) );
  buffer buf_n4180( .i (n4179), .o (n4180) );
  buffer buf_n4181( .i (n4180), .o (n4181) );
  buffer buf_n4182( .i (n4181), .o (n4182) );
  buffer buf_n4183( .i (n4182), .o (n4183) );
  buffer buf_n4184( .i (n4183), .o (n4184) );
  buffer buf_n4185( .i (n4184), .o (n4185) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n1247( .i (n1246), .o (n1247) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n3161( .i (n3160), .o (n3161) );
  buffer buf_n3162( .i (n3161), .o (n3162) );
  assign n6987 = n3918 & n6787 ;
  buffer buf_n6988( .i (n6987), .o (n6988) );
  assign n6989 = n3162 & ~n6988 ;
  assign n6990 = ~n3162 & n6988 ;
  assign n6991 = n6989 | n6990 ;
  buffer buf_n6992( .i (n6991), .o (n6992) );
  buffer buf_n6993( .i (n6992), .o (n6993) );
  buffer buf_n6994( .i (n6993), .o (n6994) );
  buffer buf_n6995( .i (n6994), .o (n6995) );
  buffer buf_n6996( .i (n6995), .o (n6996) );
  buffer buf_n6997( .i (n6996), .o (n6997) );
  buffer buf_n6998( .i (n6997), .o (n6998) );
  buffer buf_n6999( .i (n6998), .o (n6999) );
  buffer buf_n7000( .i (n6999), .o (n7000) );
  buffer buf_n7001( .i (n7000), .o (n7001) );
  buffer buf_n7002( .i (n7001), .o (n7002) );
  buffer buf_n7003( .i (n7002), .o (n7003) );
  buffer buf_n7004( .i (n7003), .o (n7004) );
  buffer buf_n7005( .i (n7004), .o (n7005) );
  buffer buf_n7006( .i (n7005), .o (n7006) );
  buffer buf_n7007( .i (n7006), .o (n7007) );
  buffer buf_n7008( .i (n7007), .o (n7008) );
  buffer buf_n7009( .i (n7008), .o (n7009) );
  buffer buf_n7010( .i (n7009), .o (n7010) );
  buffer buf_n7011( .i (n7010), .o (n7011) );
  buffer buf_n7012( .i (n7011), .o (n7012) );
  buffer buf_n7013( .i (n7012), .o (n7013) );
  buffer buf_n7014( .i (n7013), .o (n7014) );
  buffer buf_n7015( .i (n7014), .o (n7015) );
  buffer buf_n7016( .i (n7015), .o (n7016) );
  buffer buf_n7017( .i (n7016), .o (n7017) );
  buffer buf_n7018( .i (n7017), .o (n7018) );
  buffer buf_n7019( .i (n7018), .o (n7019) );
  buffer buf_n7020( .i (n7019), .o (n7020) );
  buffer buf_n7021( .i (n7020), .o (n7021) );
  buffer buf_n7022( .i (n7021), .o (n7022) );
  buffer buf_n7023( .i (n7022), .o (n7023) );
  buffer buf_n7024( .i (n7023), .o (n7024) );
  buffer buf_n7025( .i (n7024), .o (n7025) );
  buffer buf_n7026( .i (n7025), .o (n7026) );
  buffer buf_n7027( .i (n7026), .o (n7027) );
  buffer buf_n7028( .i (n7027), .o (n7028) );
  buffer buf_n7029( .i (n7028), .o (n7029) );
  buffer buf_n7030( .i (n7029), .o (n7030) );
  buffer buf_n7031( .i (n7030), .o (n7031) );
  buffer buf_n7032( .i (n7031), .o (n7032) );
  buffer buf_n7033( .i (n7032), .o (n7033) );
  buffer buf_n7034( .i (n7033), .o (n7034) );
  buffer buf_n7035( .i (n7034), .o (n7035) );
  buffer buf_n7036( .i (n7035), .o (n7036) );
  buffer buf_n7037( .i (n7036), .o (n7037) );
  buffer buf_n7038( .i (n7037), .o (n7038) );
  buffer buf_n7039( .i (n7038), .o (n7039) );
  buffer buf_n7040( .i (n7039), .o (n7040) );
  buffer buf_n7041( .i (n7040), .o (n7041) );
  buffer buf_n7042( .i (n7041), .o (n7042) );
  buffer buf_n7043( .i (n7042), .o (n7043) );
  buffer buf_n7044( .i (n7043), .o (n7044) );
  buffer buf_n7045( .i (n7044), .o (n7045) );
  buffer buf_n7046( .i (n7045), .o (n7046) );
  buffer buf_n7047( .i (n7046), .o (n7047) );
  buffer buf_n7048( .i (n7047), .o (n7048) );
  buffer buf_n7049( .i (n7048), .o (n7049) );
  buffer buf_n7050( .i (n7049), .o (n7050) );
  buffer buf_n7051( .i (n7050), .o (n7051) );
  buffer buf_n7052( .i (n7051), .o (n7052) );
  buffer buf_n7053( .i (n7052), .o (n7053) );
  buffer buf_n7054( .i (n7053), .o (n7054) );
  buffer buf_n7055( .i (n7054), .o (n7055) );
  buffer buf_n7056( .i (n7055), .o (n7056) );
  buffer buf_n7057( .i (n7056), .o (n7057) );
  buffer buf_n7058( .i (n7057), .o (n7058) );
  buffer buf_n7059( .i (n7058), .o (n7059) );
  buffer buf_n7060( .i (n7059), .o (n7060) );
  buffer buf_n7061( .i (n7060), .o (n7061) );
  buffer buf_n3781( .i (n3780), .o (n3781) );
  buffer buf_n3782( .i (n3781), .o (n3782) );
  buffer buf_n3783( .i (n3782), .o (n3783) );
  buffer buf_n3784( .i (n3783), .o (n3784) );
  buffer buf_n3785( .i (n3784), .o (n3785) );
  buffer buf_n3786( .i (n3785), .o (n3786) );
  buffer buf_n3787( .i (n3786), .o (n3787) );
  buffer buf_n3788( .i (n3787), .o (n3788) );
  buffer buf_n3789( .i (n3788), .o (n3789) );
  buffer buf_n3790( .i (n3789), .o (n3790) );
  buffer buf_n3791( .i (n3790), .o (n3791) );
  buffer buf_n3792( .i (n3791), .o (n3792) );
  buffer buf_n3793( .i (n3792), .o (n3793) );
  buffer buf_n3794( .i (n3793), .o (n3794) );
  buffer buf_n3795( .i (n3794), .o (n3795) );
  buffer buf_n3796( .i (n3795), .o (n3796) );
  buffer buf_n3797( .i (n3796), .o (n3797) );
  buffer buf_n3798( .i (n3797), .o (n3798) );
  buffer buf_n3799( .i (n3798), .o (n3799) );
  buffer buf_n3800( .i (n3799), .o (n3800) );
  buffer buf_n3801( .i (n3800), .o (n3801) );
  buffer buf_n3802( .i (n3801), .o (n3802) );
  buffer buf_n3803( .i (n3802), .o (n3803) );
  buffer buf_n3804( .i (n3803), .o (n3804) );
  buffer buf_n3805( .i (n3804), .o (n3805) );
  buffer buf_n3806( .i (n3805), .o (n3806) );
  buffer buf_n3807( .i (n3806), .o (n3807) );
  buffer buf_n3808( .i (n3807), .o (n3808) );
  buffer buf_n3809( .i (n3808), .o (n3809) );
  buffer buf_n3810( .i (n3809), .o (n3810) );
  buffer buf_n3811( .i (n3810), .o (n3811) );
  buffer buf_n3812( .i (n3811), .o (n3812) );
  buffer buf_n3813( .i (n3812), .o (n3813) );
  buffer buf_n3814( .i (n3813), .o (n3814) );
  buffer buf_n3815( .i (n3814), .o (n3815) );
  buffer buf_n3816( .i (n3815), .o (n3816) );
  buffer buf_n3817( .i (n3816), .o (n3817) );
  buffer buf_n3818( .i (n3817), .o (n3818) );
  buffer buf_n3819( .i (n3818), .o (n3819) );
  buffer buf_n3820( .i (n3819), .o (n3820) );
  buffer buf_n3821( .i (n3820), .o (n3821) );
  buffer buf_n3822( .i (n3821), .o (n3822) );
  buffer buf_n3823( .i (n3822), .o (n3823) );
  buffer buf_n3824( .i (n3823), .o (n3824) );
  buffer buf_n3825( .i (n3824), .o (n3825) );
  buffer buf_n3826( .i (n3825), .o (n3826) );
  buffer buf_n3827( .i (n3826), .o (n3827) );
  buffer buf_n3828( .i (n3827), .o (n3828) );
  buffer buf_n3829( .i (n3828), .o (n3829) );
  buffer buf_n3830( .i (n3829), .o (n3830) );
  buffer buf_n3831( .i (n3830), .o (n3831) );
  buffer buf_n3832( .i (n3831), .o (n3832) );
  buffer buf_n3833( .i (n3832), .o (n3833) );
  buffer buf_n3834( .i (n3833), .o (n3834) );
  buffer buf_n3835( .i (n3834), .o (n3835) );
  buffer buf_n3836( .i (n3835), .o (n3836) );
  buffer buf_n3837( .i (n3836), .o (n3837) );
  buffer buf_n3838( .i (n3837), .o (n3838) );
  buffer buf_n3839( .i (n3838), .o (n3839) );
  buffer buf_n3840( .i (n3839), .o (n3840) );
  buffer buf_n3841( .i (n3840), .o (n3841) );
  buffer buf_n3842( .i (n3841), .o (n3842) );
  buffer buf_n3843( .i (n3842), .o (n3843) );
  buffer buf_n3844( .i (n3843), .o (n3844) );
  buffer buf_n3845( .i (n3844), .o (n3845) );
  buffer buf_n3846( .i (n3845), .o (n3846) );
  buffer buf_n3847( .i (n3846), .o (n3847) );
  buffer buf_n3848( .i (n3847), .o (n3848) );
  buffer buf_n3849( .i (n3848), .o (n3849) );
  buffer buf_n3850( .i (n3849), .o (n3850) );
  buffer buf_n3851( .i (n3850), .o (n3851) );
  buffer buf_n3852( .i (n3851), .o (n3852) );
  buffer buf_n3853( .i (n3852), .o (n3853) );
  buffer buf_n3854( .i (n3853), .o (n3854) );
  buffer buf_n3855( .i (n3854), .o (n3855) );
  buffer buf_n3856( .i (n3855), .o (n3856) );
  buffer buf_n3857( .i (n3856), .o (n3857) );
  buffer buf_n3858( .i (n3857), .o (n3858) );
  buffer buf_n3859( .i (n3858), .o (n3859) );
  buffer buf_n3860( .i (n3859), .o (n3860) );
  buffer buf_n3861( .i (n3860), .o (n3861) );
  buffer buf_n3862( .i (n3861), .o (n3862) );
  buffer buf_n3863( .i (n3862), .o (n3863) );
  buffer buf_n3864( .i (n3863), .o (n3864) );
  buffer buf_n3865( .i (n3864), .o (n3865) );
  buffer buf_n3866( .i (n3865), .o (n3866) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  assign n7064 = n3916 & n6785 ;
  buffer buf_n7065( .i (n7064), .o (n7065) );
  assign n7066 = n1642 & n7065 ;
  assign n7067 = n1642 | n7065 ;
  assign n7068 = ~n7066 & n7067 ;
  buffer buf_n7069( .i (n7068), .o (n7069) );
  buffer buf_n7070( .i (n7069), .o (n7070) );
  buffer buf_n7071( .i (n7070), .o (n7071) );
  buffer buf_n7072( .i (n7071), .o (n7072) );
  buffer buf_n7073( .i (n7072), .o (n7073) );
  buffer buf_n7074( .i (n7073), .o (n7074) );
  buffer buf_n7075( .i (n7074), .o (n7075) );
  buffer buf_n7076( .i (n7075), .o (n7076) );
  buffer buf_n7077( .i (n7076), .o (n7077) );
  buffer buf_n7078( .i (n7077), .o (n7078) );
  buffer buf_n7079( .i (n7078), .o (n7079) );
  buffer buf_n7080( .i (n7079), .o (n7080) );
  buffer buf_n7081( .i (n7080), .o (n7081) );
  buffer buf_n7082( .i (n7081), .o (n7082) );
  buffer buf_n7083( .i (n7082), .o (n7083) );
  buffer buf_n7084( .i (n7083), .o (n7084) );
  buffer buf_n7085( .i (n7084), .o (n7085) );
  buffer buf_n7086( .i (n7085), .o (n7086) );
  buffer buf_n7087( .i (n7086), .o (n7087) );
  buffer buf_n7088( .i (n7087), .o (n7088) );
  buffer buf_n7089( .i (n7088), .o (n7089) );
  buffer buf_n7090( .i (n7089), .o (n7090) );
  buffer buf_n7091( .i (n7090), .o (n7091) );
  buffer buf_n7092( .i (n7091), .o (n7092) );
  buffer buf_n7093( .i (n7092), .o (n7093) );
  buffer buf_n7094( .i (n7093), .o (n7094) );
  buffer buf_n7095( .i (n7094), .o (n7095) );
  buffer buf_n7096( .i (n7095), .o (n7096) );
  buffer buf_n7097( .i (n7096), .o (n7097) );
  buffer buf_n7098( .i (n7097), .o (n7098) );
  buffer buf_n7099( .i (n7098), .o (n7099) );
  buffer buf_n7100( .i (n7099), .o (n7100) );
  buffer buf_n7101( .i (n7100), .o (n7101) );
  buffer buf_n7102( .i (n7101), .o (n7102) );
  buffer buf_n7103( .i (n7102), .o (n7103) );
  buffer buf_n7104( .i (n7103), .o (n7104) );
  buffer buf_n7105( .i (n7104), .o (n7105) );
  buffer buf_n7106( .i (n7105), .o (n7106) );
  buffer buf_n7107( .i (n7106), .o (n7107) );
  buffer buf_n7108( .i (n7107), .o (n7108) );
  buffer buf_n7109( .i (n7108), .o (n7109) );
  buffer buf_n7110( .i (n7109), .o (n7110) );
  buffer buf_n7111( .i (n7110), .o (n7111) );
  buffer buf_n7112( .i (n7111), .o (n7112) );
  buffer buf_n7113( .i (n7112), .o (n7113) );
  buffer buf_n7114( .i (n7113), .o (n7114) );
  buffer buf_n7115( .i (n7114), .o (n7115) );
  buffer buf_n7116( .i (n7115), .o (n7116) );
  buffer buf_n7117( .i (n7116), .o (n7117) );
  buffer buf_n7118( .i (n7117), .o (n7118) );
  buffer buf_n7119( .i (n7118), .o (n7119) );
  buffer buf_n7120( .i (n7119), .o (n7120) );
  buffer buf_n7121( .i (n7120), .o (n7121) );
  buffer buf_n7122( .i (n7121), .o (n7122) );
  buffer buf_n7123( .i (n7122), .o (n7123) );
  buffer buf_n7124( .i (n7123), .o (n7124) );
  buffer buf_n7125( .i (n7124), .o (n7125) );
  buffer buf_n7126( .i (n7125), .o (n7126) );
  buffer buf_n7127( .i (n7126), .o (n7127) );
  buffer buf_n7128( .i (n7127), .o (n7128) );
  buffer buf_n7129( .i (n7128), .o (n7129) );
  buffer buf_n7130( .i (n7129), .o (n7130) );
  buffer buf_n7131( .i (n7130), .o (n7131) );
  buffer buf_n7132( .i (n7131), .o (n7132) );
  buffer buf_n7133( .i (n7132), .o (n7133) );
  buffer buf_n7134( .i (n7133), .o (n7134) );
  buffer buf_n7135( .i (n7134), .o (n7135) );
  buffer buf_n1971( .i (n1970), .o (n1971) );
  buffer buf_n1972( .i (n1971), .o (n1972) );
  buffer buf_n1973( .i (n1972), .o (n1973) );
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  buffer buf_n1983( .i (n1982), .o (n1983) );
  buffer buf_n1984( .i (n1983), .o (n1984) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n1986( .i (n1985), .o (n1986) );
  buffer buf_n1987( .i (n1986), .o (n1987) );
  buffer buf_n1988( .i (n1987), .o (n1988) );
  buffer buf_n1989( .i (n1988), .o (n1989) );
  buffer buf_n1990( .i (n1989), .o (n1990) );
  buffer buf_n1991( .i (n1990), .o (n1991) );
  buffer buf_n1992( .i (n1991), .o (n1992) );
  buffer buf_n1993( .i (n1992), .o (n1993) );
  buffer buf_n1994( .i (n1993), .o (n1994) );
  buffer buf_n1995( .i (n1994), .o (n1995) );
  buffer buf_n1996( .i (n1995), .o (n1996) );
  buffer buf_n1997( .i (n1996), .o (n1997) );
  buffer buf_n1998( .i (n1997), .o (n1998) );
  buffer buf_n1999( .i (n1998), .o (n1999) );
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n2001( .i (n2000), .o (n2001) );
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n2003), .o (n2004) );
  buffer buf_n2005( .i (n2004), .o (n2005) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n2007( .i (n2006), .o (n2007) );
  buffer buf_n2008( .i (n2007), .o (n2008) );
  buffer buf_n2009( .i (n2008), .o (n2009) );
  buffer buf_n2010( .i (n2009), .o (n2010) );
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n2012( .i (n2011), .o (n2012) );
  buffer buf_n2013( .i (n2012), .o (n2013) );
  buffer buf_n2014( .i (n2013), .o (n2014) );
  buffer buf_n2015( .i (n2014), .o (n2015) );
  buffer buf_n2016( .i (n2015), .o (n2016) );
  buffer buf_n2017( .i (n2016), .o (n2017) );
  buffer buf_n2018( .i (n2017), .o (n2018) );
  buffer buf_n2019( .i (n2018), .o (n2019) );
  buffer buf_n2020( .i (n2019), .o (n2020) );
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2028( .i (n2027), .o (n2028) );
  buffer buf_n2029( .i (n2028), .o (n2029) );
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n2031( .i (n2030), .o (n2031) );
  buffer buf_n2032( .i (n2031), .o (n2032) );
  buffer buf_n2033( .i (n2032), .o (n2033) );
  buffer buf_n2034( .i (n2033), .o (n2034) );
  buffer buf_n2035( .i (n2034), .o (n2035) );
  buffer buf_n2036( .i (n2035), .o (n2036) );
  buffer buf_n2037( .i (n2036), .o (n2037) );
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n5471( .i (n5470), .o (n5471) );
  assign n7138 = n5473 & n5546 ;
  assign n7139 = n5471 | n7138 ;
  buffer buf_n7140( .i (n7139), .o (n7140) );
  assign n7141 = n2052 & n7140 ;
  buffer buf_n7142( .i (n7141), .o (n7142) );
  assign n7143 = n7135 | n7142 ;
  assign n7144 = n2052 | n7140 ;
  buffer buf_n7145( .i (n7144), .o (n7145) );
  buffer buf_n7146( .i (n7145), .o (n7146) );
  assign n7147 = n7143 & n7146 ;
  buffer buf_n7148( .i (n7147), .o (n7148) );
  assign n7149 = n3866 | n7148 ;
  buffer buf_n7150( .i (n7149), .o (n7150) );
  assign n7151 = n7061 & n7150 ;
  assign n7152 = n3866 & n7148 ;
  buffer buf_n7153( .i (n7152), .o (n7153) );
  buffer buf_n7154( .i (n7153), .o (n7154) );
  assign n7155 = n7151 | n7154 ;
  buffer buf_n7156( .i (n7155), .o (n7156) );
  assign n7157 = n1270 & n7156 ;
  buffer buf_n7158( .i (n7157), .o (n7158) );
  buffer buf_n7159( .i (n7158), .o (n7159) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  assign n7160 = n3920 & n6789 ;
  buffer buf_n7161( .i (n7160), .o (n7161) );
  assign n7162 = ~n1027 & n7161 ;
  assign n7163 = n1027 & ~n7161 ;
  assign n7164 = n7162 | n7163 ;
  buffer buf_n7165( .i (n7164), .o (n7165) );
  buffer buf_n7166( .i (n7165), .o (n7166) );
  buffer buf_n7167( .i (n7166), .o (n7167) );
  buffer buf_n7168( .i (n7167), .o (n7168) );
  buffer buf_n7169( .i (n7168), .o (n7169) );
  buffer buf_n7170( .i (n7169), .o (n7170) );
  buffer buf_n7171( .i (n7170), .o (n7171) );
  buffer buf_n7172( .i (n7171), .o (n7172) );
  buffer buf_n7173( .i (n7172), .o (n7173) );
  buffer buf_n7174( .i (n7173), .o (n7174) );
  buffer buf_n7175( .i (n7174), .o (n7175) );
  buffer buf_n7176( .i (n7175), .o (n7176) );
  buffer buf_n7177( .i (n7176), .o (n7177) );
  buffer buf_n7178( .i (n7177), .o (n7178) );
  buffer buf_n7179( .i (n7178), .o (n7179) );
  buffer buf_n7180( .i (n7179), .o (n7180) );
  buffer buf_n7181( .i (n7180), .o (n7181) );
  buffer buf_n7182( .i (n7181), .o (n7182) );
  buffer buf_n7183( .i (n7182), .o (n7183) );
  buffer buf_n7184( .i (n7183), .o (n7184) );
  buffer buf_n7185( .i (n7184), .o (n7185) );
  buffer buf_n7186( .i (n7185), .o (n7186) );
  buffer buf_n7187( .i (n7186), .o (n7187) );
  buffer buf_n7188( .i (n7187), .o (n7188) );
  buffer buf_n7189( .i (n7188), .o (n7189) );
  buffer buf_n7190( .i (n7189), .o (n7190) );
  buffer buf_n7191( .i (n7190), .o (n7191) );
  buffer buf_n7192( .i (n7191), .o (n7192) );
  buffer buf_n7193( .i (n7192), .o (n7193) );
  buffer buf_n7194( .i (n7193), .o (n7194) );
  buffer buf_n7195( .i (n7194), .o (n7195) );
  buffer buf_n7196( .i (n7195), .o (n7196) );
  buffer buf_n7197( .i (n7196), .o (n7197) );
  buffer buf_n7198( .i (n7197), .o (n7198) );
  buffer buf_n7199( .i (n7198), .o (n7199) );
  buffer buf_n7200( .i (n7199), .o (n7200) );
  buffer buf_n7201( .i (n7200), .o (n7201) );
  buffer buf_n7202( .i (n7201), .o (n7202) );
  buffer buf_n7203( .i (n7202), .o (n7203) );
  buffer buf_n7204( .i (n7203), .o (n7204) );
  buffer buf_n7205( .i (n7204), .o (n7205) );
  buffer buf_n7206( .i (n7205), .o (n7206) );
  buffer buf_n7207( .i (n7206), .o (n7207) );
  buffer buf_n7208( .i (n7207), .o (n7208) );
  buffer buf_n7209( .i (n7208), .o (n7209) );
  buffer buf_n7210( .i (n7209), .o (n7210) );
  buffer buf_n7211( .i (n7210), .o (n7211) );
  buffer buf_n7212( .i (n7211), .o (n7212) );
  buffer buf_n7213( .i (n7212), .o (n7213) );
  buffer buf_n7214( .i (n7213), .o (n7214) );
  buffer buf_n7215( .i (n7214), .o (n7215) );
  buffer buf_n7216( .i (n7215), .o (n7216) );
  buffer buf_n7217( .i (n7216), .o (n7217) );
  buffer buf_n7218( .i (n7217), .o (n7218) );
  buffer buf_n7219( .i (n7218), .o (n7219) );
  buffer buf_n7220( .i (n7219), .o (n7220) );
  buffer buf_n7221( .i (n7220), .o (n7221) );
  buffer buf_n7222( .i (n7221), .o (n7222) );
  buffer buf_n7223( .i (n7222), .o (n7223) );
  buffer buf_n7224( .i (n7223), .o (n7224) );
  buffer buf_n7225( .i (n7224), .o (n7225) );
  buffer buf_n7226( .i (n7225), .o (n7226) );
  buffer buf_n7227( .i (n7226), .o (n7227) );
  buffer buf_n7228( .i (n7227), .o (n7228) );
  buffer buf_n7229( .i (n7228), .o (n7229) );
  buffer buf_n7230( .i (n7229), .o (n7230) );
  buffer buf_n7231( .i (n7230), .o (n7231) );
  buffer buf_n7232( .i (n7231), .o (n7232) );
  buffer buf_n7233( .i (n7232), .o (n7233) );
  buffer buf_n7234( .i (n7233), .o (n7234) );
  buffer buf_n7235( .i (n7234), .o (n7235) );
  buffer buf_n7236( .i (n7235), .o (n7236) );
  buffer buf_n7237( .i (n7236), .o (n7237) );
  assign n7240 = n1270 | n7156 ;
  buffer buf_n7241( .i (n7240), .o (n7241) );
  assign n7242 = n7237 & n7241 ;
  assign n7243 = n7159 | n7242 ;
  buffer buf_n7244( .i (n7243), .o (n7244) );
  assign n7245 = n4185 | n7244 ;
  buffer buf_n7246( .i (n7245), .o (n7246) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  assign n7247 = n3922 & n6791 ;
  buffer buf_n7248( .i (n7247), .o (n7248) );
  assign n7249 = n289 | n7248 ;
  assign n7250 = n289 & n7248 ;
  assign n7251 = n7249 & ~n7250 ;
  buffer buf_n7252( .i (n7251), .o (n7252) );
  buffer buf_n7253( .i (n7252), .o (n7253) );
  buffer buf_n7254( .i (n7253), .o (n7254) );
  buffer buf_n7255( .i (n7254), .o (n7255) );
  buffer buf_n7256( .i (n7255), .o (n7256) );
  buffer buf_n7257( .i (n7256), .o (n7257) );
  buffer buf_n7258( .i (n7257), .o (n7258) );
  buffer buf_n7259( .i (n7258), .o (n7259) );
  buffer buf_n7260( .i (n7259), .o (n7260) );
  buffer buf_n7261( .i (n7260), .o (n7261) );
  buffer buf_n7262( .i (n7261), .o (n7262) );
  buffer buf_n7263( .i (n7262), .o (n7263) );
  buffer buf_n7264( .i (n7263), .o (n7264) );
  buffer buf_n7265( .i (n7264), .o (n7265) );
  buffer buf_n7266( .i (n7265), .o (n7266) );
  buffer buf_n7267( .i (n7266), .o (n7267) );
  buffer buf_n7268( .i (n7267), .o (n7268) );
  buffer buf_n7269( .i (n7268), .o (n7269) );
  buffer buf_n7270( .i (n7269), .o (n7270) );
  buffer buf_n7271( .i (n7270), .o (n7271) );
  buffer buf_n7272( .i (n7271), .o (n7272) );
  buffer buf_n7273( .i (n7272), .o (n7273) );
  buffer buf_n7274( .i (n7273), .o (n7274) );
  buffer buf_n7275( .i (n7274), .o (n7275) );
  buffer buf_n7276( .i (n7275), .o (n7276) );
  buffer buf_n7277( .i (n7276), .o (n7277) );
  buffer buf_n7278( .i (n7277), .o (n7278) );
  buffer buf_n7279( .i (n7278), .o (n7279) );
  buffer buf_n7280( .i (n7279), .o (n7280) );
  buffer buf_n7281( .i (n7280), .o (n7281) );
  buffer buf_n7282( .i (n7281), .o (n7282) );
  buffer buf_n7283( .i (n7282), .o (n7283) );
  buffer buf_n7284( .i (n7283), .o (n7284) );
  buffer buf_n7285( .i (n7284), .o (n7285) );
  buffer buf_n7286( .i (n7285), .o (n7286) );
  buffer buf_n7287( .i (n7286), .o (n7287) );
  buffer buf_n7288( .i (n7287), .o (n7288) );
  buffer buf_n7289( .i (n7288), .o (n7289) );
  buffer buf_n7290( .i (n7289), .o (n7290) );
  buffer buf_n7291( .i (n7290), .o (n7291) );
  buffer buf_n7292( .i (n7291), .o (n7292) );
  buffer buf_n7293( .i (n7292), .o (n7293) );
  buffer buf_n7294( .i (n7293), .o (n7294) );
  buffer buf_n7295( .i (n7294), .o (n7295) );
  buffer buf_n7296( .i (n7295), .o (n7296) );
  buffer buf_n7297( .i (n7296), .o (n7297) );
  buffer buf_n7298( .i (n7297), .o (n7298) );
  buffer buf_n7299( .i (n7298), .o (n7299) );
  buffer buf_n7300( .i (n7299), .o (n7300) );
  buffer buf_n7301( .i (n7300), .o (n7301) );
  buffer buf_n7302( .i (n7301), .o (n7302) );
  buffer buf_n7303( .i (n7302), .o (n7303) );
  buffer buf_n7304( .i (n7303), .o (n7304) );
  buffer buf_n7305( .i (n7304), .o (n7305) );
  buffer buf_n7306( .i (n7305), .o (n7306) );
  buffer buf_n7307( .i (n7306), .o (n7307) );
  buffer buf_n7308( .i (n7307), .o (n7308) );
  buffer buf_n7309( .i (n7308), .o (n7309) );
  buffer buf_n7310( .i (n7309), .o (n7310) );
  buffer buf_n7311( .i (n7310), .o (n7311) );
  buffer buf_n7312( .i (n7311), .o (n7312) );
  buffer buf_n7313( .i (n7312), .o (n7313) );
  buffer buf_n7314( .i (n7313), .o (n7314) );
  buffer buf_n7315( .i (n7314), .o (n7315) );
  buffer buf_n7316( .i (n7315), .o (n7316) );
  buffer buf_n7317( .i (n7316), .o (n7317) );
  buffer buf_n7318( .i (n7317), .o (n7318) );
  buffer buf_n7319( .i (n7318), .o (n7319) );
  buffer buf_n7320( .i (n7319), .o (n7320) );
  buffer buf_n7321( .i (n7320), .o (n7321) );
  buffer buf_n7322( .i (n7321), .o (n7322) );
  buffer buf_n7323( .i (n7322), .o (n7323) );
  buffer buf_n7324( .i (n7323), .o (n7324) );
  buffer buf_n7325( .i (n7324), .o (n7325) );
  buffer buf_n7326( .i (n7325), .o (n7326) );
  buffer buf_n7327( .i (n7326), .o (n7327) );
  assign n7330 = n7246 & n7327 ;
  assign n7331 = n4185 & n7244 ;
  buffer buf_n7332( .i (n7331), .o (n7332) );
  buffer buf_n7333( .i (n7332), .o (n7333) );
  assign n7334 = n7330 | n7333 ;
  buffer buf_n7335( .i (n7334), .o (n7335) );
  assign n7336 = n3703 | n7335 ;
  buffer buf_n7337( .i (n7336), .o (n7337) );
  buffer buf_n7338( .i (n7337), .o (n7338) );
  buffer buf_n7339( .i (n7338), .o (n7339) );
  assign n7340 = n3703 & n7335 ;
  buffer buf_n7341( .i (n7340), .o (n7341) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  assign n7343 = n3924 & n6793 ;
  buffer buf_n7344( .i (n7343), .o (n7344) );
  assign n7345 = n910 & ~n7344 ;
  assign n7346 = ~n910 & n7344 ;
  assign n7347 = n7345 | n7346 ;
  buffer buf_n7348( .i (n7347), .o (n7348) );
  buffer buf_n7349( .i (n7348), .o (n7349) );
  buffer buf_n7350( .i (n7349), .o (n7350) );
  buffer buf_n7351( .i (n7350), .o (n7351) );
  buffer buf_n7352( .i (n7351), .o (n7352) );
  buffer buf_n7353( .i (n7352), .o (n7353) );
  buffer buf_n7354( .i (n7353), .o (n7354) );
  buffer buf_n7355( .i (n7354), .o (n7355) );
  buffer buf_n7356( .i (n7355), .o (n7356) );
  buffer buf_n7357( .i (n7356), .o (n7357) );
  buffer buf_n7358( .i (n7357), .o (n7358) );
  buffer buf_n7359( .i (n7358), .o (n7359) );
  buffer buf_n7360( .i (n7359), .o (n7360) );
  buffer buf_n7361( .i (n7360), .o (n7361) );
  buffer buf_n7362( .i (n7361), .o (n7362) );
  buffer buf_n7363( .i (n7362), .o (n7363) );
  buffer buf_n7364( .i (n7363), .o (n7364) );
  buffer buf_n7365( .i (n7364), .o (n7365) );
  buffer buf_n7366( .i (n7365), .o (n7366) );
  buffer buf_n7367( .i (n7366), .o (n7367) );
  buffer buf_n7368( .i (n7367), .o (n7368) );
  buffer buf_n7369( .i (n7368), .o (n7369) );
  buffer buf_n7370( .i (n7369), .o (n7370) );
  buffer buf_n7371( .i (n7370), .o (n7371) );
  buffer buf_n7372( .i (n7371), .o (n7372) );
  buffer buf_n7373( .i (n7372), .o (n7373) );
  buffer buf_n7374( .i (n7373), .o (n7374) );
  buffer buf_n7375( .i (n7374), .o (n7375) );
  buffer buf_n7376( .i (n7375), .o (n7376) );
  buffer buf_n7377( .i (n7376), .o (n7377) );
  buffer buf_n7378( .i (n7377), .o (n7378) );
  buffer buf_n7379( .i (n7378), .o (n7379) );
  buffer buf_n7380( .i (n7379), .o (n7380) );
  buffer buf_n7381( .i (n7380), .o (n7381) );
  buffer buf_n7382( .i (n7381), .o (n7382) );
  buffer buf_n7383( .i (n7382), .o (n7383) );
  buffer buf_n7384( .i (n7383), .o (n7384) );
  buffer buf_n7385( .i (n7384), .o (n7385) );
  buffer buf_n7386( .i (n7385), .o (n7386) );
  buffer buf_n7387( .i (n7386), .o (n7387) );
  buffer buf_n7388( .i (n7387), .o (n7388) );
  buffer buf_n7389( .i (n7388), .o (n7389) );
  buffer buf_n7390( .i (n7389), .o (n7390) );
  buffer buf_n7391( .i (n7390), .o (n7391) );
  buffer buf_n7392( .i (n7391), .o (n7392) );
  buffer buf_n7393( .i (n7392), .o (n7393) );
  buffer buf_n7394( .i (n7393), .o (n7394) );
  buffer buf_n7395( .i (n7394), .o (n7395) );
  buffer buf_n7396( .i (n7395), .o (n7396) );
  buffer buf_n7397( .i (n7396), .o (n7397) );
  buffer buf_n7398( .i (n7397), .o (n7398) );
  buffer buf_n7399( .i (n7398), .o (n7399) );
  buffer buf_n7400( .i (n7399), .o (n7400) );
  buffer buf_n7401( .i (n7400), .o (n7401) );
  buffer buf_n7402( .i (n7401), .o (n7402) );
  buffer buf_n7403( .i (n7402), .o (n7403) );
  buffer buf_n7404( .i (n7403), .o (n7404) );
  buffer buf_n7405( .i (n7404), .o (n7405) );
  buffer buf_n7406( .i (n7405), .o (n7406) );
  buffer buf_n7407( .i (n7406), .o (n7407) );
  buffer buf_n7408( .i (n7407), .o (n7408) );
  buffer buf_n7409( .i (n7408), .o (n7409) );
  buffer buf_n7410( .i (n7409), .o (n7410) );
  buffer buf_n7411( .i (n7410), .o (n7411) );
  buffer buf_n7412( .i (n7411), .o (n7412) );
  buffer buf_n7413( .i (n7412), .o (n7413) );
  buffer buf_n7414( .i (n7413), .o (n7414) );
  buffer buf_n7415( .i (n7414), .o (n7415) );
  buffer buf_n7416( .i (n7415), .o (n7416) );
  buffer buf_n7417( .i (n7416), .o (n7417) );
  buffer buf_n7418( .i (n7417), .o (n7418) );
  buffer buf_n7419( .i (n7418), .o (n7419) );
  buffer buf_n7420( .i (n7419), .o (n7420) );
  buffer buf_n7421( .i (n7420), .o (n7421) );
  buffer buf_n7422( .i (n7421), .o (n7422) );
  buffer buf_n7423( .i (n7422), .o (n7423) );
  buffer buf_n7424( .i (n7423), .o (n7424) );
  buffer buf_n7425( .i (n7424), .o (n7425) );
  buffer buf_n7426( .i (n7425), .o (n7426) );
  assign n7429 = n7341 | n7426 ;
  buffer buf_n7430( .i (n7429), .o (n7430) );
  assign n7431 = n7339 & n7430 ;
  buffer buf_n7432( .i (n7431), .o (n7432) );
  assign n7433 = n2416 | n7432 ;
  buffer buf_n7434( .i (n7433), .o (n7434) );
  assign n7436 = n6984 & n7434 ;
  buffer buf_n7437( .i (n7436), .o (n7437) );
  assign n7438 = n2416 & n7432 ;
  buffer buf_n7439( .i (n7438), .o (n7439) );
  buffer buf_n7440( .i (n7439), .o (n7440) );
  buffer buf_n7441( .i (n7440), .o (n7441) );
  assign n7442 = n7437 | n7441 ;
  buffer buf_n7443( .i (n7442), .o (n7443) );
  assign n7444 = n3108 & n7443 ;
  buffer buf_n7445( .i (n7444), .o (n7445) );
  assign n7446 = n2720 & n6800 ;
  buffer buf_n7447( .i (n7446), .o (n7447) );
  assign n7448 = n6802 & ~n7447 ;
  buffer buf_n7449( .i (n7448), .o (n7449) );
  buffer buf_n7450( .i (n7449), .o (n7450) );
  buffer buf_n7451( .i (n7450), .o (n7451) );
  buffer buf_n7452( .i (n7451), .o (n7452) );
  buffer buf_n7453( .i (n7452), .o (n7453) );
  buffer buf_n7454( .i (n7453), .o (n7454) );
  buffer buf_n7455( .i (n7454), .o (n7455) );
  buffer buf_n7456( .i (n7455), .o (n7456) );
  buffer buf_n7457( .i (n7456), .o (n7457) );
  buffer buf_n7458( .i (n7457), .o (n7458) );
  buffer buf_n7459( .i (n7458), .o (n7459) );
  buffer buf_n7460( .i (n7459), .o (n7460) );
  buffer buf_n7461( .i (n7460), .o (n7461) );
  buffer buf_n7462( .i (n7461), .o (n7462) );
  buffer buf_n7463( .i (n7462), .o (n7463) );
  buffer buf_n7464( .i (n7463), .o (n7464) );
  buffer buf_n7465( .i (n7464), .o (n7465) );
  buffer buf_n7466( .i (n7465), .o (n7466) );
  buffer buf_n7467( .i (n7466), .o (n7467) );
  buffer buf_n7468( .i (n7467), .o (n7468) );
  buffer buf_n7469( .i (n7468), .o (n7469) );
  buffer buf_n7470( .i (n7469), .o (n7470) );
  buffer buf_n7471( .i (n7470), .o (n7471) );
  buffer buf_n7472( .i (n7471), .o (n7472) );
  buffer buf_n7473( .i (n7472), .o (n7473) );
  buffer buf_n7474( .i (n7473), .o (n7474) );
  buffer buf_n7475( .i (n7474), .o (n7475) );
  buffer buf_n7476( .i (n7475), .o (n7476) );
  buffer buf_n7477( .i (n7476), .o (n7477) );
  buffer buf_n7478( .i (n7477), .o (n7478) );
  buffer buf_n7479( .i (n7478), .o (n7479) );
  buffer buf_n7480( .i (n7479), .o (n7480) );
  buffer buf_n7481( .i (n7480), .o (n7481) );
  buffer buf_n7482( .i (n7481), .o (n7482) );
  buffer buf_n7483( .i (n7482), .o (n7483) );
  buffer buf_n7484( .i (n7483), .o (n7484) );
  buffer buf_n7485( .i (n7484), .o (n7485) );
  buffer buf_n7486( .i (n7485), .o (n7486) );
  buffer buf_n7487( .i (n7486), .o (n7487) );
  buffer buf_n7488( .i (n7487), .o (n7488) );
  buffer buf_n7489( .i (n7488), .o (n7489) );
  buffer buf_n7490( .i (n7489), .o (n7490) );
  buffer buf_n7491( .i (n7490), .o (n7491) );
  buffer buf_n7492( .i (n7491), .o (n7492) );
  buffer buf_n7493( .i (n7492), .o (n7493) );
  buffer buf_n7494( .i (n7493), .o (n7494) );
  buffer buf_n7495( .i (n7494), .o (n7495) );
  buffer buf_n7496( .i (n7495), .o (n7496) );
  buffer buf_n7497( .i (n7496), .o (n7497) );
  buffer buf_n7498( .i (n7497), .o (n7498) );
  buffer buf_n7499( .i (n7498), .o (n7499) );
  buffer buf_n7500( .i (n7499), .o (n7500) );
  buffer buf_n7501( .i (n7500), .o (n7501) );
  buffer buf_n7502( .i (n7501), .o (n7502) );
  buffer buf_n7503( .i (n7502), .o (n7503) );
  buffer buf_n7504( .i (n7503), .o (n7504) );
  buffer buf_n7505( .i (n7504), .o (n7505) );
  buffer buf_n7506( .i (n7505), .o (n7506) );
  buffer buf_n7507( .i (n7506), .o (n7507) );
  buffer buf_n7508( .i (n7507), .o (n7508) );
  buffer buf_n7509( .i (n7508), .o (n7509) );
  buffer buf_n7510( .i (n7509), .o (n7510) );
  buffer buf_n7511( .i (n7510), .o (n7511) );
  buffer buf_n7512( .i (n7511), .o (n7512) );
  buffer buf_n7513( .i (n7512), .o (n7513) );
  buffer buf_n7514( .i (n7513), .o (n7514) );
  buffer buf_n7515( .i (n7514), .o (n7515) );
  buffer buf_n7516( .i (n7515), .o (n7516) );
  buffer buf_n7517( .i (n7516), .o (n7517) );
  buffer buf_n7518( .i (n7517), .o (n7518) );
  buffer buf_n7519( .i (n7518), .o (n7519) );
  buffer buf_n7520( .i (n7519), .o (n7520) );
  buffer buf_n7521( .i (n7520), .o (n7521) );
  buffer buf_n7522( .i (n7521), .o (n7522) );
  buffer buf_n7523( .i (n7522), .o (n7523) );
  buffer buf_n7524( .i (n7523), .o (n7524) );
  buffer buf_n7525( .i (n7524), .o (n7525) );
  buffer buf_n7526( .i (n7525), .o (n7526) );
  buffer buf_n7527( .i (n7526), .o (n7527) );
  buffer buf_n7528( .i (n7527), .o (n7528) );
  buffer buf_n7529( .i (n7528), .o (n7529) );
  buffer buf_n7530( .i (n7529), .o (n7530) );
  buffer buf_n7531( .i (n7530), .o (n7531) );
  buffer buf_n7532( .i (n7531), .o (n7532) );
  buffer buf_n7533( .i (n7532), .o (n7533) );
  assign n7536 = n7445 | n7533 ;
  assign n7537 = n3108 | n7443 ;
  buffer buf_n7538( .i (n7537), .o (n7538) );
  buffer buf_n7539( .i (n7538), .o (n7539) );
  assign n7540 = n7536 & n7539 ;
  buffer buf_n7541( .i (n7540), .o (n7541) );
  assign n7542 = n3434 & n7541 ;
  buffer buf_n7543( .i (n7542), .o (n7543) );
  buffer buf_n7544( .i (n7543), .o (n7544) );
  buffer buf_n7545( .i (n7544), .o (n7545) );
  assign n7546 = n3434 | n7541 ;
  buffer buf_n7547( .i (n7546), .o (n7547) );
  buffer buf_n3231( .i (n3230), .o (n3231) );
  assign n7549 = n3231 & n6804 ;
  assign n7550 = n3231 | n6804 ;
  assign n7551 = ~n7549 & n7550 ;
  buffer buf_n7552( .i (n7551), .o (n7552) );
  buffer buf_n7553( .i (n7552), .o (n7553) );
  buffer buf_n7554( .i (n7553), .o (n7554) );
  buffer buf_n7555( .i (n7554), .o (n7555) );
  buffer buf_n7556( .i (n7555), .o (n7556) );
  buffer buf_n7557( .i (n7556), .o (n7557) );
  buffer buf_n7558( .i (n7557), .o (n7558) );
  buffer buf_n7559( .i (n7558), .o (n7559) );
  buffer buf_n7560( .i (n7559), .o (n7560) );
  buffer buf_n7561( .i (n7560), .o (n7561) );
  buffer buf_n7562( .i (n7561), .o (n7562) );
  buffer buf_n7563( .i (n7562), .o (n7563) );
  buffer buf_n7564( .i (n7563), .o (n7564) );
  buffer buf_n7565( .i (n7564), .o (n7565) );
  buffer buf_n7566( .i (n7565), .o (n7566) );
  buffer buf_n7567( .i (n7566), .o (n7567) );
  buffer buf_n7568( .i (n7567), .o (n7568) );
  buffer buf_n7569( .i (n7568), .o (n7569) );
  buffer buf_n7570( .i (n7569), .o (n7570) );
  buffer buf_n7571( .i (n7570), .o (n7571) );
  buffer buf_n7572( .i (n7571), .o (n7572) );
  buffer buf_n7573( .i (n7572), .o (n7573) );
  buffer buf_n7574( .i (n7573), .o (n7574) );
  buffer buf_n7575( .i (n7574), .o (n7575) );
  buffer buf_n7576( .i (n7575), .o (n7576) );
  buffer buf_n7577( .i (n7576), .o (n7577) );
  buffer buf_n7578( .i (n7577), .o (n7578) );
  buffer buf_n7579( .i (n7578), .o (n7579) );
  buffer buf_n7580( .i (n7579), .o (n7580) );
  buffer buf_n7581( .i (n7580), .o (n7581) );
  buffer buf_n7582( .i (n7581), .o (n7582) );
  buffer buf_n7583( .i (n7582), .o (n7583) );
  buffer buf_n7584( .i (n7583), .o (n7584) );
  buffer buf_n7585( .i (n7584), .o (n7585) );
  buffer buf_n7586( .i (n7585), .o (n7586) );
  buffer buf_n7587( .i (n7586), .o (n7587) );
  buffer buf_n7588( .i (n7587), .o (n7588) );
  buffer buf_n7589( .i (n7588), .o (n7589) );
  buffer buf_n7590( .i (n7589), .o (n7590) );
  buffer buf_n7591( .i (n7590), .o (n7591) );
  buffer buf_n7592( .i (n7591), .o (n7592) );
  buffer buf_n7593( .i (n7592), .o (n7593) );
  buffer buf_n7594( .i (n7593), .o (n7594) );
  buffer buf_n7595( .i (n7594), .o (n7595) );
  buffer buf_n7596( .i (n7595), .o (n7596) );
  buffer buf_n7597( .i (n7596), .o (n7597) );
  buffer buf_n7598( .i (n7597), .o (n7598) );
  buffer buf_n7599( .i (n7598), .o (n7599) );
  buffer buf_n7600( .i (n7599), .o (n7600) );
  buffer buf_n7601( .i (n7600), .o (n7601) );
  buffer buf_n7602( .i (n7601), .o (n7602) );
  buffer buf_n7603( .i (n7602), .o (n7603) );
  buffer buf_n7604( .i (n7603), .o (n7604) );
  buffer buf_n7605( .i (n7604), .o (n7605) );
  buffer buf_n7606( .i (n7605), .o (n7606) );
  buffer buf_n7607( .i (n7606), .o (n7607) );
  buffer buf_n7608( .i (n7607), .o (n7608) );
  buffer buf_n7609( .i (n7608), .o (n7609) );
  buffer buf_n7610( .i (n7609), .o (n7610) );
  buffer buf_n7611( .i (n7610), .o (n7611) );
  buffer buf_n7612( .i (n7611), .o (n7612) );
  buffer buf_n7613( .i (n7612), .o (n7613) );
  buffer buf_n7614( .i (n7613), .o (n7614) );
  buffer buf_n7615( .i (n7614), .o (n7615) );
  buffer buf_n7616( .i (n7615), .o (n7616) );
  buffer buf_n7617( .i (n7616), .o (n7617) );
  buffer buf_n7618( .i (n7617), .o (n7618) );
  buffer buf_n7619( .i (n7618), .o (n7619) );
  buffer buf_n7620( .i (n7619), .o (n7620) );
  buffer buf_n7621( .i (n7620), .o (n7621) );
  buffer buf_n7622( .i (n7621), .o (n7622) );
  buffer buf_n7623( .i (n7622), .o (n7623) );
  buffer buf_n7624( .i (n7623), .o (n7624) );
  buffer buf_n7625( .i (n7624), .o (n7625) );
  buffer buf_n7626( .i (n7625), .o (n7626) );
  buffer buf_n7627( .i (n7626), .o (n7627) );
  buffer buf_n7628( .i (n7627), .o (n7628) );
  buffer buf_n7629( .i (n7628), .o (n7629) );
  buffer buf_n7630( .i (n7629), .o (n7630) );
  buffer buf_n7631( .i (n7630), .o (n7631) );
  buffer buf_n7632( .i (n7631), .o (n7632) );
  buffer buf_n7633( .i (n7632), .o (n7633) );
  buffer buf_n7634( .i (n7633), .o (n7634) );
  buffer buf_n7635( .i (n7634), .o (n7635) );
  buffer buf_n7636( .i (n7635), .o (n7636) );
  buffer buf_n7637( .i (n7636), .o (n7637) );
  buffer buf_n7638( .i (n7637), .o (n7638) );
  assign n7641 = n7547 & n7638 ;
  buffer buf_n7642( .i (n7641), .o (n7642) );
  assign n7643 = n7545 | n7642 ;
  buffer buf_n7644( .i (n7643), .o (n7644) );
  assign n7645 = n6898 | n7644 ;
  assign n7646 = n2529 | n6810 ;
  buffer buf_n7647( .i (n7646), .o (n7647) );
  buffer buf_n7648( .i (n7647), .o (n7648) );
  buffer buf_n7649( .i (n7648), .o (n7649) );
  buffer buf_n7650( .i (n7649), .o (n7650) );
  buffer buf_n7651( .i (n7650), .o (n7651) );
  buffer buf_n7652( .i (n7651), .o (n7652) );
  buffer buf_n7653( .i (n7652), .o (n7653) );
  buffer buf_n7654( .i (n7653), .o (n7654) );
  buffer buf_n7655( .i (n7654), .o (n7655) );
  buffer buf_n7656( .i (n7655), .o (n7656) );
  buffer buf_n7657( .i (n7656), .o (n7657) );
  buffer buf_n7658( .i (n7657), .o (n7658) );
  buffer buf_n7659( .i (n7658), .o (n7659) );
  buffer buf_n7660( .i (n7659), .o (n7660) );
  buffer buf_n7661( .i (n7660), .o (n7661) );
  buffer buf_n7662( .i (n7661), .o (n7662) );
  buffer buf_n7663( .i (n7662), .o (n7663) );
  buffer buf_n7664( .i (n7663), .o (n7664) );
  buffer buf_n7665( .i (n7664), .o (n7665) );
  buffer buf_n7666( .i (n7665), .o (n7666) );
  buffer buf_n7667( .i (n7666), .o (n7667) );
  buffer buf_n7668( .i (n7667), .o (n7668) );
  buffer buf_n7669( .i (n7668), .o (n7669) );
  buffer buf_n7670( .i (n7669), .o (n7670) );
  buffer buf_n7671( .i (n7670), .o (n7671) );
  buffer buf_n7672( .i (n7671), .o (n7672) );
  buffer buf_n7673( .i (n7672), .o (n7673) );
  buffer buf_n7674( .i (n7673), .o (n7674) );
  buffer buf_n7675( .i (n7674), .o (n7675) );
  buffer buf_n7676( .i (n7675), .o (n7676) );
  buffer buf_n7677( .i (n7676), .o (n7677) );
  buffer buf_n7678( .i (n7677), .o (n7678) );
  buffer buf_n7679( .i (n7678), .o (n7679) );
  buffer buf_n7680( .i (n7679), .o (n7680) );
  buffer buf_n7681( .i (n7680), .o (n7681) );
  buffer buf_n7682( .i (n7681), .o (n7682) );
  buffer buf_n7683( .i (n7682), .o (n7683) );
  buffer buf_n7684( .i (n7683), .o (n7684) );
  buffer buf_n7685( .i (n7684), .o (n7685) );
  buffer buf_n7686( .i (n7685), .o (n7686) );
  buffer buf_n7687( .i (n7686), .o (n7687) );
  buffer buf_n7688( .i (n7687), .o (n7688) );
  buffer buf_n7689( .i (n7688), .o (n7689) );
  buffer buf_n7690( .i (n7689), .o (n7690) );
  buffer buf_n7691( .i (n7690), .o (n7691) );
  buffer buf_n7692( .i (n7691), .o (n7692) );
  buffer buf_n7693( .i (n7692), .o (n7693) );
  buffer buf_n7694( .i (n7693), .o (n7694) );
  buffer buf_n7695( .i (n7694), .o (n7695) );
  buffer buf_n7696( .i (n7695), .o (n7696) );
  buffer buf_n7697( .i (n7696), .o (n7697) );
  buffer buf_n7698( .i (n7697), .o (n7698) );
  buffer buf_n7699( .i (n7698), .o (n7699) );
  buffer buf_n7700( .i (n7699), .o (n7700) );
  buffer buf_n7701( .i (n7700), .o (n7701) );
  buffer buf_n7702( .i (n7701), .o (n7702) );
  buffer buf_n7703( .i (n7702), .o (n7703) );
  buffer buf_n7704( .i (n7703), .o (n7704) );
  buffer buf_n7705( .i (n7704), .o (n7705) );
  buffer buf_n7706( .i (n7705), .o (n7706) );
  buffer buf_n7707( .i (n7706), .o (n7707) );
  buffer buf_n7708( .i (n7707), .o (n7708) );
  buffer buf_n7709( .i (n7708), .o (n7709) );
  buffer buf_n7710( .i (n7709), .o (n7710) );
  buffer buf_n7711( .i (n7710), .o (n7711) );
  buffer buf_n7712( .i (n7711), .o (n7712) );
  buffer buf_n7713( .i (n7712), .o (n7713) );
  buffer buf_n7714( .i (n7713), .o (n7714) );
  buffer buf_n7715( .i (n7714), .o (n7715) );
  buffer buf_n7716( .i (n7715), .o (n7716) );
  buffer buf_n7717( .i (n7716), .o (n7717) );
  buffer buf_n7718( .i (n7717), .o (n7718) );
  buffer buf_n7719( .i (n7718), .o (n7719) );
  buffer buf_n7720( .i (n7719), .o (n7720) );
  buffer buf_n7721( .i (n7720), .o (n7721) );
  buffer buf_n7722( .i (n7721), .o (n7722) );
  buffer buf_n7723( .i (n7722), .o (n7723) );
  buffer buf_n7724( .i (n7723), .o (n7724) );
  buffer buf_n7725( .i (n7724), .o (n7725) );
  buffer buf_n7726( .i (n7725), .o (n7726) );
  buffer buf_n7727( .i (n7726), .o (n7727) );
  buffer buf_n7728( .i (n7727), .o (n7728) );
  buffer buf_n7729( .i (n7728), .o (n7729) );
  buffer buf_n7730( .i (n7729), .o (n7730) );
  buffer buf_n7731( .i (n7730), .o (n7731) );
  buffer buf_n7732( .i (n7731), .o (n7732) );
  buffer buf_n7733( .i (n7732), .o (n7733) );
  buffer buf_n7734( .i (n7733), .o (n7734) );
  assign n7735 = n7645 & n7734 ;
  buffer buf_n7736( .i (n7735), .o (n7736) );
  buffer buf_n7737( .i (n7736), .o (n7737) );
  buffer buf_n7738( .i (n7737), .o (n7738) );
  buffer buf_n7739( .i (n7738), .o (n7739) );
  buffer buf_n7740( .i (n7739), .o (n7740) );
  buffer buf_n7741( .i (n7740), .o (n7741) );
  buffer buf_n5373( .i (n5372), .o (n5373) );
  buffer buf_n5374( .i (n5373), .o (n5374) );
  assign n7742 = ~n5315 & n5318 ;
  buffer buf_n7743( .i (n7742), .o (n7743) );
  assign n7744 = ~n5374 & n7743 ;
  assign n7745 = n5374 & ~n7743 ;
  assign n7746 = n7744 | n7745 ;
  buffer buf_n7747( .i (n7746), .o (n7747) );
  buffer buf_n7748( .i (n7747), .o (n7748) );
  buffer buf_n7749( .i (n7748), .o (n7749) );
  buffer buf_n7750( .i (n7749), .o (n7750) );
  buffer buf_n7751( .i (n7750), .o (n7751) );
  buffer buf_n7752( .i (n7751), .o (n7752) );
  buffer buf_n7753( .i (n7752), .o (n7753) );
  buffer buf_n7754( .i (n7753), .o (n7754) );
  buffer buf_n7755( .i (n7754), .o (n7755) );
  buffer buf_n7756( .i (n7755), .o (n7756) );
  buffer buf_n7757( .i (n7756), .o (n7757) );
  buffer buf_n7758( .i (n7757), .o (n7758) );
  buffer buf_n7759( .i (n7758), .o (n7759) );
  buffer buf_n7760( .i (n7759), .o (n7760) );
  buffer buf_n7761( .i (n7760), .o (n7761) );
  buffer buf_n7762( .i (n7761), .o (n7762) );
  buffer buf_n7763( .i (n7762), .o (n7763) );
  buffer buf_n7764( .i (n7763), .o (n7764) );
  buffer buf_n7765( .i (n7764), .o (n7765) );
  buffer buf_n7766( .i (n7765), .o (n7766) );
  buffer buf_n7767( .i (n7766), .o (n7767) );
  buffer buf_n7768( .i (n7767), .o (n7768) );
  buffer buf_n7769( .i (n7768), .o (n7769) );
  buffer buf_n7770( .i (n7769), .o (n7770) );
  buffer buf_n7771( .i (n7770), .o (n7771) );
  buffer buf_n7772( .i (n7771), .o (n7772) );
  buffer buf_n7773( .i (n7772), .o (n7773) );
  buffer buf_n7774( .i (n7773), .o (n7774) );
  buffer buf_n7775( .i (n7774), .o (n7775) );
  buffer buf_n7776( .i (n7775), .o (n7776) );
  buffer buf_n7777( .i (n7776), .o (n7777) );
  buffer buf_n7778( .i (n7777), .o (n7778) );
  buffer buf_n7779( .i (n7778), .o (n7779) );
  buffer buf_n7780( .i (n7779), .o (n7780) );
  buffer buf_n7781( .i (n7780), .o (n7781) );
  buffer buf_n7782( .i (n7781), .o (n7782) );
  buffer buf_n7783( .i (n7782), .o (n7783) );
  buffer buf_n7784( .i (n7783), .o (n7784) );
  buffer buf_n7785( .i (n7784), .o (n7785) );
  buffer buf_n7786( .i (n7785), .o (n7786) );
  buffer buf_n7787( .i (n7786), .o (n7787) );
  buffer buf_n7788( .i (n7787), .o (n7788) );
  buffer buf_n7789( .i (n7788), .o (n7789) );
  buffer buf_n7790( .i (n7789), .o (n7790) );
  buffer buf_n7791( .i (n7790), .o (n7791) );
  buffer buf_n7792( .i (n7791), .o (n7792) );
  buffer buf_n7793( .i (n7792), .o (n7793) );
  buffer buf_n7794( .i (n7793), .o (n7794) );
  buffer buf_n7795( .i (n7794), .o (n7795) );
  buffer buf_n7796( .i (n7795), .o (n7796) );
  buffer buf_n7797( .i (n7796), .o (n7797) );
  buffer buf_n7798( .i (n7797), .o (n7798) );
  buffer buf_n7799( .i (n7798), .o (n7799) );
  buffer buf_n7800( .i (n7799), .o (n7800) );
  buffer buf_n7801( .i (n7800), .o (n7801) );
  buffer buf_n7802( .i (n7801), .o (n7802) );
  buffer buf_n7803( .i (n7802), .o (n7803) );
  buffer buf_n7804( .i (n7803), .o (n7804) );
  buffer buf_n7805( .i (n7804), .o (n7805) );
  buffer buf_n7806( .i (n7805), .o (n7806) );
  buffer buf_n7807( .i (n7806), .o (n7807) );
  buffer buf_n7808( .i (n7807), .o (n7808) );
  buffer buf_n7809( .i (n7808), .o (n7809) );
  buffer buf_n7810( .i (n7809), .o (n7810) );
  buffer buf_n7811( .i (n7810), .o (n7811) );
  buffer buf_n7812( .i (n7811), .o (n7812) );
  buffer buf_n7813( .i (n7812), .o (n7813) );
  buffer buf_n7814( .i (n7813), .o (n7814) );
  buffer buf_n7815( .i (n7814), .o (n7815) );
  buffer buf_n7816( .i (n7815), .o (n7816) );
  buffer buf_n7817( .i (n7816), .o (n7817) );
  buffer buf_n7818( .i (n7817), .o (n7818) );
  buffer buf_n7819( .i (n7818), .o (n7819) );
  buffer buf_n7820( .i (n7819), .o (n7820) );
  buffer buf_n7821( .i (n7820), .o (n7821) );
  buffer buf_n7328( .i (n7327), .o (n7328) );
  buffer buf_n7329( .i (n7328), .o (n7329) );
  assign n7822 = n7246 & ~n7332 ;
  buffer buf_n7823( .i (n7822), .o (n7823) );
  assign n7824 = n7329 & ~n7823 ;
  assign n7825 = ~n7329 & n7823 ;
  assign n7826 = n7824 | n7825 ;
  buffer buf_n7827( .i (n7826), .o (n7827) );
  buffer buf_n7828( .i (n7827), .o (n7828) );
  buffer buf_n7829( .i (n7828), .o (n7829) );
  buffer buf_n7830( .i (n7829), .o (n7830) );
  buffer buf_n7831( .i (n7830), .o (n7831) );
  buffer buf_n7832( .i (n7831), .o (n7832) );
  buffer buf_n7833( .i (n7832), .o (n7833) );
  buffer buf_n7834( .i (n7833), .o (n7834) );
  buffer buf_n7835( .i (n7834), .o (n7835) );
  buffer buf_n7836( .i (n7835), .o (n7836) );
  buffer buf_n7837( .i (n7836), .o (n7837) );
  buffer buf_n7838( .i (n7837), .o (n7838) );
  buffer buf_n7839( .i (n7838), .o (n7839) );
  buffer buf_n7840( .i (n7839), .o (n7840) );
  buffer buf_n7841( .i (n7840), .o (n7841) );
  buffer buf_n7842( .i (n7841), .o (n7842) );
  buffer buf_n7843( .i (n7842), .o (n7843) );
  buffer buf_n7844( .i (n7843), .o (n7844) );
  buffer buf_n7845( .i (n7844), .o (n7845) );
  buffer buf_n7846( .i (n7845), .o (n7846) );
  buffer buf_n7847( .i (n7846), .o (n7847) );
  buffer buf_n7848( .i (n7847), .o (n7848) );
  buffer buf_n7849( .i (n7848), .o (n7849) );
  buffer buf_n7850( .i (n7849), .o (n7850) );
  buffer buf_n7851( .i (n7850), .o (n7851) );
  buffer buf_n7852( .i (n7851), .o (n7852) );
  buffer buf_n7853( .i (n7852), .o (n7853) );
  buffer buf_n7854( .i (n7853), .o (n7854) );
  buffer buf_n7855( .i (n7854), .o (n7855) );
  buffer buf_n7856( .i (n7855), .o (n7856) );
  buffer buf_n4844( .i (n4843), .o (n4844) );
  buffer buf_n4845( .i (n4844), .o (n4845) );
  assign n7857 = n4835 & ~n4838 ;
  buffer buf_n7858( .i (n7857), .o (n7858) );
  assign n7859 = n4845 & n7858 ;
  assign n7860 = n4845 | n7858 ;
  assign n7861 = ~n7859 & n7860 ;
  buffer buf_n7862( .i (n7861), .o (n7862) );
  buffer buf_n7863( .i (n7862), .o (n7863) );
  buffer buf_n7864( .i (n7863), .o (n7864) );
  buffer buf_n7865( .i (n7864), .o (n7865) );
  buffer buf_n7866( .i (n7865), .o (n7866) );
  buffer buf_n7867( .i (n7866), .o (n7867) );
  buffer buf_n7868( .i (n7867), .o (n7868) );
  buffer buf_n7869( .i (n7868), .o (n7869) );
  buffer buf_n7870( .i (n7869), .o (n7870) );
  buffer buf_n7871( .i (n7870), .o (n7871) );
  buffer buf_n7872( .i (n7871), .o (n7872) );
  buffer buf_n7873( .i (n7872), .o (n7873) );
  buffer buf_n7874( .i (n7873), .o (n7874) );
  buffer buf_n7875( .i (n7874), .o (n7875) );
  buffer buf_n7876( .i (n7875), .o (n7876) );
  buffer buf_n7877( .i (n7876), .o (n7877) );
  buffer buf_n7878( .i (n7877), .o (n7878) );
  buffer buf_n7879( .i (n7878), .o (n7879) );
  buffer buf_n7880( .i (n7879), .o (n7880) );
  buffer buf_n7881( .i (n7880), .o (n7881) );
  buffer buf_n7882( .i (n7881), .o (n7882) );
  buffer buf_n7883( .i (n7882), .o (n7883) );
  buffer buf_n7884( .i (n7883), .o (n7884) );
  buffer buf_n7885( .i (n7884), .o (n7885) );
  buffer buf_n7886( .i (n7885), .o (n7886) );
  buffer buf_n7887( .i (n7886), .o (n7887) );
  buffer buf_n7888( .i (n7887), .o (n7888) );
  buffer buf_n7889( .i (n7888), .o (n7889) );
  buffer buf_n7890( .i (n7889), .o (n7890) );
  buffer buf_n7891( .i (n7890), .o (n7891) );
  buffer buf_n7892( .i (n7891), .o (n7892) );
  buffer buf_n7893( .i (n7892), .o (n7893) );
  buffer buf_n7894( .i (n7893), .o (n7894) );
  buffer buf_n7895( .i (n7894), .o (n7895) );
  buffer buf_n7896( .i (n7895), .o (n7896) );
  buffer buf_n7897( .i (n7896), .o (n7897) );
  buffer buf_n7898( .i (n7897), .o (n7898) );
  buffer buf_n7899( .i (n7898), .o (n7899) );
  buffer buf_n7900( .i (n7899), .o (n7900) );
  buffer buf_n7901( .i (n7900), .o (n7901) );
  buffer buf_n7902( .i (n7901), .o (n7902) );
  buffer buf_n7903( .i (n7902), .o (n7903) );
  buffer buf_n7904( .i (n7903), .o (n7904) );
  buffer buf_n7905( .i (n7904), .o (n7905) );
  buffer buf_n7906( .i (n7905), .o (n7906) );
  buffer buf_n7907( .i (n7906), .o (n7907) );
  buffer buf_n7908( .i (n7907), .o (n7908) );
  buffer buf_n7909( .i (n7908), .o (n7909) );
  buffer buf_n7910( .i (n7909), .o (n7910) );
  buffer buf_n7911( .i (n7910), .o (n7911) );
  buffer buf_n7912( .i (n7911), .o (n7912) );
  buffer buf_n7913( .i (n7912), .o (n7913) );
  buffer buf_n7914( .i (n7913), .o (n7914) );
  buffer buf_n7915( .i (n7914), .o (n7915) );
  buffer buf_n7916( .i (n7915), .o (n7916) );
  buffer buf_n7917( .i (n7916), .o (n7917) );
  buffer buf_n7918( .i (n7917), .o (n7918) );
  buffer buf_n7919( .i (n7918), .o (n7919) );
  buffer buf_n7920( .i (n7919), .o (n7920) );
  buffer buf_n7921( .i (n7920), .o (n7921) );
  buffer buf_n7922( .i (n7921), .o (n7922) );
  buffer buf_n7923( .i (n7922), .o (n7923) );
  buffer buf_n7924( .i (n7923), .o (n7924) );
  buffer buf_n7925( .i (n7924), .o (n7925) );
  buffer buf_n7926( .i (n7925), .o (n7926) );
  buffer buf_n7927( .i (n7926), .o (n7927) );
  buffer buf_n7928( .i (n7927), .o (n7928) );
  buffer buf_n7929( .i (n7928), .o (n7929) );
  buffer buf_n7930( .i (n7929), .o (n7930) );
  buffer buf_n7931( .i (n7930), .o (n7931) );
  buffer buf_n7932( .i (n7931), .o (n7932) );
  buffer buf_n7933( .i (n7932), .o (n7933) );
  buffer buf_n7934( .i (n7933), .o (n7934) );
  buffer buf_n7935( .i (n7934), .o (n7935) );
  buffer buf_n7936( .i (n7935), .o (n7936) );
  buffer buf_n7937( .i (n7936), .o (n7937) );
  buffer buf_n7938( .i (n7937), .o (n7938) );
  buffer buf_n7939( .i (n7938), .o (n7939) );
  buffer buf_n7940( .i (n7939), .o (n7940) );
  buffer buf_n7941( .i (n7940), .o (n7941) );
  buffer buf_n7942( .i (n7941), .o (n7942) );
  buffer buf_n7943( .i (n7942), .o (n7943) );
  buffer buf_n7944( .i (n7943), .o (n7944) );
  buffer buf_n7945( .i (n7944), .o (n7945) );
  buffer buf_n7946( .i (n7945), .o (n7946) );
  buffer buf_n7947( .i (n7946), .o (n7947) );
  buffer buf_n7948( .i (n7947), .o (n7948) );
  buffer buf_n7949( .i (n7948), .o (n7949) );
  buffer buf_n7950( .i (n7949), .o (n7950) );
  buffer buf_n7951( .i (n7950), .o (n7951) );
  buffer buf_n7952( .i (n7951), .o (n7952) );
  buffer buf_n7953( .i (n7952), .o (n7953) );
  buffer buf_n7954( .i (n7953), .o (n7954) );
  buffer buf_n7955( .i (n7954), .o (n7955) );
  buffer buf_n7956( .i (n7955), .o (n7956) );
  buffer buf_n7957( .i (n7956), .o (n7957) );
  buffer buf_n7958( .i (n7957), .o (n7958) );
  buffer buf_n7959( .i (n7958), .o (n7959) );
  buffer buf_n7960( .i (n7959), .o (n7960) );
  buffer buf_n7961( .i (n7960), .o (n7961) );
  buffer buf_n7962( .i (n7961), .o (n7962) );
  buffer buf_n7963( .i (n7962), .o (n7963) );
  buffer buf_n7964( .i (n7963), .o (n7964) );
  buffer buf_n7965( .i (n7964), .o (n7965) );
  buffer buf_n7966( .i (n7965), .o (n7966) );
  buffer buf_n7967( .i (n7966), .o (n7967) );
  buffer buf_n7968( .i (n7967), .o (n7968) );
  buffer buf_n7969( .i (n7968), .o (n7969) );
  buffer buf_n7970( .i (n7969), .o (n7970) );
  buffer buf_n7971( .i (n7970), .o (n7971) );
  buffer buf_n7972( .i (n7971), .o (n7972) );
  buffer buf_n7973( .i (n7972), .o (n7973) );
  buffer buf_n7974( .i (n7973), .o (n7974) );
  buffer buf_n7975( .i (n7974), .o (n7975) );
  buffer buf_n7976( .i (n7975), .o (n7976) );
  buffer buf_n7977( .i (n7976), .o (n7977) );
  buffer buf_n7978( .i (n7977), .o (n7978) );
  buffer buf_n7979( .i (n7978), .o (n7979) );
  buffer buf_n7980( .i (n7979), .o (n7980) );
  buffer buf_n7981( .i (n7980), .o (n7981) );
  buffer buf_n7982( .i (n7981), .o (n7982) );
  buffer buf_n7983( .i (n7982), .o (n7983) );
  buffer buf_n7984( .i (n7983), .o (n7984) );
  buffer buf_n7985( .i (n7984), .o (n7985) );
  buffer buf_n7986( .i (n7985), .o (n7986) );
  buffer buf_n7987( .i (n7986), .o (n7987) );
  buffer buf_n7988( .i (n7987), .o (n7988) );
  buffer buf_n7989( .i (n7988), .o (n7989) );
  buffer buf_n7990( .i (n7989), .o (n7990) );
  buffer buf_n7991( .i (n7990), .o (n7991) );
  buffer buf_n7992( .i (n7991), .o (n7992) );
  buffer buf_n7993( .i (n7992), .o (n7993) );
  buffer buf_n7994( .i (n7993), .o (n7994) );
  buffer buf_n7995( .i (n7994), .o (n7995) );
  buffer buf_n7996( .i (n7995), .o (n7996) );
  buffer buf_n7997( .i (n7996), .o (n7997) );
  buffer buf_n7998( .i (n7997), .o (n7998) );
  buffer buf_n7999( .i (n7998), .o (n7999) );
  buffer buf_n8000( .i (n7999), .o (n8000) );
  buffer buf_n8001( .i (n8000), .o (n8001) );
  buffer buf_n8002( .i (n8001), .o (n8002) );
  buffer buf_n8003( .i (n8002), .o (n8003) );
  buffer buf_n8004( .i (n8003), .o (n8004) );
  buffer buf_n8005( .i (n8004), .o (n8005) );
  buffer buf_n8006( .i (n8005), .o (n8006) );
  buffer buf_n8007( .i (n8006), .o (n8007) );
  buffer buf_n8008( .i (n8007), .o (n8008) );
  buffer buf_n8009( .i (n8008), .o (n8009) );
  buffer buf_n8010( .i (n8009), .o (n8010) );
  buffer buf_n8011( .i (n8010), .o (n8011) );
  buffer buf_n8012( .i (n8011), .o (n8012) );
  buffer buf_n8013( .i (n8012), .o (n8013) );
  buffer buf_n8014( .i (n8013), .o (n8014) );
  buffer buf_n8015( .i (n8014), .o (n8015) );
  buffer buf_n8016( .i (n8015), .o (n8016) );
  buffer buf_n8017( .i (n8016), .o (n8017) );
  buffer buf_n8018( .i (n8017), .o (n8018) );
  buffer buf_n7136( .i (n7135), .o (n7136) );
  buffer buf_n7137( .i (n7136), .o (n7137) );
  assign n8019 = ~n7142 & n7145 ;
  buffer buf_n8020( .i (n8019), .o (n8020) );
  assign n8021 = ~n7137 & n8020 ;
  assign n8022 = n7137 & ~n8020 ;
  assign n8023 = n8021 | n8022 ;
  buffer buf_n8024( .i (n8023), .o (n8024) );
  buffer buf_n8025( .i (n8024), .o (n8025) );
  buffer buf_n8026( .i (n8025), .o (n8026) );
  buffer buf_n8027( .i (n8026), .o (n8027) );
  buffer buf_n8028( .i (n8027), .o (n8028) );
  buffer buf_n8029( .i (n8028), .o (n8029) );
  buffer buf_n8030( .i (n8029), .o (n8030) );
  buffer buf_n8031( .i (n8030), .o (n8031) );
  buffer buf_n8032( .i (n8031), .o (n8032) );
  buffer buf_n8033( .i (n8032), .o (n8033) );
  buffer buf_n8034( .i (n8033), .o (n8034) );
  buffer buf_n8035( .i (n8034), .o (n8035) );
  buffer buf_n8036( .i (n8035), .o (n8036) );
  buffer buf_n8037( .i (n8036), .o (n8037) );
  buffer buf_n8038( .i (n8037), .o (n8038) );
  buffer buf_n8039( .i (n8038), .o (n8039) );
  buffer buf_n8040( .i (n8039), .o (n8040) );
  buffer buf_n8041( .i (n8040), .o (n8041) );
  buffer buf_n8042( .i (n8041), .o (n8042) );
  buffer buf_n8043( .i (n8042), .o (n8043) );
  buffer buf_n8044( .i (n8043), .o (n8044) );
  buffer buf_n8045( .i (n8044), .o (n8045) );
  buffer buf_n8046( .i (n8045), .o (n8046) );
  buffer buf_n8047( .i (n8046), .o (n8047) );
  buffer buf_n8048( .i (n8047), .o (n8048) );
  buffer buf_n8049( .i (n8048), .o (n8049) );
  buffer buf_n8050( .i (n8049), .o (n8050) );
  buffer buf_n8051( .i (n8050), .o (n8051) );
  buffer buf_n8052( .i (n8051), .o (n8052) );
  buffer buf_n8053( .i (n8052), .o (n8053) );
  buffer buf_n8054( .i (n8053), .o (n8054) );
  buffer buf_n8055( .i (n8054), .o (n8055) );
  buffer buf_n8056( .i (n8055), .o (n8056) );
  buffer buf_n8057( .i (n8056), .o (n8057) );
  buffer buf_n8058( .i (n8057), .o (n8058) );
  buffer buf_n8059( .i (n8058), .o (n8059) );
  buffer buf_n8060( .i (n8059), .o (n8060) );
  buffer buf_n8061( .i (n8060), .o (n8061) );
  buffer buf_n8062( .i (n8061), .o (n8062) );
  buffer buf_n8063( .i (n8062), .o (n8063) );
  buffer buf_n8064( .i (n8063), .o (n8064) );
  buffer buf_n8065( .i (n8064), .o (n8065) );
  buffer buf_n8066( .i (n8065), .o (n8066) );
  buffer buf_n8067( .i (n8066), .o (n8067) );
  buffer buf_n8068( .i (n8067), .o (n8068) );
  assign n8069 = n2996 & ~n5912 ;
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  assign n8070 = n1309 & n5912 ;
  assign n8071 = n8069 | n8070 ;
  buffer buf_n8072( .i (n8071), .o (n8072) );
  buffer buf_n8073( .i (n8072), .o (n8073) );
  buffer buf_n8074( .i (n6215), .o (n8074) );
  assign n8075 = ~n6542 & n8074 ;
  buffer buf_n8076( .i (n8075), .o (n8076) );
  assign n8077 = n8073 & n8076 ;
  buffer buf_n8078( .i (n8077), .o (n8078) );
  buffer buf_n4358( .i (n4357), .o (n4358) );
  buffer buf_n4359( .i (n4358), .o (n4359) );
  buffer buf_n4360( .i (n4359), .o (n4360) );
  buffer buf_n4361( .i (n4360), .o (n4361) );
  buffer buf_n4362( .i (n4361), .o (n4362) );
  buffer buf_n4363( .i (n4362), .o (n4363) );
  buffer buf_n4364( .i (n4363), .o (n4364) );
  buffer buf_n4365( .i (n4364), .o (n4365) );
  buffer buf_n4366( .i (n4365), .o (n4366) );
  buffer buf_n4367( .i (n4366), .o (n4367) );
  buffer buf_n4368( .i (n4367), .o (n4368) );
  buffer buf_n4369( .i (n4368), .o (n4369) );
  buffer buf_n4370( .i (n4369), .o (n4370) );
  buffer buf_n4371( .i (n4370), .o (n4371) );
  buffer buf_n4372( .i (n4371), .o (n4372) );
  buffer buf_n4373( .i (n4372), .o (n4373) );
  buffer buf_n4374( .i (n4373), .o (n4374) );
  buffer buf_n4375( .i (n4374), .o (n4375) );
  buffer buf_n4376( .i (n4375), .o (n4376) );
  buffer buf_n4377( .i (n4376), .o (n4377) );
  buffer buf_n4378( .i (n4377), .o (n4378) );
  buffer buf_n4379( .i (n4378), .o (n4379) );
  buffer buf_n4380( .i (n4379), .o (n4380) );
  buffer buf_n4381( .i (n4380), .o (n4381) );
  buffer buf_n4382( .i (n4381), .o (n4382) );
  buffer buf_n4383( .i (n4382), .o (n4383) );
  buffer buf_n4384( .i (n4383), .o (n4384) );
  buffer buf_n4385( .i (n4384), .o (n4385) );
  buffer buf_n4386( .i (n4385), .o (n4386) );
  buffer buf_n4387( .i (n4386), .o (n4387) );
  buffer buf_n4388( .i (n4387), .o (n4388) );
  buffer buf_n4389( .i (n4388), .o (n4389) );
  buffer buf_n4390( .i (n4389), .o (n4390) );
  buffer buf_n4391( .i (n4390), .o (n4391) );
  buffer buf_n4392( .i (n4391), .o (n4392) );
  assign n8079 = n3318 & ~n5913 ;
  buffer buf_n2954( .i (n2953), .o (n2954) );
  buffer buf_n2955( .i (n2954), .o (n2955) );
  buffer buf_n2956( .i (n2955), .o (n2956) );
  buffer buf_n2957( .i (n2956), .o (n2957) );
  assign n8080 = n2957 & n5913 ;
  assign n8081 = n8079 | n8080 ;
  buffer buf_n8082( .i (n8081), .o (n8082) );
  assign n8083 = ~n4392 & n8082 ;
  buffer buf_n8084( .i (n3560), .o (n8084) );
  assign n8085 = n8083 | n8084 ;
  assign n8086 = n8078 | n8085 ;
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n2571( .i (n2570), .o (n2571) );
  assign n8087 = n2310 & ~n5912 ;
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n8088( .i (n5911), .o (n8088) );
  assign n8089 = n487 & n8088 ;
  assign n8090 = n8087 | n8089 ;
  buffer buf_n8091( .i (n8090), .o (n8091) );
  assign n8092 = ~n2571 & n8091 ;
  buffer buf_n4048( .i (n4047), .o (n4048) );
  buffer buf_n4049( .i (n4048), .o (n4049) );
  buffer buf_n8093( .i (n6577), .o (n8093) );
  assign n8094 = n4049 & n8093 ;
  assign n8095 = n3602 & ~n8093 ;
  assign n8096 = n8094 | n8095 ;
  buffer buf_n8097( .i (n8096), .o (n8097) );
  buffer buf_n8098( .i (n8097), .o (n8098) );
  assign n8099 = n2571 & n8098 ;
  assign n8100 = n8092 | n8099 ;
  buffer buf_n8101( .i (n8100), .o (n8101) );
  assign n8102 = n45 & n8101 ;
  assign n8103 = n8086 | n8102 ;
  buffer buf_n8104( .i (n8103), .o (n8104) );
  assign n8105 = n44 & n6589 ;
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  assign n8106 = n756 & n8093 ;
  assign n8107 = n4089 & ~n8093 ;
  assign n8108 = n8106 | n8107 ;
  buffer buf_n8109( .i (n8108), .o (n8109) );
  assign n8110 = ~n8074 & n8109 ;
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n8111( .i (n6577), .o (n8111) );
  assign n8112 = n718 & n8111 ;
  assign n8113 = n1179 & ~n8111 ;
  assign n8114 = n8112 | n8113 ;
  buffer buf_n8115( .i (n8114), .o (n8115) );
  assign n8116 = n8074 & n8115 ;
  assign n8117 = n8110 | n8116 ;
  buffer buf_n8118( .i (n8117), .o (n8118) );
  buffer buf_n8119( .i (n6630), .o (n8119) );
  buffer buf_n8120( .i (n8119), .o (n8120) );
  assign n8121 = n8118 & ~n8120 ;
  assign n8122 = n8105 | n8121 ;
  buffer buf_n8123( .i (n8122), .o (n8123) );
  assign n8124 = n3564 & ~n8123 ;
  assign n8125 = n8104 & ~n8124 ;
  buffer buf_n8126( .i (n6557), .o (n8126) );
  assign n8127 = n8125 & ~n8126 ;
  assign n8128 = n6226 & n8126 ;
  assign n8129 = n8127 | n8128 ;
  assign n8130 = ~n6641 & n8129 ;
  buffer buf_n8131( .i (n8130), .o (n8131) );
  assign n8132 = n6146 & n8126 ;
  buffer buf_n6285( .i (n6284), .o (n6285) );
  assign n8133 = n6285 & ~n8126 ;
  assign n8134 = n8132 | n8133 ;
  buffer buf_n8135( .i (n8134), .o (n8135) );
  assign n8136 = n135 & n8135 ;
  assign n8137 = n8131 | n8136 ;
  buffer buf_n8138( .i (n8137), .o (n8138) );
  assign n8139 = n5928 & ~n8138 ;
  assign n8140 = n5885 & ~n8139 ;
  assign n8141 = n38 & n2955 ;
  buffer buf_n8142( .i (n8141), .o (n8142) );
  buffer buf_n8143( .i (n8142), .o (n8143) );
  assign n8144 = n6058 & ~n8143 ;
  assign n8145 = n6089 | n8144 ;
  buffer buf_n6059( .i (n6058), .o (n6059) );
  assign n8146 = n39 & n6067 ;
  assign n8147 = n2957 | n8146 ;
  assign n8148 = n6080 & n8142 ;
  assign n8149 = n8147 & ~n8148 ;
  assign n8150 = n6059 | n8149 ;
  assign n8151 = ~n8145 & n8150 ;
  buffer buf_n8152( .i (n8151), .o (n8152) );
  buffer buf_n8153( .i (n8152), .o (n8153) );
  assign n8154 = n5919 | n8153 ;
  buffer buf_n8155( .i (n8154), .o (n8155) );
  buffer buf_n8156( .i (n8155), .o (n8156) );
  buffer buf_n8157( .i (n8156), .o (n8157) );
  buffer buf_n8158( .i (n8157), .o (n8158) );
  buffer buf_n8159( .i (n8158), .o (n8159) );
  buffer buf_n8160( .i (n8159), .o (n8160) );
  buffer buf_n8161( .i (n8160), .o (n8161) );
  buffer buf_n8162( .i (n8161), .o (n8162) );
  assign n8163 = n5971 & ~n6557 ;
  assign n8164 = n6150 | n8163 ;
  buffer buf_n8165( .i (n8164), .o (n8165) );
  assign n8166 = ~n6641 & n8165 ;
  assign n8167 = n5950 | n8166 ;
  buffer buf_n8168( .i (n8167), .o (n8168) );
  assign n8170 = n6101 & n8168 ;
  assign n8171 = n8162 | n8170 ;
  buffer buf_n8172( .i (n8171), .o (n8172) );
  assign n8173 = n8140 & n8172 ;
  assign n8174 = ~n5632 & n7905 ;
  assign n8175 = n8173 | n8174 ;
  buffer buf_n8176( .i (n8175), .o (n8176) );
  buffer buf_n8177( .i (n8176), .o (n8177) );
  buffer buf_n8178( .i (n8177), .o (n8178) );
  buffer buf_n8179( .i (n8178), .o (n8179) );
  buffer buf_n8180( .i (n8179), .o (n8180) );
  buffer buf_n8181( .i (n8180), .o (n8181) );
  buffer buf_n8182( .i (n8181), .o (n8182) );
  buffer buf_n8183( .i (n8182), .o (n8183) );
  buffer buf_n8184( .i (n8183), .o (n8184) );
  buffer buf_n8185( .i (n8184), .o (n8185) );
  buffer buf_n8186( .i (n8185), .o (n8186) );
  buffer buf_n8187( .i (n8186), .o (n8187) );
  buffer buf_n8188( .i (n8187), .o (n8188) );
  buffer buf_n8189( .i (n8188), .o (n8189) );
  buffer buf_n8190( .i (n8189), .o (n8190) );
  buffer buf_n8191( .i (n8190), .o (n8191) );
  buffer buf_n8192( .i (n8191), .o (n8192) );
  buffer buf_n8193( .i (n8192), .o (n8193) );
  buffer buf_n8194( .i (n8193), .o (n8194) );
  buffer buf_n8195( .i (n8194), .o (n8195) );
  buffer buf_n8196( .i (n8195), .o (n8196) );
  buffer buf_n8197( .i (n8196), .o (n8197) );
  buffer buf_n8198( .i (n8197), .o (n8198) );
  buffer buf_n8199( .i (n8198), .o (n8199) );
  buffer buf_n8200( .i (n8199), .o (n8200) );
  buffer buf_n8201( .i (n8200), .o (n8201) );
  buffer buf_n8202( .i (n8201), .o (n8202) );
  buffer buf_n8203( .i (n8202), .o (n8203) );
  buffer buf_n8204( .i (n8203), .o (n8204) );
  buffer buf_n8205( .i (n8204), .o (n8205) );
  buffer buf_n8206( .i (n8205), .o (n8206) );
  buffer buf_n8207( .i (n8206), .o (n8207) );
  buffer buf_n8208( .i (n8207), .o (n8208) );
  buffer buf_n8209( .i (n8208), .o (n8209) );
  buffer buf_n8210( .i (n8209), .o (n8210) );
  buffer buf_n8211( .i (n8210), .o (n8211) );
  buffer buf_n8212( .i (n8211), .o (n8212) );
  buffer buf_n8213( .i (n8212), .o (n8213) );
  buffer buf_n8214( .i (n8213), .o (n8214) );
  buffer buf_n8215( .i (n8214), .o (n8215) );
  buffer buf_n8216( .i (n8215), .o (n8216) );
  buffer buf_n8217( .i (n8216), .o (n8217) );
  buffer buf_n8218( .i (n8217), .o (n8218) );
  buffer buf_n8219( .i (n8218), .o (n8219) );
  buffer buf_n8220( .i (n8219), .o (n8220) );
  buffer buf_n8221( .i (n8220), .o (n8221) );
  buffer buf_n8222( .i (n8221), .o (n8222) );
  buffer buf_n8223( .i (n8222), .o (n8223) );
  buffer buf_n8224( .i (n8223), .o (n8224) );
  buffer buf_n8225( .i (n8224), .o (n8225) );
  buffer buf_n8226( .i (n8225), .o (n8226) );
  buffer buf_n8227( .i (n8226), .o (n8227) );
  buffer buf_n8228( .i (n8227), .o (n8228) );
  buffer buf_n8229( .i (n8228), .o (n8229) );
  buffer buf_n8230( .i (n8229), .o (n8230) );
  buffer buf_n8231( .i (n8230), .o (n8231) );
  buffer buf_n8232( .i (n8231), .o (n8232) );
  buffer buf_n8233( .i (n8232), .o (n8233) );
  buffer buf_n8234( .i (n8233), .o (n8234) );
  buffer buf_n8235( .i (n8234), .o (n8235) );
  buffer buf_n8236( .i (n8235), .o (n8236) );
  buffer buf_n8237( .i (n8236), .o (n8237) );
  buffer buf_n8238( .i (n8237), .o (n8238) );
  buffer buf_n8239( .i (n8238), .o (n8239) );
  buffer buf_n8240( .i (n8239), .o (n8240) );
  buffer buf_n8241( .i (n8240), .o (n8241) );
  buffer buf_n8242( .i (n8241), .o (n8242) );
  buffer buf_n8243( .i (n8242), .o (n8243) );
  buffer buf_n8244( .i (n8243), .o (n8244) );
  buffer buf_n8245( .i (n8244), .o (n8245) );
  buffer buf_n8246( .i (n8245), .o (n8246) );
  buffer buf_n8247( .i (n8246), .o (n8247) );
  buffer buf_n8248( .i (n8247), .o (n8248) );
  buffer buf_n8249( .i (n8248), .o (n8249) );
  buffer buf_n8250( .i (n8249), .o (n8250) );
  buffer buf_n8251( .i (n8250), .o (n8251) );
  buffer buf_n8252( .i (n8251), .o (n8252) );
  buffer buf_n8253( .i (n8252), .o (n8253) );
  buffer buf_n8254( .i (n8253), .o (n8254) );
  buffer buf_n8255( .i (n8254), .o (n8255) );
  buffer buf_n8256( .i (n8255), .o (n8256) );
  buffer buf_n8257( .i (n8256), .o (n8257) );
  buffer buf_n8258( .i (n8257), .o (n8258) );
  buffer buf_n8259( .i (n8258), .o (n8259) );
  buffer buf_n8260( .i (n8259), .o (n8260) );
  buffer buf_n8261( .i (n8260), .o (n8261) );
  buffer buf_n8262( .i (n8261), .o (n8262) );
  buffer buf_n8263( .i (n8262), .o (n8263) );
  buffer buf_n8264( .i (n8263), .o (n8264) );
  buffer buf_n8265( .i (n8264), .o (n8265) );
  buffer buf_n8266( .i (n8265), .o (n8266) );
  buffer buf_n8267( .i (n8266), .o (n8267) );
  buffer buf_n8268( .i (n8267), .o (n8268) );
  buffer buf_n8269( .i (n8268), .o (n8269) );
  buffer buf_n8270( .i (n8269), .o (n8270) );
  buffer buf_n8271( .i (n8270), .o (n8271) );
  buffer buf_n8272( .i (n8271), .o (n8272) );
  buffer buf_n8273( .i (n8272), .o (n8273) );
  buffer buf_n8274( .i (n8273), .o (n8274) );
  buffer buf_n8275( .i (n8274), .o (n8275) );
  buffer buf_n8276( .i (n8275), .o (n8276) );
  buffer buf_n8277( .i (n8276), .o (n8277) );
  buffer buf_n8278( .i (n8277), .o (n8278) );
  buffer buf_n8279( .i (n8278), .o (n8279) );
  buffer buf_n8280( .i (n8279), .o (n8280) );
  buffer buf_n8281( .i (n8280), .o (n8281) );
  buffer buf_n8282( .i (n8281), .o (n8282) );
  buffer buf_n8283( .i (n8282), .o (n8283) );
  buffer buf_n8284( .i (n8283), .o (n8284) );
  buffer buf_n8285( .i (n8284), .o (n8285) );
  buffer buf_n8286( .i (n8285), .o (n8286) );
  buffer buf_n4990( .i (n4989), .o (n4990) );
  buffer buf_n4991( .i (n4990), .o (n4991) );
  assign n8287 = ~n4965 & n4994 ;
  buffer buf_n8288( .i (n8287), .o (n8288) );
  assign n8289 = n4991 & n8288 ;
  assign n8290 = n4991 | n8288 ;
  assign n8291 = ~n8289 & n8290 ;
  buffer buf_n8292( .i (n8291), .o (n8292) );
  buffer buf_n8293( .i (n8292), .o (n8293) );
  buffer buf_n8294( .i (n8293), .o (n8294) );
  buffer buf_n8295( .i (n8294), .o (n8295) );
  buffer buf_n8296( .i (n8295), .o (n8296) );
  buffer buf_n8297( .i (n8296), .o (n8297) );
  buffer buf_n8298( .i (n8297), .o (n8298) );
  buffer buf_n8299( .i (n8298), .o (n8299) );
  buffer buf_n8300( .i (n8299), .o (n8300) );
  buffer buf_n8301( .i (n8300), .o (n8301) );
  buffer buf_n8302( .i (n8301), .o (n8302) );
  buffer buf_n8303( .i (n8302), .o (n8303) );
  buffer buf_n8304( .i (n8303), .o (n8304) );
  buffer buf_n8305( .i (n8304), .o (n8305) );
  buffer buf_n8306( .i (n8305), .o (n8306) );
  buffer buf_n8307( .i (n8306), .o (n8307) );
  buffer buf_n8308( .i (n8307), .o (n8308) );
  buffer buf_n8309( .i (n8308), .o (n8309) );
  buffer buf_n8310( .i (n8309), .o (n8310) );
  buffer buf_n8311( .i (n8310), .o (n8311) );
  buffer buf_n8312( .i (n8311), .o (n8312) );
  buffer buf_n8313( .i (n8312), .o (n8313) );
  buffer buf_n8314( .i (n8313), .o (n8314) );
  buffer buf_n8315( .i (n8314), .o (n8315) );
  buffer buf_n8316( .i (n8315), .o (n8316) );
  buffer buf_n8317( .i (n8316), .o (n8317) );
  buffer buf_n8318( .i (n8317), .o (n8318) );
  buffer buf_n8319( .i (n8318), .o (n8319) );
  buffer buf_n8320( .i (n8319), .o (n8320) );
  buffer buf_n8321( .i (n8320), .o (n8321) );
  buffer buf_n8322( .i (n8321), .o (n8322) );
  buffer buf_n8323( .i (n8322), .o (n8323) );
  buffer buf_n8324( .i (n8323), .o (n8324) );
  buffer buf_n8325( .i (n8324), .o (n8325) );
  buffer buf_n8326( .i (n8325), .o (n8326) );
  buffer buf_n8327( .i (n8326), .o (n8327) );
  buffer buf_n8328( .i (n8327), .o (n8328) );
  buffer buf_n8329( .i (n8328), .o (n8329) );
  buffer buf_n8330( .i (n8329), .o (n8330) );
  buffer buf_n8331( .i (n8330), .o (n8331) );
  buffer buf_n8332( .i (n8331), .o (n8332) );
  buffer buf_n8333( .i (n8332), .o (n8333) );
  buffer buf_n8334( .i (n8333), .o (n8334) );
  buffer buf_n8335( .i (n8334), .o (n8335) );
  buffer buf_n8336( .i (n8335), .o (n8336) );
  buffer buf_n8337( .i (n8336), .o (n8337) );
  buffer buf_n8338( .i (n8337), .o (n8338) );
  buffer buf_n8339( .i (n8338), .o (n8339) );
  buffer buf_n8340( .i (n8339), .o (n8340) );
  buffer buf_n8341( .i (n8340), .o (n8341) );
  buffer buf_n8342( .i (n8341), .o (n8342) );
  buffer buf_n8343( .i (n8342), .o (n8343) );
  buffer buf_n8344( .i (n8343), .o (n8344) );
  buffer buf_n8345( .i (n8344), .o (n8345) );
  buffer buf_n8346( .i (n8345), .o (n8346) );
  buffer buf_n8347( .i (n8346), .o (n8347) );
  buffer buf_n8348( .i (n8347), .o (n8348) );
  buffer buf_n8349( .i (n8348), .o (n8349) );
  buffer buf_n8350( .i (n8349), .o (n8350) );
  buffer buf_n8351( .i (n8350), .o (n8351) );
  buffer buf_n8352( .i (n8351), .o (n8352) );
  buffer buf_n8353( .i (n8352), .o (n8353) );
  buffer buf_n8354( .i (n8353), .o (n8354) );
  buffer buf_n8355( .i (n8354), .o (n8355) );
  buffer buf_n8356( .i (n8355), .o (n8356) );
  buffer buf_n8357( .i (n8356), .o (n8357) );
  buffer buf_n8358( .i (n8357), .o (n8358) );
  buffer buf_n8359( .i (n8358), .o (n8359) );
  buffer buf_n8360( .i (n8359), .o (n8360) );
  buffer buf_n8361( .i (n8360), .o (n8361) );
  buffer buf_n8362( .i (n8361), .o (n8362) );
  buffer buf_n8363( .i (n8362), .o (n8363) );
  buffer buf_n8364( .i (n8363), .o (n8364) );
  buffer buf_n8365( .i (n8364), .o (n8365) );
  buffer buf_n8366( .i (n8365), .o (n8366) );
  buffer buf_n8367( .i (n8366), .o (n8367) );
  buffer buf_n8368( .i (n8367), .o (n8368) );
  buffer buf_n8369( .i (n8368), .o (n8369) );
  buffer buf_n8370( .i (n8369), .o (n8370) );
  buffer buf_n8371( .i (n8370), .o (n8371) );
  buffer buf_n8372( .i (n8371), .o (n8372) );
  buffer buf_n8373( .i (n8372), .o (n8373) );
  buffer buf_n8374( .i (n8373), .o (n8374) );
  buffer buf_n8375( .i (n8374), .o (n8375) );
  buffer buf_n8376( .i (n8375), .o (n8376) );
  buffer buf_n8377( .i (n8376), .o (n8377) );
  buffer buf_n8378( .i (n8377), .o (n8378) );
  buffer buf_n8379( .i (n8378), .o (n8379) );
  buffer buf_n8380( .i (n8379), .o (n8380) );
  buffer buf_n8381( .i (n8380), .o (n8381) );
  buffer buf_n8382( .i (n8381), .o (n8382) );
  buffer buf_n8383( .i (n8382), .o (n8383) );
  buffer buf_n8384( .i (n8383), .o (n8384) );
  buffer buf_n8385( .i (n8384), .o (n8385) );
  buffer buf_n8386( .i (n8385), .o (n8386) );
  buffer buf_n8387( .i (n8386), .o (n8387) );
  buffer buf_n8388( .i (n8387), .o (n8388) );
  buffer buf_n8389( .i (n8388), .o (n8389) );
  buffer buf_n8390( .i (n8389), .o (n8390) );
  buffer buf_n8391( .i (n8390), .o (n8391) );
  buffer buf_n8392( .i (n8391), .o (n8392) );
  buffer buf_n8393( .i (n8392), .o (n8393) );
  buffer buf_n8394( .i (n8393), .o (n8394) );
  buffer buf_n8395( .i (n8394), .o (n8395) );
  buffer buf_n8396( .i (n8395), .o (n8396) );
  buffer buf_n8397( .i (n8396), .o (n8397) );
  buffer buf_n8398( .i (n8397), .o (n8398) );
  buffer buf_n8399( .i (n8398), .o (n8399) );
  buffer buf_n8400( .i (n8399), .o (n8400) );
  buffer buf_n8401( .i (n8400), .o (n8401) );
  buffer buf_n8402( .i (n8401), .o (n8402) );
  buffer buf_n8403( .i (n8402), .o (n8403) );
  buffer buf_n8404( .i (n8403), .o (n8404) );
  buffer buf_n8405( .i (n8404), .o (n8405) );
  buffer buf_n8406( .i (n8405), .o (n8406) );
  buffer buf_n8407( .i (n8406), .o (n8407) );
  buffer buf_n8408( .i (n8407), .o (n8408) );
  buffer buf_n8409( .i (n8408), .o (n8409) );
  buffer buf_n8410( .i (n8409), .o (n8410) );
  buffer buf_n8411( .i (n8410), .o (n8411) );
  buffer buf_n8412( .i (n8411), .o (n8412) );
  buffer buf_n8413( .i (n8412), .o (n8413) );
  buffer buf_n4804( .i (n4803), .o (n4804) );
  buffer buf_n4805( .i (n4804), .o (n4805) );
  buffer buf_n4806( .i (n4805), .o (n4806) );
  buffer buf_n4807( .i (n4806), .o (n4807) );
  buffer buf_n4808( .i (n4807), .o (n4808) );
  buffer buf_n4809( .i (n4808), .o (n4809) );
  buffer buf_n4810( .i (n4809), .o (n4810) );
  buffer buf_n4811( .i (n4810), .o (n4811) );
  buffer buf_n4812( .i (n4811), .o (n4812) );
  buffer buf_n4813( .i (n4812), .o (n4813) );
  buffer buf_n4814( .i (n4813), .o (n4814) );
  buffer buf_n4815( .i (n4814), .o (n4815) );
  buffer buf_n4816( .i (n4815), .o (n4816) );
  buffer buf_n4817( .i (n4816), .o (n4817) );
  buffer buf_n4818( .i (n4817), .o (n4818) );
  buffer buf_n4819( .i (n4818), .o (n4819) );
  buffer buf_n4820( .i (n4819), .o (n4820) );
  buffer buf_n4821( .i (n4820), .o (n4821) );
  buffer buf_n4822( .i (n4821), .o (n4822) );
  buffer buf_n4823( .i (n4822), .o (n4823) );
  buffer buf_n4824( .i (n4823), .o (n4824) );
  buffer buf_n4825( .i (n4824), .o (n4825) );
  buffer buf_n4826( .i (n4825), .o (n4826) );
  buffer buf_n4827( .i (n4826), .o (n4827) );
  buffer buf_n4828( .i (n4827), .o (n4828) );
  buffer buf_n4829( .i (n4828), .o (n4829) );
  buffer buf_n4830( .i (n4829), .o (n4830) );
  buffer buf_n4831( .i (n4830), .o (n4831) );
  assign n8414 = n2187 | n2562 ;
  buffer buf_n8415( .i (n8414), .o (n8415) );
  assign n8416 = ~n4831 & n8415 ;
  buffer buf_n8417( .i (n8416), .o (n8417) );
  buffer buf_n8418( .i (n8417), .o (n8418) );
  buffer buf_n8419( .i (n8418), .o (n8419) );
  buffer buf_n8420( .i (n8419), .o (n8420) );
  buffer buf_n8421( .i (n8420), .o (n8421) );
  buffer buf_n8422( .i (n8421), .o (n8422) );
  buffer buf_n8423( .i (n8422), .o (n8423) );
  buffer buf_n8424( .i (n8423), .o (n8424) );
  buffer buf_n8425( .i (n8424), .o (n8425) );
  buffer buf_n8426( .i (n8425), .o (n8426) );
  buffer buf_n8427( .i (n8426), .o (n8427) );
  buffer buf_n8428( .i (n8427), .o (n8428) );
  buffer buf_n8429( .i (n8428), .o (n8429) );
  buffer buf_n8430( .i (n8429), .o (n8430) );
  buffer buf_n8431( .i (n8430), .o (n8431) );
  buffer buf_n8432( .i (n8431), .o (n8432) );
  buffer buf_n8433( .i (n8432), .o (n8433) );
  buffer buf_n8434( .i (n8433), .o (n8434) );
  buffer buf_n8435( .i (n8434), .o (n8435) );
  buffer buf_n8436( .i (n8435), .o (n8436) );
  buffer buf_n8437( .i (n8436), .o (n8437) );
  buffer buf_n8438( .i (n8437), .o (n8438) );
  buffer buf_n8439( .i (n8438), .o (n8439) );
  buffer buf_n8440( .i (n8439), .o (n8440) );
  buffer buf_n8441( .i (n8440), .o (n8441) );
  buffer buf_n8442( .i (n8441), .o (n8442) );
  buffer buf_n8443( .i (n8442), .o (n8443) );
  buffer buf_n8444( .i (n8443), .o (n8444) );
  buffer buf_n8445( .i (n8444), .o (n8445) );
  buffer buf_n8446( .i (n8445), .o (n8446) );
  buffer buf_n8447( .i (n8446), .o (n8447) );
  buffer buf_n8448( .i (n8447), .o (n8448) );
  buffer buf_n8449( .i (n8448), .o (n8449) );
  buffer buf_n8450( .i (n8449), .o (n8450) );
  buffer buf_n8451( .i (n8450), .o (n8451) );
  buffer buf_n8452( .i (n8451), .o (n8452) );
  buffer buf_n8453( .i (n8452), .o (n8453) );
  buffer buf_n8454( .i (n8453), .o (n8454) );
  buffer buf_n8455( .i (n8454), .o (n8455) );
  buffer buf_n8456( .i (n8455), .o (n8456) );
  buffer buf_n8457( .i (n8456), .o (n8457) );
  buffer buf_n8458( .i (n8457), .o (n8458) );
  buffer buf_n8459( .i (n8458), .o (n8459) );
  buffer buf_n8460( .i (n8459), .o (n8460) );
  buffer buf_n8461( .i (n8460), .o (n8461) );
  buffer buf_n8462( .i (n8461), .o (n8462) );
  buffer buf_n8463( .i (n8462), .o (n8463) );
  buffer buf_n8464( .i (n8463), .o (n8464) );
  buffer buf_n8465( .i (n8464), .o (n8465) );
  buffer buf_n8466( .i (n8465), .o (n8466) );
  buffer buf_n8467( .i (n8466), .o (n8467) );
  buffer buf_n8468( .i (n8467), .o (n8468) );
  buffer buf_n8469( .i (n8468), .o (n8469) );
  buffer buf_n8470( .i (n8469), .o (n8470) );
  buffer buf_n8471( .i (n8470), .o (n8471) );
  buffer buf_n8472( .i (n8471), .o (n8472) );
  buffer buf_n8473( .i (n8472), .o (n8473) );
  buffer buf_n8474( .i (n8473), .o (n8474) );
  buffer buf_n8475( .i (n8474), .o (n8475) );
  buffer buf_n8476( .i (n8475), .o (n8476) );
  buffer buf_n8477( .i (n8476), .o (n8477) );
  buffer buf_n8478( .i (n8477), .o (n8478) );
  buffer buf_n8479( .i (n8478), .o (n8479) );
  buffer buf_n8480( .i (n8479), .o (n8480) );
  buffer buf_n8481( .i (n8480), .o (n8481) );
  buffer buf_n8482( .i (n8481), .o (n8482) );
  buffer buf_n8483( .i (n8482), .o (n8483) );
  buffer buf_n8484( .i (n8483), .o (n8484) );
  buffer buf_n8485( .i (n8484), .o (n8485) );
  buffer buf_n8486( .i (n8485), .o (n8486) );
  buffer buf_n8487( .i (n8486), .o (n8487) );
  buffer buf_n8488( .i (n8487), .o (n8488) );
  buffer buf_n8489( .i (n8488), .o (n8489) );
  buffer buf_n8490( .i (n8489), .o (n8490) );
  buffer buf_n8491( .i (n8490), .o (n8491) );
  buffer buf_n8492( .i (n8491), .o (n8492) );
  buffer buf_n8493( .i (n8492), .o (n8493) );
  buffer buf_n8494( .i (n8493), .o (n8494) );
  buffer buf_n8495( .i (n8494), .o (n8495) );
  buffer buf_n8496( .i (n8495), .o (n8496) );
  buffer buf_n8497( .i (n8496), .o (n8497) );
  buffer buf_n8498( .i (n8497), .o (n8498) );
  buffer buf_n8499( .i (n8498), .o (n8499) );
  buffer buf_n8500( .i (n8499), .o (n8500) );
  buffer buf_n8501( .i (n8500), .o (n8501) );
  buffer buf_n8502( .i (n8501), .o (n8502) );
  buffer buf_n8503( .i (n8502), .o (n8503) );
  buffer buf_n8504( .i (n8503), .o (n8504) );
  buffer buf_n8505( .i (n8504), .o (n8505) );
  buffer buf_n8506( .i (n8505), .o (n8506) );
  buffer buf_n8507( .i (n8506), .o (n8507) );
  buffer buf_n8508( .i (n8507), .o (n8508) );
  buffer buf_n8509( .i (n8508), .o (n8509) );
  buffer buf_n8510( .i (n8509), .o (n8510) );
  buffer buf_n8511( .i (n8510), .o (n8511) );
  buffer buf_n8512( .i (n8511), .o (n8512) );
  buffer buf_n8513( .i (n8512), .o (n8513) );
  buffer buf_n8514( .i (n8513), .o (n8514) );
  buffer buf_n8515( .i (n8514), .o (n8515) );
  buffer buf_n8516( .i (n8515), .o (n8516) );
  buffer buf_n8517( .i (n8516), .o (n8517) );
  buffer buf_n8518( .i (n8517), .o (n8518) );
  buffer buf_n8519( .i (n8518), .o (n8519) );
  buffer buf_n8520( .i (n8519), .o (n8520) );
  buffer buf_n8521( .i (n8520), .o (n8521) );
  buffer buf_n8522( .i (n8521), .o (n8522) );
  buffer buf_n8523( .i (n8522), .o (n8523) );
  buffer buf_n8524( .i (n8523), .o (n8524) );
  buffer buf_n8525( .i (n8524), .o (n8525) );
  buffer buf_n8526( .i (n8525), .o (n8526) );
  buffer buf_n8527( .i (n8526), .o (n8527) );
  buffer buf_n8528( .i (n8527), .o (n8528) );
  buffer buf_n8529( .i (n8528), .o (n8529) );
  buffer buf_n8530( .i (n8529), .o (n8530) );
  buffer buf_n8531( .i (n8530), .o (n8531) );
  buffer buf_n8532( .i (n8531), .o (n8532) );
  buffer buf_n8533( .i (n8532), .o (n8533) );
  buffer buf_n8534( .i (n8533), .o (n8534) );
  buffer buf_n8535( .i (n8534), .o (n8535) );
  buffer buf_n8536( .i (n8535), .o (n8536) );
  buffer buf_n8537( .i (n8536), .o (n8537) );
  buffer buf_n8538( .i (n8537), .o (n8538) );
  buffer buf_n8539( .i (n8538), .o (n8539) );
  buffer buf_n8540( .i (n8539), .o (n8540) );
  buffer buf_n8541( .i (n8540), .o (n8541) );
  buffer buf_n8542( .i (n8541), .o (n8542) );
  buffer buf_n8543( .i (n8542), .o (n8543) );
  buffer buf_n8544( .i (n8543), .o (n8544) );
  buffer buf_n8545( .i (n8544), .o (n8545) );
  buffer buf_n8546( .i (n8545), .o (n8546) );
  buffer buf_n8547( .i (n8546), .o (n8547) );
  buffer buf_n8548( .i (n8547), .o (n8548) );
  buffer buf_n8549( .i (n8548), .o (n8549) );
  buffer buf_n8550( .i (n8549), .o (n8550) );
  buffer buf_n6426( .i (n6425), .o (n6426) );
  buffer buf_n6427( .i (n6426), .o (n6427) );
  buffer buf_n6428( .i (n6427), .o (n6428) );
  buffer buf_n6429( .i (n6428), .o (n6429) );
  buffer buf_n6430( .i (n6429), .o (n6430) );
  buffer buf_n6431( .i (n6430), .o (n6431) );
  buffer buf_n6432( .i (n6431), .o (n6432) );
  buffer buf_n6433( .i (n6432), .o (n6433) );
  buffer buf_n6434( .i (n6433), .o (n6434) );
  buffer buf_n6435( .i (n6434), .o (n6435) );
  buffer buf_n6436( .i (n6435), .o (n6436) );
  buffer buf_n6437( .i (n6436), .o (n6437) );
  buffer buf_n6438( .i (n6437), .o (n6438) );
  buffer buf_n6439( .i (n6438), .o (n6439) );
  buffer buf_n6440( .i (n6439), .o (n6440) );
  buffer buf_n6441( .i (n6440), .o (n6441) );
  buffer buf_n6442( .i (n6441), .o (n6442) );
  buffer buf_n6443( .i (n6442), .o (n6443) );
  buffer buf_n6444( .i (n6443), .o (n6444) );
  buffer buf_n6445( .i (n6444), .o (n6445) );
  buffer buf_n6446( .i (n6445), .o (n6446) );
  buffer buf_n6447( .i (n6446), .o (n6447) );
  buffer buf_n6448( .i (n6447), .o (n6448) );
  buffer buf_n6449( .i (n6448), .o (n6449) );
  buffer buf_n6450( .i (n6449), .o (n6450) );
  buffer buf_n6451( .i (n6450), .o (n6451) );
  buffer buf_n6452( .i (n6451), .o (n6452) );
  buffer buf_n6453( .i (n6452), .o (n6453) );
  buffer buf_n6454( .i (n6453), .o (n6454) );
  buffer buf_n6455( .i (n6454), .o (n6455) );
  buffer buf_n6456( .i (n6455), .o (n6456) );
  buffer buf_n6457( .i (n6456), .o (n6457) );
  buffer buf_n6458( .i (n6457), .o (n6458) );
  buffer buf_n6459( .i (n6458), .o (n6459) );
  buffer buf_n6460( .i (n6459), .o (n6460) );
  buffer buf_n6461( .i (n6460), .o (n6461) );
  buffer buf_n6462( .i (n6461), .o (n6462) );
  buffer buf_n6463( .i (n6462), .o (n6463) );
  buffer buf_n6464( .i (n6463), .o (n6464) );
  buffer buf_n6465( .i (n6464), .o (n6465) );
  buffer buf_n6466( .i (n6465), .o (n6466) );
  buffer buf_n6467( .i (n6466), .o (n6467) );
  buffer buf_n6468( .i (n6467), .o (n6468) );
  buffer buf_n6469( .i (n6468), .o (n6469) );
  buffer buf_n6470( .i (n6469), .o (n6470) );
  buffer buf_n6471( .i (n6470), .o (n6471) );
  buffer buf_n6472( .i (n6471), .o (n6472) );
  buffer buf_n6473( .i (n6472), .o (n6473) );
  buffer buf_n6474( .i (n6473), .o (n6474) );
  buffer buf_n6475( .i (n6474), .o (n6475) );
  buffer buf_n6476( .i (n6475), .o (n6476) );
  buffer buf_n6477( .i (n6476), .o (n6477) );
  buffer buf_n6478( .i (n6477), .o (n6478) );
  buffer buf_n6479( .i (n6478), .o (n6479) );
  buffer buf_n6480( .i (n6479), .o (n6480) );
  buffer buf_n6481( .i (n6480), .o (n6481) );
  buffer buf_n6482( .i (n6481), .o (n6482) );
  buffer buf_n6483( .i (n6482), .o (n6483) );
  buffer buf_n6484( .i (n6483), .o (n6484) );
  buffer buf_n6485( .i (n6484), .o (n6485) );
  buffer buf_n6486( .i (n6485), .o (n6486) );
  buffer buf_n6487( .i (n6486), .o (n6487) );
  buffer buf_n6488( .i (n6487), .o (n6488) );
  buffer buf_n6489( .i (n6488), .o (n6489) );
  buffer buf_n6490( .i (n6489), .o (n6490) );
  buffer buf_n6491( .i (n6490), .o (n6491) );
  buffer buf_n6492( .i (n6491), .o (n6492) );
  buffer buf_n6493( .i (n6492), .o (n6493) );
  buffer buf_n6494( .i (n6493), .o (n6494) );
  buffer buf_n6495( .i (n6494), .o (n6495) );
  buffer buf_n6496( .i (n6495), .o (n6496) );
  buffer buf_n6497( .i (n6496), .o (n6497) );
  buffer buf_n6498( .i (n6497), .o (n6498) );
  buffer buf_n6499( .i (n6498), .o (n6499) );
  buffer buf_n6500( .i (n6499), .o (n6500) );
  buffer buf_n6501( .i (n6500), .o (n6501) );
  buffer buf_n6502( .i (n6501), .o (n6502) );
  buffer buf_n6503( .i (n6502), .o (n6503) );
  buffer buf_n6504( .i (n6503), .o (n6504) );
  buffer buf_n6505( .i (n6504), .o (n6505) );
  buffer buf_n6506( .i (n6505), .o (n6506) );
  buffer buf_n6507( .i (n6506), .o (n6507) );
  buffer buf_n6508( .i (n6507), .o (n6508) );
  buffer buf_n6509( .i (n6508), .o (n6509) );
  buffer buf_n6510( .i (n6509), .o (n6510) );
  buffer buf_n6511( .i (n6510), .o (n6511) );
  buffer buf_n6512( .i (n6511), .o (n6512) );
  buffer buf_n6513( .i (n6512), .o (n6513) );
  buffer buf_n6514( .i (n6513), .o (n6514) );
  buffer buf_n6515( .i (n6514), .o (n6515) );
  buffer buf_n6516( .i (n6515), .o (n6516) );
  buffer buf_n6517( .i (n6516), .o (n6517) );
  buffer buf_n6518( .i (n6517), .o (n6518) );
  buffer buf_n6519( .i (n6518), .o (n6519) );
  buffer buf_n6520( .i (n6519), .o (n6520) );
  buffer buf_n6521( .i (n6520), .o (n6521) );
  buffer buf_n6522( .i (n6521), .o (n6522) );
  buffer buf_n6523( .i (n6522), .o (n6523) );
  buffer buf_n6524( .i (n6523), .o (n6524) );
  buffer buf_n6525( .i (n6524), .o (n6525) );
  buffer buf_n6526( .i (n6525), .o (n6526) );
  buffer buf_n6527( .i (n6526), .o (n6527) );
  buffer buf_n6528( .i (n6527), .o (n6528) );
  buffer buf_n6529( .i (n6528), .o (n6529) );
  buffer buf_n6530( .i (n6529), .o (n6530) );
  buffer buf_n6531( .i (n6530), .o (n6531) );
  buffer buf_n6532( .i (n6531), .o (n6532) );
  buffer buf_n6533( .i (n6532), .o (n6533) );
  buffer buf_n6534( .i (n6533), .o (n6534) );
  buffer buf_n6535( .i (n6534), .o (n6535) );
  buffer buf_n6536( .i (n6535), .o (n6536) );
  buffer buf_n6537( .i (n6536), .o (n6537) );
  buffer buf_n6538( .i (n6537), .o (n6538) );
  buffer buf_n6539( .i (n6538), .o (n6539) );
  buffer buf_n5246( .i (n5245), .o (n5246) );
  buffer buf_n5247( .i (n5246), .o (n5247) );
  assign n8551 = ~n5198 & n5250 ;
  buffer buf_n8552( .i (n8551), .o (n8552) );
  assign n8553 = ~n5247 & n8552 ;
  assign n8554 = n5247 & ~n8552 ;
  assign n8555 = n8553 | n8554 ;
  buffer buf_n8556( .i (n8555), .o (n8556) );
  assign n8641 = ~n5661 & n8556 ;
  buffer buf_n8642( .i (n1863), .o (n8642) );
  assign n8643 = n6637 & n8642 ;
  assign n8644 = n6247 & ~n6269 ;
  buffer buf_n8645( .i (n6135), .o (n8645) );
  assign n8646 = n6268 & n8645 ;
  assign n8647 = n8644 | n8646 ;
  buffer buf_n8648( .i (n8647), .o (n8648) );
  assign n8649 = ~n6630 & n8648 ;
  buffer buf_n8650( .i (n40), .o (n8650) );
  buffer buf_n8651( .i (n8650), .o (n8651) );
  assign n8652 = n5986 & n8651 ;
  assign n8653 = n8649 | n8652 ;
  buffer buf_n8654( .i (n8653), .o (n8654) );
  assign n8655 = n6552 & n8654 ;
  assign n8656 = n6231 & ~n8645 ;
  assign n8657 = n6254 & n8645 ;
  assign n8658 = n8656 | n8657 ;
  buffer buf_n8659( .i (n8658), .o (n8659) );
  assign n8660 = n8651 & n8659 ;
  assign n8661 = n6194 & ~n8645 ;
  buffer buf_n8662( .i (n2566), .o (n8662) );
  buffer buf_n8663( .i (n8662), .o (n8663) );
  assign n8664 = n6237 & n8663 ;
  assign n8665 = n8661 | n8664 ;
  buffer buf_n8666( .i (n8665), .o (n8666) );
  assign n8668 = ~n8651 & n8666 ;
  assign n8669 = n8660 | n8668 ;
  buffer buf_n8670( .i (n8669), .o (n8670) );
  buffer buf_n8672( .i (n8084), .o (n8672) );
  assign n8673 = n8670 & ~n8672 ;
  assign n8674 = n8655 | n8673 ;
  buffer buf_n8675( .i (n8674), .o (n8675) );
  assign n8677 = ~n8642 & n8675 ;
  assign n8678 = n8643 | n8677 ;
  buffer buf_n8679( .i (n8678), .o (n8679) );
  assign n8680 = ~n6641 & n8679 ;
  buffer buf_n8681( .i (n5949), .o (n8681) );
  assign n8682 = n8680 | n8681 ;
  buffer buf_n8683( .i (n8682), .o (n8683) );
  assign n8684 = n6101 & n8683 ;
  buffer buf_n2234( .i (n2233), .o (n2234) );
  assign n8685 = n2234 & n6078 ;
  assign n8686 = n1346 & ~n6053 ;
  buffer buf_n8687( .i (n8686), .o (n8687) );
  buffer buf_n8688( .i (n8687), .o (n8688) );
  assign n8689 = ~n8685 & n8688 ;
  assign n8690 = n1348 | n6066 ;
  assign n8691 = n2234 & ~n8687 ;
  assign n8692 = n8690 & n8691 ;
  assign n8693 = n8689 | n8692 ;
  buffer buf_n8694( .i (n8693), .o (n8694) );
  buffer buf_n8695( .i (n8694), .o (n8695) );
  assign n8696 = ~n6090 & n8695 ;
  buffer buf_n8697( .i (n8696), .o (n8697) );
  buffer buf_n8698( .i (n8697), .o (n8698) );
  buffer buf_n8699( .i (n5918), .o (n8699) );
  assign n8700 = n8698 | n8699 ;
  buffer buf_n8701( .i (n8700), .o (n8701) );
  buffer buf_n8702( .i (n8701), .o (n8702) );
  buffer buf_n8703( .i (n8702), .o (n8703) );
  buffer buf_n8704( .i (n8703), .o (n8704) );
  buffer buf_n8705( .i (n8704), .o (n8705) );
  buffer buf_n8706( .i (n8705), .o (n8706) );
  buffer buf_n8707( .i (n8706), .o (n8707) );
  buffer buf_n8708( .i (n8707), .o (n8708) );
  assign n8709 = n8684 | n8708 ;
  buffer buf_n6556( .i (n6555), .o (n6556) );
  buffer buf_n8710( .i (n8642), .o (n8710) );
  assign n8711 = ~n6556 & n8710 ;
  buffer buf_n8712( .i (n8711), .o (n8712) );
  assign n8713 = n6617 | n8710 ;
  assign n8714 = ~n133 & n8713 ;
  assign n8715 = ~n8712 & n8714 ;
  buffer buf_n5936( .i (n5935), .o (n5936) );
  buffer buf_n4430( .i (n4429), .o (n4430) );
  buffer buf_n4431( .i (n4430), .o (n4431) );
  buffer buf_n4432( .i (n4431), .o (n4432) );
  buffer buf_n4433( .i (n4432), .o (n4433) );
  buffer buf_n4434( .i (n4433), .o (n4434) );
  buffer buf_n4435( .i (n4434), .o (n4435) );
  buffer buf_n4436( .i (n4435), .o (n4436) );
  buffer buf_n4437( .i (n4436), .o (n4437) );
  buffer buf_n4438( .i (n4437), .o (n4438) );
  buffer buf_n4439( .i (n4438), .o (n4439) );
  buffer buf_n4440( .i (n4439), .o (n4440) );
  buffer buf_n4441( .i (n4440), .o (n4441) );
  buffer buf_n4442( .i (n4441), .o (n4442) );
  buffer buf_n4443( .i (n4442), .o (n4443) );
  buffer buf_n4444( .i (n4443), .o (n4444) );
  buffer buf_n4445( .i (n4444), .o (n4445) );
  buffer buf_n4446( .i (n4445), .o (n4446) );
  buffer buf_n4447( .i (n4446), .o (n4447) );
  assign n8716 = ~n3903 & n4447 ;
  assign n8717 = n121 & ~n8716 ;
  buffer buf_n8718( .i (n8717), .o (n8718) );
  buffer buf_n8719( .i (n8718), .o (n8719) );
  buffer buf_n8720( .i (n8719), .o (n8720) );
  buffer buf_n8721( .i (n8720), .o (n8721) );
  assign n8722 = n5936 & n8721 ;
  buffer buf_n8723( .i (n8722), .o (n8723) );
  buffer buf_n8724( .i (n8723), .o (n8724) );
  buffer buf_n8725( .i (n8724), .o (n8725) );
  buffer buf_n8726( .i (n8725), .o (n8726) );
  buffer buf_n8727( .i (n8726), .o (n8727) );
  buffer buf_n8728( .i (n8727), .o (n8728) );
  buffer buf_n8729( .i (n8728), .o (n8729) );
  buffer buf_n8730( .i (n8729), .o (n8730) );
  assign n8731 = n8715 | n8730 ;
  buffer buf_n8732( .i (n8731), .o (n8732) );
  assign n8733 = n5927 & ~n8732 ;
  assign n8734 = n5884 & ~n8733 ;
  assign n8735 = n8709 & n8734 ;
  buffer buf_n8736( .i (n8735), .o (n8736) );
  buffer buf_n8737( .i (n8736), .o (n8737) );
  buffer buf_n8738( .i (n8737), .o (n8738) );
  buffer buf_n8739( .i (n8738), .o (n8739) );
  buffer buf_n8740( .i (n8739), .o (n8740) );
  buffer buf_n8741( .i (n8740), .o (n8741) );
  buffer buf_n8742( .i (n8741), .o (n8742) );
  buffer buf_n8743( .i (n8742), .o (n8743) );
  buffer buf_n8744( .i (n8743), .o (n8744) );
  buffer buf_n8745( .i (n8744), .o (n8745) );
  buffer buf_n8746( .i (n8745), .o (n8746) );
  buffer buf_n8747( .i (n8746), .o (n8747) );
  buffer buf_n8748( .i (n8747), .o (n8748) );
  buffer buf_n8749( .i (n8748), .o (n8749) );
  buffer buf_n8750( .i (n8749), .o (n8750) );
  buffer buf_n8751( .i (n8750), .o (n8751) );
  buffer buf_n8752( .i (n8751), .o (n8752) );
  buffer buf_n8753( .i (n8752), .o (n8753) );
  buffer buf_n8754( .i (n8753), .o (n8754) );
  buffer buf_n8755( .i (n8754), .o (n8755) );
  buffer buf_n8756( .i (n8755), .o (n8756) );
  buffer buf_n8757( .i (n8756), .o (n8757) );
  buffer buf_n8758( .i (n8757), .o (n8758) );
  buffer buf_n8759( .i (n8758), .o (n8759) );
  buffer buf_n8760( .i (n8759), .o (n8760) );
  buffer buf_n8761( .i (n8760), .o (n8761) );
  buffer buf_n8762( .i (n8761), .o (n8762) );
  buffer buf_n8763( .i (n8762), .o (n8763) );
  buffer buf_n8764( .i (n8763), .o (n8764) );
  buffer buf_n8765( .i (n8764), .o (n8765) );
  assign n8766 = n8641 | n8765 ;
  buffer buf_n8767( .i (n8766), .o (n8767) );
  buffer buf_n8768( .i (n8767), .o (n8768) );
  buffer buf_n8769( .i (n8768), .o (n8769) );
  buffer buf_n8770( .i (n8769), .o (n8770) );
  buffer buf_n8771( .i (n8770), .o (n8771) );
  buffer buf_n8772( .i (n8771), .o (n8772) );
  buffer buf_n8773( .i (n8772), .o (n8773) );
  buffer buf_n8774( .i (n8773), .o (n8774) );
  buffer buf_n8775( .i (n8774), .o (n8775) );
  buffer buf_n8776( .i (n8775), .o (n8776) );
  buffer buf_n8777( .i (n8776), .o (n8777) );
  buffer buf_n8778( .i (n8777), .o (n8778) );
  buffer buf_n8779( .i (n8778), .o (n8779) );
  buffer buf_n8780( .i (n8779), .o (n8780) );
  buffer buf_n8781( .i (n8780), .o (n8781) );
  buffer buf_n8782( .i (n8781), .o (n8782) );
  buffer buf_n8783( .i (n8782), .o (n8783) );
  buffer buf_n8784( .i (n8783), .o (n8784) );
  buffer buf_n8785( .i (n8784), .o (n8785) );
  buffer buf_n8786( .i (n8785), .o (n8786) );
  buffer buf_n8787( .i (n8786), .o (n8787) );
  buffer buf_n8788( .i (n8787), .o (n8788) );
  buffer buf_n8789( .i (n8788), .o (n8789) );
  buffer buf_n8790( .i (n8789), .o (n8790) );
  buffer buf_n8791( .i (n8790), .o (n8791) );
  buffer buf_n8792( .i (n8791), .o (n8792) );
  buffer buf_n8793( .i (n8792), .o (n8793) );
  buffer buf_n8794( .i (n8793), .o (n8794) );
  buffer buf_n8795( .i (n8794), .o (n8795) );
  buffer buf_n8796( .i (n8795), .o (n8796) );
  buffer buf_n8797( .i (n8796), .o (n8797) );
  buffer buf_n8798( .i (n8797), .o (n8798) );
  buffer buf_n8799( .i (n8798), .o (n8799) );
  buffer buf_n8800( .i (n8799), .o (n8800) );
  buffer buf_n8801( .i (n8800), .o (n8801) );
  buffer buf_n8802( .i (n8801), .o (n8802) );
  buffer buf_n8803( .i (n8802), .o (n8803) );
  buffer buf_n8804( .i (n8803), .o (n8804) );
  buffer buf_n8805( .i (n8804), .o (n8805) );
  buffer buf_n8806( .i (n8805), .o (n8806) );
  buffer buf_n8807( .i (n8806), .o (n8807) );
  buffer buf_n8808( .i (n8807), .o (n8808) );
  buffer buf_n8809( .i (n8808), .o (n8809) );
  buffer buf_n8810( .i (n8809), .o (n8810) );
  buffer buf_n8811( .i (n8810), .o (n8811) );
  buffer buf_n8812( .i (n8811), .o (n8812) );
  buffer buf_n8813( .i (n8812), .o (n8813) );
  buffer buf_n8814( .i (n8813), .o (n8814) );
  buffer buf_n8815( .i (n8814), .o (n8815) );
  buffer buf_n8816( .i (n8815), .o (n8816) );
  buffer buf_n8817( .i (n8816), .o (n8817) );
  buffer buf_n8818( .i (n8817), .o (n8818) );
  buffer buf_n8819( .i (n8818), .o (n8819) );
  buffer buf_n8820( .i (n8819), .o (n8820) );
  buffer buf_n8821( .i (n8820), .o (n8821) );
  buffer buf_n8822( .i (n8821), .o (n8822) );
  buffer buf_n8823( .i (n8822), .o (n8823) );
  buffer buf_n8824( .i (n8823), .o (n8824) );
  buffer buf_n8825( .i (n8824), .o (n8825) );
  buffer buf_n8826( .i (n8825), .o (n8826) );
  buffer buf_n8827( .i (n8826), .o (n8827) );
  buffer buf_n8828( .i (n8827), .o (n8828) );
  buffer buf_n8829( .i (n8828), .o (n8829) );
  buffer buf_n8830( .i (n8829), .o (n8830) );
  buffer buf_n8831( .i (n8830), .o (n8831) );
  buffer buf_n8832( .i (n8831), .o (n8832) );
  buffer buf_n8833( .i (n8832), .o (n8833) );
  buffer buf_n8834( .i (n8833), .o (n8834) );
  buffer buf_n8835( .i (n8834), .o (n8835) );
  buffer buf_n8836( .i (n8835), .o (n8836) );
  buffer buf_n8837( .i (n8836), .o (n8837) );
  buffer buf_n8838( .i (n8837), .o (n8838) );
  buffer buf_n8839( .i (n8838), .o (n8839) );
  buffer buf_n8840( .i (n8839), .o (n8840) );
  buffer buf_n8841( .i (n8840), .o (n8841) );
  buffer buf_n8842( .i (n8841), .o (n8842) );
  buffer buf_n8843( .i (n8842), .o (n8843) );
  buffer buf_n8844( .i (n8843), .o (n8844) );
  buffer buf_n8845( .i (n8844), .o (n8845) );
  buffer buf_n8846( .i (n8845), .o (n8846) );
  buffer buf_n8847( .i (n8846), .o (n8847) );
  buffer buf_n8848( .i (n8847), .o (n8848) );
  buffer buf_n5697( .i (n5696), .o (n5697) );
  buffer buf_n5698( .i (n5697), .o (n5698) );
  buffer buf_n5699( .i (n5698), .o (n5699) );
  buffer buf_n5700( .i (n5699), .o (n5700) );
  buffer buf_n5701( .i (n5700), .o (n5701) );
  buffer buf_n5702( .i (n5701), .o (n5702) );
  buffer buf_n5703( .i (n5702), .o (n5703) );
  buffer buf_n5704( .i (n5703), .o (n5704) );
  buffer buf_n5705( .i (n5704), .o (n5705) );
  buffer buf_n5706( .i (n5705), .o (n5706) );
  buffer buf_n5707( .i (n5706), .o (n5707) );
  buffer buf_n5708( .i (n5707), .o (n5708) );
  buffer buf_n5709( .i (n5708), .o (n5709) );
  buffer buf_n5710( .i (n5709), .o (n5710) );
  buffer buf_n5711( .i (n5710), .o (n5711) );
  buffer buf_n5712( .i (n5711), .o (n5712) );
  buffer buf_n5713( .i (n5712), .o (n5713) );
  buffer buf_n5714( .i (n5713), .o (n5714) );
  buffer buf_n5715( .i (n5714), .o (n5715) );
  buffer buf_n5716( .i (n5715), .o (n5716) );
  buffer buf_n5717( .i (n5716), .o (n5717) );
  buffer buf_n5718( .i (n5717), .o (n5718) );
  buffer buf_n5719( .i (n5718), .o (n5719) );
  buffer buf_n5720( .i (n5719), .o (n5720) );
  buffer buf_n5721( .i (n5720), .o (n5721) );
  buffer buf_n5722( .i (n5721), .o (n5722) );
  buffer buf_n5723( .i (n5722), .o (n5723) );
  buffer buf_n5724( .i (n5723), .o (n5724) );
  buffer buf_n5725( .i (n5724), .o (n5725) );
  buffer buf_n5726( .i (n5725), .o (n5726) );
  buffer buf_n5727( .i (n5726), .o (n5727) );
  buffer buf_n5728( .i (n5727), .o (n5728) );
  buffer buf_n5729( .i (n5728), .o (n5729) );
  buffer buf_n5730( .i (n5729), .o (n5730) );
  buffer buf_n5731( .i (n5730), .o (n5731) );
  buffer buf_n5732( .i (n5731), .o (n5732) );
  buffer buf_n5733( .i (n5732), .o (n5733) );
  buffer buf_n5734( .i (n5733), .o (n5734) );
  buffer buf_n5735( .i (n5734), .o (n5735) );
  buffer buf_n5736( .i (n5735), .o (n5736) );
  buffer buf_n5737( .i (n5736), .o (n5737) );
  buffer buf_n5738( .i (n5737), .o (n5738) );
  buffer buf_n5739( .i (n5738), .o (n5739) );
  buffer buf_n5740( .i (n5739), .o (n5740) );
  assign n8849 = ~n6896 & n7731 ;
  buffer buf_n8850( .i (n8849), .o (n8850) );
  assign n8851 = n7644 & ~n8850 ;
  assign n8852 = ~n7644 & n8850 ;
  assign n8853 = n8851 | n8852 ;
  buffer buf_n8854( .i (n8853), .o (n8854) );
  assign n8860 = ~n5740 & n8854 ;
  buffer buf_n8861( .i (n133), .o (n8861) );
  assign n8862 = n8679 & n8861 ;
  assign n8863 = n6164 & n6215 ;
  assign n8864 = ~n6215 & n6580 ;
  assign n8865 = n8863 | n8864 ;
  buffer buf_n8866( .i (n8865), .o (n8866) );
  assign n8868 = ~n8119 & n8866 ;
  buffer buf_n8869( .i (n8663), .o (n8869) );
  assign n8870 = n6158 & ~n8869 ;
  assign n8871 = n6180 & n8869 ;
  assign n8872 = n8870 | n8871 ;
  buffer buf_n8873( .i (n8872), .o (n8873) );
  assign n8874 = n8119 & n8873 ;
  assign n8875 = n8868 | n8874 ;
  buffer buf_n8876( .i (n8875), .o (n8876) );
  assign n8878 = ~n6223 & n8876 ;
  assign n8879 = n6209 & n8869 ;
  assign n8880 = n6174 & ~n8869 ;
  assign n8881 = n8879 | n8880 ;
  buffer buf_n8882( .i (n8881), .o (n8882) );
  assign n8883 = ~n8119 & n8882 ;
  buffer buf_n8884( .i (n8663), .o (n8884) );
  assign n8885 = n6214 & ~n8884 ;
  assign n8886 = n6200 & n8884 ;
  assign n8887 = n8885 | n8886 ;
  buffer buf_n8888( .i (n8887), .o (n8888) );
  buffer buf_n8889( .i (n8651), .o (n8889) );
  assign n8890 = n8888 & n8889 ;
  assign n8891 = n8883 | n8890 ;
  buffer buf_n8892( .i (n8891), .o (n8892) );
  buffer buf_n8893( .i (n8672), .o (n8893) );
  assign n8894 = n8892 & n8893 ;
  assign n8895 = n8878 | n8894 ;
  buffer buf_n8896( .i (n8895), .o (n8896) );
  assign n8897 = n8710 & n8896 ;
  buffer buf_n2191( .i (n2190), .o (n2191) );
  buffer buf_n2192( .i (n2191), .o (n2192) );
  buffer buf_n2193( .i (n2192), .o (n2193) );
  buffer buf_n2194( .i (n2193), .o (n2194) );
  buffer buf_n2195( .i (n2194), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  assign n8898 = ~n2196 & n5915 ;
  assign n8899 = n2496 | n5914 ;
  assign n8900 = ~n4391 & n8899 ;
  assign n8901 = ~n8898 & n8900 ;
  assign n8902 = n8084 | n8901 ;
  buffer buf_n8903( .i (n8902), .o (n8903) );
  buffer buf_n8904( .i (n8903), .o (n8904) );
  assign n8905 = n8076 & n8082 ;
  buffer buf_n8906( .i (n8905), .o (n8906) );
  buffer buf_n8907( .i (n8906), .o (n8907) );
  assign n8908 = ~n2571 & n8072 ;
  assign n8909 = n2571 & n8091 ;
  assign n8910 = n8908 | n8909 ;
  buffer buf_n8911( .i (n8910), .o (n8911) );
  assign n8912 = n45 & n8911 ;
  assign n8913 = n8907 | n8912 ;
  assign n8914 = n8904 | n8913 ;
  assign n8915 = n6586 & n8074 ;
  buffer buf_n8916( .i (n8884), .o (n8916) );
  assign n8917 = n8115 & ~n8916 ;
  assign n8918 = n8915 | n8917 ;
  buffer buf_n8919( .i (n8918), .o (n8919) );
  assign n8920 = n8120 & n8919 ;
  assign n8921 = n8097 & ~n8916 ;
  assign n8922 = n8109 & n8916 ;
  assign n8923 = n8921 | n8922 ;
  buffer buf_n8924( .i (n8923), .o (n8924) );
  assign n8925 = ~n8120 & n8924 ;
  assign n8926 = n8920 | n8925 ;
  buffer buf_n8927( .i (n8926), .o (n8927) );
  assign n8928 = n3564 & ~n8927 ;
  assign n8929 = n8914 & ~n8928 ;
  assign n8930 = ~n8710 & n8929 ;
  assign n8931 = n8897 | n8930 ;
  assign n8932 = ~n8861 & n8931 ;
  assign n8933 = n8862 | n8932 ;
  buffer buf_n8934( .i (n8933), .o (n8934) );
  buffer buf_n8935( .i (n6100), .o (n8935) );
  assign n8936 = n8934 & n8935 ;
  assign n8937 = n2496 & ~n6081 ;
  assign n8938 = n2494 & ~n2759 ;
  buffer buf_n8939( .i (n8938), .o (n8939) );
  assign n8940 = ~n2493 & n2758 ;
  buffer buf_n8941( .i (n8940), .o (n8941) );
  assign n8943 = n6068 & n8941 ;
  assign n8944 = n8939 | n8943 ;
  assign n8945 = n8937 | n8944 ;
  assign n8946 = n2494 & n2759 ;
  assign n8947 = n6057 & ~n8946 ;
  buffer buf_n8948( .i (n8947), .o (n8948) );
  assign n8949 = n6089 | n8948 ;
  assign n8950 = n8945 & ~n8949 ;
  buffer buf_n8951( .i (n8950), .o (n8951) );
  buffer buf_n8952( .i (n8951), .o (n8952) );
  assign n8953 = n8699 | n8952 ;
  buffer buf_n8954( .i (n8953), .o (n8954) );
  buffer buf_n8955( .i (n8954), .o (n8955) );
  buffer buf_n8956( .i (n8955), .o (n8956) );
  buffer buf_n8957( .i (n8956), .o (n8957) );
  buffer buf_n8958( .i (n8957), .o (n8958) );
  buffer buf_n8959( .i (n8958), .o (n8959) );
  buffer buf_n8960( .i (n8959), .o (n8960) );
  buffer buf_n8961( .i (n8960), .o (n8961) );
  assign n8962 = n8936 | n8961 ;
  buffer buf_n4460( .i (n4459), .o (n4460) );
  buffer buf_n4461( .i (n4460), .o (n4461) );
  buffer buf_n4462( .i (n4461), .o (n4462) );
  buffer buf_n4463( .i (n4462), .o (n4463) );
  buffer buf_n4464( .i (n4463), .o (n4464) );
  buffer buf_n4465( .i (n4464), .o (n4465) );
  buffer buf_n4466( .i (n4465), .o (n4466) );
  buffer buf_n4467( .i (n4466), .o (n4467) );
  buffer buf_n4468( .i (n4467), .o (n4468) );
  buffer buf_n4469( .i (n4468), .o (n4469) );
  buffer buf_n4470( .i (n4469), .o (n4470) );
  buffer buf_n4471( .i (n4470), .o (n4471) );
  buffer buf_n4472( .i (n4471), .o (n4472) );
  assign n8963 = ~n3903 & n4472 ;
  buffer buf_n8964( .i (n8963), .o (n8964) );
  buffer buf_n8965( .i (n8964), .o (n8965) );
  buffer buf_n8966( .i (n8965), .o (n8966) );
  buffer buf_n8967( .i (n8966), .o (n8967) );
  buffer buf_n8968( .i (n8967), .o (n8968) );
  assign n8969 = n5936 & ~n8968 ;
  buffer buf_n8970( .i (n8969), .o (n8970) );
  buffer buf_n8971( .i (n8970), .o (n8971) );
  assign n8972 = n8699 & ~n8971 ;
  assign n8973 = n5876 & ~n8972 ;
  buffer buf_n8974( .i (n8973), .o (n8974) );
  buffer buf_n8975( .i (n8974), .o (n8975) );
  buffer buf_n8976( .i (n8975), .o (n8976) );
  buffer buf_n8977( .i (n8976), .o (n8977) );
  buffer buf_n8978( .i (n8977), .o (n8978) );
  buffer buf_n8979( .i (n8978), .o (n8979) );
  buffer buf_n8980( .i (n8979), .o (n8980) );
  buffer buf_n8981( .i (n8980), .o (n8981) );
  assign n8982 = n8962 & n8981 ;
  buffer buf_n8983( .i (n8982), .o (n8983) );
  buffer buf_n8984( .i (n8983), .o (n8984) );
  buffer buf_n8985( .i (n8984), .o (n8985) );
  buffer buf_n8986( .i (n8985), .o (n8986) );
  buffer buf_n8987( .i (n8986), .o (n8987) );
  buffer buf_n8988( .i (n8987), .o (n8988) );
  buffer buf_n8989( .i (n8988), .o (n8989) );
  buffer buf_n8990( .i (n8989), .o (n8990) );
  buffer buf_n8991( .i (n8990), .o (n8991) );
  buffer buf_n8992( .i (n8991), .o (n8992) );
  buffer buf_n8993( .i (n8992), .o (n8993) );
  buffer buf_n8994( .i (n8993), .o (n8994) );
  buffer buf_n8995( .i (n8994), .o (n8995) );
  buffer buf_n8996( .i (n8995), .o (n8996) );
  buffer buf_n8997( .i (n8996), .o (n8997) );
  buffer buf_n8998( .i (n8997), .o (n8998) );
  buffer buf_n8999( .i (n8998), .o (n8999) );
  buffer buf_n9000( .i (n8999), .o (n9000) );
  buffer buf_n9001( .i (n9000), .o (n9001) );
  buffer buf_n9002( .i (n9001), .o (n9002) );
  buffer buf_n9003( .i (n9002), .o (n9003) );
  buffer buf_n9004( .i (n9003), .o (n9004) );
  buffer buf_n9005( .i (n9004), .o (n9005) );
  buffer buf_n9006( .i (n9005), .o (n9006) );
  buffer buf_n9007( .i (n9006), .o (n9007) );
  buffer buf_n9008( .i (n9007), .o (n9008) );
  buffer buf_n9009( .i (n9008), .o (n9009) );
  buffer buf_n9010( .i (n9009), .o (n9010) );
  buffer buf_n9011( .i (n9010), .o (n9011) );
  buffer buf_n9012( .i (n9011), .o (n9012) );
  buffer buf_n9013( .i (n9012), .o (n9013) );
  buffer buf_n9014( .i (n9013), .o (n9014) );
  buffer buf_n9015( .i (n9014), .o (n9015) );
  buffer buf_n9016( .i (n9015), .o (n9016) );
  buffer buf_n9017( .i (n9016), .o (n9017) );
  buffer buf_n9018( .i (n9017), .o (n9018) );
  buffer buf_n9019( .i (n9018), .o (n9019) );
  buffer buf_n9020( .i (n9019), .o (n9020) );
  buffer buf_n9021( .i (n9020), .o (n9021) );
  buffer buf_n9022( .i (n9021), .o (n9022) );
  buffer buf_n9023( .i (n9022), .o (n9023) );
  buffer buf_n9024( .i (n9023), .o (n9024) );
  buffer buf_n9025( .i (n9024), .o (n9025) );
  buffer buf_n9026( .i (n9025), .o (n9026) );
  buffer buf_n9027( .i (n9026), .o (n9027) );
  buffer buf_n9028( .i (n9027), .o (n9028) );
  buffer buf_n9029( .i (n9028), .o (n9029) );
  buffer buf_n9030( .i (n9029), .o (n9030) );
  buffer buf_n9031( .i (n9030), .o (n9031) );
  buffer buf_n9032( .i (n9031), .o (n9032) );
  buffer buf_n9033( .i (n9032), .o (n9033) );
  buffer buf_n9034( .i (n9033), .o (n9034) );
  buffer buf_n9035( .i (n9034), .o (n9035) );
  buffer buf_n9036( .i (n9035), .o (n9036) );
  buffer buf_n9037( .i (n9036), .o (n9037) );
  buffer buf_n9038( .i (n9037), .o (n9038) );
  buffer buf_n9039( .i (n9038), .o (n9039) );
  buffer buf_n9040( .i (n9039), .o (n9040) );
  buffer buf_n9041( .i (n9040), .o (n9041) );
  buffer buf_n9042( .i (n9041), .o (n9042) );
  buffer buf_n9043( .i (n9042), .o (n9043) );
  buffer buf_n9044( .i (n9043), .o (n9044) );
  buffer buf_n9045( .i (n9044), .o (n9045) );
  buffer buf_n9046( .i (n9045), .o (n9046) );
  buffer buf_n9047( .i (n9046), .o (n9047) );
  buffer buf_n9048( .i (n9047), .o (n9048) );
  buffer buf_n9049( .i (n9048), .o (n9049) );
  buffer buf_n9050( .i (n9049), .o (n9050) );
  buffer buf_n9051( .i (n9050), .o (n9051) );
  buffer buf_n9052( .i (n9051), .o (n9052) );
  buffer buf_n9053( .i (n9052), .o (n9053) );
  buffer buf_n9054( .i (n9053), .o (n9054) );
  buffer buf_n9055( .i (n9054), .o (n9055) );
  buffer buf_n9056( .i (n9055), .o (n9056) );
  buffer buf_n9057( .i (n9056), .o (n9057) );
  buffer buf_n9058( .i (n9057), .o (n9058) );
  buffer buf_n9059( .i (n9058), .o (n9059) );
  buffer buf_n9060( .i (n9059), .o (n9060) );
  buffer buf_n9061( .i (n9060), .o (n9061) );
  buffer buf_n9062( .i (n9061), .o (n9062) );
  buffer buf_n9063( .i (n9062), .o (n9063) );
  buffer buf_n9064( .i (n9063), .o (n9064) );
  buffer buf_n9065( .i (n9064), .o (n9065) );
  buffer buf_n9066( .i (n9065), .o (n9066) );
  buffer buf_n9067( .i (n9066), .o (n9067) );
  buffer buf_n9068( .i (n9067), .o (n9068) );
  buffer buf_n9069( .i (n9068), .o (n9069) );
  buffer buf_n9070( .i (n9069), .o (n9070) );
  buffer buf_n9071( .i (n9070), .o (n9071) );
  buffer buf_n9072( .i (n9071), .o (n9072) );
  buffer buf_n9073( .i (n9072), .o (n9073) );
  buffer buf_n9074( .i (n9073), .o (n9074) );
  buffer buf_n9075( .i (n9074), .o (n9075) );
  buffer buf_n9076( .i (n9075), .o (n9076) );
  buffer buf_n9077( .i (n9076), .o (n9077) );
  buffer buf_n9078( .i (n9077), .o (n9078) );
  buffer buf_n9079( .i (n9078), .o (n9079) );
  buffer buf_n9080( .i (n9079), .o (n9080) );
  buffer buf_n9081( .i (n9080), .o (n9081) );
  buffer buf_n9082( .i (n9081), .o (n9082) );
  buffer buf_n9083( .i (n9082), .o (n9083) );
  buffer buf_n9084( .i (n9083), .o (n9084) );
  buffer buf_n9085( .i (n9084), .o (n9085) );
  buffer buf_n9086( .i (n9085), .o (n9086) );
  buffer buf_n9087( .i (n9086), .o (n9087) );
  buffer buf_n9088( .i (n9087), .o (n9088) );
  buffer buf_n9089( .i (n9088), .o (n9089) );
  buffer buf_n9090( .i (n9089), .o (n9090) );
  buffer buf_n9091( .i (n9090), .o (n9091) );
  assign n9092 = n8860 | n9091 ;
  buffer buf_n9093( .i (n9092), .o (n9093) );
  buffer buf_n9094( .i (n9093), .o (n9094) );
  buffer buf_n9095( .i (n9094), .o (n9095) );
  buffer buf_n4787( .i (n4786), .o (n4787) );
  buffer buf_n4788( .i (n4787), .o (n4788) );
  assign n9096 = ~n5036 & n5039 ;
  buffer buf_n9097( .i (n9096), .o (n9097) );
  assign n9098 = n4788 | n9097 ;
  assign n9099 = n4788 & n9097 ;
  assign n9100 = n9098 & ~n9099 ;
  buffer buf_n9101( .i (n9100), .o (n9101) );
  buffer buf_n9102( .i (n9101), .o (n9102) );
  buffer buf_n9103( .i (n9102), .o (n9103) );
  buffer buf_n9104( .i (n9103), .o (n9104) );
  buffer buf_n9105( .i (n9104), .o (n9105) );
  buffer buf_n9106( .i (n9105), .o (n9106) );
  buffer buf_n9107( .i (n9106), .o (n9107) );
  buffer buf_n9108( .i (n9107), .o (n9108) );
  buffer buf_n9109( .i (n9108), .o (n9109) );
  buffer buf_n9110( .i (n9109), .o (n9110) );
  buffer buf_n9111( .i (n9110), .o (n9111) );
  buffer buf_n9112( .i (n9111), .o (n9112) );
  buffer buf_n9113( .i (n9112), .o (n9113) );
  buffer buf_n9114( .i (n9113), .o (n9114) );
  buffer buf_n9115( .i (n9114), .o (n9115) );
  buffer buf_n9116( .i (n9115), .o (n9116) );
  buffer buf_n9117( .i (n9116), .o (n9117) );
  buffer buf_n9118( .i (n9117), .o (n9118) );
  buffer buf_n9119( .i (n9118), .o (n9119) );
  buffer buf_n9120( .i (n9119), .o (n9120) );
  buffer buf_n9121( .i (n9120), .o (n9121) );
  buffer buf_n9122( .i (n9121), .o (n9122) );
  buffer buf_n9123( .i (n9122), .o (n9123) );
  buffer buf_n9124( .i (n9123), .o (n9124) );
  buffer buf_n9125( .i (n9124), .o (n9125) );
  buffer buf_n9126( .i (n9125), .o (n9126) );
  buffer buf_n9127( .i (n9126), .o (n9127) );
  buffer buf_n9128( .i (n9127), .o (n9128) );
  buffer buf_n9129( .i (n9128), .o (n9129) );
  buffer buf_n9130( .i (n9129), .o (n9130) );
  buffer buf_n9131( .i (n9130), .o (n9131) );
  buffer buf_n9132( .i (n9131), .o (n9132) );
  buffer buf_n9133( .i (n9132), .o (n9133) );
  buffer buf_n9134( .i (n9133), .o (n9134) );
  buffer buf_n9135( .i (n9134), .o (n9135) );
  buffer buf_n9136( .i (n9135), .o (n9136) );
  buffer buf_n9137( .i (n9136), .o (n9137) );
  buffer buf_n9138( .i (n9137), .o (n9138) );
  buffer buf_n9139( .i (n9138), .o (n9139) );
  buffer buf_n9140( .i (n9139), .o (n9140) );
  buffer buf_n9141( .i (n9140), .o (n9141) );
  buffer buf_n9142( .i (n9141), .o (n9142) );
  buffer buf_n9143( .i (n9142), .o (n9143) );
  buffer buf_n9144( .i (n9143), .o (n9144) );
  buffer buf_n9145( .i (n9144), .o (n9145) );
  buffer buf_n9146( .i (n9145), .o (n9146) );
  buffer buf_n9147( .i (n9146), .o (n9147) );
  buffer buf_n9148( .i (n9147), .o (n9148) );
  buffer buf_n9149( .i (n9148), .o (n9149) );
  buffer buf_n9150( .i (n9149), .o (n9150) );
  buffer buf_n9151( .i (n9150), .o (n9151) );
  buffer buf_n9152( .i (n9151), .o (n9152) );
  buffer buf_n9153( .i (n9152), .o (n9153) );
  buffer buf_n9154( .i (n9153), .o (n9154) );
  buffer buf_n9155( .i (n9154), .o (n9155) );
  buffer buf_n9156( .i (n9155), .o (n9156) );
  buffer buf_n9157( .i (n9156), .o (n9157) );
  buffer buf_n9158( .i (n9157), .o (n9158) );
  buffer buf_n9159( .i (n9158), .o (n9159) );
  buffer buf_n9160( .i (n9159), .o (n9160) );
  buffer buf_n9161( .i (n9160), .o (n9161) );
  buffer buf_n9162( .i (n9161), .o (n9162) );
  buffer buf_n9163( .i (n9162), .o (n9163) );
  buffer buf_n9164( .i (n9163), .o (n9164) );
  buffer buf_n9165( .i (n9164), .o (n9165) );
  buffer buf_n9166( .i (n9165), .o (n9166) );
  buffer buf_n9167( .i (n9166), .o (n9167) );
  buffer buf_n9168( .i (n9167), .o (n9168) );
  buffer buf_n9169( .i (n9168), .o (n9169) );
  buffer buf_n9170( .i (n9169), .o (n9170) );
  buffer buf_n9171( .i (n9170), .o (n9171) );
  buffer buf_n9172( .i (n9171), .o (n9172) );
  buffer buf_n9173( .i (n9172), .o (n9173) );
  buffer buf_n9174( .i (n9173), .o (n9174) );
  buffer buf_n9175( .i (n9174), .o (n9175) );
  buffer buf_n9176( .i (n9175), .o (n9176) );
  buffer buf_n9177( .i (n9176), .o (n9177) );
  buffer buf_n9178( .i (n9177), .o (n9178) );
  buffer buf_n9179( .i (n9178), .o (n9179) );
  buffer buf_n9180( .i (n9179), .o (n9180) );
  buffer buf_n9181( .i (n9180), .o (n9181) );
  buffer buf_n9182( .i (n9181), .o (n9182) );
  buffer buf_n9183( .i (n9182), .o (n9183) );
  buffer buf_n9184( .i (n9183), .o (n9184) );
  buffer buf_n9185( .i (n9184), .o (n9185) );
  buffer buf_n9186( .i (n9185), .o (n9186) );
  buffer buf_n9187( .i (n9186), .o (n9187) );
  buffer buf_n9188( .i (n9187), .o (n9188) );
  buffer buf_n9189( .i (n9188), .o (n9189) );
  buffer buf_n9190( .i (n9189), .o (n9190) );
  buffer buf_n9191( .i (n9190), .o (n9191) );
  buffer buf_n9192( .i (n9191), .o (n9192) );
  buffer buf_n9193( .i (n9192), .o (n9193) );
  buffer buf_n9194( .i (n9193), .o (n9194) );
  buffer buf_n9195( .i (n9194), .o (n9195) );
  buffer buf_n9196( .i (n9195), .o (n9196) );
  buffer buf_n9197( .i (n9196), .o (n9197) );
  buffer buf_n9198( .i (n9197), .o (n9198) );
  buffer buf_n9199( .i (n9198), .o (n9199) );
  buffer buf_n9200( .i (n9199), .o (n9200) );
  buffer buf_n9201( .i (n9200), .o (n9201) );
  buffer buf_n9202( .i (n9201), .o (n9202) );
  buffer buf_n9203( .i (n9202), .o (n9203) );
  buffer buf_n9204( .i (n9203), .o (n9204) );
  buffer buf_n9205( .i (n9204), .o (n9205) );
  buffer buf_n9206( .i (n9205), .o (n9206) );
  buffer buf_n9207( .i (n9206), .o (n9207) );
  buffer buf_n9208( .i (n9207), .o (n9208) );
  buffer buf_n9209( .i (n9208), .o (n9209) );
  buffer buf_n9210( .i (n9209), .o (n9210) );
  buffer buf_n9211( .i (n9210), .o (n9211) );
  buffer buf_n9212( .i (n9211), .o (n9212) );
  assign n9213 = n1009 & n1179 ;
  buffer buf_n9214( .i (n9213), .o (n9214) );
  assign n9216 = n6080 & n9214 ;
  assign n9217 = n1010 & n6067 ;
  assign n9218 = n1181 | n9217 ;
  assign n9219 = ~n9216 & n9218 ;
  assign n9220 = n6059 | n9219 ;
  buffer buf_n9215( .i (n9214), .o (n9215) );
  assign n9221 = n6058 & ~n9215 ;
  assign n9222 = n6089 | n9221 ;
  assign n9223 = n9220 & ~n9222 ;
  buffer buf_n9224( .i (n9223), .o (n9224) );
  buffer buf_n9225( .i (n9224), .o (n9225) );
  assign n9226 = n8699 | n9225 ;
  buffer buf_n9227( .i (n9226), .o (n9227) );
  buffer buf_n9228( .i (n9227), .o (n9228) );
  buffer buf_n9229( .i (n9228), .o (n9229) );
  buffer buf_n9230( .i (n9229), .o (n9230) );
  buffer buf_n9231( .i (n9230), .o (n9231) );
  buffer buf_n9232( .i (n9231), .o (n9232) );
  buffer buf_n9233( .i (n9232), .o (n9233) );
  buffer buf_n9234( .i (n9233), .o (n9234) );
  assign n9235 = n6044 & n8861 ;
  assign n9236 = n8888 & ~n8889 ;
  buffer buf_n8667( .i (n8666), .o (n8667) );
  assign n9237 = n8667 & n8889 ;
  assign n9238 = n9236 | n9237 ;
  buffer buf_n9239( .i (n9238), .o (n9239) );
  assign n9240 = ~n8893 & n9239 ;
  buffer buf_n9241( .i (n8650), .o (n9241) );
  assign n9242 = n8648 & n9241 ;
  assign n9243 = n8659 & ~n9241 ;
  assign n9244 = n9242 | n9243 ;
  buffer buf_n9245( .i (n9244), .o (n9245) );
  buffer buf_n9246( .i (n9245), .o (n9246) );
  assign n9247 = n8893 & n9246 ;
  assign n9248 = n9240 | n9247 ;
  buffer buf_n9249( .i (n9248), .o (n9249) );
  buffer buf_n9250( .i (n8642), .o (n9250) );
  assign n9251 = ~n9249 & n9250 ;
  assign n9252 = n8882 & n8889 ;
  buffer buf_n9253( .i (n9241), .o (n9253) );
  assign n9254 = n8873 & ~n9253 ;
  assign n9255 = n9252 | n9254 ;
  buffer buf_n9256( .i (n9255), .o (n9256) );
  buffer buf_n9257( .i (n9256), .o (n9257) );
  buffer buf_n9258( .i (n8893), .o (n9258) );
  assign n9259 = ~n9257 & n9258 ;
  buffer buf_n8867( .i (n8866), .o (n8867) );
  assign n9260 = n8120 & n8867 ;
  buffer buf_n9261( .i (n9253), .o (n9261) );
  assign n9262 = n8919 & ~n9261 ;
  assign n9263 = n9260 | n9262 ;
  buffer buf_n9264( .i (n9263), .o (n9264) );
  assign n9265 = n9258 | n9264 ;
  assign n9266 = ~n9259 & n9265 ;
  assign n9267 = n9250 | n9266 ;
  assign n9268 = ~n9251 & n9267 ;
  assign n9269 = ~n8861 & n9268 ;
  assign n9270 = n9235 | n9269 ;
  buffer buf_n9271( .i (n9270), .o (n9271) );
  assign n9272 = n8935 & n9271 ;
  assign n9273 = n9234 | n9272 ;
  buffer buf_n9274( .i (n9273), .o (n9274) );
  buffer buf_n5951( .i (n5950), .o (n5951) );
  assign n9275 = ~n135 & n6153 ;
  assign n9276 = n5951 | n9275 ;
  buffer buf_n9277( .i (n9276), .o (n9277) );
  assign n9278 = n5928 & ~n9277 ;
  assign n9279 = n5885 & ~n9278 ;
  assign n9280 = n9274 & n9279 ;
  buffer buf_n9281( .i (n9280), .o (n9281) );
  buffer buf_n9282( .i (n9281), .o (n9282) );
  buffer buf_n9283( .i (n9282), .o (n9283) );
  buffer buf_n9284( .i (n9283), .o (n9284) );
  buffer buf_n9285( .i (n9284), .o (n9285) );
  buffer buf_n9286( .i (n9285), .o (n9286) );
  buffer buf_n9287( .i (n9286), .o (n9287) );
  buffer buf_n9288( .i (n9287), .o (n9288) );
  buffer buf_n9289( .i (n9288), .o (n9289) );
  buffer buf_n9290( .i (n9289), .o (n9290) );
  buffer buf_n9291( .i (n9290), .o (n9291) );
  buffer buf_n9292( .i (n9291), .o (n9292) );
  buffer buf_n9293( .i (n9292), .o (n9293) );
  buffer buf_n9294( .i (n9293), .o (n9294) );
  buffer buf_n9295( .i (n9294), .o (n9295) );
  buffer buf_n9296( .i (n9295), .o (n9296) );
  buffer buf_n9297( .i (n9296), .o (n9297) );
  buffer buf_n9298( .i (n9297), .o (n9298) );
  buffer buf_n9299( .i (n9298), .o (n9299) );
  buffer buf_n9300( .i (n9299), .o (n9300) );
  buffer buf_n9301( .i (n9300), .o (n9301) );
  buffer buf_n9302( .i (n9301), .o (n9302) );
  buffer buf_n9303( .i (n9302), .o (n9303) );
  buffer buf_n9304( .i (n9303), .o (n9304) );
  buffer buf_n9305( .i (n9304), .o (n9305) );
  buffer buf_n9306( .i (n9305), .o (n9306) );
  buffer buf_n9307( .i (n9306), .o (n9307) );
  buffer buf_n9308( .i (n9307), .o (n9308) );
  buffer buf_n9309( .i (n9308), .o (n9309) );
  buffer buf_n9310( .i (n9309), .o (n9310) );
  buffer buf_n9311( .i (n9310), .o (n9311) );
  buffer buf_n9312( .i (n9311), .o (n9312) );
  buffer buf_n9313( .i (n9312), .o (n9313) );
  buffer buf_n9314( .i (n9313), .o (n9314) );
  buffer buf_n9315( .i (n9314), .o (n9315) );
  buffer buf_n9316( .i (n9315), .o (n9316) );
  buffer buf_n9317( .i (n9316), .o (n9317) );
  buffer buf_n9318( .i (n9317), .o (n9318) );
  buffer buf_n9319( .i (n9318), .o (n9319) );
  buffer buf_n9320( .i (n9319), .o (n9320) );
  buffer buf_n9321( .i (n9320), .o (n9321) );
  buffer buf_n9322( .i (n9321), .o (n9322) );
  buffer buf_n9323( .i (n9322), .o (n9323) );
  buffer buf_n9324( .i (n9323), .o (n9324) );
  buffer buf_n9325( .i (n9324), .o (n9325) );
  buffer buf_n9326( .i (n9325), .o (n9326) );
  buffer buf_n9327( .i (n9326), .o (n9327) );
  buffer buf_n9328( .i (n9327), .o (n9328) );
  buffer buf_n9329( .i (n9328), .o (n9329) );
  buffer buf_n9330( .i (n9329), .o (n9330) );
  buffer buf_n9331( .i (n9330), .o (n9331) );
  buffer buf_n9332( .i (n9331), .o (n9332) );
  buffer buf_n9333( .i (n9332), .o (n9333) );
  buffer buf_n9334( .i (n9333), .o (n9334) );
  buffer buf_n9335( .i (n9334), .o (n9335) );
  buffer buf_n9336( .i (n9335), .o (n9336) );
  buffer buf_n9337( .i (n9336), .o (n9337) );
  buffer buf_n9338( .i (n9337), .o (n9338) );
  buffer buf_n9339( .i (n9338), .o (n9339) );
  buffer buf_n9340( .i (n9339), .o (n9340) );
  buffer buf_n9341( .i (n9340), .o (n9341) );
  buffer buf_n9342( .i (n9341), .o (n9342) );
  buffer buf_n9343( .i (n9342), .o (n9343) );
  buffer buf_n9344( .i (n9343), .o (n9344) );
  buffer buf_n9345( .i (n9344), .o (n9345) );
  buffer buf_n9346( .i (n9345), .o (n9346) );
  buffer buf_n9347( .i (n9346), .o (n9347) );
  buffer buf_n9348( .i (n9347), .o (n9348) );
  buffer buf_n9349( .i (n9348), .o (n9349) );
  buffer buf_n9350( .i (n9349), .o (n9350) );
  buffer buf_n9351( .i (n9350), .o (n9351) );
  buffer buf_n9352( .i (n9351), .o (n9352) );
  buffer buf_n9353( .i (n9352), .o (n9353) );
  buffer buf_n9354( .i (n9353), .o (n9354) );
  buffer buf_n9355( .i (n9354), .o (n9355) );
  buffer buf_n9356( .i (n9355), .o (n9356) );
  buffer buf_n9357( .i (n9356), .o (n9357) );
  buffer buf_n9358( .i (n9357), .o (n9358) );
  buffer buf_n9359( .i (n9358), .o (n9359) );
  buffer buf_n7238( .i (n7237), .o (n7238) );
  buffer buf_n7239( .i (n7238), .o (n7239) );
  assign n9360 = ~n7158 & n7241 ;
  buffer buf_n9361( .i (n9360), .o (n9361) );
  assign n9362 = n7239 | n9361 ;
  assign n9363 = n7239 & n9361 ;
  assign n9364 = n9362 & ~n9363 ;
  buffer buf_n9365( .i (n9364), .o (n9365) );
  assign n9400 = ~n5711 & n9365 ;
  assign n9401 = n9359 | n9400 ;
  buffer buf_n9402( .i (n9401), .o (n9402) );
  buffer buf_n9403( .i (n9402), .o (n9403) );
  buffer buf_n9404( .i (n9403), .o (n9404) );
  buffer buf_n9405( .i (n9404), .o (n9405) );
  buffer buf_n9406( .i (n9405), .o (n9406) );
  buffer buf_n9407( .i (n9406), .o (n9407) );
  buffer buf_n9408( .i (n9407), .o (n9408) );
  buffer buf_n9409( .i (n9408), .o (n9409) );
  buffer buf_n9410( .i (n9409), .o (n9410) );
  buffer buf_n9411( .i (n9410), .o (n9411) );
  buffer buf_n9412( .i (n9411), .o (n9412) );
  buffer buf_n9413( .i (n9412), .o (n9413) );
  buffer buf_n9414( .i (n9413), .o (n9414) );
  buffer buf_n9415( .i (n9414), .o (n9415) );
  buffer buf_n9416( .i (n9415), .o (n9416) );
  buffer buf_n9417( .i (n9416), .o (n9417) );
  buffer buf_n9418( .i (n9417), .o (n9418) );
  buffer buf_n9419( .i (n9418), .o (n9419) );
  buffer buf_n9420( .i (n9419), .o (n9420) );
  buffer buf_n9421( .i (n9420), .o (n9421) );
  buffer buf_n9422( .i (n9421), .o (n9422) );
  buffer buf_n9423( .i (n9422), .o (n9423) );
  buffer buf_n9424( .i (n9423), .o (n9424) );
  buffer buf_n9425( .i (n9424), .o (n9425) );
  buffer buf_n9426( .i (n9425), .o (n9426) );
  buffer buf_n9427( .i (n9426), .o (n9427) );
  buffer buf_n9428( .i (n9427), .o (n9428) );
  buffer buf_n9429( .i (n9428), .o (n9429) );
  buffer buf_n9430( .i (n9429), .o (n9430) );
  buffer buf_n9431( .i (n9430), .o (n9431) );
  buffer buf_n9432( .i (n9431), .o (n9432) );
  buffer buf_n9433( .i (n9432), .o (n9433) );
  assign n9434 = ~n5634 & n9101 ;
  buffer buf_n3962( .i (n3961), .o (n3962) );
  buffer buf_n3963( .i (n3962), .o (n3963) );
  buffer buf_n3964( .i (n3963), .o (n3964) );
  buffer buf_n3965( .i (n3964), .o (n3965) );
  buffer buf_n3966( .i (n3965), .o (n3966) );
  buffer buf_n3967( .i (n3966), .o (n3967) );
  buffer buf_n3968( .i (n3967), .o (n3968) );
  buffer buf_n3969( .i (n3968), .o (n3969) );
  buffer buf_n3970( .i (n3969), .o (n3970) );
  buffer buf_n3971( .i (n3970), .o (n3971) );
  buffer buf_n3972( .i (n3971), .o (n3972) );
  assign n9435 = n3972 & n6078 ;
  assign n9436 = n4221 & ~n6053 ;
  buffer buf_n9437( .i (n9436), .o (n9437) );
  buffer buf_n9438( .i (n9437), .o (n9438) );
  assign n9439 = ~n9435 & n9438 ;
  assign n9440 = n3972 & ~n9437 ;
  assign n9441 = n4223 | n6066 ;
  assign n9442 = n9440 & n9441 ;
  assign n9443 = n9439 | n9442 ;
  buffer buf_n9444( .i (n9443), .o (n9444) );
  buffer buf_n9445( .i (n9444), .o (n9445) );
  assign n9446 = ~n6090 & n9445 ;
  buffer buf_n9447( .i (n9446), .o (n9447) );
  buffer buf_n9448( .i (n9447), .o (n9448) );
  buffer buf_n9449( .i (n5918), .o (n9449) );
  assign n9450 = n9448 | n9449 ;
  buffer buf_n9451( .i (n9450), .o (n9451) );
  buffer buf_n9452( .i (n9451), .o (n9452) );
  buffer buf_n9453( .i (n9452), .o (n9453) );
  buffer buf_n9454( .i (n9453), .o (n9454) );
  buffer buf_n9455( .i (n9454), .o (n9455) );
  buffer buf_n9456( .i (n9455), .o (n9456) );
  buffer buf_n9457( .i (n9456), .o (n9457) );
  buffer buf_n9458( .i (n9457), .o (n9458) );
  buffer buf_n9459( .i (n9458), .o (n9459) );
  buffer buf_n5969( .i (n5968), .o (n5969) );
  buffer buf_n9460( .i (n8672), .o (n9460) );
  assign n9461 = n6143 & ~n9460 ;
  assign n9462 = n5969 | n9461 ;
  buffer buf_n9463( .i (n9462), .o (n9463) );
  assign n9464 = n9250 & ~n9463 ;
  buffer buf_n6281( .i (n6280), .o (n6281) );
  assign n9465 = n6281 & ~n9460 ;
  assign n9466 = n6129 & n9460 ;
  assign n9467 = n9465 | n9466 ;
  buffer buf_n9468( .i (n9467), .o (n9468) );
  assign n9469 = n9250 | n9468 ;
  assign n9470 = ~n9464 & n9469 ;
  buffer buf_n9471( .i (n9470), .o (n9471) );
  assign n9472 = ~n135 & n9471 ;
  assign n9473 = n5951 | n9472 ;
  buffer buf_n9474( .i (n9473), .o (n9474) );
  assign n9475 = n6102 & n9474 ;
  assign n9476 = n9459 | n9475 ;
  assign n9477 = n6003 & n8672 ;
  buffer buf_n9478( .i (n8084), .o (n9478) );
  assign n9479 = n9245 & ~n9478 ;
  assign n9480 = n9477 | n9479 ;
  buffer buf_n9481( .i (n9480), .o (n9481) );
  buffer buf_n9482( .i (n1863), .o (n9482) );
  assign n9483 = n9481 & n9482 ;
  assign n9484 = n132 | n9483 ;
  assign n9485 = n9256 & ~n9460 ;
  buffer buf_n9486( .i (n9478), .o (n9486) );
  assign n9487 = n9239 & n9486 ;
  assign n9488 = n9485 | n9487 ;
  buffer buf_n9489( .i (n9488), .o (n9489) );
  buffer buf_n9490( .i (n9482), .o (n9490) );
  assign n9491 = n9489 & ~n9490 ;
  assign n9492 = n9484 | n9491 ;
  buffer buf_n9493( .i (n9492), .o (n9493) );
  assign n9494 = ~n5965 & n9478 ;
  assign n9495 = n6037 | n9478 ;
  assign n9496 = ~n9494 & n9495 ;
  buffer buf_n9497( .i (n9496), .o (n9497) );
  assign n9498 = ~n9482 & n9497 ;
  assign n9499 = n6150 | n9498 ;
  buffer buf_n9500( .i (n9499), .o (n9500) );
  buffer buf_n9501( .i (n132), .o (n9501) );
  buffer buf_n9502( .i (n9501), .o (n9502) );
  assign n9503 = ~n9500 & n9502 ;
  assign n9504 = n9493 & ~n9503 ;
  buffer buf_n9505( .i (n9504), .o (n9505) );
  assign n9506 = n5927 & ~n9505 ;
  assign n9507 = n5884 & ~n9506 ;
  buffer buf_n9508( .i (n9507), .o (n9508) );
  assign n9509 = n9476 & n9508 ;
  buffer buf_n9510( .i (n9509), .o (n9510) );
  buffer buf_n9511( .i (n9510), .o (n9511) );
  assign n9512 = n9434 | n9511 ;
  buffer buf_n9513( .i (n9512), .o (n9513) );
  buffer buf_n9514( .i (n9513), .o (n9514) );
  buffer buf_n9515( .i (n9514), .o (n9515) );
  buffer buf_n9516( .i (n9515), .o (n9516) );
  buffer buf_n9517( .i (n9516), .o (n9517) );
  buffer buf_n9518( .i (n9517), .o (n9518) );
  buffer buf_n9519( .i (n9518), .o (n9519) );
  buffer buf_n9520( .i (n9519), .o (n9520) );
  buffer buf_n9521( .i (n9520), .o (n9521) );
  buffer buf_n9522( .i (n9521), .o (n9522) );
  buffer buf_n9523( .i (n9522), .o (n9523) );
  buffer buf_n9524( .i (n9523), .o (n9524) );
  buffer buf_n9525( .i (n9524), .o (n9525) );
  buffer buf_n9526( .i (n9525), .o (n9526) );
  buffer buf_n9527( .i (n9526), .o (n9527) );
  buffer buf_n9528( .i (n9527), .o (n9528) );
  buffer buf_n9529( .i (n9528), .o (n9529) );
  buffer buf_n9530( .i (n9529), .o (n9530) );
  buffer buf_n9531( .i (n9530), .o (n9531) );
  buffer buf_n9532( .i (n9531), .o (n9532) );
  buffer buf_n9533( .i (n9532), .o (n9533) );
  buffer buf_n9534( .i (n9533), .o (n9534) );
  buffer buf_n9535( .i (n9534), .o (n9535) );
  buffer buf_n9536( .i (n9535), .o (n9536) );
  buffer buf_n9537( .i (n9536), .o (n9537) );
  buffer buf_n9538( .i (n9537), .o (n9538) );
  buffer buf_n9539( .i (n9538), .o (n9539) );
  buffer buf_n9540( .i (n9539), .o (n9540) );
  buffer buf_n9541( .i (n9540), .o (n9541) );
  buffer buf_n9542( .i (n9541), .o (n9542) );
  buffer buf_n9543( .i (n9542), .o (n9543) );
  buffer buf_n9544( .i (n9543), .o (n9544) );
  buffer buf_n9545( .i (n9544), .o (n9545) );
  buffer buf_n9546( .i (n9545), .o (n9546) );
  buffer buf_n9547( .i (n9546), .o (n9547) );
  buffer buf_n9548( .i (n9547), .o (n9548) );
  buffer buf_n9549( .i (n9548), .o (n9549) );
  buffer buf_n9550( .i (n9549), .o (n9550) );
  buffer buf_n9551( .i (n9550), .o (n9551) );
  buffer buf_n9552( .i (n9551), .o (n9552) );
  buffer buf_n9553( .i (n9552), .o (n9553) );
  buffer buf_n9554( .i (n9553), .o (n9554) );
  buffer buf_n9555( .i (n9554), .o (n9555) );
  buffer buf_n9556( .i (n9555), .o (n9556) );
  buffer buf_n9557( .i (n9556), .o (n9557) );
  buffer buf_n9558( .i (n9557), .o (n9558) );
  buffer buf_n9559( .i (n9558), .o (n9559) );
  buffer buf_n9560( .i (n9559), .o (n9560) );
  buffer buf_n9561( .i (n9560), .o (n9561) );
  buffer buf_n9562( .i (n9561), .o (n9562) );
  buffer buf_n9563( .i (n9562), .o (n9563) );
  buffer buf_n9564( .i (n9563), .o (n9564) );
  buffer buf_n9565( .i (n9564), .o (n9565) );
  buffer buf_n9566( .i (n9565), .o (n9566) );
  buffer buf_n9567( .i (n9566), .o (n9567) );
  buffer buf_n9568( .i (n9567), .o (n9568) );
  buffer buf_n9569( .i (n9568), .o (n9569) );
  buffer buf_n9570( .i (n9569), .o (n9570) );
  buffer buf_n9571( .i (n9570), .o (n9571) );
  buffer buf_n9572( .i (n9571), .o (n9572) );
  buffer buf_n9573( .i (n9572), .o (n9573) );
  buffer buf_n9574( .i (n9573), .o (n9574) );
  buffer buf_n9575( .i (n9574), .o (n9575) );
  buffer buf_n9576( .i (n9575), .o (n9576) );
  buffer buf_n9577( .i (n9576), .o (n9577) );
  buffer buf_n9578( .i (n9577), .o (n9578) );
  buffer buf_n9579( .i (n9578), .o (n9579) );
  buffer buf_n9580( .i (n9579), .o (n9580) );
  buffer buf_n9581( .i (n9580), .o (n9581) );
  buffer buf_n9582( .i (n9581), .o (n9582) );
  buffer buf_n9583( .i (n9582), .o (n9583) );
  buffer buf_n9584( .i (n9583), .o (n9584) );
  buffer buf_n9585( .i (n9584), .o (n9585) );
  buffer buf_n9586( .i (n9585), .o (n9586) );
  buffer buf_n9587( .i (n9586), .o (n9587) );
  buffer buf_n9588( .i (n9587), .o (n9588) );
  buffer buf_n9589( .i (n9588), .o (n9589) );
  buffer buf_n9590( .i (n9589), .o (n9590) );
  buffer buf_n9591( .i (n9590), .o (n9591) );
  buffer buf_n9592( .i (n9591), .o (n9592) );
  buffer buf_n9593( .i (n9592), .o (n9593) );
  buffer buf_n9594( .i (n9593), .o (n9594) );
  buffer buf_n9595( .i (n9594), .o (n9595) );
  buffer buf_n9596( .i (n9595), .o (n9596) );
  buffer buf_n9597( .i (n9596), .o (n9597) );
  buffer buf_n9598( .i (n9597), .o (n9598) );
  buffer buf_n9599( .i (n9598), .o (n9599) );
  buffer buf_n9600( .i (n9599), .o (n9600) );
  buffer buf_n9601( .i (n9600), .o (n9601) );
  buffer buf_n9602( .i (n9601), .o (n9602) );
  buffer buf_n9603( .i (n9602), .o (n9603) );
  buffer buf_n9604( .i (n9603), .o (n9604) );
  buffer buf_n9605( .i (n9604), .o (n9605) );
  buffer buf_n9606( .i (n9605), .o (n9606) );
  buffer buf_n9607( .i (n9606), .o (n9607) );
  buffer buf_n9608( .i (n9607), .o (n9608) );
  buffer buf_n9609( .i (n9608), .o (n9609) );
  buffer buf_n9610( .i (n9609), .o (n9610) );
  buffer buf_n9611( .i (n9610), .o (n9611) );
  buffer buf_n9612( .i (n9611), .o (n9612) );
  buffer buf_n9613( .i (n9612), .o (n9613) );
  buffer buf_n9614( .i (n9613), .o (n9614) );
  buffer buf_n9615( .i (n9614), .o (n9615) );
  buffer buf_n9616( .i (n9615), .o (n9616) );
  buffer buf_n9617( .i (n9616), .o (n9617) );
  buffer buf_n9618( .i (n9617), .o (n9618) );
  buffer buf_n9619( .i (n9618), .o (n9619) );
  buffer buf_n9620( .i (n9619), .o (n9620) );
  buffer buf_n9621( .i (n9620), .o (n9621) );
  buffer buf_n9622( .i (n9502), .o (n9622) );
  assign n9623 = n8135 & ~n9622 ;
  assign n9624 = n5951 | n9623 ;
  buffer buf_n9625( .i (n9624), .o (n9625) );
  assign n9626 = n6102 & n9625 ;
  buffer buf_n447( .i (n446), .o (n447) );
  assign n9627 = n447 & n1063 ;
  buffer buf_n9628( .i (n9627), .o (n9628) );
  assign n9630 = n6078 & n9628 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n9631 = n448 & n6065 ;
  assign n9632 = n1065 | n9631 ;
  assign n9633 = ~n9630 & n9632 ;
  assign n9634 = n6057 | n9633 ;
  buffer buf_n9629( .i (n9628), .o (n9629) );
  assign n9635 = n6056 & ~n9629 ;
  assign n9636 = n6087 | n9635 ;
  assign n9637 = n9634 & ~n9636 ;
  buffer buf_n9638( .i (n9637), .o (n9638) );
  buffer buf_n9639( .i (n9638), .o (n9639) );
  buffer buf_n9640( .i (n9639), .o (n9640) );
  buffer buf_n9641( .i (n9640), .o (n9641) );
  assign n9642 = n9449 | n9641 ;
  buffer buf_n9643( .i (n9642), .o (n9643) );
  buffer buf_n9644( .i (n9643), .o (n9644) );
  buffer buf_n9645( .i (n9644), .o (n9645) );
  buffer buf_n9646( .i (n9645), .o (n9646) );
  buffer buf_n9647( .i (n9646), .o (n9647) );
  buffer buf_n9648( .i (n9647), .o (n9648) );
  buffer buf_n9649( .i (n9648), .o (n9649) );
  buffer buf_n9650( .i (n9649), .o (n9650) );
  buffer buf_n9651( .i (n9650), .o (n9651) );
  assign n9652 = n9626 | n9651 ;
  assign n9653 = n8165 & n9502 ;
  buffer buf_n6041( .i (n6040), .o (n6041) );
  assign n9654 = ~n6041 & n9490 ;
  assign n9655 = n9249 | n9490 ;
  assign n9656 = ~n9654 & n9655 ;
  assign n9657 = ~n9502 & n9656 ;
  assign n9658 = n9653 | n9657 ;
  buffer buf_n9659( .i (n9658), .o (n9659) );
  buffer buf_n9660( .i (n5926), .o (n9660) );
  assign n9661 = ~n9659 & n9660 ;
  buffer buf_n9662( .i (n5883), .o (n9662) );
  assign n9663 = ~n9661 & n9662 ;
  buffer buf_n9664( .i (n9663), .o (n9664) );
  assign n9665 = n9652 & n9664 ;
  buffer buf_n9666( .i (n9665), .o (n9666) );
  buffer buf_n9667( .i (n9666), .o (n9667) );
  buffer buf_n9668( .i (n9667), .o (n9668) );
  buffer buf_n9669( .i (n9668), .o (n9669) );
  buffer buf_n9670( .i (n9669), .o (n9670) );
  buffer buf_n9671( .i (n9670), .o (n9671) );
  buffer buf_n9672( .i (n9671), .o (n9672) );
  buffer buf_n9673( .i (n9672), .o (n9673) );
  buffer buf_n9674( .i (n9673), .o (n9674) );
  buffer buf_n9675( .i (n9674), .o (n9675) );
  buffer buf_n9676( .i (n9675), .o (n9676) );
  buffer buf_n9677( .i (n9676), .o (n9677) );
  buffer buf_n9678( .i (n9677), .o (n9678) );
  buffer buf_n9679( .i (n9678), .o (n9679) );
  buffer buf_n9680( .i (n9679), .o (n9680) );
  buffer buf_n9681( .i (n9680), .o (n9681) );
  buffer buf_n9682( .i (n9681), .o (n9682) );
  buffer buf_n9683( .i (n9682), .o (n9683) );
  buffer buf_n9684( .i (n9683), .o (n9684) );
  buffer buf_n9685( .i (n9684), .o (n9685) );
  buffer buf_n9686( .i (n9685), .o (n9686) );
  buffer buf_n9687( .i (n9686), .o (n9687) );
  buffer buf_n9688( .i (n9687), .o (n9688) );
  buffer buf_n9689( .i (n9688), .o (n9689) );
  buffer buf_n4755( .i (n4754), .o (n4755) );
  buffer buf_n4756( .i (n4755), .o (n4756) );
  assign n9690 = ~n5190 & n5193 ;
  buffer buf_n9691( .i (n9690), .o (n9691) );
  assign n9692 = n4756 | n9691 ;
  assign n9693 = n4756 & n9691 ;
  assign n9694 = n9692 & ~n9693 ;
  buffer buf_n9695( .i (n9694), .o (n9695) );
  assign n9785 = ~n5656 & n9695 ;
  assign n9786 = n9689 | n9785 ;
  buffer buf_n9787( .i (n9786), .o (n9787) );
  buffer buf_n9788( .i (n9787), .o (n9788) );
  buffer buf_n9789( .i (n9788), .o (n9789) );
  buffer buf_n9790( .i (n9789), .o (n9790) );
  buffer buf_n9791( .i (n9790), .o (n9791) );
  buffer buf_n9792( .i (n9791), .o (n9792) );
  buffer buf_n9793( .i (n9792), .o (n9793) );
  buffer buf_n9794( .i (n9793), .o (n9794) );
  buffer buf_n9795( .i (n9794), .o (n9795) );
  buffer buf_n9796( .i (n9795), .o (n9796) );
  buffer buf_n9797( .i (n9796), .o (n9797) );
  buffer buf_n9798( .i (n9797), .o (n9798) );
  buffer buf_n9799( .i (n9798), .o (n9799) );
  buffer buf_n9800( .i (n9799), .o (n9800) );
  buffer buf_n9801( .i (n9800), .o (n9801) );
  buffer buf_n9802( .i (n9801), .o (n9802) );
  buffer buf_n9803( .i (n9802), .o (n9803) );
  buffer buf_n9804( .i (n9803), .o (n9804) );
  buffer buf_n9805( .i (n9804), .o (n9805) );
  buffer buf_n9806( .i (n9805), .o (n9806) );
  buffer buf_n9807( .i (n9806), .o (n9807) );
  buffer buf_n9808( .i (n9807), .o (n9808) );
  buffer buf_n9809( .i (n9808), .o (n9809) );
  buffer buf_n9810( .i (n9809), .o (n9810) );
  buffer buf_n9811( .i (n9810), .o (n9811) );
  buffer buf_n9812( .i (n9811), .o (n9812) );
  buffer buf_n9813( .i (n9812), .o (n9813) );
  buffer buf_n9814( .i (n9813), .o (n9814) );
  buffer buf_n9815( .i (n9814), .o (n9815) );
  buffer buf_n9816( .i (n9815), .o (n9816) );
  buffer buf_n9817( .i (n9816), .o (n9817) );
  buffer buf_n9818( .i (n9817), .o (n9818) );
  buffer buf_n9819( .i (n9818), .o (n9819) );
  buffer buf_n9820( .i (n9819), .o (n9820) );
  buffer buf_n9821( .i (n9820), .o (n9821) );
  buffer buf_n9822( .i (n9821), .o (n9822) );
  buffer buf_n9823( .i (n9822), .o (n9823) );
  buffer buf_n9824( .i (n9823), .o (n9824) );
  buffer buf_n9825( .i (n9824), .o (n9825) );
  buffer buf_n9826( .i (n9825), .o (n9826) );
  buffer buf_n9827( .i (n9826), .o (n9827) );
  buffer buf_n9828( .i (n9827), .o (n9828) );
  buffer buf_n9829( .i (n9828), .o (n9829) );
  buffer buf_n9830( .i (n9829), .o (n9830) );
  buffer buf_n9831( .i (n9830), .o (n9831) );
  buffer buf_n9832( .i (n9831), .o (n9832) );
  buffer buf_n9833( .i (n9832), .o (n9833) );
  buffer buf_n9834( .i (n9833), .o (n9834) );
  buffer buf_n9835( .i (n9834), .o (n9835) );
  buffer buf_n9836( .i (n9835), .o (n9836) );
  buffer buf_n9837( .i (n9836), .o (n9837) );
  buffer buf_n9838( .i (n9837), .o (n9838) );
  buffer buf_n9839( .i (n9838), .o (n9839) );
  buffer buf_n9840( .i (n9839), .o (n9840) );
  buffer buf_n9841( .i (n9840), .o (n9841) );
  buffer buf_n9842( .i (n9841), .o (n9842) );
  buffer buf_n9843( .i (n9842), .o (n9843) );
  buffer buf_n9844( .i (n9843), .o (n9844) );
  buffer buf_n9845( .i (n9844), .o (n9845) );
  buffer buf_n9846( .i (n9845), .o (n9846) );
  buffer buf_n9847( .i (n9846), .o (n9847) );
  buffer buf_n9848( .i (n9847), .o (n9848) );
  buffer buf_n9849( .i (n9848), .o (n9849) );
  buffer buf_n9850( .i (n9849), .o (n9850) );
  buffer buf_n9851( .i (n9850), .o (n9851) );
  buffer buf_n9852( .i (n9851), .o (n9852) );
  buffer buf_n9853( .i (n9852), .o (n9853) );
  buffer buf_n9854( .i (n9853), .o (n9854) );
  buffer buf_n9855( .i (n9854), .o (n9855) );
  buffer buf_n9856( .i (n9855), .o (n9856) );
  buffer buf_n9857( .i (n9856), .o (n9857) );
  buffer buf_n9858( .i (n9857), .o (n9858) );
  buffer buf_n9859( .i (n9858), .o (n9859) );
  buffer buf_n9860( .i (n9859), .o (n9860) );
  buffer buf_n9861( .i (n9860), .o (n9861) );
  buffer buf_n9862( .i (n9861), .o (n9862) );
  buffer buf_n9863( .i (n9862), .o (n9863) );
  buffer buf_n9864( .i (n9863), .o (n9864) );
  buffer buf_n9865( .i (n9864), .o (n9865) );
  buffer buf_n9866( .i (n9865), .o (n9866) );
  buffer buf_n9867( .i (n9866), .o (n9867) );
  buffer buf_n9868( .i (n9867), .o (n9868) );
  buffer buf_n9869( .i (n9868), .o (n9869) );
  buffer buf_n9870( .i (n9869), .o (n9870) );
  buffer buf_n9871( .i (n9870), .o (n9871) );
  buffer buf_n9872( .i (n9871), .o (n9872) );
  buffer buf_n9873( .i (n9872), .o (n9873) );
  assign n9874 = ~n6644 & n9660 ;
  assign n9875 = n9662 & ~n9874 ;
  assign n9876 = n3146 & n3780 ;
  buffer buf_n9877( .i (n9876), .o (n9877) );
  buffer buf_n9878( .i (n9877), .o (n9878) );
  buffer buf_n9879( .i (n6057), .o (n9879) );
  assign n9880 = ~n9878 & n9879 ;
  buffer buf_n9881( .i (n6088), .o (n9881) );
  assign n9882 = n9880 | n9881 ;
  assign n9883 = n6080 & n9877 ;
  assign n9884 = n3147 & n6067 ;
  assign n9885 = n3782 | n9884 ;
  assign n9886 = ~n9883 & n9885 ;
  assign n9887 = n6059 | n9886 ;
  assign n9888 = ~n9882 & n9887 ;
  buffer buf_n9889( .i (n9888), .o (n9889) );
  buffer buf_n9890( .i (n9889), .o (n9890) );
  assign n9891 = n9449 | n9890 ;
  buffer buf_n9892( .i (n9891), .o (n9892) );
  buffer buf_n9893( .i (n9892), .o (n9893) );
  buffer buf_n9894( .i (n9893), .o (n9894) );
  buffer buf_n9895( .i (n9894), .o (n9895) );
  buffer buf_n9896( .i (n9895), .o (n9896) );
  buffer buf_n9897( .i (n9896), .o (n9897) );
  buffer buf_n9898( .i (n9897), .o (n9898) );
  buffer buf_n9899( .i (n9898), .o (n9899) );
  assign n9900 = n6622 & n8935 ;
  assign n9901 = n9899 | n9900 ;
  assign n9902 = n9875 & n9901 ;
  buffer buf_n9903( .i (n9902), .o (n9903) );
  buffer buf_n9904( .i (n9903), .o (n9904) );
  buffer buf_n9905( .i (n9904), .o (n9905) );
  buffer buf_n9906( .i (n9905), .o (n9906) );
  buffer buf_n9907( .i (n9906), .o (n9907) );
  buffer buf_n9908( .i (n9907), .o (n9908) );
  buffer buf_n9909( .i (n9908), .o (n9909) );
  buffer buf_n9910( .i (n9909), .o (n9910) );
  buffer buf_n9911( .i (n9910), .o (n9911) );
  buffer buf_n9912( .i (n9911), .o (n9912) );
  buffer buf_n9913( .i (n9912), .o (n9913) );
  buffer buf_n9914( .i (n9913), .o (n9914) );
  buffer buf_n9915( .i (n9914), .o (n9915) );
  buffer buf_n9916( .i (n9915), .o (n9916) );
  buffer buf_n9917( .i (n9916), .o (n9917) );
  buffer buf_n9918( .i (n9917), .o (n9918) );
  buffer buf_n9919( .i (n9918), .o (n9919) );
  buffer buf_n9920( .i (n9919), .o (n9920) );
  buffer buf_n9921( .i (n9920), .o (n9921) );
  buffer buf_n9922( .i (n9921), .o (n9922) );
  buffer buf_n9923( .i (n9922), .o (n9923) );
  buffer buf_n9924( .i (n9923), .o (n9924) );
  buffer buf_n9925( .i (n9924), .o (n9925) );
  buffer buf_n9926( .i (n9925), .o (n9926) );
  buffer buf_n9927( .i (n9926), .o (n9927) );
  buffer buf_n9928( .i (n9927), .o (n9928) );
  buffer buf_n9929( .i (n9928), .o (n9929) );
  buffer buf_n9930( .i (n9929), .o (n9930) );
  buffer buf_n9931( .i (n9930), .o (n9931) );
  buffer buf_n9932( .i (n9931), .o (n9932) );
  buffer buf_n9933( .i (n9932), .o (n9933) );
  buffer buf_n9934( .i (n9933), .o (n9934) );
  buffer buf_n9935( .i (n9934), .o (n9935) );
  buffer buf_n9936( .i (n9935), .o (n9936) );
  buffer buf_n9937( .i (n9936), .o (n9937) );
  buffer buf_n9938( .i (n9937), .o (n9938) );
  buffer buf_n9939( .i (n9938), .o (n9939) );
  buffer buf_n9940( .i (n9939), .o (n9940) );
  buffer buf_n9941( .i (n9940), .o (n9941) );
  buffer buf_n9942( .i (n9941), .o (n9942) );
  buffer buf_n9943( .i (n9942), .o (n9943) );
  buffer buf_n9944( .i (n9943), .o (n9944) );
  buffer buf_n9945( .i (n9944), .o (n9945) );
  buffer buf_n9946( .i (n9945), .o (n9946) );
  buffer buf_n9947( .i (n9946), .o (n9947) );
  buffer buf_n9948( .i (n9947), .o (n9948) );
  buffer buf_n9949( .i (n9948), .o (n9949) );
  buffer buf_n9950( .i (n9949), .o (n9950) );
  buffer buf_n9951( .i (n9950), .o (n9951) );
  buffer buf_n9952( .i (n9951), .o (n9952) );
  buffer buf_n9953( .i (n9952), .o (n9953) );
  buffer buf_n9954( .i (n9953), .o (n9954) );
  buffer buf_n9955( .i (n9954), .o (n9955) );
  buffer buf_n9956( .i (n9955), .o (n9956) );
  buffer buf_n9957( .i (n9956), .o (n9957) );
  buffer buf_n9958( .i (n9957), .o (n9958) );
  buffer buf_n9959( .i (n9958), .o (n9959) );
  buffer buf_n9960( .i (n9959), .o (n9960) );
  buffer buf_n9961( .i (n9960), .o (n9961) );
  buffer buf_n9962( .i (n9961), .o (n9962) );
  buffer buf_n9963( .i (n9962), .o (n9963) );
  buffer buf_n9964( .i (n9963), .o (n9964) );
  buffer buf_n9965( .i (n9964), .o (n9965) );
  buffer buf_n9966( .i (n9965), .o (n9966) );
  buffer buf_n9967( .i (n9966), .o (n9967) );
  buffer buf_n9968( .i (n9967), .o (n9968) );
  buffer buf_n9969( .i (n9968), .o (n9969) );
  buffer buf_n9970( .i (n9969), .o (n9970) );
  buffer buf_n9971( .i (n9970), .o (n9971) );
  buffer buf_n9972( .i (n9971), .o (n9972) );
  buffer buf_n9973( .i (n9972), .o (n9973) );
  buffer buf_n9974( .i (n9973), .o (n9974) );
  buffer buf_n9975( .i (n9974), .o (n9975) );
  buffer buf_n9976( .i (n9975), .o (n9976) );
  buffer buf_n9977( .i (n9976), .o (n9977) );
  buffer buf_n7062( .i (n7061), .o (n7062) );
  buffer buf_n7063( .i (n7062), .o (n7063) );
  assign n9978 = n7150 & ~n7153 ;
  buffer buf_n9979( .i (n9978), .o (n9979) );
  assign n9980 = n7063 | n9979 ;
  assign n9981 = n7063 & n9979 ;
  assign n9982 = n9980 & ~n9981 ;
  buffer buf_n9983( .i (n9982), .o (n9983) );
  assign n10023 = ~n5706 & n9983 ;
  assign n10024 = n9977 | n10023 ;
  buffer buf_n10025( .i (n10024), .o (n10025) );
  buffer buf_n10026( .i (n10025), .o (n10026) );
  buffer buf_n10027( .i (n10026), .o (n10027) );
  buffer buf_n10028( .i (n10027), .o (n10028) );
  buffer buf_n10029( .i (n10028), .o (n10029) );
  buffer buf_n10030( .i (n10029), .o (n10030) );
  buffer buf_n10031( .i (n10030), .o (n10031) );
  buffer buf_n10032( .i (n10031), .o (n10032) );
  buffer buf_n10033( .i (n10032), .o (n10033) );
  buffer buf_n10034( .i (n10033), .o (n10034) );
  buffer buf_n10035( .i (n10034), .o (n10035) );
  buffer buf_n10036( .i (n10035), .o (n10036) );
  buffer buf_n10037( .i (n10036), .o (n10037) );
  buffer buf_n10038( .i (n10037), .o (n10038) );
  buffer buf_n10039( .i (n10038), .o (n10039) );
  buffer buf_n10040( .i (n10039), .o (n10040) );
  buffer buf_n10041( .i (n10040), .o (n10041) );
  buffer buf_n10042( .i (n10041), .o (n10042) );
  buffer buf_n10043( .i (n10042), .o (n10043) );
  buffer buf_n10044( .i (n10043), .o (n10044) );
  buffer buf_n10045( .i (n10044), .o (n10045) );
  buffer buf_n10046( .i (n10045), .o (n10046) );
  buffer buf_n10047( .i (n10046), .o (n10047) );
  buffer buf_n10048( .i (n10047), .o (n10048) );
  buffer buf_n10049( .i (n10048), .o (n10049) );
  buffer buf_n10050( .i (n10049), .o (n10050) );
  buffer buf_n10051( .i (n10050), .o (n10051) );
  buffer buf_n10052( .i (n10051), .o (n10052) );
  buffer buf_n10053( .i (n10052), .o (n10053) );
  buffer buf_n10054( .i (n10053), .o (n10054) );
  buffer buf_n10055( .i (n10054), .o (n10055) );
  buffer buf_n10056( .i (n10055), .o (n10056) );
  buffer buf_n10057( .i (n10056), .o (n10057) );
  buffer buf_n10058( .i (n10057), .o (n10058) );
  buffer buf_n10059( .i (n10058), .o (n10059) );
  buffer buf_n10060( .i (n10059), .o (n10060) );
  buffer buf_n10061( .i (n10060), .o (n10061) );
  buffer buf_n4897( .i (n4896), .o (n4897) );
  buffer buf_n4898( .i (n4897), .o (n4898) );
  assign n10062 = ~n4890 & n4901 ;
  buffer buf_n10063( .i (n10062), .o (n10063) );
  assign n10064 = n4898 & ~n10063 ;
  assign n10065 = ~n4898 & n10063 ;
  assign n10066 = n10064 | n10065 ;
  buffer buf_n10067( .i (n10066), .o (n10067) );
  buffer buf_n10068( .i (n10067), .o (n10068) );
  buffer buf_n10069( .i (n10068), .o (n10069) );
  buffer buf_n10070( .i (n10069), .o (n10070) );
  buffer buf_n10071( .i (n10070), .o (n10071) );
  buffer buf_n10072( .i (n10071), .o (n10072) );
  buffer buf_n10073( .i (n10072), .o (n10073) );
  buffer buf_n10074( .i (n10073), .o (n10074) );
  buffer buf_n10075( .i (n10074), .o (n10075) );
  buffer buf_n10076( .i (n10075), .o (n10076) );
  buffer buf_n10077( .i (n10076), .o (n10077) );
  buffer buf_n10078( .i (n10077), .o (n10078) );
  buffer buf_n10079( .i (n10078), .o (n10079) );
  buffer buf_n10080( .i (n10079), .o (n10080) );
  buffer buf_n10081( .i (n10080), .o (n10081) );
  buffer buf_n10082( .i (n10081), .o (n10082) );
  buffer buf_n10083( .i (n10082), .o (n10083) );
  buffer buf_n10084( .i (n10083), .o (n10084) );
  buffer buf_n10085( .i (n10084), .o (n10085) );
  buffer buf_n10086( .i (n10085), .o (n10086) );
  buffer buf_n10087( .i (n10086), .o (n10087) );
  buffer buf_n10088( .i (n10087), .o (n10088) );
  buffer buf_n10089( .i (n10088), .o (n10089) );
  buffer buf_n10090( .i (n10089), .o (n10090) );
  buffer buf_n10091( .i (n10090), .o (n10091) );
  buffer buf_n10092( .i (n10091), .o (n10092) );
  buffer buf_n10093( .i (n10092), .o (n10093) );
  buffer buf_n10094( .i (n10093), .o (n10094) );
  buffer buf_n10095( .i (n10094), .o (n10095) );
  buffer buf_n10096( .i (n10095), .o (n10096) );
  buffer buf_n10097( .i (n10096), .o (n10097) );
  buffer buf_n10098( .i (n10097), .o (n10098) );
  buffer buf_n10099( .i (n10098), .o (n10099) );
  buffer buf_n10100( .i (n10099), .o (n10100) );
  buffer buf_n10101( .i (n10100), .o (n10101) );
  buffer buf_n10102( .i (n10101), .o (n10102) );
  buffer buf_n10103( .i (n10102), .o (n10103) );
  buffer buf_n10104( .i (n10103), .o (n10104) );
  buffer buf_n10105( .i (n10104), .o (n10105) );
  buffer buf_n10106( .i (n10105), .o (n10106) );
  buffer buf_n10107( .i (n10106), .o (n10107) );
  buffer buf_n10108( .i (n10107), .o (n10108) );
  buffer buf_n10109( .i (n10108), .o (n10109) );
  buffer buf_n10110( .i (n10109), .o (n10110) );
  buffer buf_n10111( .i (n10110), .o (n10111) );
  buffer buf_n10112( .i (n10111), .o (n10112) );
  buffer buf_n10113( .i (n10112), .o (n10113) );
  buffer buf_n10114( .i (n10113), .o (n10114) );
  buffer buf_n10115( .i (n10114), .o (n10115) );
  buffer buf_n10116( .i (n10115), .o (n10116) );
  buffer buf_n10117( .i (n10116), .o (n10117) );
  buffer buf_n10118( .i (n10117), .o (n10118) );
  buffer buf_n10119( .i (n10118), .o (n10119) );
  buffer buf_n10120( .i (n10119), .o (n10120) );
  buffer buf_n10121( .i (n10120), .o (n10121) );
  buffer buf_n10122( .i (n10121), .o (n10122) );
  buffer buf_n10123( .i (n10122), .o (n10123) );
  buffer buf_n10124( .i (n10123), .o (n10124) );
  buffer buf_n10125( .i (n10124), .o (n10125) );
  buffer buf_n10126( .i (n10125), .o (n10126) );
  buffer buf_n10127( .i (n10126), .o (n10127) );
  buffer buf_n10128( .i (n10127), .o (n10128) );
  buffer buf_n10129( .i (n10128), .o (n10129) );
  buffer buf_n10130( .i (n10129), .o (n10130) );
  buffer buf_n10131( .i (n10130), .o (n10131) );
  buffer buf_n10132( .i (n10131), .o (n10132) );
  buffer buf_n10133( .i (n10132), .o (n10133) );
  buffer buf_n10134( .i (n10133), .o (n10134) );
  buffer buf_n10135( .i (n10134), .o (n10135) );
  buffer buf_n10136( .i (n10135), .o (n10136) );
  buffer buf_n10137( .i (n10136), .o (n10137) );
  buffer buf_n10138( .i (n10137), .o (n10138) );
  buffer buf_n10139( .i (n10138), .o (n10139) );
  buffer buf_n10140( .i (n10139), .o (n10140) );
  buffer buf_n10141( .i (n10140), .o (n10141) );
  buffer buf_n10142( .i (n10141), .o (n10142) );
  buffer buf_n10143( .i (n10142), .o (n10143) );
  buffer buf_n10144( .i (n10143), .o (n10144) );
  buffer buf_n10145( .i (n10144), .o (n10145) );
  buffer buf_n10146( .i (n10145), .o (n10146) );
  buffer buf_n10147( .i (n10146), .o (n10147) );
  buffer buf_n10148( .i (n10147), .o (n10148) );
  buffer buf_n10149( .i (n10148), .o (n10149) );
  buffer buf_n10150( .i (n10149), .o (n10150) );
  buffer buf_n10151( .i (n10150), .o (n10151) );
  buffer buf_n10152( .i (n10151), .o (n10152) );
  buffer buf_n10153( .i (n10152), .o (n10153) );
  buffer buf_n10154( .i (n10153), .o (n10154) );
  buffer buf_n10155( .i (n10154), .o (n10155) );
  buffer buf_n10156( .i (n10155), .o (n10156) );
  buffer buf_n10157( .i (n10156), .o (n10157) );
  buffer buf_n10158( .i (n10157), .o (n10158) );
  buffer buf_n10159( .i (n10158), .o (n10159) );
  buffer buf_n10160( .i (n10159), .o (n10160) );
  buffer buf_n10161( .i (n10160), .o (n10161) );
  buffer buf_n10162( .i (n10161), .o (n10162) );
  buffer buf_n10163( .i (n10162), .o (n10163) );
  buffer buf_n10164( .i (n10163), .o (n10164) );
  buffer buf_n10165( .i (n10164), .o (n10165) );
  buffer buf_n10166( .i (n10165), .o (n10166) );
  buffer buf_n10167( .i (n10166), .o (n10167) );
  buffer buf_n10168( .i (n10167), .o (n10168) );
  buffer buf_n10169( .i (n10168), .o (n10169) );
  buffer buf_n10170( .i (n10169), .o (n10170) );
  buffer buf_n10171( .i (n10170), .o (n10171) );
  buffer buf_n10172( .i (n10171), .o (n10172) );
  buffer buf_n10173( .i (n10172), .o (n10173) );
  buffer buf_n10174( .i (n10173), .o (n10174) );
  buffer buf_n10175( .i (n10174), .o (n10175) );
  buffer buf_n10176( .i (n10175), .o (n10176) );
  buffer buf_n10177( .i (n10176), .o (n10177) );
  buffer buf_n10178( .i (n10177), .o (n10178) );
  buffer buf_n10179( .i (n10178), .o (n10179) );
  buffer buf_n10180( .i (n10179), .o (n10180) );
  buffer buf_n10181( .i (n10180), .o (n10181) );
  buffer buf_n10182( .i (n10181), .o (n10182) );
  buffer buf_n10183( .i (n10182), .o (n10183) );
  buffer buf_n10184( .i (n10183), .o (n10184) );
  buffer buf_n10185( .i (n10184), .o (n10185) );
  buffer buf_n10186( .i (n10185), .o (n10186) );
  buffer buf_n10187( .i (n10186), .o (n10187) );
  buffer buf_n10188( .i (n10187), .o (n10188) );
  buffer buf_n10189( .i (n10188), .o (n10189) );
  buffer buf_n10190( .i (n10189), .o (n10190) );
  buffer buf_n10191( .i (n10190), .o (n10191) );
  buffer buf_n10192( .i (n10191), .o (n10192) );
  buffer buf_n10193( .i (n10192), .o (n10193) );
  buffer buf_n10194( .i (n10193), .o (n10194) );
  buffer buf_n10195( .i (n10194), .o (n10195) );
  buffer buf_n10196( .i (n10195), .o (n10196) );
  buffer buf_n10197( .i (n10196), .o (n10197) );
  buffer buf_n10198( .i (n10197), .o (n10198) );
  buffer buf_n10199( .i (n10198), .o (n10199) );
  buffer buf_n10200( .i (n10199), .o (n10200) );
  buffer buf_n10201( .i (n10200), .o (n10201) );
  buffer buf_n10202( .i (n10201), .o (n10202) );
  buffer buf_n10203( .i (n10202), .o (n10203) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n10204( .i (n6065), .o (n10204) );
  assign n10205 = n2129 | n10204 ;
  assign n10206 = n363 & n10205 ;
  assign n10207 = n2129 & ~n6055 ;
  buffer buf_n10208( .i (n10207), .o (n10208) );
  assign n10209 = n10206 | n10208 ;
  buffer buf_n10210( .i (n10209), .o (n10210) );
  assign n10211 = n363 & n6079 ;
  assign n10212 = n10208 & n10211 ;
  assign n10213 = n6088 | n10212 ;
  assign n10214 = n10210 & ~n10213 ;
  buffer buf_n10215( .i (n10214), .o (n10215) );
  buffer buf_n10216( .i (n10215), .o (n10216) );
  buffer buf_n10217( .i (n10216), .o (n10217) );
  assign n10218 = n9449 | n10217 ;
  buffer buf_n10219( .i (n10218), .o (n10219) );
  buffer buf_n10220( .i (n10219), .o (n10220) );
  buffer buf_n10221( .i (n10220), .o (n10221) );
  buffer buf_n10222( .i (n10221), .o (n10222) );
  buffer buf_n10223( .i (n10222), .o (n10223) );
  buffer buf_n10224( .i (n10223), .o (n10224) );
  buffer buf_n10225( .i (n10224), .o (n10225) );
  buffer buf_n10226( .i (n10225), .o (n10226) );
  buffer buf_n10227( .i (n3560), .o (n10227) );
  buffer buf_n10228( .i (n10227), .o (n10228) );
  assign n10229 = n6613 & ~n10228 ;
  assign n10230 = n6551 & n10228 ;
  assign n10231 = n10229 | n10230 ;
  buffer buf_n10232( .i (n10231), .o (n10232) );
  assign n10233 = ~n9482 & n10232 ;
  buffer buf_n5937( .i (n5936), .o (n5937) );
  assign n10234 = ~n3909 & n4392 ;
  assign n10235 = n5937 & ~n10234 ;
  assign n10236 = n10228 & ~n10235 ;
  assign n10237 = n6546 | n10228 ;
  assign n10238 = ~n10236 & n10237 ;
  buffer buf_n10239( .i (n10238), .o (n10239) );
  buffer buf_n10240( .i (n1862), .o (n10240) );
  buffer buf_n10241( .i (n10240), .o (n10241) );
  assign n10242 = n10239 & n10241 ;
  assign n10243 = n10233 | n10242 ;
  buffer buf_n10244( .i (n10243), .o (n10244) );
  buffer buf_n10245( .i (n9501), .o (n10245) );
  assign n10246 = n10244 & ~n10245 ;
  assign n10247 = n8681 | n10246 ;
  buffer buf_n10248( .i (n10247), .o (n10248) );
  assign n10249 = n8935 & n10248 ;
  assign n10250 = n10226 | n10249 ;
  assign n10251 = n8892 & ~n9486 ;
  buffer buf_n8671( .i (n8670), .o (n8671) );
  assign n10252 = n8671 & n9486 ;
  assign n10253 = n10251 | n10252 ;
  buffer buf_n10254( .i (n10253), .o (n10254) );
  assign n10255 = n9490 | n10254 ;
  buffer buf_n10256( .i (n10227), .o (n10256) );
  assign n10257 = n8654 & ~n10256 ;
  assign n10258 = n6634 & n10256 ;
  assign n10259 = n10257 | n10258 ;
  buffer buf_n10260( .i (n10259), .o (n10260) );
  buffer buf_n10261( .i (n10260), .o (n10261) );
  buffer buf_n10262( .i (n10241), .o (n10262) );
  assign n10263 = ~n10261 & n10262 ;
  assign n10264 = n10255 & ~n10263 ;
  assign n10265 = ~n10245 & n10264 ;
  assign n10266 = n6628 & ~n10256 ;
  assign n10267 = n5968 | n10266 ;
  buffer buf_n10268( .i (n10267), .o (n10268) );
  assign n10269 = ~n10241 & n10268 ;
  buffer buf_n10270( .i (n6149), .o (n10270) );
  assign n10271 = n10269 | n10270 ;
  buffer buf_n10272( .i (n10271), .o (n10272) );
  assign n10273 = n10245 & n10272 ;
  assign n10274 = n10265 | n10273 ;
  buffer buf_n10275( .i (n10274), .o (n10275) );
  assign n10276 = n9660 & ~n10275 ;
  assign n10277 = n9662 & ~n10276 ;
  assign n10278 = n10250 & n10277 ;
  buffer buf_n10279( .i (n10278), .o (n10279) );
  buffer buf_n10280( .i (n10279), .o (n10280) );
  buffer buf_n10281( .i (n10280), .o (n10281) );
  buffer buf_n10282( .i (n10281), .o (n10282) );
  buffer buf_n10283( .i (n10282), .o (n10283) );
  buffer buf_n10284( .i (n10283), .o (n10284) );
  buffer buf_n10285( .i (n10284), .o (n10285) );
  buffer buf_n10286( .i (n10285), .o (n10286) );
  buffer buf_n10287( .i (n10286), .o (n10287) );
  buffer buf_n10288( .i (n10287), .o (n10288) );
  buffer buf_n10289( .i (n10288), .o (n10289) );
  buffer buf_n10290( .i (n10289), .o (n10290) );
  buffer buf_n10291( .i (n10290), .o (n10291) );
  buffer buf_n10292( .i (n10291), .o (n10292) );
  buffer buf_n5128( .i (n5127), .o (n5128) );
  buffer buf_n5129( .i (n5128), .o (n5129) );
  assign n10293 = ~n5090 & n5132 ;
  buffer buf_n10294( .i (n10293), .o (n10294) );
  assign n10295 = n5129 | n10294 ;
  assign n10296 = n5129 & n10294 ;
  assign n10297 = n10295 & ~n10296 ;
  buffer buf_n10298( .i (n10297), .o (n10298) );
  assign n10399 = ~n5645 & n10298 ;
  assign n10400 = n10292 | n10399 ;
  buffer buf_n10401( .i (n10400), .o (n10401) );
  buffer buf_n10402( .i (n10401), .o (n10402) );
  buffer buf_n10403( .i (n10402), .o (n10403) );
  buffer buf_n10404( .i (n10403), .o (n10404) );
  buffer buf_n10405( .i (n10404), .o (n10405) );
  buffer buf_n10406( .i (n10405), .o (n10406) );
  buffer buf_n10407( .i (n10406), .o (n10407) );
  buffer buf_n10408( .i (n10407), .o (n10408) );
  buffer buf_n10409( .i (n10408), .o (n10409) );
  buffer buf_n10410( .i (n10409), .o (n10410) );
  buffer buf_n10411( .i (n10410), .o (n10411) );
  buffer buf_n10412( .i (n10411), .o (n10412) );
  buffer buf_n10413( .i (n10412), .o (n10413) );
  buffer buf_n10414( .i (n10413), .o (n10414) );
  buffer buf_n10415( .i (n10414), .o (n10415) );
  buffer buf_n10416( .i (n10415), .o (n10416) );
  buffer buf_n10417( .i (n10416), .o (n10417) );
  buffer buf_n10418( .i (n10417), .o (n10418) );
  buffer buf_n10419( .i (n10418), .o (n10419) );
  buffer buf_n10420( .i (n10419), .o (n10420) );
  buffer buf_n10421( .i (n10420), .o (n10421) );
  buffer buf_n10422( .i (n10421), .o (n10422) );
  buffer buf_n10423( .i (n10422), .o (n10423) );
  buffer buf_n10424( .i (n10423), .o (n10424) );
  buffer buf_n10425( .i (n10424), .o (n10425) );
  buffer buf_n10426( .i (n10425), .o (n10426) );
  buffer buf_n10427( .i (n10426), .o (n10427) );
  buffer buf_n10428( .i (n10427), .o (n10428) );
  buffer buf_n10429( .i (n10428), .o (n10429) );
  buffer buf_n10430( .i (n10429), .o (n10430) );
  buffer buf_n10431( .i (n10430), .o (n10431) );
  buffer buf_n10432( .i (n10431), .o (n10432) );
  buffer buf_n10433( .i (n10432), .o (n10433) );
  buffer buf_n10434( .i (n10433), .o (n10434) );
  buffer buf_n10435( .i (n10434), .o (n10435) );
  buffer buf_n10436( .i (n10435), .o (n10436) );
  buffer buf_n10437( .i (n10436), .o (n10437) );
  buffer buf_n10438( .i (n10437), .o (n10438) );
  buffer buf_n10439( .i (n10438), .o (n10439) );
  buffer buf_n10440( .i (n10439), .o (n10440) );
  buffer buf_n10441( .i (n10440), .o (n10441) );
  buffer buf_n10442( .i (n10441), .o (n10442) );
  buffer buf_n10443( .i (n10442), .o (n10443) );
  buffer buf_n10444( .i (n10443), .o (n10444) );
  buffer buf_n10445( .i (n10444), .o (n10445) );
  buffer buf_n10446( .i (n10445), .o (n10446) );
  buffer buf_n10447( .i (n10446), .o (n10447) );
  buffer buf_n10448( .i (n10447), .o (n10448) );
  buffer buf_n10449( .i (n10448), .o (n10449) );
  buffer buf_n10450( .i (n10449), .o (n10450) );
  buffer buf_n10451( .i (n10450), .o (n10451) );
  buffer buf_n10452( .i (n10451), .o (n10452) );
  buffer buf_n10453( .i (n10452), .o (n10453) );
  buffer buf_n10454( .i (n10453), .o (n10454) );
  buffer buf_n10455( .i (n10454), .o (n10455) );
  buffer buf_n10456( .i (n10455), .o (n10456) );
  buffer buf_n10457( .i (n10456), .o (n10457) );
  buffer buf_n10458( .i (n10457), .o (n10458) );
  buffer buf_n10459( .i (n10458), .o (n10459) );
  buffer buf_n10460( .i (n10459), .o (n10460) );
  buffer buf_n10461( .i (n10460), .o (n10461) );
  buffer buf_n10462( .i (n10461), .o (n10462) );
  buffer buf_n10463( .i (n10462), .o (n10463) );
  buffer buf_n10464( .i (n10463), .o (n10464) );
  buffer buf_n10465( .i (n10464), .o (n10465) );
  buffer buf_n10466( .i (n10465), .o (n10466) );
  buffer buf_n10467( .i (n10466), .o (n10467) );
  buffer buf_n10468( .i (n10467), .o (n10468) );
  buffer buf_n10469( .i (n10468), .o (n10469) );
  buffer buf_n10470( .i (n10469), .o (n10470) );
  buffer buf_n10471( .i (n10470), .o (n10471) );
  buffer buf_n10472( .i (n10471), .o (n10472) );
  buffer buf_n10473( .i (n10472), .o (n10473) );
  buffer buf_n10474( .i (n10473), .o (n10474) );
  buffer buf_n10475( .i (n10474), .o (n10475) );
  buffer buf_n10476( .i (n10475), .o (n10476) );
  buffer buf_n10477( .i (n10476), .o (n10477) );
  buffer buf_n10478( .i (n10477), .o (n10478) );
  buffer buf_n10479( .i (n10478), .o (n10479) );
  buffer buf_n10480( .i (n10479), .o (n10480) );
  buffer buf_n10481( .i (n10480), .o (n10481) );
  buffer buf_n10482( .i (n10481), .o (n10482) );
  buffer buf_n10483( .i (n10482), .o (n10483) );
  buffer buf_n10484( .i (n10483), .o (n10484) );
  buffer buf_n10485( .i (n10484), .o (n10485) );
  buffer buf_n10486( .i (n10485), .o (n10486) );
  buffer buf_n10487( .i (n10486), .o (n10487) );
  buffer buf_n10488( .i (n10487), .o (n10488) );
  buffer buf_n10489( .i (n10488), .o (n10489) );
  buffer buf_n10490( .i (n10489), .o (n10490) );
  buffer buf_n10491( .i (n10490), .o (n10491) );
  buffer buf_n10492( .i (n10491), .o (n10492) );
  buffer buf_n10493( .i (n10492), .o (n10493) );
  buffer buf_n10494( .i (n10493), .o (n10494) );
  buffer buf_n10495( .i (n10494), .o (n10495) );
  buffer buf_n10496( .i (n10495), .o (n10496) );
  buffer buf_n10497( .i (n10496), .o (n10497) );
  buffer buf_n10498( .i (n10497), .o (n10498) );
  buffer buf_n5028( .i (n5027), .o (n5028) );
  buffer buf_n5029( .i (n5028), .o (n5029) );
  assign n10499 = n4999 & ~n5031 ;
  buffer buf_n10500( .i (n10499), .o (n10500) );
  assign n10501 = ~n5029 & n10500 ;
  assign n10502 = n5029 & ~n10500 ;
  assign n10503 = n10501 | n10502 ;
  buffer buf_n10504( .i (n10503), .o (n10504) );
  buffer buf_n10505( .i (n10504), .o (n10505) );
  buffer buf_n10506( .i (n10505), .o (n10506) );
  buffer buf_n10507( .i (n10506), .o (n10507) );
  buffer buf_n10508( .i (n10507), .o (n10508) );
  buffer buf_n10509( .i (n10508), .o (n10509) );
  buffer buf_n10510( .i (n10509), .o (n10510) );
  buffer buf_n10511( .i (n10510), .o (n10511) );
  buffer buf_n10512( .i (n10511), .o (n10512) );
  buffer buf_n10513( .i (n10512), .o (n10513) );
  buffer buf_n10514( .i (n10513), .o (n10514) );
  buffer buf_n10515( .i (n10514), .o (n10515) );
  buffer buf_n10516( .i (n10515), .o (n10516) );
  buffer buf_n10517( .i (n10516), .o (n10517) );
  buffer buf_n10518( .i (n10517), .o (n10518) );
  buffer buf_n10519( .i (n10518), .o (n10519) );
  buffer buf_n10520( .i (n10519), .o (n10520) );
  buffer buf_n10521( .i (n10520), .o (n10521) );
  buffer buf_n10522( .i (n10521), .o (n10522) );
  buffer buf_n10523( .i (n10522), .o (n10523) );
  buffer buf_n10524( .i (n10523), .o (n10524) );
  buffer buf_n10525( .i (n10524), .o (n10525) );
  buffer buf_n10526( .i (n10525), .o (n10526) );
  buffer buf_n10527( .i (n10526), .o (n10527) );
  buffer buf_n10528( .i (n10527), .o (n10528) );
  buffer buf_n10529( .i (n10528), .o (n10529) );
  buffer buf_n10530( .i (n10529), .o (n10530) );
  buffer buf_n10531( .i (n10530), .o (n10531) );
  buffer buf_n10532( .i (n10531), .o (n10532) );
  buffer buf_n10533( .i (n10532), .o (n10533) );
  buffer buf_n10534( .i (n10533), .o (n10534) );
  buffer buf_n10535( .i (n10534), .o (n10535) );
  buffer buf_n10536( .i (n10535), .o (n10536) );
  buffer buf_n10537( .i (n10536), .o (n10537) );
  buffer buf_n10538( .i (n10537), .o (n10538) );
  buffer buf_n10539( .i (n10538), .o (n10539) );
  buffer buf_n10540( .i (n10539), .o (n10540) );
  buffer buf_n10541( .i (n10540), .o (n10541) );
  buffer buf_n10542( .i (n10541), .o (n10542) );
  buffer buf_n10543( .i (n10542), .o (n10543) );
  buffer buf_n10544( .i (n10543), .o (n10544) );
  buffer buf_n10545( .i (n10544), .o (n10545) );
  buffer buf_n10546( .i (n10545), .o (n10546) );
  buffer buf_n10547( .i (n10546), .o (n10547) );
  buffer buf_n10548( .i (n10547), .o (n10548) );
  buffer buf_n10549( .i (n10548), .o (n10549) );
  buffer buf_n10550( .i (n10549), .o (n10550) );
  buffer buf_n10551( .i (n10550), .o (n10551) );
  buffer buf_n10552( .i (n10551), .o (n10552) );
  buffer buf_n10553( .i (n10552), .o (n10553) );
  buffer buf_n10554( .i (n10553), .o (n10554) );
  buffer buf_n10555( .i (n10554), .o (n10555) );
  buffer buf_n10556( .i (n10555), .o (n10556) );
  buffer buf_n10557( .i (n10556), .o (n10557) );
  buffer buf_n10558( .i (n10557), .o (n10558) );
  buffer buf_n10559( .i (n10558), .o (n10559) );
  buffer buf_n10560( .i (n10559), .o (n10560) );
  buffer buf_n10561( .i (n10560), .o (n10561) );
  buffer buf_n10562( .i (n10561), .o (n10562) );
  buffer buf_n10563( .i (n10562), .o (n10563) );
  buffer buf_n10564( .i (n10563), .o (n10564) );
  buffer buf_n10565( .i (n10564), .o (n10565) );
  buffer buf_n10566( .i (n10565), .o (n10566) );
  buffer buf_n10567( .i (n10566), .o (n10567) );
  buffer buf_n10568( .i (n10567), .o (n10568) );
  buffer buf_n10569( .i (n10568), .o (n10569) );
  buffer buf_n10570( .i (n10569), .o (n10570) );
  buffer buf_n10571( .i (n10570), .o (n10571) );
  buffer buf_n10572( .i (n10571), .o (n10572) );
  buffer buf_n10573( .i (n10572), .o (n10573) );
  buffer buf_n10574( .i (n10573), .o (n10574) );
  buffer buf_n10575( .i (n10574), .o (n10575) );
  buffer buf_n10576( .i (n10575), .o (n10576) );
  buffer buf_n10577( .i (n10576), .o (n10577) );
  buffer buf_n10578( .i (n10577), .o (n10578) );
  buffer buf_n10579( .i (n10578), .o (n10579) );
  buffer buf_n10580( .i (n10579), .o (n10580) );
  buffer buf_n10581( .i (n10580), .o (n10581) );
  buffer buf_n10582( .i (n10581), .o (n10582) );
  buffer buf_n10583( .i (n10582), .o (n10583) );
  buffer buf_n10584( .i (n10583), .o (n10584) );
  buffer buf_n10585( .i (n10584), .o (n10585) );
  buffer buf_n10586( .i (n10585), .o (n10586) );
  buffer buf_n10587( .i (n10586), .o (n10587) );
  buffer buf_n10588( .i (n10587), .o (n10588) );
  buffer buf_n10589( .i (n10588), .o (n10589) );
  buffer buf_n10590( .i (n10589), .o (n10590) );
  buffer buf_n10591( .i (n10590), .o (n10591) );
  buffer buf_n10592( .i (n10591), .o (n10592) );
  buffer buf_n10593( .i (n10592), .o (n10593) );
  buffer buf_n10594( .i (n10593), .o (n10594) );
  buffer buf_n10595( .i (n10594), .o (n10595) );
  buffer buf_n10596( .i (n10595), .o (n10596) );
  buffer buf_n10597( .i (n10596), .o (n10597) );
  buffer buf_n10598( .i (n10597), .o (n10598) );
  buffer buf_n10599( .i (n10598), .o (n10599) );
  buffer buf_n10600( .i (n10599), .o (n10600) );
  buffer buf_n10601( .i (n10600), .o (n10601) );
  buffer buf_n10602( .i (n10601), .o (n10602) );
  buffer buf_n10603( .i (n10602), .o (n10603) );
  buffer buf_n10604( .i (n10603), .o (n10604) );
  buffer buf_n10605( .i (n10604), .o (n10605) );
  buffer buf_n10606( .i (n10605), .o (n10606) );
  buffer buf_n10607( .i (n10606), .o (n10607) );
  buffer buf_n10608( .i (n10607), .o (n10608) );
  buffer buf_n10609( .i (n10608), .o (n10609) );
  buffer buf_n10610( .i (n10609), .o (n10610) );
  buffer buf_n10611( .i (n10610), .o (n10611) );
  buffer buf_n10612( .i (n10611), .o (n10612) );
  buffer buf_n10613( .i (n10612), .o (n10613) );
  buffer buf_n10614( .i (n10613), .o (n10614) );
  buffer buf_n10615( .i (n10614), .o (n10615) );
  buffer buf_n10616( .i (n10615), .o (n10616) );
  buffer buf_n10617( .i (n10616), .o (n10617) );
  buffer buf_n10618( .i (n10617), .o (n10618) );
  buffer buf_n10619( .i (n10618), .o (n10619) );
  buffer buf_n10620( .i (n10619), .o (n10620) );
  assign n10621 = ~n7545 & n7642 ;
  buffer buf_n7639( .i (n7638), .o (n7639) );
  buffer buf_n7640( .i (n7639), .o (n7640) );
  buffer buf_n7548( .i (n7547), .o (n7548) );
  assign n10622 = ~n7544 & n7548 ;
  assign n10623 = n7640 | n10622 ;
  assign n10624 = ~n10621 & n10623 ;
  buffer buf_n10625( .i (n10624), .o (n10625) );
  buffer buf_n10626( .i (n10625), .o (n10626) );
  buffer buf_n10627( .i (n10626), .o (n10627) );
  buffer buf_n10628( .i (n10627), .o (n10628) );
  buffer buf_n10629( .i (n10628), .o (n10629) );
  buffer buf_n10630( .i (n10629), .o (n10630) );
  buffer buf_n10631( .i (n10630), .o (n10631) );
  buffer buf_n10632( .i (n10631), .o (n10632) );
  buffer buf_n10299( .i (n10298), .o (n10299) );
  buffer buf_n10300( .i (n10299), .o (n10300) );
  buffer buf_n10301( .i (n10300), .o (n10301) );
  buffer buf_n10302( .i (n10301), .o (n10302) );
  buffer buf_n10303( .i (n10302), .o (n10303) );
  buffer buf_n10304( .i (n10303), .o (n10304) );
  buffer buf_n10305( .i (n10304), .o (n10305) );
  buffer buf_n10306( .i (n10305), .o (n10306) );
  buffer buf_n10307( .i (n10306), .o (n10307) );
  buffer buf_n10308( .i (n10307), .o (n10308) );
  buffer buf_n10309( .i (n10308), .o (n10309) );
  buffer buf_n10310( .i (n10309), .o (n10310) );
  buffer buf_n10311( .i (n10310), .o (n10311) );
  buffer buf_n10312( .i (n10311), .o (n10312) );
  buffer buf_n10313( .i (n10312), .o (n10313) );
  buffer buf_n10314( .i (n10313), .o (n10314) );
  buffer buf_n10315( .i (n10314), .o (n10315) );
  buffer buf_n10316( .i (n10315), .o (n10316) );
  buffer buf_n10317( .i (n10316), .o (n10317) );
  buffer buf_n10318( .i (n10317), .o (n10318) );
  buffer buf_n10319( .i (n10318), .o (n10319) );
  buffer buf_n10320( .i (n10319), .o (n10320) );
  buffer buf_n10321( .i (n10320), .o (n10321) );
  buffer buf_n10322( .i (n10321), .o (n10322) );
  buffer buf_n10323( .i (n10322), .o (n10323) );
  buffer buf_n10324( .i (n10323), .o (n10324) );
  buffer buf_n10325( .i (n10324), .o (n10325) );
  buffer buf_n10326( .i (n10325), .o (n10326) );
  buffer buf_n10327( .i (n10326), .o (n10327) );
  buffer buf_n10328( .i (n10327), .o (n10328) );
  buffer buf_n10329( .i (n10328), .o (n10329) );
  buffer buf_n10330( .i (n10329), .o (n10330) );
  buffer buf_n10331( .i (n10330), .o (n10331) );
  buffer buf_n10332( .i (n10331), .o (n10332) );
  buffer buf_n10333( .i (n10332), .o (n10333) );
  buffer buf_n10334( .i (n10333), .o (n10334) );
  buffer buf_n10335( .i (n10334), .o (n10335) );
  buffer buf_n10336( .i (n10335), .o (n10336) );
  buffer buf_n10337( .i (n10336), .o (n10337) );
  buffer buf_n10338( .i (n10337), .o (n10338) );
  buffer buf_n10339( .i (n10338), .o (n10339) );
  buffer buf_n10340( .i (n10339), .o (n10340) );
  buffer buf_n10341( .i (n10340), .o (n10341) );
  buffer buf_n10342( .i (n10341), .o (n10342) );
  buffer buf_n10343( .i (n10342), .o (n10343) );
  buffer buf_n10344( .i (n10343), .o (n10344) );
  buffer buf_n10345( .i (n10344), .o (n10345) );
  buffer buf_n10346( .i (n10345), .o (n10346) );
  buffer buf_n10347( .i (n10346), .o (n10347) );
  buffer buf_n10348( .i (n10347), .o (n10348) );
  buffer buf_n10349( .i (n10348), .o (n10349) );
  buffer buf_n10350( .i (n10349), .o (n10350) );
  buffer buf_n10351( .i (n10350), .o (n10351) );
  buffer buf_n10352( .i (n10351), .o (n10352) );
  buffer buf_n10353( .i (n10352), .o (n10353) );
  buffer buf_n10354( .i (n10353), .o (n10354) );
  buffer buf_n10355( .i (n10354), .o (n10355) );
  buffer buf_n10356( .i (n10355), .o (n10356) );
  buffer buf_n10357( .i (n10356), .o (n10357) );
  buffer buf_n10358( .i (n10357), .o (n10358) );
  buffer buf_n10359( .i (n10358), .o (n10359) );
  buffer buf_n10360( .i (n10359), .o (n10360) );
  buffer buf_n10361( .i (n10360), .o (n10361) );
  buffer buf_n10362( .i (n10361), .o (n10362) );
  buffer buf_n10363( .i (n10362), .o (n10363) );
  buffer buf_n10364( .i (n10363), .o (n10364) );
  buffer buf_n10365( .i (n10364), .o (n10365) );
  buffer buf_n10366( .i (n10365), .o (n10366) );
  buffer buf_n10367( .i (n10366), .o (n10367) );
  buffer buf_n10368( .i (n10367), .o (n10368) );
  buffer buf_n10369( .i (n10368), .o (n10369) );
  buffer buf_n10370( .i (n10369), .o (n10370) );
  buffer buf_n10371( .i (n10370), .o (n10371) );
  buffer buf_n10372( .i (n10371), .o (n10372) );
  buffer buf_n10373( .i (n10372), .o (n10373) );
  buffer buf_n10374( .i (n10373), .o (n10374) );
  buffer buf_n10375( .i (n10374), .o (n10375) );
  buffer buf_n10376( .i (n10375), .o (n10376) );
  buffer buf_n10377( .i (n10376), .o (n10377) );
  buffer buf_n10378( .i (n10377), .o (n10378) );
  buffer buf_n10379( .i (n10378), .o (n10379) );
  buffer buf_n10380( .i (n10379), .o (n10380) );
  buffer buf_n10381( .i (n10380), .o (n10381) );
  buffer buf_n10382( .i (n10381), .o (n10382) );
  buffer buf_n10383( .i (n10382), .o (n10383) );
  buffer buf_n10384( .i (n10383), .o (n10384) );
  buffer buf_n10385( .i (n10384), .o (n10385) );
  buffer buf_n10386( .i (n10385), .o (n10386) );
  buffer buf_n10387( .i (n10386), .o (n10387) );
  buffer buf_n10388( .i (n10387), .o (n10388) );
  buffer buf_n10389( .i (n10388), .o (n10389) );
  buffer buf_n10390( .i (n10389), .o (n10390) );
  buffer buf_n10391( .i (n10390), .o (n10391) );
  buffer buf_n10392( .i (n10391), .o (n10392) );
  buffer buf_n10393( .i (n10392), .o (n10393) );
  buffer buf_n10394( .i (n10393), .o (n10394) );
  buffer buf_n10395( .i (n10394), .o (n10395) );
  buffer buf_n10396( .i (n10395), .o (n10396) );
  buffer buf_n10397( .i (n10396), .o (n10397) );
  buffer buf_n10398( .i (n10397), .o (n10398) );
  buffer buf_n5180( .i (n5179), .o (n5180) );
  buffer buf_n5181( .i (n5180), .o (n5181) );
  buffer buf_n5184( .i (n5183), .o (n5184) );
  assign n10633 = n5138 & ~n5184 ;
  assign n10634 = n5181 & ~n10633 ;
  assign n10635 = n5139 & ~n5186 ;
  assign n10636 = n10634 | n10635 ;
  buffer buf_n10637( .i (n10636), .o (n10637) );
  buffer buf_n10638( .i (n10637), .o (n10638) );
  buffer buf_n10639( .i (n10638), .o (n10639) );
  buffer buf_n10640( .i (n10639), .o (n10640) );
  buffer buf_n10641( .i (n10640), .o (n10641) );
  buffer buf_n10642( .i (n10641), .o (n10642) );
  buffer buf_n10643( .i (n10642), .o (n10643) );
  buffer buf_n10644( .i (n10643), .o (n10644) );
  buffer buf_n10645( .i (n10644), .o (n10645) );
  buffer buf_n10646( .i (n10645), .o (n10646) );
  buffer buf_n10647( .i (n10646), .o (n10647) );
  buffer buf_n10648( .i (n10647), .o (n10648) );
  buffer buf_n10649( .i (n10648), .o (n10649) );
  buffer buf_n10650( .i (n10649), .o (n10650) );
  buffer buf_n10651( .i (n10650), .o (n10651) );
  buffer buf_n10652( .i (n10651), .o (n10652) );
  buffer buf_n10653( .i (n10652), .o (n10653) );
  buffer buf_n10654( .i (n10653), .o (n10654) );
  buffer buf_n10655( .i (n10654), .o (n10655) );
  buffer buf_n10656( .i (n10655), .o (n10656) );
  buffer buf_n10657( .i (n10656), .o (n10657) );
  buffer buf_n10658( .i (n10657), .o (n10658) );
  buffer buf_n10659( .i (n10658), .o (n10659) );
  buffer buf_n10660( .i (n10659), .o (n10660) );
  buffer buf_n10661( .i (n10660), .o (n10661) );
  buffer buf_n10662( .i (n10661), .o (n10662) );
  buffer buf_n10663( .i (n10662), .o (n10663) );
  buffer buf_n10664( .i (n10663), .o (n10664) );
  buffer buf_n10665( .i (n10664), .o (n10665) );
  buffer buf_n10666( .i (n10665), .o (n10666) );
  buffer buf_n10667( .i (n10666), .o (n10667) );
  buffer buf_n10668( .i (n10667), .o (n10668) );
  buffer buf_n10669( .i (n10668), .o (n10669) );
  buffer buf_n10670( .i (n10669), .o (n10670) );
  buffer buf_n10671( .i (n10670), .o (n10671) );
  buffer buf_n10672( .i (n10671), .o (n10672) );
  buffer buf_n10673( .i (n10672), .o (n10673) );
  buffer buf_n10674( .i (n10673), .o (n10674) );
  buffer buf_n10675( .i (n10674), .o (n10675) );
  buffer buf_n10676( .i (n10675), .o (n10676) );
  buffer buf_n10677( .i (n10676), .o (n10677) );
  buffer buf_n10678( .i (n10677), .o (n10678) );
  buffer buf_n10679( .i (n10678), .o (n10679) );
  buffer buf_n10680( .i (n10679), .o (n10680) );
  buffer buf_n10681( .i (n10680), .o (n10681) );
  buffer buf_n10682( .i (n10681), .o (n10682) );
  buffer buf_n10683( .i (n10682), .o (n10683) );
  buffer buf_n10684( .i (n10683), .o (n10684) );
  buffer buf_n10685( .i (n10684), .o (n10685) );
  buffer buf_n10686( .i (n10685), .o (n10686) );
  buffer buf_n10687( .i (n10686), .o (n10687) );
  buffer buf_n10688( .i (n10687), .o (n10688) );
  buffer buf_n10689( .i (n10688), .o (n10689) );
  buffer buf_n10690( .i (n10689), .o (n10690) );
  buffer buf_n10691( .i (n10690), .o (n10691) );
  buffer buf_n10692( .i (n10691), .o (n10692) );
  buffer buf_n10693( .i (n10692), .o (n10693) );
  buffer buf_n10694( .i (n10693), .o (n10694) );
  buffer buf_n10695( .i (n10694), .o (n10695) );
  buffer buf_n10696( .i (n10695), .o (n10696) );
  buffer buf_n10697( .i (n10696), .o (n10697) );
  buffer buf_n10698( .i (n10697), .o (n10698) );
  buffer buf_n10699( .i (n10698), .o (n10699) );
  buffer buf_n10700( .i (n10699), .o (n10700) );
  buffer buf_n10701( .i (n10700), .o (n10701) );
  buffer buf_n10702( .i (n10701), .o (n10702) );
  buffer buf_n10703( .i (n10702), .o (n10703) );
  buffer buf_n10704( .i (n10703), .o (n10704) );
  buffer buf_n10705( .i (n10704), .o (n10705) );
  buffer buf_n10706( .i (n10705), .o (n10706) );
  buffer buf_n10707( .i (n10706), .o (n10707) );
  buffer buf_n10708( .i (n10707), .o (n10708) );
  buffer buf_n10709( .i (n10708), .o (n10709) );
  buffer buf_n10710( .i (n10709), .o (n10710) );
  buffer buf_n10711( .i (n10710), .o (n10711) );
  buffer buf_n10712( .i (n10711), .o (n10712) );
  buffer buf_n10713( .i (n10712), .o (n10713) );
  buffer buf_n10714( .i (n10713), .o (n10714) );
  buffer buf_n10715( .i (n10714), .o (n10715) );
  buffer buf_n10716( .i (n10715), .o (n10716) );
  buffer buf_n10717( .i (n10716), .o (n10717) );
  buffer buf_n10718( .i (n10717), .o (n10718) );
  buffer buf_n10719( .i (n10718), .o (n10719) );
  buffer buf_n10720( .i (n10719), .o (n10720) );
  buffer buf_n10721( .i (n10720), .o (n10721) );
  buffer buf_n10722( .i (n10721), .o (n10722) );
  buffer buf_n10723( .i (n10722), .o (n10723) );
  buffer buf_n10724( .i (n10723), .o (n10724) );
  buffer buf_n10725( .i (n10724), .o (n10725) );
  buffer buf_n10726( .i (n10725), .o (n10726) );
  buffer buf_n10727( .i (n10726), .o (n10727) );
  buffer buf_n10728( .i (n10727), .o (n10728) );
  buffer buf_n10729( .i (n10728), .o (n10729) );
  buffer buf_n10730( .i (n10729), .o (n10730) );
  buffer buf_n10731( .i (n10730), .o (n10731) );
  buffer buf_n10732( .i (n10731), .o (n10732) );
  assign n10733 = ~n9468 & n10262 ;
  buffer buf_n6262( .i (n6261), .o (n6262) );
  assign n10734 = n6262 & n9486 ;
  buffer buf_n10735( .i (n10256), .o (n10735) );
  assign n10736 = n6221 & ~n10735 ;
  assign n10737 = n10734 | n10736 ;
  buffer buf_n10738( .i (n10737), .o (n10738) );
  assign n10739 = n10262 | n10738 ;
  assign n10740 = ~n10733 & n10739 ;
  assign n10741 = ~n10245 & n10740 ;
  buffer buf_n10742( .i (n10741), .o (n10742) );
  assign n10743 = n9463 & ~n10262 ;
  assign n10744 = n6151 | n10743 ;
  buffer buf_n10745( .i (n10744), .o (n10745) );
  assign n10746 = n9622 & n10745 ;
  assign n10747 = n10742 | n10746 ;
  buffer buf_n10748( .i (n10747), .o (n10748) );
  assign n10749 = n5928 & ~n10748 ;
  assign n10750 = n5885 & ~n10749 ;
  assign n10751 = n9481 & ~n10241 ;
  buffer buf_n10752( .i (n10240), .o (n10752) );
  assign n10753 = n9497 & n10752 ;
  assign n10754 = n10751 | n10753 ;
  buffer buf_n10755( .i (n10754), .o (n10755) );
  buffer buf_n10756( .i (n9501), .o (n10756) );
  assign n10757 = n10755 & ~n10756 ;
  assign n10758 = n8681 | n10757 ;
  buffer buf_n10759( .i (n10758), .o (n10759) );
  buffer buf_n10761( .i (n6100), .o (n10761) );
  assign n10762 = n10759 & n10761 ;
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2089( .i (n2088), .o (n2089) );
  buffer buf_n2090( .i (n2089), .o (n2090) );
  buffer buf_n2091( .i (n2090), .o (n2091) );
  assign n10763 = n2091 & n6079 ;
  assign n10764 = n1903 & ~n6055 ;
  buffer buf_n10765( .i (n10764), .o (n10765) );
  assign n10766 = n10763 & n10765 ;
  buffer buf_n10767( .i (n6087), .o (n10767) );
  assign n10768 = n10766 | n10767 ;
  assign n10769 = n1903 | n10204 ;
  assign n10770 = n2091 & n10769 ;
  assign n10771 = n10765 | n10770 ;
  buffer buf_n10772( .i (n10771), .o (n10772) );
  assign n10773 = ~n10768 & n10772 ;
  buffer buf_n10774( .i (n10773), .o (n10774) );
  buffer buf_n10775( .i (n10774), .o (n10775) );
  buffer buf_n10776( .i (n10775), .o (n10776) );
  buffer buf_n10777( .i (n5918), .o (n10777) );
  assign n10778 = n10776 | n10777 ;
  buffer buf_n10779( .i (n10778), .o (n10779) );
  buffer buf_n10780( .i (n10779), .o (n10780) );
  buffer buf_n10781( .i (n10780), .o (n10781) );
  buffer buf_n10782( .i (n10781), .o (n10782) );
  buffer buf_n10783( .i (n10782), .o (n10783) );
  buffer buf_n10784( .i (n10783), .o (n10784) );
  buffer buf_n10785( .i (n10784), .o (n10785) );
  buffer buf_n10786( .i (n10785), .o (n10786) );
  assign n10787 = n10762 | n10786 ;
  buffer buf_n10788( .i (n10787), .o (n10788) );
  assign n10789 = n10750 & n10788 ;
  buffer buf_n10790( .i (n10789), .o (n10790) );
  buffer buf_n10791( .i (n10790), .o (n10791) );
  buffer buf_n10792( .i (n10791), .o (n10792) );
  buffer buf_n10793( .i (n10792), .o (n10793) );
  buffer buf_n10794( .i (n10793), .o (n10794) );
  buffer buf_n10795( .i (n10794), .o (n10795) );
  buffer buf_n10796( .i (n10795), .o (n10796) );
  buffer buf_n10797( .i (n10796), .o (n10797) );
  buffer buf_n10798( .i (n10797), .o (n10798) );
  buffer buf_n10799( .i (n10798), .o (n10799) );
  buffer buf_n10800( .i (n10799), .o (n10800) );
  buffer buf_n10801( .i (n10800), .o (n10801) );
  buffer buf_n10802( .i (n10801), .o (n10802) );
  buffer buf_n10803( .i (n10802), .o (n10803) );
  buffer buf_n10804( .i (n10803), .o (n10804) );
  buffer buf_n10805( .i (n10804), .o (n10805) );
  buffer buf_n10806( .i (n10805), .o (n10806) );
  buffer buf_n10807( .i (n10806), .o (n10807) );
  assign n10808 = ~n5650 & n10637 ;
  assign n10809 = n10807 | n10808 ;
  buffer buf_n10810( .i (n10809), .o (n10810) );
  buffer buf_n10811( .i (n10810), .o (n10811) );
  buffer buf_n10812( .i (n10811), .o (n10812) );
  buffer buf_n10813( .i (n10812), .o (n10813) );
  buffer buf_n10814( .i (n10813), .o (n10814) );
  buffer buf_n10815( .i (n10814), .o (n10815) );
  buffer buf_n10816( .i (n10815), .o (n10816) );
  buffer buf_n10817( .i (n10816), .o (n10817) );
  buffer buf_n10818( .i (n10817), .o (n10818) );
  buffer buf_n10819( .i (n10818), .o (n10819) );
  buffer buf_n10820( .i (n10819), .o (n10820) );
  buffer buf_n10821( .i (n10820), .o (n10821) );
  buffer buf_n10822( .i (n10821), .o (n10822) );
  buffer buf_n10823( .i (n10822), .o (n10823) );
  buffer buf_n10824( .i (n10823), .o (n10824) );
  buffer buf_n10825( .i (n10824), .o (n10825) );
  buffer buf_n10826( .i (n10825), .o (n10826) );
  buffer buf_n10827( .i (n10826), .o (n10827) );
  buffer buf_n10828( .i (n10827), .o (n10828) );
  buffer buf_n10829( .i (n10828), .o (n10829) );
  buffer buf_n10830( .i (n10829), .o (n10830) );
  buffer buf_n10831( .i (n10830), .o (n10831) );
  buffer buf_n10832( .i (n10831), .o (n10832) );
  buffer buf_n10833( .i (n10832), .o (n10833) );
  buffer buf_n10834( .i (n10833), .o (n10834) );
  buffer buf_n10835( .i (n10834), .o (n10835) );
  buffer buf_n10836( .i (n10835), .o (n10836) );
  buffer buf_n10837( .i (n10836), .o (n10837) );
  buffer buf_n10838( .i (n10837), .o (n10838) );
  buffer buf_n10839( .i (n10838), .o (n10839) );
  buffer buf_n10840( .i (n10839), .o (n10840) );
  buffer buf_n10841( .i (n10840), .o (n10841) );
  buffer buf_n10842( .i (n10841), .o (n10842) );
  buffer buf_n10843( .i (n10842), .o (n10843) );
  buffer buf_n10844( .i (n10843), .o (n10844) );
  buffer buf_n10845( .i (n10844), .o (n10845) );
  buffer buf_n10846( .i (n10845), .o (n10846) );
  buffer buf_n10847( .i (n10846), .o (n10847) );
  buffer buf_n10848( .i (n10847), .o (n10848) );
  buffer buf_n10849( .i (n10848), .o (n10849) );
  buffer buf_n10850( .i (n10849), .o (n10850) );
  buffer buf_n10851( .i (n10850), .o (n10851) );
  buffer buf_n10852( .i (n10851), .o (n10852) );
  buffer buf_n10853( .i (n10852), .o (n10853) );
  buffer buf_n10854( .i (n10853), .o (n10854) );
  buffer buf_n10855( .i (n10854), .o (n10855) );
  buffer buf_n10856( .i (n10855), .o (n10856) );
  buffer buf_n10857( .i (n10856), .o (n10857) );
  buffer buf_n10858( .i (n10857), .o (n10858) );
  buffer buf_n10859( .i (n10858), .o (n10859) );
  buffer buf_n10860( .i (n10859), .o (n10860) );
  buffer buf_n10861( .i (n10860), .o (n10861) );
  buffer buf_n10862( .i (n10861), .o (n10862) );
  buffer buf_n10863( .i (n10862), .o (n10863) );
  buffer buf_n10864( .i (n10863), .o (n10864) );
  buffer buf_n10865( .i (n10864), .o (n10865) );
  buffer buf_n10866( .i (n10865), .o (n10866) );
  buffer buf_n10867( .i (n10866), .o (n10867) );
  buffer buf_n10868( .i (n10867), .o (n10868) );
  buffer buf_n10869( .i (n10868), .o (n10869) );
  buffer buf_n10870( .i (n10869), .o (n10870) );
  buffer buf_n10871( .i (n10870), .o (n10871) );
  buffer buf_n10872( .i (n10871), .o (n10872) );
  buffer buf_n10873( .i (n10872), .o (n10873) );
  buffer buf_n10874( .i (n10873), .o (n10874) );
  buffer buf_n10875( .i (n10874), .o (n10875) );
  buffer buf_n10876( .i (n10875), .o (n10876) );
  buffer buf_n10877( .i (n10876), .o (n10877) );
  buffer buf_n10878( .i (n10877), .o (n10878) );
  buffer buf_n10879( .i (n10878), .o (n10879) );
  buffer buf_n10880( .i (n10879), .o (n10880) );
  buffer buf_n10881( .i (n10880), .o (n10881) );
  buffer buf_n10882( .i (n10881), .o (n10882) );
  buffer buf_n10883( .i (n10882), .o (n10883) );
  buffer buf_n10884( .i (n10883), .o (n10884) );
  buffer buf_n10885( .i (n10884), .o (n10885) );
  buffer buf_n10886( .i (n10885), .o (n10886) );
  buffer buf_n10887( .i (n10886), .o (n10887) );
  buffer buf_n10888( .i (n10887), .o (n10888) );
  buffer buf_n10889( .i (n10888), .o (n10889) );
  buffer buf_n10890( .i (n10889), .o (n10890) );
  buffer buf_n10891( .i (n10890), .o (n10891) );
  buffer buf_n10892( .i (n10891), .o (n10892) );
  buffer buf_n10893( .i (n10892), .o (n10893) );
  buffer buf_n10894( .i (n10893), .o (n10894) );
  buffer buf_n10895( .i (n10894), .o (n10895) );
  buffer buf_n10896( .i (n10895), .o (n10896) );
  buffer buf_n10897( .i (n10896), .o (n10897) );
  buffer buf_n10898( .i (n10897), .o (n10898) );
  buffer buf_n10899( .i (n10898), .o (n10899) );
  buffer buf_n10900( .i (n10899), .o (n10900) );
  buffer buf_n10901( .i (n10900), .o (n10901) );
  buffer buf_n10902( .i (n10901), .o (n10902) );
  buffer buf_n10903( .i (n9660), .o (n10903) );
  assign n10904 = ~n9474 & n10903 ;
  buffer buf_n10905( .i (n9662), .o (n10905) );
  assign n10906 = ~n10904 & n10905 ;
  assign n10907 = n9505 & n10761 ;
  buffer buf_n10908( .i (n10204), .o (n10908) );
  assign n10909 = n402 & n10908 ;
  assign n10910 = n1521 | n10909 ;
  assign n10911 = n401 & n1519 ;
  buffer buf_n10912( .i (n10911), .o (n10912) );
  buffer buf_n10914( .i (n6077), .o (n10914) );
  buffer buf_n10915( .i (n10914), .o (n10915) );
  buffer buf_n10916( .i (n10915), .o (n10916) );
  assign n10917 = n10912 & n10916 ;
  assign n10918 = n10910 & ~n10917 ;
  assign n10919 = n6059 | n10918 ;
  buffer buf_n10913( .i (n10912), .o (n10913) );
  assign n10920 = n9879 & ~n10913 ;
  assign n10921 = n9881 | n10920 ;
  assign n10922 = n10919 & ~n10921 ;
  buffer buf_n10923( .i (n10922), .o (n10923) );
  buffer buf_n10924( .i (n10923), .o (n10924) );
  assign n10925 = n10777 | n10924 ;
  buffer buf_n10926( .i (n10925), .o (n10926) );
  buffer buf_n10927( .i (n10926), .o (n10927) );
  buffer buf_n10928( .i (n10927), .o (n10928) );
  buffer buf_n10929( .i (n10928), .o (n10929) );
  buffer buf_n10930( .i (n10929), .o (n10930) );
  buffer buf_n10931( .i (n10930), .o (n10931) );
  buffer buf_n10932( .i (n10931), .o (n10932) );
  buffer buf_n10933( .i (n10932), .o (n10933) );
  assign n10934 = n10907 | n10933 ;
  buffer buf_n10935( .i (n10934), .o (n10935) );
  assign n10936 = n10906 & n10935 ;
  buffer buf_n10937( .i (n10936), .o (n10937) );
  buffer buf_n10938( .i (n10937), .o (n10938) );
  buffer buf_n10939( .i (n10938), .o (n10939) );
  buffer buf_n10940( .i (n10939), .o (n10940) );
  buffer buf_n10941( .i (n10940), .o (n10941) );
  buffer buf_n10942( .i (n10941), .o (n10942) );
  buffer buf_n10943( .i (n10942), .o (n10943) );
  buffer buf_n10944( .i (n10943), .o (n10944) );
  buffer buf_n10945( .i (n10944), .o (n10945) );
  buffer buf_n10946( .i (n10945), .o (n10946) );
  buffer buf_n10947( .i (n10946), .o (n10947) );
  buffer buf_n10948( .i (n10947), .o (n10948) );
  buffer buf_n10949( .i (n10948), .o (n10949) );
  buffer buf_n10950( .i (n10949), .o (n10950) );
  buffer buf_n10951( .i (n10950), .o (n10951) );
  buffer buf_n10952( .i (n10951), .o (n10952) );
  buffer buf_n10953( .i (n10952), .o (n10953) );
  buffer buf_n10954( .i (n10953), .o (n10954) );
  buffer buf_n10955( .i (n10954), .o (n10955) );
  buffer buf_n10956( .i (n10955), .o (n10956) );
  buffer buf_n10957( .i (n10956), .o (n10957) );
  buffer buf_n10958( .i (n10957), .o (n10958) );
  buffer buf_n10959( .i (n10958), .o (n10959) );
  buffer buf_n10960( .i (n10959), .o (n10960) );
  buffer buf_n10961( .i (n10960), .o (n10961) );
  buffer buf_n10962( .i (n10961), .o (n10962) );
  buffer buf_n10963( .i (n10962), .o (n10963) );
  buffer buf_n10964( .i (n10963), .o (n10964) );
  buffer buf_n10965( .i (n10964), .o (n10965) );
  buffer buf_n10966( .i (n10965), .o (n10966) );
  buffer buf_n10967( .i (n10966), .o (n10967) );
  buffer buf_n10968( .i (n10967), .o (n10968) );
  buffer buf_n10969( .i (n10968), .o (n10969) );
  buffer buf_n10970( .i (n10969), .o (n10970) );
  buffer buf_n10971( .i (n10970), .o (n10971) );
  buffer buf_n10972( .i (n10971), .o (n10972) );
  buffer buf_n10973( .i (n10972), .o (n10973) );
  buffer buf_n10974( .i (n10973), .o (n10974) );
  buffer buf_n10975( .i (n10974), .o (n10975) );
  buffer buf_n10976( .i (n10975), .o (n10976) );
  buffer buf_n10977( .i (n10976), .o (n10977) );
  buffer buf_n10978( .i (n10977), .o (n10978) );
  buffer buf_n10979( .i (n10978), .o (n10979) );
  buffer buf_n10980( .i (n10979), .o (n10980) );
  buffer buf_n10981( .i (n10980), .o (n10981) );
  buffer buf_n10982( .i (n10981), .o (n10982) );
  buffer buf_n10983( .i (n10982), .o (n10983) );
  buffer buf_n10984( .i (n10983), .o (n10984) );
  buffer buf_n10985( .i (n10984), .o (n10985) );
  buffer buf_n10986( .i (n10985), .o (n10986) );
  buffer buf_n10987( .i (n10986), .o (n10987) );
  buffer buf_n10988( .i (n10987), .o (n10988) );
  buffer buf_n10989( .i (n10988), .o (n10989) );
  buffer buf_n10990( .i (n10989), .o (n10990) );
  buffer buf_n10991( .i (n10990), .o (n10991) );
  buffer buf_n10992( .i (n10991), .o (n10992) );
  buffer buf_n10993( .i (n10992), .o (n10993) );
  buffer buf_n10994( .i (n10993), .o (n10994) );
  buffer buf_n10995( .i (n10994), .o (n10995) );
  buffer buf_n4582( .i (n4581), .o (n4582) );
  buffer buf_n4583( .i (n4582), .o (n4583) );
  assign n10996 = ~n5462 & n5465 ;
  buffer buf_n10997( .i (n10996), .o (n10997) );
  assign n10998 = n4583 & ~n10997 ;
  assign n10999 = ~n4583 & n10997 ;
  assign n11000 = n10998 | n10999 ;
  buffer buf_n11001( .i (n11000), .o (n11001) );
  assign n11056 = ~n5691 & n11001 ;
  assign n11057 = n10995 | n11056 ;
  buffer buf_n11058( .i (n11057), .o (n11058) );
  buffer buf_n11059( .i (n11058), .o (n11059) );
  buffer buf_n11060( .i (n11059), .o (n11060) );
  buffer buf_n11061( .i (n11060), .o (n11061) );
  buffer buf_n11062( .i (n11061), .o (n11062) );
  buffer buf_n11063( .i (n11062), .o (n11063) );
  buffer buf_n11064( .i (n11063), .o (n11064) );
  buffer buf_n11065( .i (n11064), .o (n11065) );
  buffer buf_n11066( .i (n11065), .o (n11066) );
  buffer buf_n11067( .i (n11066), .o (n11067) );
  buffer buf_n11068( .i (n11067), .o (n11068) );
  buffer buf_n11069( .i (n11068), .o (n11069) );
  buffer buf_n11070( .i (n11069), .o (n11070) );
  buffer buf_n11071( .i (n11070), .o (n11071) );
  buffer buf_n11072( .i (n11071), .o (n11072) );
  buffer buf_n11073( .i (n11072), .o (n11073) );
  buffer buf_n11074( .i (n11073), .o (n11074) );
  buffer buf_n11075( .i (n11074), .o (n11075) );
  buffer buf_n11076( .i (n11075), .o (n11076) );
  buffer buf_n11077( .i (n11076), .o (n11077) );
  buffer buf_n11078( .i (n11077), .o (n11078) );
  buffer buf_n11079( .i (n11078), .o (n11079) );
  buffer buf_n11080( .i (n11079), .o (n11080) );
  buffer buf_n11081( .i (n11080), .o (n11081) );
  buffer buf_n11082( .i (n11081), .o (n11082) );
  buffer buf_n11083( .i (n11082), .o (n11083) );
  buffer buf_n11084( .i (n11083), .o (n11084) );
  buffer buf_n11085( .i (n11084), .o (n11085) );
  buffer buf_n11086( .i (n11085), .o (n11086) );
  buffer buf_n11087( .i (n11086), .o (n11087) );
  buffer buf_n11088( .i (n11087), .o (n11088) );
  buffer buf_n11089( .i (n11088), .o (n11089) );
  buffer buf_n11090( .i (n11089), .o (n11090) );
  buffer buf_n11091( .i (n11090), .o (n11091) );
  buffer buf_n11092( .i (n11091), .o (n11092) );
  buffer buf_n11093( .i (n11092), .o (n11093) );
  buffer buf_n11094( .i (n11093), .o (n11094) );
  buffer buf_n11095( .i (n11094), .o (n11095) );
  buffer buf_n11096( .i (n11095), .o (n11096) );
  buffer buf_n11097( .i (n11096), .o (n11097) );
  buffer buf_n11098( .i (n11097), .o (n11098) );
  buffer buf_n11099( .i (n11098), .o (n11099) );
  buffer buf_n11100( .i (n11099), .o (n11100) );
  buffer buf_n11101( .i (n11100), .o (n11101) );
  buffer buf_n11102( .i (n11101), .o (n11102) );
  buffer buf_n11103( .i (n11102), .o (n11103) );
  buffer buf_n11104( .i (n11103), .o (n11104) );
  buffer buf_n11105( .i (n11104), .o (n11105) );
  buffer buf_n11106( .i (n11105), .o (n11106) );
  buffer buf_n11107( .i (n11106), .o (n11107) );
  buffer buf_n11108( .i (n11107), .o (n11108) );
  buffer buf_n11109( .i (n11108), .o (n11109) );
  buffer buf_n5306( .i (n5305), .o (n5306) );
  buffer buf_n5307( .i (n5306), .o (n5307) );
  assign n11110 = n5255 & ~n5310 ;
  buffer buf_n11111( .i (n11110), .o (n11111) );
  assign n11112 = n5307 & n11111 ;
  assign n11113 = n5307 | n11111 ;
  assign n11114 = ~n11112 & n11113 ;
  buffer buf_n11115( .i (n11114), .o (n11115) );
  buffer buf_n11116( .i (n11115), .o (n11116) );
  buffer buf_n11117( .i (n11116), .o (n11117) );
  buffer buf_n11118( .i (n11117), .o (n11118) );
  buffer buf_n11119( .i (n11118), .o (n11119) );
  buffer buf_n11120( .i (n11119), .o (n11120) );
  buffer buf_n11121( .i (n11120), .o (n11121) );
  buffer buf_n11122( .i (n11121), .o (n11122) );
  buffer buf_n11123( .i (n11122), .o (n11123) );
  buffer buf_n11124( .i (n11123), .o (n11124) );
  buffer buf_n11125( .i (n11124), .o (n11125) );
  buffer buf_n11126( .i (n11125), .o (n11126) );
  buffer buf_n11127( .i (n11126), .o (n11127) );
  buffer buf_n11128( .i (n11127), .o (n11128) );
  buffer buf_n11129( .i (n11128), .o (n11129) );
  buffer buf_n11130( .i (n11129), .o (n11130) );
  buffer buf_n11131( .i (n11130), .o (n11131) );
  buffer buf_n11132( .i (n11131), .o (n11132) );
  buffer buf_n11133( .i (n11132), .o (n11133) );
  buffer buf_n11134( .i (n11133), .o (n11134) );
  buffer buf_n11135( .i (n11134), .o (n11135) );
  buffer buf_n11136( .i (n11135), .o (n11136) );
  buffer buf_n11137( .i (n11136), .o (n11137) );
  buffer buf_n11138( .i (n11137), .o (n11138) );
  buffer buf_n11139( .i (n11138), .o (n11139) );
  buffer buf_n11140( .i (n11139), .o (n11140) );
  buffer buf_n11141( .i (n11140), .o (n11141) );
  buffer buf_n11142( .i (n11141), .o (n11142) );
  buffer buf_n11143( .i (n11142), .o (n11143) );
  buffer buf_n11144( .i (n11143), .o (n11144) );
  buffer buf_n11145( .i (n11144), .o (n11145) );
  buffer buf_n11146( .i (n11145), .o (n11146) );
  buffer buf_n11147( .i (n11146), .o (n11147) );
  buffer buf_n11148( .i (n11147), .o (n11148) );
  buffer buf_n11149( .i (n11148), .o (n11149) );
  buffer buf_n11150( .i (n11149), .o (n11150) );
  buffer buf_n11151( .i (n11150), .o (n11151) );
  buffer buf_n11152( .i (n11151), .o (n11152) );
  buffer buf_n11153( .i (n11152), .o (n11153) );
  buffer buf_n11154( .i (n11153), .o (n11154) );
  buffer buf_n11155( .i (n11154), .o (n11155) );
  buffer buf_n11156( .i (n11155), .o (n11156) );
  buffer buf_n11157( .i (n11156), .o (n11157) );
  buffer buf_n11158( .i (n11157), .o (n11158) );
  buffer buf_n11159( .i (n11158), .o (n11159) );
  buffer buf_n11160( .i (n11159), .o (n11160) );
  buffer buf_n11161( .i (n11160), .o (n11161) );
  buffer buf_n11162( .i (n11161), .o (n11162) );
  buffer buf_n11163( .i (n11162), .o (n11163) );
  buffer buf_n11164( .i (n11163), .o (n11164) );
  buffer buf_n11165( .i (n11164), .o (n11165) );
  buffer buf_n11166( .i (n11165), .o (n11166) );
  buffer buf_n11167( .i (n11166), .o (n11167) );
  buffer buf_n11168( .i (n11167), .o (n11168) );
  buffer buf_n11169( .i (n11168), .o (n11169) );
  buffer buf_n11170( .i (n11169), .o (n11170) );
  buffer buf_n11171( .i (n11170), .o (n11171) );
  buffer buf_n11172( .i (n11171), .o (n11172) );
  buffer buf_n11173( .i (n11172), .o (n11173) );
  buffer buf_n11174( .i (n11173), .o (n11174) );
  buffer buf_n11175( .i (n11174), .o (n11175) );
  buffer buf_n11176( .i (n11175), .o (n11176) );
  buffer buf_n11177( .i (n11176), .o (n11177) );
  buffer buf_n11178( .i (n11177), .o (n11178) );
  buffer buf_n11179( .i (n11178), .o (n11179) );
  buffer buf_n11180( .i (n11179), .o (n11180) );
  buffer buf_n11181( .i (n11180), .o (n11181) );
  buffer buf_n11182( .i (n11181), .o (n11182) );
  buffer buf_n11183( .i (n11182), .o (n11183) );
  buffer buf_n11184( .i (n11183), .o (n11184) );
  buffer buf_n11185( .i (n11184), .o (n11185) );
  buffer buf_n11186( .i (n11185), .o (n11186) );
  buffer buf_n11187( .i (n11186), .o (n11187) );
  buffer buf_n11188( .i (n11187), .o (n11188) );
  buffer buf_n11189( .i (n11188), .o (n11189) );
  buffer buf_n11190( .i (n11189), .o (n11190) );
  buffer buf_n11191( .i (n11190), .o (n11191) );
  buffer buf_n11192( .i (n11191), .o (n11192) );
  buffer buf_n11193( .i (n11192), .o (n11193) );
  buffer buf_n11194( .i (n11193), .o (n11194) );
  buffer buf_n8169( .i (n8168), .o (n8169) );
  assign n11195 = ~n8169 & n10903 ;
  assign n11196 = n10905 & ~n11195 ;
  assign n11197 = n3204 & n6082 ;
  buffer buf_n11198( .i (n6056), .o (n11198) );
  assign n11199 = n3318 & ~n11198 ;
  buffer buf_n11200( .i (n11199), .o (n11200) );
  buffer buf_n11201( .i (n11200), .o (n11201) );
  assign n11202 = ~n11197 & n11201 ;
  buffer buf_n6070( .i (n6069), .o (n6070) );
  assign n11203 = n3320 | n6070 ;
  assign n11204 = n3204 & ~n11200 ;
  assign n11205 = n11203 & n11204 ;
  assign n11206 = n11202 | n11205 ;
  assign n11207 = ~n6092 & n11206 ;
  assign n11208 = n10777 | n11207 ;
  buffer buf_n11209( .i (n11208), .o (n11209) );
  buffer buf_n11210( .i (n11209), .o (n11210) );
  buffer buf_n11211( .i (n11210), .o (n11211) );
  buffer buf_n11212( .i (n11211), .o (n11212) );
  buffer buf_n11213( .i (n11212), .o (n11213) );
  buffer buf_n11214( .i (n11213), .o (n11214) );
  buffer buf_n11215( .i (n11214), .o (n11215) );
  buffer buf_n11216( .i (n11215), .o (n11216) );
  buffer buf_n11217( .i (n11216), .o (n11217) );
  assign n11218 = n6102 & n8138 ;
  assign n11219 = n11217 | n11218 ;
  assign n11220 = n11196 & n11219 ;
  buffer buf_n11221( .i (n11220), .o (n11221) );
  buffer buf_n11222( .i (n11221), .o (n11222) );
  buffer buf_n11223( .i (n11222), .o (n11223) );
  buffer buf_n11224( .i (n11223), .o (n11224) );
  buffer buf_n11225( .i (n11224), .o (n11225) );
  buffer buf_n11226( .i (n11225), .o (n11226) );
  buffer buf_n11227( .i (n11226), .o (n11227) );
  buffer buf_n11228( .i (n11227), .o (n11228) );
  buffer buf_n11229( .i (n11228), .o (n11229) );
  buffer buf_n11230( .i (n11229), .o (n11230) );
  buffer buf_n11231( .i (n11230), .o (n11231) );
  buffer buf_n11232( .i (n11231), .o (n11232) );
  buffer buf_n11233( .i (n11232), .o (n11233) );
  buffer buf_n11234( .i (n11233), .o (n11234) );
  buffer buf_n11235( .i (n11234), .o (n11235) );
  buffer buf_n11236( .i (n11235), .o (n11236) );
  buffer buf_n11237( .i (n11236), .o (n11237) );
  buffer buf_n11238( .i (n11237), .o (n11238) );
  buffer buf_n11239( .i (n11238), .o (n11239) );
  buffer buf_n11240( .i (n11239), .o (n11240) );
  buffer buf_n11241( .i (n11240), .o (n11241) );
  buffer buf_n11242( .i (n11241), .o (n11242) );
  buffer buf_n11243( .i (n11242), .o (n11243) );
  buffer buf_n11244( .i (n11243), .o (n11244) );
  buffer buf_n11245( .i (n11244), .o (n11245) );
  buffer buf_n11246( .i (n11245), .o (n11246) );
  buffer buf_n11247( .i (n11246), .o (n11247) );
  buffer buf_n11248( .i (n11247), .o (n11248) );
  buffer buf_n11249( .i (n11248), .o (n11249) );
  buffer buf_n11250( .i (n11249), .o (n11250) );
  buffer buf_n11251( .i (n11250), .o (n11251) );
  buffer buf_n11252( .i (n11251), .o (n11252) );
  buffer buf_n11253( .i (n11252), .o (n11253) );
  buffer buf_n11254( .i (n11253), .o (n11254) );
  buffer buf_n11255( .i (n11254), .o (n11255) );
  buffer buf_n11256( .i (n11255), .o (n11256) );
  buffer buf_n11257( .i (n11256), .o (n11257) );
  buffer buf_n11258( .i (n11257), .o (n11258) );
  buffer buf_n11259( .i (n11258), .o (n11259) );
  buffer buf_n11260( .i (n11259), .o (n11260) );
  buffer buf_n11261( .i (n11260), .o (n11261) );
  buffer buf_n11262( .i (n11261), .o (n11262) );
  buffer buf_n11263( .i (n11262), .o (n11263) );
  buffer buf_n11264( .i (n11263), .o (n11264) );
  buffer buf_n11265( .i (n11264), .o (n11265) );
  buffer buf_n11266( .i (n11265), .o (n11266) );
  buffer buf_n11267( .i (n11266), .o (n11267) );
  buffer buf_n11268( .i (n11267), .o (n11268) );
  buffer buf_n11269( .i (n11268), .o (n11269) );
  buffer buf_n11270( .i (n11269), .o (n11270) );
  buffer buf_n11271( .i (n11270), .o (n11271) );
  buffer buf_n11272( .i (n11271), .o (n11272) );
  buffer buf_n11273( .i (n11272), .o (n11273) );
  buffer buf_n11274( .i (n11273), .o (n11274) );
  buffer buf_n11275( .i (n11274), .o (n11275) );
  buffer buf_n11276( .i (n11275), .o (n11276) );
  buffer buf_n11277( .i (n11276), .o (n11277) );
  buffer buf_n11278( .i (n11277), .o (n11278) );
  buffer buf_n11279( .i (n11278), .o (n11279) );
  buffer buf_n11280( .i (n11279), .o (n11280) );
  buffer buf_n11281( .i (n11280), .o (n11281) );
  buffer buf_n11282( .i (n11281), .o (n11282) );
  buffer buf_n11283( .i (n11282), .o (n11283) );
  buffer buf_n11284( .i (n11283), .o (n11284) );
  buffer buf_n11285( .i (n11284), .o (n11285) );
  buffer buf_n11286( .i (n11285), .o (n11286) );
  buffer buf_n11287( .i (n11286), .o (n11287) );
  buffer buf_n11288( .i (n11287), .o (n11288) );
  buffer buf_n11289( .i (n11288), .o (n11289) );
  buffer buf_n11290( .i (n11289), .o (n11290) );
  buffer buf_n11291( .i (n11290), .o (n11291) );
  buffer buf_n11292( .i (n11291), .o (n11292) );
  buffer buf_n11293( .i (n11292), .o (n11293) );
  buffer buf_n11294( .i (n11293), .o (n11294) );
  buffer buf_n11295( .i (n11294), .o (n11295) );
  buffer buf_n11296( .i (n11295), .o (n11296) );
  buffer buf_n11297( .i (n11296), .o (n11297) );
  buffer buf_n11298( .i (n11297), .o (n11298) );
  buffer buf_n11299( .i (n11298), .o (n11299) );
  buffer buf_n11300( .i (n11299), .o (n11300) );
  buffer buf_n11301( .i (n11300), .o (n11301) );
  buffer buf_n11302( .i (n11301), .o (n11302) );
  buffer buf_n11303( .i (n11302), .o (n11303) );
  buffer buf_n11304( .i (n11303), .o (n11304) );
  buffer buf_n11305( .i (n11304), .o (n11305) );
  buffer buf_n11306( .i (n11305), .o (n11306) );
  buffer buf_n11307( .i (n11306), .o (n11307) );
  buffer buf_n11308( .i (n11307), .o (n11308) );
  buffer buf_n11309( .i (n11308), .o (n11309) );
  buffer buf_n11310( .i (n11309), .o (n11310) );
  buffer buf_n11311( .i (n11310), .o (n11311) );
  buffer buf_n11312( .i (n11311), .o (n11312) );
  buffer buf_n11313( .i (n11312), .o (n11313) );
  buffer buf_n11314( .i (n11313), .o (n11314) );
  buffer buf_n11315( .i (n11314), .o (n11315) );
  buffer buf_n11316( .i (n11315), .o (n11316) );
  buffer buf_n11317( .i (n11316), .o (n11317) );
  buffer buf_n11318( .i (n11317), .o (n11318) );
  buffer buf_n11319( .i (n11318), .o (n11319) );
  buffer buf_n11320( .i (n11319), .o (n11320) );
  buffer buf_n11321( .i (n11320), .o (n11321) );
  buffer buf_n11322( .i (n11321), .o (n11322) );
  buffer buf_n11323( .i (n11322), .o (n11323) );
  buffer buf_n11324( .i (n11323), .o (n11324) );
  buffer buf_n11325( .i (n11324), .o (n11325) );
  buffer buf_n11326( .i (n11325), .o (n11326) );
  assign n11327 = ~n5738 & n10625 ;
  assign n11328 = n11326 | n11327 ;
  buffer buf_n11329( .i (n11328), .o (n11329) );
  buffer buf_n11330( .i (n11329), .o (n11330) );
  buffer buf_n11331( .i (n11330), .o (n11331) );
  buffer buf_n11332( .i (n11331), .o (n11332) );
  buffer buf_n11333( .i (n11332), .o (n11333) );
  buffer buf_n4800( .i (n4799), .o (n4800) );
  buffer buf_n4801( .i (n4800), .o (n4801) );
  assign n11334 = ~n4850 & n4853 ;
  buffer buf_n11335( .i (n11334), .o (n11335) );
  assign n11336 = ~n4801 & n11335 ;
  assign n11337 = n4801 & ~n11335 ;
  assign n11338 = n11336 | n11337 ;
  buffer buf_n11339( .i (n11338), .o (n11339) );
  buffer buf_n11340( .i (n11339), .o (n11340) );
  buffer buf_n11341( .i (n11340), .o (n11341) );
  buffer buf_n11342( .i (n11341), .o (n11342) );
  buffer buf_n11343( .i (n11342), .o (n11343) );
  buffer buf_n11344( .i (n11343), .o (n11344) );
  buffer buf_n11345( .i (n11344), .o (n11345) );
  buffer buf_n11346( .i (n11345), .o (n11346) );
  buffer buf_n11347( .i (n11346), .o (n11347) );
  buffer buf_n11348( .i (n11347), .o (n11348) );
  buffer buf_n11349( .i (n11348), .o (n11349) );
  buffer buf_n11350( .i (n11349), .o (n11350) );
  buffer buf_n11351( .i (n11350), .o (n11351) );
  buffer buf_n11352( .i (n11351), .o (n11352) );
  buffer buf_n11353( .i (n11352), .o (n11353) );
  buffer buf_n11354( .i (n11353), .o (n11354) );
  buffer buf_n11355( .i (n11354), .o (n11355) );
  buffer buf_n11356( .i (n11355), .o (n11356) );
  buffer buf_n11357( .i (n11356), .o (n11357) );
  buffer buf_n11358( .i (n11357), .o (n11358) );
  buffer buf_n11359( .i (n11358), .o (n11359) );
  buffer buf_n11360( .i (n11359), .o (n11360) );
  buffer buf_n11361( .i (n11360), .o (n11361) );
  buffer buf_n11362( .i (n11361), .o (n11362) );
  buffer buf_n11363( .i (n11362), .o (n11363) );
  buffer buf_n11364( .i (n11363), .o (n11364) );
  buffer buf_n11365( .i (n11364), .o (n11365) );
  buffer buf_n11366( .i (n11365), .o (n11366) );
  buffer buf_n11367( .i (n11366), .o (n11367) );
  buffer buf_n11368( .i (n11367), .o (n11368) );
  buffer buf_n11369( .i (n11368), .o (n11369) );
  buffer buf_n11370( .i (n11369), .o (n11370) );
  buffer buf_n11371( .i (n11370), .o (n11371) );
  buffer buf_n11372( .i (n11371), .o (n11372) );
  buffer buf_n11373( .i (n11372), .o (n11373) );
  buffer buf_n11374( .i (n11373), .o (n11374) );
  buffer buf_n11375( .i (n11374), .o (n11375) );
  buffer buf_n11376( .i (n11375), .o (n11376) );
  buffer buf_n11377( .i (n11376), .o (n11377) );
  buffer buf_n11378( .i (n11377), .o (n11378) );
  buffer buf_n11379( .i (n11378), .o (n11379) );
  buffer buf_n11380( .i (n11379), .o (n11380) );
  buffer buf_n11381( .i (n11380), .o (n11381) );
  buffer buf_n11382( .i (n11381), .o (n11382) );
  buffer buf_n11383( .i (n11382), .o (n11383) );
  buffer buf_n11384( .i (n11383), .o (n11384) );
  buffer buf_n11385( .i (n11384), .o (n11385) );
  buffer buf_n11386( .i (n11385), .o (n11386) );
  buffer buf_n11387( .i (n11386), .o (n11387) );
  buffer buf_n11388( .i (n11387), .o (n11388) );
  buffer buf_n11389( .i (n11388), .o (n11389) );
  buffer buf_n11390( .i (n11389), .o (n11390) );
  buffer buf_n11391( .i (n11390), .o (n11391) );
  buffer buf_n11392( .i (n11391), .o (n11392) );
  buffer buf_n11393( .i (n11392), .o (n11393) );
  buffer buf_n11394( .i (n11393), .o (n11394) );
  buffer buf_n11395( .i (n11394), .o (n11395) );
  buffer buf_n11396( .i (n11395), .o (n11396) );
  buffer buf_n11397( .i (n11396), .o (n11397) );
  buffer buf_n11398( .i (n11397), .o (n11398) );
  buffer buf_n11399( .i (n11398), .o (n11399) );
  buffer buf_n11400( .i (n11399), .o (n11400) );
  buffer buf_n11401( .i (n11400), .o (n11401) );
  buffer buf_n11402( .i (n11401), .o (n11402) );
  buffer buf_n11403( .i (n11402), .o (n11403) );
  buffer buf_n11404( .i (n11403), .o (n11404) );
  buffer buf_n11405( .i (n11404), .o (n11405) );
  buffer buf_n11406( .i (n11405), .o (n11406) );
  buffer buf_n11407( .i (n11406), .o (n11407) );
  buffer buf_n11408( .i (n11407), .o (n11408) );
  buffer buf_n11409( .i (n11408), .o (n11409) );
  buffer buf_n11410( .i (n11409), .o (n11410) );
  buffer buf_n11411( .i (n11410), .o (n11411) );
  buffer buf_n11412( .i (n11411), .o (n11412) );
  buffer buf_n11413( .i (n11412), .o (n11413) );
  buffer buf_n11414( .i (n11413), .o (n11414) );
  buffer buf_n11415( .i (n11414), .o (n11415) );
  buffer buf_n11416( .i (n11415), .o (n11416) );
  buffer buf_n11417( .i (n11416), .o (n11417) );
  buffer buf_n11418( .i (n11417), .o (n11418) );
  buffer buf_n11419( .i (n11418), .o (n11419) );
  buffer buf_n11420( .i (n11419), .o (n11420) );
  buffer buf_n11421( .i (n11420), .o (n11421) );
  buffer buf_n11422( .i (n11421), .o (n11422) );
  buffer buf_n11423( .i (n11422), .o (n11423) );
  buffer buf_n11424( .i (n11423), .o (n11424) );
  buffer buf_n11425( .i (n11424), .o (n11425) );
  buffer buf_n11426( .i (n11425), .o (n11426) );
  buffer buf_n11427( .i (n11426), .o (n11427) );
  buffer buf_n11428( .i (n11427), .o (n11428) );
  buffer buf_n11429( .i (n11428), .o (n11429) );
  buffer buf_n11430( .i (n11429), .o (n11430) );
  buffer buf_n11431( .i (n11430), .o (n11431) );
  buffer buf_n11432( .i (n11431), .o (n11432) );
  buffer buf_n11433( .i (n11432), .o (n11433) );
  buffer buf_n11434( .i (n11433), .o (n11434) );
  buffer buf_n11435( .i (n11434), .o (n11435) );
  buffer buf_n11436( .i (n11435), .o (n11436) );
  buffer buf_n11437( .i (n11436), .o (n11437) );
  buffer buf_n11438( .i (n11437), .o (n11438) );
  buffer buf_n11439( .i (n11438), .o (n11439) );
  buffer buf_n11440( .i (n11439), .o (n11440) );
  buffer buf_n11441( .i (n11440), .o (n11441) );
  buffer buf_n11442( .i (n11441), .o (n11442) );
  buffer buf_n11443( .i (n11442), .o (n11443) );
  buffer buf_n11444( .i (n11443), .o (n11444) );
  buffer buf_n11445( .i (n11444), .o (n11445) );
  buffer buf_n11446( .i (n11445), .o (n11446) );
  buffer buf_n11447( .i (n11446), .o (n11447) );
  buffer buf_n11448( .i (n11447), .o (n11448) );
  buffer buf_n11449( .i (n11448), .o (n11449) );
  buffer buf_n11450( .i (n11449), .o (n11450) );
  buffer buf_n11451( .i (n11450), .o (n11451) );
  buffer buf_n11452( .i (n11451), .o (n11452) );
  buffer buf_n11453( .i (n11452), .o (n11453) );
  buffer buf_n11454( .i (n11453), .o (n11454) );
  buffer buf_n11455( .i (n11454), .o (n11455) );
  buffer buf_n11456( .i (n11455), .o (n11456) );
  buffer buf_n11457( .i (n11456), .o (n11457) );
  buffer buf_n11458( .i (n11457), .o (n11458) );
  buffer buf_n11459( .i (n11458), .o (n11459) );
  buffer buf_n11460( .i (n11459), .o (n11460) );
  buffer buf_n11461( .i (n11460), .o (n11461) );
  buffer buf_n11462( .i (n11461), .o (n11462) );
  buffer buf_n11463( .i (n11462), .o (n11463) );
  buffer buf_n11464( .i (n11463), .o (n11464) );
  buffer buf_n11465( .i (n11464), .o (n11465) );
  buffer buf_n11466( .i (n11465), .o (n11466) );
  buffer buf_n11467( .i (n11466), .o (n11467) );
  buffer buf_n11468( .i (n11467), .o (n11468) );
  buffer buf_n11469( .i (n11468), .o (n11469) );
  buffer buf_n11470( .i (n11469), .o (n11470) );
  buffer buf_n11471( .i (n11470), .o (n11471) );
  buffer buf_n11472( .i (n11471), .o (n11472) );
  buffer buf_n11473( .i (n11472), .o (n11473) );
  buffer buf_n11474( .i (n11473), .o (n11474) );
  buffer buf_n11475( .i (n11474), .o (n11475) );
  buffer buf_n11476( .i (n11475), .o (n11476) );
  buffer buf_n11477( .i (n11476), .o (n11477) );
  buffer buf_n11478( .i (n11477), .o (n11478) );
  buffer buf_n11479( .i (n11478), .o (n11479) );
  buffer buf_n11480( .i (n11479), .o (n11480) );
  buffer buf_n11481( .i (n11480), .o (n11481) );
  buffer buf_n11482( .i (n11481), .o (n11482) );
  buffer buf_n11483( .i (n11482), .o (n11483) );
  buffer buf_n11484( .i (n11483), .o (n11484) );
  buffer buf_n11485( .i (n11484), .o (n11485) );
  buffer buf_n11486( .i (n11485), .o (n11486) );
  buffer buf_n11487( .i (n11486), .o (n11487) );
  buffer buf_n11488( .i (n11487), .o (n11488) );
  buffer buf_n11489( .i (n11488), .o (n11489) );
  buffer buf_n11490( .i (n11489), .o (n11490) );
  assign n11491 = ~n5632 & n11377 ;
  assign n11492 = n9258 & ~n9264 ;
  assign n11493 = n8924 & n9261 ;
  buffer buf_n11494( .i (n10227), .o (n11494) );
  assign n11495 = n11493 | n11494 ;
  assign n11496 = ~n45 & n8911 ;
  assign n11497 = n11495 | n11496 ;
  buffer buf_n11498( .i (n11497), .o (n11498) );
  assign n11499 = ~n11492 & n11498 ;
  buffer buf_n11500( .i (n10752), .o (n11500) );
  assign n11501 = n11499 & ~n11500 ;
  buffer buf_n11502( .i (n11501), .o (n11502) );
  assign n11503 = n9489 & n11500 ;
  assign n11504 = n9501 | n11503 ;
  assign n11505 = n11502 | n11504 ;
  assign n11506 = ~n10755 & n10756 ;
  assign n11507 = n11505 & ~n11506 ;
  buffer buf_n11508( .i (n11507), .o (n11508) );
  buffer buf_n11509( .i (n5926), .o (n11509) );
  assign n11510 = ~n11508 & n11509 ;
  buffer buf_n11511( .i (n5883), .o (n11511) );
  assign n11512 = ~n11510 & n11511 ;
  buffer buf_n11513( .i (n11512), .o (n11513) );
  assign n11514 = n1308 & n3555 ;
  buffer buf_n11515( .i (n11514), .o (n11515) );
  buffer buf_n11516( .i (n11515), .o (n11516) );
  assign n11517 = n9879 & ~n11516 ;
  assign n11518 = n9881 | n11517 ;
  assign n11519 = n10916 & n11515 ;
  buffer buf_n1310( .i (n1309), .o (n1310) );
  assign n11520 = n3556 & n10908 ;
  assign n11521 = n1310 | n11520 ;
  assign n11522 = ~n11519 & n11521 ;
  buffer buf_n11523( .i (n9879), .o (n11523) );
  assign n11524 = n11522 | n11523 ;
  assign n11525 = ~n11518 & n11524 ;
  buffer buf_n11526( .i (n11525), .o (n11526) );
  buffer buf_n11527( .i (n11526), .o (n11527) );
  assign n11528 = n10777 | n11527 ;
  buffer buf_n11529( .i (n11528), .o (n11529) );
  buffer buf_n11530( .i (n11529), .o (n11530) );
  buffer buf_n11531( .i (n11530), .o (n11531) );
  buffer buf_n11532( .i (n11531), .o (n11532) );
  buffer buf_n11533( .i (n11532), .o (n11533) );
  buffer buf_n11534( .i (n11533), .o (n11534) );
  buffer buf_n11535( .i (n11534), .o (n11535) );
  buffer buf_n11536( .i (n11535), .o (n11536) );
  buffer buf_n11537( .i (n11536), .o (n11537) );
  assign n11538 = ~n9622 & n10745 ;
  assign n11539 = n5951 | n11538 ;
  buffer buf_n11540( .i (n11539), .o (n11540) );
  buffer buf_n11541( .i (n10761), .o (n11541) );
  assign n11542 = n11540 & n11541 ;
  assign n11543 = n11537 | n11542 ;
  assign n11544 = n11513 & n11543 ;
  assign n11545 = n11491 | n11544 ;
  buffer buf_n11546( .i (n11545), .o (n11546) );
  buffer buf_n11547( .i (n11546), .o (n11547) );
  buffer buf_n11548( .i (n11547), .o (n11548) );
  buffer buf_n11549( .i (n11548), .o (n11549) );
  buffer buf_n11550( .i (n11549), .o (n11550) );
  buffer buf_n11551( .i (n11550), .o (n11551) );
  buffer buf_n11552( .i (n11551), .o (n11552) );
  buffer buf_n11553( .i (n11552), .o (n11553) );
  buffer buf_n11554( .i (n11553), .o (n11554) );
  buffer buf_n11555( .i (n11554), .o (n11555) );
  buffer buf_n11556( .i (n11555), .o (n11556) );
  buffer buf_n11557( .i (n11556), .o (n11557) );
  buffer buf_n11558( .i (n11557), .o (n11558) );
  buffer buf_n11559( .i (n11558), .o (n11559) );
  buffer buf_n11560( .i (n11559), .o (n11560) );
  buffer buf_n11561( .i (n11560), .o (n11561) );
  buffer buf_n11562( .i (n11561), .o (n11562) );
  buffer buf_n11563( .i (n11562), .o (n11563) );
  buffer buf_n11564( .i (n11563), .o (n11564) );
  buffer buf_n11565( .i (n11564), .o (n11565) );
  buffer buf_n11566( .i (n11565), .o (n11566) );
  buffer buf_n11567( .i (n11566), .o (n11567) );
  buffer buf_n11568( .i (n11567), .o (n11568) );
  buffer buf_n11569( .i (n11568), .o (n11569) );
  buffer buf_n11570( .i (n11569), .o (n11570) );
  buffer buf_n11571( .i (n11570), .o (n11571) );
  buffer buf_n11572( .i (n11571), .o (n11572) );
  buffer buf_n11573( .i (n11572), .o (n11573) );
  buffer buf_n11574( .i (n11573), .o (n11574) );
  buffer buf_n11575( .i (n11574), .o (n11575) );
  buffer buf_n11576( .i (n11575), .o (n11576) );
  buffer buf_n11577( .i (n11576), .o (n11577) );
  buffer buf_n11578( .i (n11577), .o (n11578) );
  buffer buf_n11579( .i (n11578), .o (n11579) );
  buffer buf_n11580( .i (n11579), .o (n11580) );
  buffer buf_n11581( .i (n11580), .o (n11581) );
  buffer buf_n11582( .i (n11581), .o (n11582) );
  buffer buf_n11583( .i (n11582), .o (n11583) );
  buffer buf_n11584( .i (n11583), .o (n11584) );
  buffer buf_n11585( .i (n11584), .o (n11585) );
  buffer buf_n11586( .i (n11585), .o (n11586) );
  buffer buf_n11587( .i (n11586), .o (n11587) );
  buffer buf_n11588( .i (n11587), .o (n11588) );
  buffer buf_n11589( .i (n11588), .o (n11589) );
  buffer buf_n11590( .i (n11589), .o (n11590) );
  buffer buf_n11591( .i (n11590), .o (n11591) );
  buffer buf_n11592( .i (n11591), .o (n11592) );
  buffer buf_n11593( .i (n11592), .o (n11593) );
  buffer buf_n11594( .i (n11593), .o (n11594) );
  buffer buf_n11595( .i (n11594), .o (n11595) );
  buffer buf_n11596( .i (n11595), .o (n11596) );
  buffer buf_n11597( .i (n11596), .o (n11597) );
  buffer buf_n11598( .i (n11597), .o (n11598) );
  buffer buf_n11599( .i (n11598), .o (n11599) );
  buffer buf_n11600( .i (n11599), .o (n11600) );
  buffer buf_n11601( .i (n11600), .o (n11601) );
  buffer buf_n11602( .i (n11601), .o (n11602) );
  buffer buf_n11603( .i (n11602), .o (n11603) );
  buffer buf_n11604( .i (n11603), .o (n11604) );
  buffer buf_n11605( .i (n11604), .o (n11605) );
  buffer buf_n11606( .i (n11605), .o (n11606) );
  buffer buf_n11607( .i (n11606), .o (n11607) );
  buffer buf_n11608( .i (n11607), .o (n11608) );
  buffer buf_n11609( .i (n11608), .o (n11609) );
  buffer buf_n11610( .i (n11609), .o (n11610) );
  buffer buf_n11611( .i (n11610), .o (n11611) );
  buffer buf_n11612( .i (n11611), .o (n11612) );
  buffer buf_n11613( .i (n11612), .o (n11613) );
  buffer buf_n11614( .i (n11613), .o (n11614) );
  buffer buf_n11615( .i (n11614), .o (n11615) );
  buffer buf_n11616( .i (n11615), .o (n11616) );
  buffer buf_n11617( .i (n11616), .o (n11617) );
  buffer buf_n11618( .i (n11617), .o (n11618) );
  buffer buf_n11619( .i (n11618), .o (n11619) );
  buffer buf_n11620( .i (n11619), .o (n11620) );
  buffer buf_n11621( .i (n11620), .o (n11621) );
  buffer buf_n11622( .i (n11621), .o (n11622) );
  buffer buf_n11623( .i (n11622), .o (n11623) );
  buffer buf_n11624( .i (n11623), .o (n11624) );
  buffer buf_n11625( .i (n11624), .o (n11625) );
  buffer buf_n11626( .i (n11625), .o (n11626) );
  buffer buf_n11627( .i (n11626), .o (n11627) );
  buffer buf_n11628( .i (n11627), .o (n11628) );
  buffer buf_n11629( .i (n11628), .o (n11629) );
  buffer buf_n11630( .i (n11629), .o (n11630) );
  buffer buf_n11631( .i (n11630), .o (n11631) );
  buffer buf_n11632( .i (n11631), .o (n11632) );
  buffer buf_n11633( .i (n11632), .o (n11633) );
  buffer buf_n11634( .i (n11633), .o (n11634) );
  buffer buf_n11635( .i (n11634), .o (n11635) );
  buffer buf_n11636( .i (n11635), .o (n11636) );
  buffer buf_n11637( .i (n11636), .o (n11637) );
  buffer buf_n11638( .i (n11637), .o (n11638) );
  buffer buf_n11639( .i (n11638), .o (n11639) );
  buffer buf_n11640( .i (n11639), .o (n11640) );
  buffer buf_n11641( .i (n11640), .o (n11641) );
  buffer buf_n11642( .i (n11641), .o (n11642) );
  buffer buf_n11643( .i (n11642), .o (n11643) );
  buffer buf_n11644( .i (n11643), .o (n11644) );
  buffer buf_n11645( .i (n11644), .o (n11645) );
  buffer buf_n11646( .i (n11645), .o (n11646) );
  buffer buf_n11647( .i (n11646), .o (n11647) );
  buffer buf_n11648( .i (n11647), .o (n11648) );
  buffer buf_n11649( .i (n11648), .o (n11649) );
  buffer buf_n11650( .i (n11649), .o (n11650) );
  buffer buf_n11651( .i (n11650), .o (n11651) );
  buffer buf_n11652( .i (n11651), .o (n11652) );
  buffer buf_n11653( .i (n11652), .o (n11653) );
  buffer buf_n11654( .i (n11653), .o (n11654) );
  buffer buf_n11655( .i (n11654), .o (n11655) );
  buffer buf_n11656( .i (n11655), .o (n11656) );
  buffer buf_n8855( .i (n8854), .o (n8855) );
  buffer buf_n8856( .i (n8855), .o (n8856) );
  buffer buf_n8857( .i (n8856), .o (n8857) );
  buffer buf_n8858( .i (n8857), .o (n8858) );
  buffer buf_n8859( .i (n8858), .o (n8859) );
  buffer buf_n9696( .i (n9695), .o (n9696) );
  buffer buf_n9697( .i (n9696), .o (n9697) );
  buffer buf_n9698( .i (n9697), .o (n9698) );
  buffer buf_n9699( .i (n9698), .o (n9699) );
  buffer buf_n9700( .i (n9699), .o (n9700) );
  buffer buf_n9701( .i (n9700), .o (n9701) );
  buffer buf_n9702( .i (n9701), .o (n9702) );
  buffer buf_n9703( .i (n9702), .o (n9703) );
  buffer buf_n9704( .i (n9703), .o (n9704) );
  buffer buf_n9705( .i (n9704), .o (n9705) );
  buffer buf_n9706( .i (n9705), .o (n9706) );
  buffer buf_n9707( .i (n9706), .o (n9707) );
  buffer buf_n9708( .i (n9707), .o (n9708) );
  buffer buf_n9709( .i (n9708), .o (n9709) );
  buffer buf_n9710( .i (n9709), .o (n9710) );
  buffer buf_n9711( .i (n9710), .o (n9711) );
  buffer buf_n9712( .i (n9711), .o (n9712) );
  buffer buf_n9713( .i (n9712), .o (n9713) );
  buffer buf_n9714( .i (n9713), .o (n9714) );
  buffer buf_n9715( .i (n9714), .o (n9715) );
  buffer buf_n9716( .i (n9715), .o (n9716) );
  buffer buf_n9717( .i (n9716), .o (n9717) );
  buffer buf_n9718( .i (n9717), .o (n9718) );
  buffer buf_n9719( .i (n9718), .o (n9719) );
  buffer buf_n9720( .i (n9719), .o (n9720) );
  buffer buf_n9721( .i (n9720), .o (n9721) );
  buffer buf_n9722( .i (n9721), .o (n9722) );
  buffer buf_n9723( .i (n9722), .o (n9723) );
  buffer buf_n9724( .i (n9723), .o (n9724) );
  buffer buf_n9725( .i (n9724), .o (n9725) );
  buffer buf_n9726( .i (n9725), .o (n9726) );
  buffer buf_n9727( .i (n9726), .o (n9727) );
  buffer buf_n9728( .i (n9727), .o (n9728) );
  buffer buf_n9729( .i (n9728), .o (n9729) );
  buffer buf_n9730( .i (n9729), .o (n9730) );
  buffer buf_n9731( .i (n9730), .o (n9731) );
  buffer buf_n9732( .i (n9731), .o (n9732) );
  buffer buf_n9733( .i (n9732), .o (n9733) );
  buffer buf_n9734( .i (n9733), .o (n9734) );
  buffer buf_n9735( .i (n9734), .o (n9735) );
  buffer buf_n9736( .i (n9735), .o (n9736) );
  buffer buf_n9737( .i (n9736), .o (n9737) );
  buffer buf_n9738( .i (n9737), .o (n9738) );
  buffer buf_n9739( .i (n9738), .o (n9739) );
  buffer buf_n9740( .i (n9739), .o (n9740) );
  buffer buf_n9741( .i (n9740), .o (n9741) );
  buffer buf_n9742( .i (n9741), .o (n9742) );
  buffer buf_n9743( .i (n9742), .o (n9743) );
  buffer buf_n9744( .i (n9743), .o (n9744) );
  buffer buf_n9745( .i (n9744), .o (n9745) );
  buffer buf_n9746( .i (n9745), .o (n9746) );
  buffer buf_n9747( .i (n9746), .o (n9747) );
  buffer buf_n9748( .i (n9747), .o (n9748) );
  buffer buf_n9749( .i (n9748), .o (n9749) );
  buffer buf_n9750( .i (n9749), .o (n9750) );
  buffer buf_n9751( .i (n9750), .o (n9751) );
  buffer buf_n9752( .i (n9751), .o (n9752) );
  buffer buf_n9753( .i (n9752), .o (n9753) );
  buffer buf_n9754( .i (n9753), .o (n9754) );
  buffer buf_n9755( .i (n9754), .o (n9755) );
  buffer buf_n9756( .i (n9755), .o (n9756) );
  buffer buf_n9757( .i (n9756), .o (n9757) );
  buffer buf_n9758( .i (n9757), .o (n9758) );
  buffer buf_n9759( .i (n9758), .o (n9759) );
  buffer buf_n9760( .i (n9759), .o (n9760) );
  buffer buf_n9761( .i (n9760), .o (n9761) );
  buffer buf_n9762( .i (n9761), .o (n9762) );
  buffer buf_n9763( .i (n9762), .o (n9763) );
  buffer buf_n9764( .i (n9763), .o (n9764) );
  buffer buf_n9765( .i (n9764), .o (n9765) );
  buffer buf_n9766( .i (n9765), .o (n9766) );
  buffer buf_n9767( .i (n9766), .o (n9767) );
  buffer buf_n9768( .i (n9767), .o (n9768) );
  buffer buf_n9769( .i (n9768), .o (n9769) );
  buffer buf_n9770( .i (n9769), .o (n9770) );
  buffer buf_n9771( .i (n9770), .o (n9771) );
  buffer buf_n9772( .i (n9771), .o (n9772) );
  buffer buf_n9773( .i (n9772), .o (n9773) );
  buffer buf_n9774( .i (n9773), .o (n9774) );
  buffer buf_n9775( .i (n9774), .o (n9775) );
  buffer buf_n9776( .i (n9775), .o (n9776) );
  buffer buf_n9777( .i (n9776), .o (n9777) );
  buffer buf_n9778( .i (n9777), .o (n9778) );
  buffer buf_n9779( .i (n9778), .o (n9779) );
  buffer buf_n9780( .i (n9779), .o (n9780) );
  buffer buf_n9781( .i (n9780), .o (n9781) );
  buffer buf_n9782( .i (n9781), .o (n9782) );
  buffer buf_n9783( .i (n9782), .o (n9783) );
  buffer buf_n9784( .i (n9783), .o (n9784) );
  assign n11657 = ~n5716 & n7827 ;
  buffer buf_n11658( .i (n11198), .o (n11658) );
  assign n11659 = n4092 & ~n11658 ;
  buffer buf_n11660( .i (n11659), .o (n11660) );
  assign n11661 = n4092 | n6069 ;
  assign n11662 = n273 & n11661 ;
  assign n11663 = n11660 | n11662 ;
  buffer buf_n11664( .i (n11663), .o (n11664) );
  assign n11665 = n273 & n6082 ;
  assign n11666 = n11660 & n11665 ;
  assign n11667 = n6091 | n11666 ;
  assign n11668 = n11664 & ~n11667 ;
  buffer buf_n11669( .i (n5917), .o (n11669) );
  buffer buf_n11670( .i (n11669), .o (n11670) );
  assign n11671 = n11668 | n11670 ;
  buffer buf_n11672( .i (n11671), .o (n11672) );
  buffer buf_n11673( .i (n11672), .o (n11673) );
  buffer buf_n11674( .i (n11673), .o (n11674) );
  buffer buf_n11675( .i (n11674), .o (n11675) );
  buffer buf_n11676( .i (n11675), .o (n11676) );
  buffer buf_n11677( .i (n11676), .o (n11677) );
  buffer buf_n11678( .i (n11677), .o (n11678) );
  buffer buf_n11679( .i (n11678), .o (n11679) );
  buffer buf_n11680( .i (n11679), .o (n11680) );
  assign n11681 = n9471 & n9622 ;
  assign n11682 = n8123 | n9258 ;
  buffer buf_n6188( .i (n6187), .o (n6188) );
  buffer buf_n11683( .i (n10735), .o (n11683) );
  assign n11684 = ~n6188 & n11683 ;
  assign n11685 = n11682 & ~n11684 ;
  assign n11686 = n11500 | n11685 ;
  assign n11687 = ~n10738 & n11500 ;
  assign n11688 = n11686 & ~n11687 ;
  assign n11689 = ~n10756 & n11688 ;
  buffer buf_n11690( .i (n11689), .o (n11690) );
  assign n11691 = n11681 | n11690 ;
  buffer buf_n11692( .i (n11691), .o (n11692) );
  assign n11693 = n11541 & n11692 ;
  assign n11694 = n11680 | n11693 ;
  assign n11695 = n9500 & ~n10756 ;
  assign n11696 = n8681 | n11695 ;
  buffer buf_n11697( .i (n11696), .o (n11697) );
  buffer buf_n11698( .i (n11697), .o (n11698) );
  assign n11699 = n10903 & ~n11698 ;
  assign n11700 = n10905 & ~n11699 ;
  assign n11701 = n11694 & n11700 ;
  buffer buf_n11702( .i (n11701), .o (n11702) );
  buffer buf_n11703( .i (n11702), .o (n11703) );
  buffer buf_n11704( .i (n11703), .o (n11704) );
  buffer buf_n11705( .i (n11704), .o (n11705) );
  buffer buf_n11706( .i (n11705), .o (n11706) );
  buffer buf_n11707( .i (n11706), .o (n11707) );
  buffer buf_n11708( .i (n11707), .o (n11708) );
  buffer buf_n11709( .i (n11708), .o (n11709) );
  buffer buf_n11710( .i (n11709), .o (n11710) );
  buffer buf_n11711( .i (n11710), .o (n11711) );
  buffer buf_n11712( .i (n11711), .o (n11712) );
  buffer buf_n11713( .i (n11712), .o (n11713) );
  buffer buf_n11714( .i (n11713), .o (n11714) );
  buffer buf_n11715( .i (n11714), .o (n11715) );
  buffer buf_n11716( .i (n11715), .o (n11716) );
  buffer buf_n11717( .i (n11716), .o (n11717) );
  buffer buf_n11718( .i (n11717), .o (n11718) );
  buffer buf_n11719( .i (n11718), .o (n11719) );
  buffer buf_n11720( .i (n11719), .o (n11720) );
  buffer buf_n11721( .i (n11720), .o (n11721) );
  buffer buf_n11722( .i (n11721), .o (n11722) );
  buffer buf_n11723( .i (n11722), .o (n11723) );
  buffer buf_n11724( .i (n11723), .o (n11724) );
  buffer buf_n11725( .i (n11724), .o (n11725) );
  buffer buf_n11726( .i (n11725), .o (n11726) );
  buffer buf_n11727( .i (n11726), .o (n11727) );
  buffer buf_n11728( .i (n11727), .o (n11728) );
  buffer buf_n11729( .i (n11728), .o (n11729) );
  buffer buf_n11730( .i (n11729), .o (n11730) );
  buffer buf_n11731( .i (n11730), .o (n11731) );
  buffer buf_n11732( .i (n11731), .o (n11732) );
  buffer buf_n11733( .i (n11732), .o (n11733) );
  buffer buf_n11734( .i (n11733), .o (n11734) );
  buffer buf_n11735( .i (n11734), .o (n11735) );
  buffer buf_n11736( .i (n11735), .o (n11736) );
  buffer buf_n11737( .i (n11736), .o (n11737) );
  buffer buf_n11738( .i (n11737), .o (n11738) );
  buffer buf_n11739( .i (n11738), .o (n11739) );
  buffer buf_n11740( .i (n11739), .o (n11740) );
  buffer buf_n11741( .i (n11740), .o (n11741) );
  buffer buf_n11742( .i (n11741), .o (n11742) );
  buffer buf_n11743( .i (n11742), .o (n11743) );
  buffer buf_n11744( .i (n11743), .o (n11744) );
  buffer buf_n11745( .i (n11744), .o (n11745) );
  buffer buf_n11746( .i (n11745), .o (n11746) );
  buffer buf_n11747( .i (n11746), .o (n11747) );
  buffer buf_n11748( .i (n11747), .o (n11748) );
  buffer buf_n11749( .i (n11748), .o (n11749) );
  buffer buf_n11750( .i (n11749), .o (n11750) );
  buffer buf_n11751( .i (n11750), .o (n11751) );
  buffer buf_n11752( .i (n11751), .o (n11752) );
  buffer buf_n11753( .i (n11752), .o (n11753) );
  buffer buf_n11754( .i (n11753), .o (n11754) );
  buffer buf_n11755( .i (n11754), .o (n11755) );
  buffer buf_n11756( .i (n11755), .o (n11756) );
  buffer buf_n11757( .i (n11756), .o (n11757) );
  buffer buf_n11758( .i (n11757), .o (n11758) );
  buffer buf_n11759( .i (n11758), .o (n11759) );
  buffer buf_n11760( .i (n11759), .o (n11760) );
  buffer buf_n11761( .i (n11760), .o (n11761) );
  buffer buf_n11762( .i (n11761), .o (n11762) );
  buffer buf_n11763( .i (n11762), .o (n11763) );
  buffer buf_n11764( .i (n11763), .o (n11764) );
  buffer buf_n11765( .i (n11764), .o (n11765) );
  buffer buf_n11766( .i (n11765), .o (n11766) );
  buffer buf_n11767( .i (n11766), .o (n11767) );
  buffer buf_n11768( .i (n11767), .o (n11768) );
  buffer buf_n11769( .i (n11768), .o (n11769) );
  buffer buf_n11770( .i (n11769), .o (n11770) );
  buffer buf_n11771( .i (n11770), .o (n11771) );
  buffer buf_n11772( .i (n11771), .o (n11772) );
  buffer buf_n11773( .i (n11772), .o (n11773) );
  buffer buf_n11774( .i (n11773), .o (n11774) );
  buffer buf_n11775( .i (n11774), .o (n11775) );
  buffer buf_n11776( .i (n11775), .o (n11776) );
  buffer buf_n11777( .i (n11776), .o (n11777) );
  buffer buf_n11778( .i (n11777), .o (n11778) );
  buffer buf_n11779( .i (n11778), .o (n11779) );
  buffer buf_n11780( .i (n11779), .o (n11780) );
  buffer buf_n11781( .i (n11780), .o (n11781) );
  buffer buf_n11782( .i (n11781), .o (n11782) );
  buffer buf_n11783( .i (n11782), .o (n11783) );
  buffer buf_n11784( .i (n11783), .o (n11784) );
  buffer buf_n11785( .i (n11784), .o (n11785) );
  assign n11786 = n11657 | n11785 ;
  buffer buf_n11787( .i (n11786), .o (n11787) );
  buffer buf_n11788( .i (n11787), .o (n11788) );
  buffer buf_n11789( .i (n11788), .o (n11789) );
  buffer buf_n11790( .i (n11789), .o (n11790) );
  buffer buf_n11791( .i (n11790), .o (n11791) );
  buffer buf_n11792( .i (n11791), .o (n11792) );
  buffer buf_n11793( .i (n11792), .o (n11793) );
  buffer buf_n11794( .i (n11793), .o (n11794) );
  buffer buf_n11795( .i (n11794), .o (n11795) );
  buffer buf_n11796( .i (n11795), .o (n11796) );
  buffer buf_n11797( .i (n11796), .o (n11797) );
  buffer buf_n11798( .i (n11797), .o (n11798) );
  buffer buf_n11799( .i (n11798), .o (n11799) );
  buffer buf_n11800( .i (n11799), .o (n11800) );
  buffer buf_n11801( .i (n11800), .o (n11801) );
  buffer buf_n11802( .i (n11801), .o (n11802) );
  buffer buf_n11803( .i (n11802), .o (n11803) );
  buffer buf_n11804( .i (n11803), .o (n11804) );
  buffer buf_n11805( .i (n11804), .o (n11805) );
  buffer buf_n11806( .i (n11805), .o (n11806) );
  buffer buf_n11807( .i (n11806), .o (n11807) );
  buffer buf_n11808( .i (n11807), .o (n11808) );
  buffer buf_n11809( .i (n11808), .o (n11809) );
  buffer buf_n11810( .i (n11809), .o (n11810) );
  buffer buf_n11811( .i (n11810), .o (n11811) );
  buffer buf_n11812( .i (n11811), .o (n11812) );
  buffer buf_n11813( .i (n11812), .o (n11813) );
  assign n11814 = ~n5671 & n7747 ;
  assign n11815 = n525 & n1139 ;
  buffer buf_n11816( .i (n11815), .o (n11816) );
  buffer buf_n11817( .i (n11816), .o (n11817) );
  assign n11818 = n11658 & ~n11817 ;
  assign n11819 = n9881 | n11818 ;
  assign n11820 = n10916 & n11816 ;
  assign n11821 = n1140 & n10908 ;
  assign n11822 = n527 | n11821 ;
  assign n11823 = ~n11820 & n11822 ;
  assign n11824 = n11523 | n11823 ;
  assign n11825 = ~n11819 & n11824 ;
  buffer buf_n11826( .i (n11825), .o (n11826) );
  buffer buf_n11827( .i (n11826), .o (n11827) );
  assign n11828 = n11670 | n11827 ;
  buffer buf_n11829( .i (n11828), .o (n11829) );
  buffer buf_n11830( .i (n11829), .o (n11830) );
  buffer buf_n11831( .i (n11830), .o (n11831) );
  buffer buf_n11832( .i (n11831), .o (n11832) );
  buffer buf_n11833( .i (n11832), .o (n11833) );
  buffer buf_n11834( .i (n11833), .o (n11834) );
  buffer buf_n11835( .i (n11834), .o (n11835) );
  buffer buf_n11836( .i (n11835), .o (n11836) );
  assign n11837 = n9659 & n10761 ;
  assign n11838 = n11836 | n11837 ;
  buffer buf_n11839( .i (n11838), .o (n11839) );
  assign n11840 = ~n9625 & n10903 ;
  assign n11841 = n10905 & ~n11840 ;
  assign n11842 = n11839 & n11841 ;
  buffer buf_n11843( .i (n11842), .o (n11843) );
  buffer buf_n11844( .i (n11843), .o (n11844) );
  buffer buf_n11845( .i (n11844), .o (n11845) );
  buffer buf_n11846( .i (n11845), .o (n11846) );
  buffer buf_n11847( .i (n11846), .o (n11847) );
  buffer buf_n11848( .i (n11847), .o (n11848) );
  buffer buf_n11849( .i (n11848), .o (n11849) );
  buffer buf_n11850( .i (n11849), .o (n11850) );
  buffer buf_n11851( .i (n11850), .o (n11851) );
  buffer buf_n11852( .i (n11851), .o (n11852) );
  buffer buf_n11853( .i (n11852), .o (n11853) );
  buffer buf_n11854( .i (n11853), .o (n11854) );
  buffer buf_n11855( .i (n11854), .o (n11855) );
  buffer buf_n11856( .i (n11855), .o (n11856) );
  buffer buf_n11857( .i (n11856), .o (n11857) );
  buffer buf_n11858( .i (n11857), .o (n11858) );
  buffer buf_n11859( .i (n11858), .o (n11859) );
  buffer buf_n11860( .i (n11859), .o (n11860) );
  buffer buf_n11861( .i (n11860), .o (n11861) );
  buffer buf_n11862( .i (n11861), .o (n11862) );
  buffer buf_n11863( .i (n11862), .o (n11863) );
  buffer buf_n11864( .i (n11863), .o (n11864) );
  buffer buf_n11865( .i (n11864), .o (n11865) );
  buffer buf_n11866( .i (n11865), .o (n11866) );
  buffer buf_n11867( .i (n11866), .o (n11867) );
  buffer buf_n11868( .i (n11867), .o (n11868) );
  buffer buf_n11869( .i (n11868), .o (n11869) );
  buffer buf_n11870( .i (n11869), .o (n11870) );
  buffer buf_n11871( .i (n11870), .o (n11871) );
  buffer buf_n11872( .i (n11871), .o (n11872) );
  buffer buf_n11873( .i (n11872), .o (n11873) );
  buffer buf_n11874( .i (n11873), .o (n11874) );
  buffer buf_n11875( .i (n11874), .o (n11875) );
  buffer buf_n11876( .i (n11875), .o (n11876) );
  buffer buf_n11877( .i (n11876), .o (n11877) );
  buffer buf_n11878( .i (n11877), .o (n11878) );
  buffer buf_n11879( .i (n11878), .o (n11879) );
  buffer buf_n11880( .i (n11879), .o (n11880) );
  buffer buf_n11881( .i (n11880), .o (n11881) );
  assign n11882 = n11814 | n11881 ;
  buffer buf_n11883( .i (n11882), .o (n11883) );
  buffer buf_n11884( .i (n11883), .o (n11884) );
  buffer buf_n11885( .i (n11884), .o (n11885) );
  buffer buf_n11886( .i (n11885), .o (n11886) );
  buffer buf_n11887( .i (n11886), .o (n11887) );
  buffer buf_n11888( .i (n11887), .o (n11888) );
  buffer buf_n11889( .i (n11888), .o (n11889) );
  buffer buf_n11890( .i (n11889), .o (n11890) );
  buffer buf_n11891( .i (n11890), .o (n11891) );
  buffer buf_n11892( .i (n11891), .o (n11892) );
  buffer buf_n11893( .i (n11892), .o (n11893) );
  buffer buf_n11894( .i (n11893), .o (n11894) );
  buffer buf_n11895( .i (n11894), .o (n11895) );
  buffer buf_n11896( .i (n11895), .o (n11896) );
  buffer buf_n11897( .i (n11896), .o (n11897) );
  buffer buf_n11898( .i (n11897), .o (n11898) );
  buffer buf_n11899( .i (n11898), .o (n11899) );
  buffer buf_n11900( .i (n11899), .o (n11900) );
  buffer buf_n11901( .i (n11900), .o (n11901) );
  buffer buf_n11902( .i (n11901), .o (n11902) );
  buffer buf_n11903( .i (n11902), .o (n11903) );
  buffer buf_n11904( .i (n11903), .o (n11904) );
  buffer buf_n11905( .i (n11904), .o (n11905) );
  buffer buf_n11906( .i (n11905), .o (n11906) );
  buffer buf_n11907( .i (n11906), .o (n11907) );
  buffer buf_n11908( .i (n11907), .o (n11908) );
  buffer buf_n11909( .i (n11908), .o (n11909) );
  buffer buf_n11910( .i (n11909), .o (n11910) );
  buffer buf_n11911( .i (n11910), .o (n11911) );
  buffer buf_n11912( .i (n11911), .o (n11912) );
  buffer buf_n11913( .i (n11912), .o (n11913) );
  buffer buf_n11914( .i (n11913), .o (n11914) );
  buffer buf_n11915( .i (n11914), .o (n11915) );
  buffer buf_n11916( .i (n11915), .o (n11916) );
  buffer buf_n11917( .i (n11916), .o (n11917) );
  buffer buf_n11918( .i (n11917), .o (n11918) );
  buffer buf_n11919( .i (n11918), .o (n11919) );
  buffer buf_n11920( .i (n11919), .o (n11920) );
  buffer buf_n11921( .i (n11920), .o (n11921) );
  buffer buf_n11922( .i (n11921), .o (n11922) );
  buffer buf_n11923( .i (n11922), .o (n11923) );
  buffer buf_n11924( .i (n11923), .o (n11924) );
  buffer buf_n11925( .i (n11924), .o (n11925) );
  buffer buf_n11926( .i (n11925), .o (n11926) );
  buffer buf_n11927( .i (n11926), .o (n11927) );
  buffer buf_n11928( .i (n11927), .o (n11928) );
  buffer buf_n11929( .i (n11928), .o (n11929) );
  buffer buf_n11930( .i (n11929), .o (n11930) );
  buffer buf_n11931( .i (n11930), .o (n11931) );
  buffer buf_n11932( .i (n11931), .o (n11932) );
  buffer buf_n11933( .i (n11932), .o (n11933) );
  buffer buf_n11934( .i (n11933), .o (n11934) );
  buffer buf_n11935( .i (n11934), .o (n11935) );
  buffer buf_n11936( .i (n11935), .o (n11936) );
  buffer buf_n11937( .i (n11936), .o (n11937) );
  buffer buf_n11938( .i (n11937), .o (n11938) );
  buffer buf_n11939( .i (n11938), .o (n11939) );
  buffer buf_n11940( .i (n11939), .o (n11940) );
  buffer buf_n11941( .i (n11940), .o (n11941) );
  buffer buf_n11942( .i (n11941), .o (n11942) );
  buffer buf_n11943( .i (n11942), .o (n11943) );
  buffer buf_n11944( .i (n11943), .o (n11944) );
  buffer buf_n11945( .i (n11944), .o (n11945) );
  buffer buf_n11946( .i (n11945), .o (n11946) );
  buffer buf_n11947( .i (n11946), .o (n11947) );
  buffer buf_n11948( .i (n11947), .o (n11948) );
  buffer buf_n11949( .i (n11948), .o (n11949) );
  buffer buf_n11950( .i (n11949), .o (n11950) );
  buffer buf_n11951( .i (n11950), .o (n11951) );
  buffer buf_n11952( .i (n11951), .o (n11952) );
  buffer buf_n11953( .i (n11952), .o (n11953) );
  buffer buf_n11954( .i (n11953), .o (n11954) );
  buffer buf_n4926( .i (n4925), .o (n4926) );
  buffer buf_n4927( .i (n4926), .o (n4927) );
  assign n11955 = ~n4906 & n4929 ;
  buffer buf_n11956( .i (n11955), .o (n11956) );
  assign n11957 = n4927 & n11956 ;
  assign n11958 = n4927 | n11956 ;
  assign n11959 = ~n11957 & n11958 ;
  buffer buf_n11960( .i (n11959), .o (n11960) );
  buffer buf_n11961( .i (n11960), .o (n11961) );
  buffer buf_n11962( .i (n11961), .o (n11962) );
  buffer buf_n11963( .i (n11962), .o (n11963) );
  buffer buf_n11964( .i (n11963), .o (n11964) );
  buffer buf_n11965( .i (n11964), .o (n11965) );
  buffer buf_n11966( .i (n11965), .o (n11966) );
  buffer buf_n11967( .i (n11966), .o (n11967) );
  buffer buf_n11968( .i (n11967), .o (n11968) );
  buffer buf_n11969( .i (n11968), .o (n11969) );
  buffer buf_n11970( .i (n11969), .o (n11970) );
  buffer buf_n11971( .i (n11970), .o (n11971) );
  buffer buf_n11972( .i (n11971), .o (n11972) );
  buffer buf_n11973( .i (n11972), .o (n11973) );
  buffer buf_n11974( .i (n11973), .o (n11974) );
  buffer buf_n11975( .i (n11974), .o (n11975) );
  buffer buf_n11976( .i (n11975), .o (n11976) );
  buffer buf_n11977( .i (n11976), .o (n11977) );
  buffer buf_n11978( .i (n11977), .o (n11978) );
  buffer buf_n11979( .i (n11978), .o (n11979) );
  buffer buf_n11980( .i (n11979), .o (n11980) );
  buffer buf_n11981( .i (n11980), .o (n11981) );
  buffer buf_n11982( .i (n11981), .o (n11982) );
  buffer buf_n11983( .i (n11982), .o (n11983) );
  buffer buf_n11984( .i (n11983), .o (n11984) );
  buffer buf_n11985( .i (n11984), .o (n11985) );
  buffer buf_n11986( .i (n11985), .o (n11986) );
  buffer buf_n11987( .i (n11986), .o (n11987) );
  buffer buf_n11988( .i (n11987), .o (n11988) );
  buffer buf_n11989( .i (n11988), .o (n11989) );
  buffer buf_n11990( .i (n11989), .o (n11990) );
  buffer buf_n11991( .i (n11990), .o (n11991) );
  buffer buf_n11992( .i (n11991), .o (n11992) );
  buffer buf_n11993( .i (n11992), .o (n11993) );
  buffer buf_n11994( .i (n11993), .o (n11994) );
  buffer buf_n11995( .i (n11994), .o (n11995) );
  buffer buf_n11996( .i (n11995), .o (n11996) );
  buffer buf_n11997( .i (n11996), .o (n11997) );
  buffer buf_n11998( .i (n11997), .o (n11998) );
  buffer buf_n11999( .i (n11998), .o (n11999) );
  buffer buf_n12000( .i (n11999), .o (n12000) );
  buffer buf_n12001( .i (n12000), .o (n12001) );
  buffer buf_n12002( .i (n12001), .o (n12002) );
  buffer buf_n12003( .i (n12002), .o (n12003) );
  buffer buf_n12004( .i (n12003), .o (n12004) );
  buffer buf_n12005( .i (n12004), .o (n12005) );
  buffer buf_n12006( .i (n12005), .o (n12006) );
  buffer buf_n12007( .i (n12006), .o (n12007) );
  buffer buf_n12008( .i (n12007), .o (n12008) );
  buffer buf_n12009( .i (n12008), .o (n12009) );
  buffer buf_n12010( .i (n12009), .o (n12010) );
  buffer buf_n12011( .i (n12010), .o (n12011) );
  buffer buf_n12012( .i (n12011), .o (n12012) );
  buffer buf_n12013( .i (n12012), .o (n12013) );
  buffer buf_n12014( .i (n12013), .o (n12014) );
  buffer buf_n12015( .i (n12014), .o (n12015) );
  buffer buf_n12016( .i (n12015), .o (n12016) );
  buffer buf_n12017( .i (n12016), .o (n12017) );
  buffer buf_n12018( .i (n12017), .o (n12018) );
  buffer buf_n12019( .i (n12018), .o (n12019) );
  buffer buf_n12020( .i (n12019), .o (n12020) );
  buffer buf_n12021( .i (n12020), .o (n12021) );
  buffer buf_n12022( .i (n12021), .o (n12022) );
  buffer buf_n12023( .i (n12022), .o (n12023) );
  buffer buf_n12024( .i (n12023), .o (n12024) );
  buffer buf_n12025( .i (n12024), .o (n12025) );
  buffer buf_n12026( .i (n12025), .o (n12026) );
  buffer buf_n12027( .i (n12026), .o (n12027) );
  buffer buf_n12028( .i (n12027), .o (n12028) );
  buffer buf_n12029( .i (n12028), .o (n12029) );
  buffer buf_n12030( .i (n12029), .o (n12030) );
  buffer buf_n12031( .i (n12030), .o (n12031) );
  buffer buf_n12032( .i (n12031), .o (n12032) );
  buffer buf_n12033( .i (n12032), .o (n12033) );
  buffer buf_n12034( .i (n12033), .o (n12034) );
  buffer buf_n12035( .i (n12034), .o (n12035) );
  buffer buf_n12036( .i (n12035), .o (n12036) );
  buffer buf_n12037( .i (n12036), .o (n12037) );
  buffer buf_n12038( .i (n12037), .o (n12038) );
  buffer buf_n12039( .i (n12038), .o (n12039) );
  buffer buf_n12040( .i (n12039), .o (n12040) );
  buffer buf_n12041( .i (n12040), .o (n12041) );
  buffer buf_n12042( .i (n12041), .o (n12042) );
  buffer buf_n12043( .i (n12042), .o (n12043) );
  buffer buf_n12044( .i (n12043), .o (n12044) );
  buffer buf_n12045( .i (n12044), .o (n12045) );
  buffer buf_n12046( .i (n12045), .o (n12046) );
  buffer buf_n12047( .i (n12046), .o (n12047) );
  buffer buf_n12048( .i (n12047), .o (n12048) );
  buffer buf_n12049( .i (n12048), .o (n12049) );
  buffer buf_n12050( .i (n12049), .o (n12050) );
  buffer buf_n12051( .i (n12050), .o (n12051) );
  buffer buf_n12052( .i (n12051), .o (n12052) );
  buffer buf_n12053( .i (n12052), .o (n12053) );
  buffer buf_n12054( .i (n12053), .o (n12054) );
  buffer buf_n12055( .i (n12054), .o (n12055) );
  buffer buf_n12056( .i (n12055), .o (n12056) );
  buffer buf_n12057( .i (n12056), .o (n12057) );
  buffer buf_n12058( .i (n12057), .o (n12058) );
  buffer buf_n12059( .i (n12058), .o (n12059) );
  buffer buf_n12060( .i (n12059), .o (n12060) );
  buffer buf_n12061( .i (n12060), .o (n12061) );
  buffer buf_n12062( .i (n12061), .o (n12062) );
  buffer buf_n12063( .i (n12062), .o (n12063) );
  buffer buf_n12064( .i (n12063), .o (n12064) );
  buffer buf_n12065( .i (n12064), .o (n12065) );
  buffer buf_n12066( .i (n12065), .o (n12066) );
  buffer buf_n12067( .i (n12066), .o (n12067) );
  buffer buf_n12068( .i (n12067), .o (n12068) );
  buffer buf_n12069( .i (n12068), .o (n12069) );
  buffer buf_n12070( .i (n12069), .o (n12070) );
  buffer buf_n12071( .i (n12070), .o (n12071) );
  buffer buf_n12072( .i (n12071), .o (n12072) );
  buffer buf_n12073( .i (n12072), .o (n12073) );
  buffer buf_n12074( .i (n12073), .o (n12074) );
  buffer buf_n12075( .i (n12074), .o (n12075) );
  buffer buf_n12076( .i (n12075), .o (n12076) );
  buffer buf_n12077( .i (n12076), .o (n12077) );
  buffer buf_n12078( .i (n12077), .o (n12078) );
  buffer buf_n12079( .i (n12078), .o (n12079) );
  buffer buf_n12080( .i (n12079), .o (n12080) );
  buffer buf_n12081( .i (n12080), .o (n12081) );
  buffer buf_n12082( .i (n12081), .o (n12082) );
  buffer buf_n12083( .i (n12082), .o (n12083) );
  buffer buf_n12084( .i (n12083), .o (n12084) );
  buffer buf_n12085( .i (n12084), .o (n12085) );
  buffer buf_n12086( .i (n12085), .o (n12086) );
  buffer buf_n12087( .i (n12086), .o (n12087) );
  buffer buf_n12088( .i (n12087), .o (n12088) );
  buffer buf_n12089( .i (n12088), .o (n12089) );
  buffer buf_n12090( .i (n12089), .o (n12090) );
  buffer buf_n12091( .i (n12090), .o (n12091) );
  buffer buf_n5440( .i (n5439), .o (n5440) );
  buffer buf_n5441( .i (n5440), .o (n5441) );
  assign n12092 = ~n5379 & n5382 ;
  buffer buf_n12093( .i (n12092), .o (n12093) );
  assign n12094 = n5441 & ~n12093 ;
  assign n12095 = ~n5441 & n12093 ;
  assign n12096 = n12094 | n12095 ;
  buffer buf_n12097( .i (n12096), .o (n12097) );
  assign n12167 = ~n5676 & n12097 ;
  buffer buf_n10760( .i (n10759), .o (n10760) );
  buffer buf_n12168( .i (n11509), .o (n12168) );
  assign n12169 = ~n10760 & n12168 ;
  buffer buf_n12170( .i (n11511), .o (n12170) );
  assign n12171 = ~n12169 & n12170 ;
  assign n12172 = n794 & n2829 ;
  buffer buf_n12173( .i (n12172), .o (n12173) );
  buffer buf_n12174( .i (n12173), .o (n12174) );
  assign n12175 = n11658 & ~n12174 ;
  buffer buf_n12176( .i (n10767), .o (n12176) );
  assign n12177 = n12175 | n12176 ;
  assign n12178 = n2830 & n10908 ;
  assign n12179 = n796 | n12178 ;
  assign n12180 = n10916 & n12173 ;
  assign n12181 = n12179 & ~n12180 ;
  assign n12182 = n11523 | n12181 ;
  assign n12183 = ~n12177 & n12182 ;
  buffer buf_n12184( .i (n12183), .o (n12184) );
  buffer buf_n12185( .i (n12184), .o (n12185) );
  assign n12186 = n11670 | n12185 ;
  buffer buf_n12187( .i (n12186), .o (n12187) );
  buffer buf_n12188( .i (n12187), .o (n12188) );
  buffer buf_n12189( .i (n12188), .o (n12189) );
  buffer buf_n12190( .i (n12189), .o (n12190) );
  buffer buf_n12191( .i (n12190), .o (n12191) );
  buffer buf_n12192( .i (n12191), .o (n12192) );
  buffer buf_n12193( .i (n12192), .o (n12193) );
  buffer buf_n12194( .i (n12193), .o (n12194) );
  buffer buf_n12195( .i (n12194), .o (n12195) );
  assign n12196 = n10748 & n11541 ;
  assign n12197 = n12195 | n12196 ;
  assign n12198 = n12171 & n12197 ;
  buffer buf_n12199( .i (n12198), .o (n12199) );
  buffer buf_n12200( .i (n12199), .o (n12200) );
  buffer buf_n12201( .i (n12200), .o (n12201) );
  buffer buf_n12202( .i (n12201), .o (n12202) );
  buffer buf_n12203( .i (n12202), .o (n12203) );
  buffer buf_n12204( .i (n12203), .o (n12204) );
  buffer buf_n12205( .i (n12204), .o (n12205) );
  buffer buf_n12206( .i (n12205), .o (n12206) );
  buffer buf_n12207( .i (n12206), .o (n12207) );
  buffer buf_n12208( .i (n12207), .o (n12208) );
  buffer buf_n12209( .i (n12208), .o (n12209) );
  buffer buf_n12210( .i (n12209), .o (n12210) );
  buffer buf_n12211( .i (n12210), .o (n12211) );
  buffer buf_n12212( .i (n12211), .o (n12212) );
  buffer buf_n12213( .i (n12212), .o (n12213) );
  buffer buf_n12214( .i (n12213), .o (n12214) );
  buffer buf_n12215( .i (n12214), .o (n12215) );
  buffer buf_n12216( .i (n12215), .o (n12216) );
  buffer buf_n12217( .i (n12216), .o (n12217) );
  buffer buf_n12218( .i (n12217), .o (n12218) );
  buffer buf_n12219( .i (n12218), .o (n12219) );
  buffer buf_n12220( .i (n12219), .o (n12220) );
  buffer buf_n12221( .i (n12220), .o (n12221) );
  buffer buf_n12222( .i (n12221), .o (n12222) );
  buffer buf_n12223( .i (n12222), .o (n12223) );
  buffer buf_n12224( .i (n12223), .o (n12224) );
  buffer buf_n12225( .i (n12224), .o (n12225) );
  buffer buf_n12226( .i (n12225), .o (n12226) );
  buffer buf_n12227( .i (n12226), .o (n12227) );
  buffer buf_n12228( .i (n12227), .o (n12228) );
  buffer buf_n12229( .i (n12228), .o (n12229) );
  buffer buf_n12230( .i (n12229), .o (n12230) );
  buffer buf_n12231( .i (n12230), .o (n12231) );
  buffer buf_n12232( .i (n12231), .o (n12232) );
  buffer buf_n12233( .i (n12232), .o (n12233) );
  buffer buf_n12234( .i (n12233), .o (n12234) );
  buffer buf_n12235( .i (n12234), .o (n12235) );
  buffer buf_n12236( .i (n12235), .o (n12236) );
  buffer buf_n12237( .i (n12236), .o (n12237) );
  buffer buf_n12238( .i (n12237), .o (n12238) );
  buffer buf_n12239( .i (n12238), .o (n12239) );
  buffer buf_n12240( .i (n12239), .o (n12240) );
  buffer buf_n12241( .i (n12240), .o (n12241) );
  buffer buf_n12242( .i (n12241), .o (n12242) );
  assign n12243 = n12167 | n12242 ;
  buffer buf_n12244( .i (n12243), .o (n12244) );
  buffer buf_n12245( .i (n12244), .o (n12245) );
  buffer buf_n12246( .i (n12245), .o (n12246) );
  buffer buf_n12247( .i (n12246), .o (n12247) );
  buffer buf_n12248( .i (n12247), .o (n12248) );
  buffer buf_n12249( .i (n12248), .o (n12249) );
  buffer buf_n12250( .i (n12249), .o (n12250) );
  buffer buf_n12251( .i (n12250), .o (n12251) );
  buffer buf_n12252( .i (n12251), .o (n12252) );
  buffer buf_n12253( .i (n12252), .o (n12253) );
  buffer buf_n12254( .i (n12253), .o (n12254) );
  buffer buf_n12255( .i (n12254), .o (n12255) );
  buffer buf_n12256( .i (n12255), .o (n12256) );
  buffer buf_n12257( .i (n12256), .o (n12257) );
  buffer buf_n12258( .i (n12257), .o (n12258) );
  buffer buf_n12259( .i (n12258), .o (n12259) );
  buffer buf_n12260( .i (n12259), .o (n12260) );
  buffer buf_n12261( .i (n12260), .o (n12261) );
  buffer buf_n12262( .i (n12261), .o (n12262) );
  buffer buf_n12263( .i (n12262), .o (n12263) );
  buffer buf_n12264( .i (n12263), .o (n12264) );
  buffer buf_n12265( .i (n12264), .o (n12265) );
  buffer buf_n12266( .i (n12265), .o (n12266) );
  buffer buf_n12267( .i (n12266), .o (n12267) );
  buffer buf_n12268( .i (n12267), .o (n12268) );
  buffer buf_n12269( .i (n12268), .o (n12269) );
  buffer buf_n12270( .i (n12269), .o (n12270) );
  buffer buf_n12271( .i (n12270), .o (n12271) );
  buffer buf_n12272( .i (n12271), .o (n12272) );
  buffer buf_n12273( .i (n12272), .o (n12273) );
  buffer buf_n12274( .i (n12273), .o (n12274) );
  buffer buf_n12275( .i (n12274), .o (n12275) );
  buffer buf_n12276( .i (n12275), .o (n12276) );
  buffer buf_n12277( .i (n12276), .o (n12277) );
  buffer buf_n12278( .i (n12277), .o (n12278) );
  buffer buf_n12279( .i (n12278), .o (n12279) );
  buffer buf_n12280( .i (n12279), .o (n12280) );
  buffer buf_n12281( .i (n12280), .o (n12281) );
  buffer buf_n12282( .i (n12281), .o (n12282) );
  buffer buf_n12283( .i (n12282), .o (n12283) );
  buffer buf_n12284( .i (n12283), .o (n12284) );
  buffer buf_n12285( .i (n12284), .o (n12285) );
  buffer buf_n12286( .i (n12285), .o (n12286) );
  buffer buf_n12287( .i (n12286), .o (n12287) );
  buffer buf_n12288( .i (n12287), .o (n12288) );
  buffer buf_n12289( .i (n12288), .o (n12289) );
  buffer buf_n12290( .i (n12289), .o (n12290) );
  buffer buf_n12291( .i (n12290), .o (n12291) );
  buffer buf_n12292( .i (n12291), .o (n12292) );
  buffer buf_n12293( .i (n12292), .o (n12293) );
  buffer buf_n12294( .i (n12293), .o (n12294) );
  buffer buf_n12295( .i (n12294), .o (n12295) );
  buffer buf_n12296( .i (n12295), .o (n12296) );
  buffer buf_n12297( .i (n12296), .o (n12297) );
  buffer buf_n12298( .i (n12297), .o (n12298) );
  buffer buf_n12299( .i (n12298), .o (n12299) );
  buffer buf_n12300( .i (n12299), .o (n12300) );
  buffer buf_n12301( .i (n12300), .o (n12301) );
  buffer buf_n12302( .i (n12301), .o (n12302) );
  buffer buf_n12303( .i (n12302), .o (n12303) );
  buffer buf_n12304( .i (n12303), .o (n12304) );
  buffer buf_n12305( .i (n12304), .o (n12305) );
  buffer buf_n12306( .i (n12305), .o (n12306) );
  buffer buf_n12307( .i (n12306), .o (n12307) );
  buffer buf_n12308( .i (n12307), .o (n12308) );
  buffer buf_n12309( .i (n12308), .o (n12309) );
  buffer buf_n12310( .i (n12309), .o (n12310) );
  buffer buf_n5741( .i (n5740), .o (n5741) );
  buffer buf_n5742( .i (n5741), .o (n5742) );
  buffer buf_n5743( .i (n5742), .o (n5743) );
  assign n12311 = n5743 | n8548 ;
  buffer buf_n5753( .i (n5752), .o (n5753) );
  buffer buf_n5754( .i (n5753), .o (n5754) );
  assign n12312 = n6092 & n8970 ;
  buffer buf_n4832( .i (n4831), .o (n4832) );
  buffer buf_n4833( .i (n4832), .o (n4833) );
  assign n12313 = n4833 & n6054 ;
  assign n12314 = ~n6052 & n8415 ;
  assign n12315 = n2189 | n6063 ;
  assign n12316 = n12314 & n12315 ;
  assign n12317 = n4832 & n6076 ;
  assign n12318 = n12316 & ~n12317 ;
  assign n12319 = n12313 | n12318 ;
  assign n12320 = ~n6086 & n12319 ;
  buffer buf_n12321( .i (n12320), .o (n12321) );
  buffer buf_n12322( .i (n12321), .o (n12322) );
  buffer buf_n12323( .i (n12322), .o (n12323) );
  assign n12324 = n5916 | n12323 ;
  buffer buf_n12325( .i (n12324), .o (n12325) );
  buffer buf_n12326( .i (n12325), .o (n12326) );
  assign n12327 = n12312 | n12326 ;
  assign n12328 = ~n5754 & n12327 ;
  buffer buf_n12329( .i (n12328), .o (n12329) );
  buffer buf_n12330( .i (n12329), .o (n12330) );
  buffer buf_n12331( .i (n12330), .o (n12331) );
  buffer buf_n12332( .i (n12331), .o (n12332) );
  buffer buf_n12333( .i (n12332), .o (n12333) );
  buffer buf_n12334( .i (n12333), .o (n12334) );
  buffer buf_n12335( .i (n12334), .o (n12335) );
  assign n12336 = ~n8934 & n11509 ;
  assign n12337 = n12335 & ~n12336 ;
  assign n12338 = n5631 & ~n12337 ;
  buffer buf_n12339( .i (n12338), .o (n12339) );
  buffer buf_n12340( .i (n12339), .o (n12340) );
  buffer buf_n12341( .i (n12340), .o (n12341) );
  buffer buf_n12342( .i (n12341), .o (n12342) );
  buffer buf_n12343( .i (n12342), .o (n12343) );
  buffer buf_n12344( .i (n12343), .o (n12344) );
  buffer buf_n12345( .i (n12344), .o (n12345) );
  buffer buf_n12346( .i (n12345), .o (n12346) );
  buffer buf_n12347( .i (n12346), .o (n12347) );
  buffer buf_n12348( .i (n12347), .o (n12348) );
  buffer buf_n12349( .i (n12348), .o (n12349) );
  buffer buf_n12350( .i (n12349), .o (n12350) );
  buffer buf_n12351( .i (n12350), .o (n12351) );
  buffer buf_n12352( .i (n12351), .o (n12352) );
  buffer buf_n12353( .i (n12352), .o (n12353) );
  buffer buf_n12354( .i (n12353), .o (n12354) );
  buffer buf_n12355( .i (n12354), .o (n12355) );
  buffer buf_n12356( .i (n12355), .o (n12356) );
  buffer buf_n12357( .i (n12356), .o (n12357) );
  buffer buf_n12358( .i (n12357), .o (n12358) );
  buffer buf_n12359( .i (n12358), .o (n12359) );
  buffer buf_n12360( .i (n12359), .o (n12360) );
  buffer buf_n12361( .i (n12360), .o (n12361) );
  buffer buf_n12362( .i (n12361), .o (n12362) );
  buffer buf_n12363( .i (n12362), .o (n12363) );
  buffer buf_n12364( .i (n12363), .o (n12364) );
  buffer buf_n12365( .i (n12364), .o (n12365) );
  buffer buf_n12366( .i (n12365), .o (n12366) );
  buffer buf_n12367( .i (n12366), .o (n12367) );
  buffer buf_n12368( .i (n12367), .o (n12368) );
  buffer buf_n12369( .i (n12368), .o (n12369) );
  buffer buf_n12370( .i (n12369), .o (n12370) );
  buffer buf_n12371( .i (n12370), .o (n12371) );
  buffer buf_n12372( .i (n12371), .o (n12372) );
  buffer buf_n12373( .i (n12372), .o (n12373) );
  buffer buf_n12374( .i (n12373), .o (n12374) );
  buffer buf_n12375( .i (n12374), .o (n12375) );
  buffer buf_n12376( .i (n12375), .o (n12376) );
  buffer buf_n12377( .i (n12376), .o (n12377) );
  buffer buf_n12378( .i (n12377), .o (n12378) );
  buffer buf_n12379( .i (n12378), .o (n12379) );
  buffer buf_n12380( .i (n12379), .o (n12380) );
  buffer buf_n12381( .i (n12380), .o (n12381) );
  buffer buf_n12382( .i (n12381), .o (n12382) );
  buffer buf_n12383( .i (n12382), .o (n12383) );
  buffer buf_n12384( .i (n12383), .o (n12384) );
  buffer buf_n12385( .i (n12384), .o (n12385) );
  buffer buf_n12386( .i (n12385), .o (n12386) );
  buffer buf_n12387( .i (n12386), .o (n12387) );
  buffer buf_n12388( .i (n12387), .o (n12388) );
  buffer buf_n12389( .i (n12388), .o (n12389) );
  buffer buf_n12390( .i (n12389), .o (n12390) );
  buffer buf_n12391( .i (n12390), .o (n12391) );
  buffer buf_n12392( .i (n12391), .o (n12392) );
  buffer buf_n12393( .i (n12392), .o (n12393) );
  buffer buf_n12394( .i (n12393), .o (n12394) );
  buffer buf_n12395( .i (n12394), .o (n12395) );
  buffer buf_n12396( .i (n12395), .o (n12396) );
  buffer buf_n12397( .i (n12396), .o (n12397) );
  buffer buf_n12398( .i (n12397), .o (n12398) );
  buffer buf_n12399( .i (n12398), .o (n12399) );
  buffer buf_n12400( .i (n12399), .o (n12400) );
  buffer buf_n12401( .i (n12400), .o (n12401) );
  buffer buf_n12402( .i (n12401), .o (n12402) );
  buffer buf_n12403( .i (n12402), .o (n12403) );
  buffer buf_n12404( .i (n12403), .o (n12404) );
  buffer buf_n12405( .i (n12404), .o (n12405) );
  buffer buf_n12406( .i (n12405), .o (n12406) );
  buffer buf_n12407( .i (n12406), .o (n12407) );
  buffer buf_n12408( .i (n12407), .o (n12408) );
  buffer buf_n12409( .i (n12408), .o (n12409) );
  buffer buf_n12410( .i (n12409), .o (n12410) );
  buffer buf_n12411( .i (n12410), .o (n12411) );
  buffer buf_n12412( .i (n12411), .o (n12412) );
  buffer buf_n12413( .i (n12412), .o (n12413) );
  buffer buf_n12414( .i (n12413), .o (n12414) );
  buffer buf_n12415( .i (n12414), .o (n12415) );
  buffer buf_n12416( .i (n12415), .o (n12416) );
  buffer buf_n12417( .i (n12416), .o (n12417) );
  buffer buf_n12418( .i (n12417), .o (n12418) );
  buffer buf_n12419( .i (n12418), .o (n12419) );
  buffer buf_n12420( .i (n12419), .o (n12420) );
  buffer buf_n12421( .i (n12420), .o (n12421) );
  buffer buf_n12422( .i (n12421), .o (n12422) );
  buffer buf_n12423( .i (n12422), .o (n12423) );
  buffer buf_n12424( .i (n12423), .o (n12424) );
  buffer buf_n12425( .i (n12424), .o (n12425) );
  buffer buf_n12426( .i (n12425), .o (n12426) );
  buffer buf_n12427( .i (n12426), .o (n12427) );
  buffer buf_n12428( .i (n12427), .o (n12428) );
  buffer buf_n12429( .i (n12428), .o (n12429) );
  buffer buf_n12430( .i (n12429), .o (n12430) );
  buffer buf_n12431( .i (n12430), .o (n12431) );
  buffer buf_n12432( .i (n12431), .o (n12432) );
  buffer buf_n12433( .i (n12432), .o (n12433) );
  buffer buf_n12434( .i (n12433), .o (n12434) );
  buffer buf_n12435( .i (n12434), .o (n12435) );
  buffer buf_n12436( .i (n12435), .o (n12436) );
  buffer buf_n12437( .i (n12436), .o (n12437) );
  buffer buf_n12438( .i (n12437), .o (n12438) );
  buffer buf_n12439( .i (n12438), .o (n12439) );
  buffer buf_n12440( .i (n12439), .o (n12440) );
  buffer buf_n12441( .i (n12440), .o (n12441) );
  buffer buf_n12442( .i (n12441), .o (n12442) );
  buffer buf_n12443( .i (n12442), .o (n12443) );
  buffer buf_n12444( .i (n12443), .o (n12444) );
  buffer buf_n12445( .i (n12444), .o (n12445) );
  buffer buf_n12446( .i (n12445), .o (n12446) );
  buffer buf_n12447( .i (n12446), .o (n12447) );
  buffer buf_n12448( .i (n12447), .o (n12448) );
  buffer buf_n12449( .i (n12448), .o (n12449) );
  buffer buf_n5755( .i (n5754), .o (n5755) );
  buffer buf_n5756( .i (n5755), .o (n5756) );
  buffer buf_n5757( .i (n5756), .o (n5757) );
  buffer buf_n5758( .i (n5757), .o (n5758) );
  buffer buf_n5759( .i (n5758), .o (n5759) );
  buffer buf_n5760( .i (n5759), .o (n5760) );
  buffer buf_n5761( .i (n5760), .o (n5761) );
  buffer buf_n5762( .i (n5761), .o (n5762) );
  buffer buf_n5763( .i (n5762), .o (n5763) );
  buffer buf_n5764( .i (n5763), .o (n5764) );
  buffer buf_n5765( .i (n5764), .o (n5765) );
  buffer buf_n5766( .i (n5765), .o (n5766) );
  buffer buf_n5767( .i (n5766), .o (n5767) );
  buffer buf_n5768( .i (n5767), .o (n5768) );
  buffer buf_n5769( .i (n5768), .o (n5769) );
  buffer buf_n5770( .i (n5769), .o (n5770) );
  buffer buf_n5771( .i (n5770), .o (n5771) );
  buffer buf_n5772( .i (n5771), .o (n5772) );
  buffer buf_n5773( .i (n5772), .o (n5773) );
  buffer buf_n5774( .i (n5773), .o (n5774) );
  buffer buf_n5775( .i (n5774), .o (n5775) );
  buffer buf_n5776( .i (n5775), .o (n5776) );
  buffer buf_n5777( .i (n5776), .o (n5777) );
  buffer buf_n5778( .i (n5777), .o (n5778) );
  buffer buf_n5779( .i (n5778), .o (n5779) );
  buffer buf_n5780( .i (n5779), .o (n5780) );
  buffer buf_n5781( .i (n5780), .o (n5781) );
  buffer buf_n5782( .i (n5781), .o (n5782) );
  buffer buf_n5783( .i (n5782), .o (n5783) );
  buffer buf_n5784( .i (n5783), .o (n5784) );
  buffer buf_n5785( .i (n5784), .o (n5785) );
  buffer buf_n5786( .i (n5785), .o (n5786) );
  buffer buf_n5787( .i (n5786), .o (n5787) );
  buffer buf_n5788( .i (n5787), .o (n5788) );
  buffer buf_n5789( .i (n5788), .o (n5789) );
  buffer buf_n5790( .i (n5789), .o (n5790) );
  buffer buf_n5791( .i (n5790), .o (n5791) );
  buffer buf_n5792( .i (n5791), .o (n5792) );
  buffer buf_n5793( .i (n5792), .o (n5793) );
  buffer buf_n5794( .i (n5793), .o (n5794) );
  buffer buf_n5795( .i (n5794), .o (n5795) );
  buffer buf_n5796( .i (n5795), .o (n5796) );
  buffer buf_n5797( .i (n5796), .o (n5797) );
  buffer buf_n5798( .i (n5797), .o (n5798) );
  buffer buf_n5799( .i (n5798), .o (n5799) );
  buffer buf_n5800( .i (n5799), .o (n5800) );
  buffer buf_n5801( .i (n5800), .o (n5801) );
  buffer buf_n5802( .i (n5801), .o (n5802) );
  buffer buf_n5803( .i (n5802), .o (n5803) );
  buffer buf_n5804( .i (n5803), .o (n5804) );
  buffer buf_n5805( .i (n5804), .o (n5805) );
  buffer buf_n5806( .i (n5805), .o (n5806) );
  buffer buf_n5807( .i (n5806), .o (n5807) );
  buffer buf_n5808( .i (n5807), .o (n5808) );
  buffer buf_n5809( .i (n5808), .o (n5809) );
  buffer buf_n5810( .i (n5809), .o (n5810) );
  buffer buf_n5811( .i (n5810), .o (n5811) );
  buffer buf_n5812( .i (n5811), .o (n5812) );
  buffer buf_n5813( .i (n5812), .o (n5813) );
  buffer buf_n5814( .i (n5813), .o (n5814) );
  buffer buf_n5815( .i (n5814), .o (n5815) );
  buffer buf_n5816( .i (n5815), .o (n5816) );
  buffer buf_n5817( .i (n5816), .o (n5817) );
  buffer buf_n5818( .i (n5817), .o (n5818) );
  buffer buf_n5819( .i (n5818), .o (n5819) );
  buffer buf_n5820( .i (n5819), .o (n5820) );
  buffer buf_n5821( .i (n5820), .o (n5821) );
  buffer buf_n5822( .i (n5821), .o (n5822) );
  buffer buf_n5823( .i (n5822), .o (n5823) );
  buffer buf_n5824( .i (n5823), .o (n5824) );
  buffer buf_n5825( .i (n5824), .o (n5825) );
  buffer buf_n5826( .i (n5825), .o (n5826) );
  buffer buf_n5827( .i (n5826), .o (n5827) );
  buffer buf_n5828( .i (n5827), .o (n5828) );
  buffer buf_n5829( .i (n5828), .o (n5829) );
  buffer buf_n5830( .i (n5829), .o (n5830) );
  buffer buf_n5831( .i (n5830), .o (n5831) );
  buffer buf_n5832( .i (n5831), .o (n5832) );
  buffer buf_n5833( .i (n5832), .o (n5833) );
  buffer buf_n5834( .i (n5833), .o (n5834) );
  buffer buf_n5835( .i (n5834), .o (n5835) );
  buffer buf_n5836( .i (n5835), .o (n5836) );
  buffer buf_n5837( .i (n5836), .o (n5837) );
  buffer buf_n5838( .i (n5837), .o (n5838) );
  buffer buf_n5839( .i (n5838), .o (n5839) );
  buffer buf_n5840( .i (n5839), .o (n5840) );
  buffer buf_n5841( .i (n5840), .o (n5841) );
  buffer buf_n5842( .i (n5841), .o (n5842) );
  buffer buf_n5843( .i (n5842), .o (n5843) );
  buffer buf_n5844( .i (n5843), .o (n5844) );
  buffer buf_n5845( .i (n5844), .o (n5845) );
  buffer buf_n5846( .i (n5845), .o (n5846) );
  buffer buf_n5847( .i (n5846), .o (n5847) );
  buffer buf_n5848( .i (n5847), .o (n5848) );
  buffer buf_n5849( .i (n5848), .o (n5849) );
  buffer buf_n5850( .i (n5849), .o (n5850) );
  buffer buf_n5851( .i (n5850), .o (n5851) );
  buffer buf_n5852( .i (n5851), .o (n5852) );
  buffer buf_n5853( .i (n5852), .o (n5853) );
  buffer buf_n5854( .i (n5853), .o (n5854) );
  buffer buf_n5855( .i (n5854), .o (n5855) );
  buffer buf_n5856( .i (n5855), .o (n5856) );
  buffer buf_n5857( .i (n5856), .o (n5857) );
  buffer buf_n5858( .i (n5857), .o (n5858) );
  buffer buf_n5859( .i (n5858), .o (n5859) );
  buffer buf_n5860( .i (n5859), .o (n5860) );
  buffer buf_n5861( .i (n5860), .o (n5861) );
  buffer buf_n5862( .i (n5861), .o (n5862) );
  buffer buf_n5863( .i (n5862), .o (n5863) );
  buffer buf_n5864( .i (n5863), .o (n5864) );
  buffer buf_n5865( .i (n5864), .o (n5865) );
  buffer buf_n5866( .i (n5865), .o (n5866) );
  buffer buf_n5867( .i (n5866), .o (n5867) );
  buffer buf_n5868( .i (n5867), .o (n5868) );
  buffer buf_n5869( .i (n5868), .o (n5869) );
  buffer buf_n5870( .i (n5869), .o (n5870) );
  buffer buf_n5871( .i (n5870), .o (n5871) );
  buffer buf_n5872( .i (n5871), .o (n5872) );
  buffer buf_n5873( .i (n5872), .o (n5873) );
  buffer buf_n5874( .i (n5873), .o (n5874) );
  buffer buf_n8942( .i (n8941), .o (n8942) );
  assign n12450 = n8939 | n8942 ;
  buffer buf_n12451( .i (n12450), .o (n12451) );
  buffer buf_n12452( .i (n12451), .o (n12452) );
  buffer buf_n12453( .i (n12452), .o (n12453) );
  buffer buf_n12454( .i (n12453), .o (n12454) );
  buffer buf_n12455( .i (n12454), .o (n12455) );
  buffer buf_n12456( .i (n12455), .o (n12456) );
  buffer buf_n12457( .i (n12456), .o (n12457) );
  buffer buf_n12458( .i (n12457), .o (n12458) );
  buffer buf_n12459( .i (n12458), .o (n12459) );
  buffer buf_n12460( .i (n12459), .o (n12460) );
  buffer buf_n12461( .i (n12460), .o (n12461) );
  buffer buf_n12462( .i (n12461), .o (n12462) );
  buffer buf_n12463( .i (n12462), .o (n12463) );
  buffer buf_n12464( .i (n12463), .o (n12464) );
  buffer buf_n12465( .i (n12464), .o (n12465) );
  buffer buf_n12466( .i (n12465), .o (n12466) );
  buffer buf_n12467( .i (n12466), .o (n12467) );
  buffer buf_n12468( .i (n12467), .o (n12468) );
  buffer buf_n12469( .i (n12468), .o (n12469) );
  buffer buf_n12470( .i (n12469), .o (n12470) );
  buffer buf_n12471( .i (n12470), .o (n12471) );
  buffer buf_n12472( .i (n12471), .o (n12472) );
  buffer buf_n12473( .i (n12472), .o (n12473) );
  buffer buf_n12474( .i (n12473), .o (n12474) );
  buffer buf_n12475( .i (n12474), .o (n12475) );
  buffer buf_n12476( .i (n12475), .o (n12476) );
  buffer buf_n12477( .i (n12476), .o (n12477) );
  buffer buf_n12478( .i (n12477), .o (n12478) );
  buffer buf_n12479( .i (n12478), .o (n12479) );
  buffer buf_n12480( .i (n12479), .o (n12480) );
  buffer buf_n12481( .i (n12480), .o (n12481) );
  buffer buf_n12482( .i (n12481), .o (n12482) );
  buffer buf_n12483( .i (n12482), .o (n12483) );
  buffer buf_n12484( .i (n12483), .o (n12484) );
  buffer buf_n12485( .i (n12484), .o (n12485) );
  buffer buf_n12486( .i (n12485), .o (n12486) );
  buffer buf_n12487( .i (n12486), .o (n12487) );
  buffer buf_n12488( .i (n12487), .o (n12488) );
  buffer buf_n12489( .i (n12488), .o (n12489) );
  buffer buf_n12490( .i (n12489), .o (n12490) );
  buffer buf_n12491( .i (n12490), .o (n12491) );
  buffer buf_n12492( .i (n12491), .o (n12492) );
  buffer buf_n12493( .i (n12492), .o (n12493) );
  buffer buf_n12494( .i (n12493), .o (n12494) );
  buffer buf_n12495( .i (n12494), .o (n12495) );
  buffer buf_n12496( .i (n12495), .o (n12496) );
  buffer buf_n12497( .i (n12496), .o (n12497) );
  buffer buf_n12498( .i (n12497), .o (n12498) );
  buffer buf_n12499( .i (n12498), .o (n12499) );
  buffer buf_n12500( .i (n12499), .o (n12500) );
  buffer buf_n12501( .i (n12500), .o (n12501) );
  buffer buf_n12502( .i (n12501), .o (n12502) );
  buffer buf_n12503( .i (n12502), .o (n12503) );
  buffer buf_n12504( .i (n12503), .o (n12504) );
  buffer buf_n12505( .i (n12504), .o (n12505) );
  buffer buf_n12506( .i (n12505), .o (n12506) );
  buffer buf_n12507( .i (n12506), .o (n12507) );
  buffer buf_n12508( .i (n12507), .o (n12508) );
  buffer buf_n12509( .i (n12508), .o (n12509) );
  buffer buf_n12510( .i (n12509), .o (n12510) );
  buffer buf_n12511( .i (n12510), .o (n12511) );
  buffer buf_n12512( .i (n12511), .o (n12512) );
  buffer buf_n12513( .i (n12512), .o (n12513) );
  buffer buf_n12514( .i (n12513), .o (n12514) );
  buffer buf_n12515( .i (n12514), .o (n12515) );
  buffer buf_n12516( .i (n12515), .o (n12516) );
  buffer buf_n12517( .i (n12516), .o (n12517) );
  buffer buf_n12518( .i (n12517), .o (n12518) );
  buffer buf_n12519( .i (n12518), .o (n12519) );
  buffer buf_n12520( .i (n12519), .o (n12520) );
  buffer buf_n12521( .i (n12520), .o (n12521) );
  buffer buf_n12522( .i (n12521), .o (n12522) );
  buffer buf_n12523( .i (n12522), .o (n12523) );
  buffer buf_n12524( .i (n12523), .o (n12524) );
  buffer buf_n12525( .i (n12524), .o (n12525) );
  buffer buf_n12526( .i (n12525), .o (n12526) );
  buffer buf_n12527( .i (n12526), .o (n12527) );
  buffer buf_n12528( .i (n12527), .o (n12528) );
  buffer buf_n12529( .i (n12528), .o (n12529) );
  buffer buf_n12530( .i (n12529), .o (n12530) );
  buffer buf_n12531( .i (n12530), .o (n12531) );
  buffer buf_n12532( .i (n12531), .o (n12532) );
  buffer buf_n12533( .i (n12532), .o (n12533) );
  buffer buf_n12534( .i (n12533), .o (n12534) );
  buffer buf_n12535( .i (n12534), .o (n12535) );
  buffer buf_n12536( .i (n12535), .o (n12536) );
  buffer buf_n12537( .i (n12536), .o (n12537) );
  buffer buf_n12538( .i (n12537), .o (n12538) );
  buffer buf_n12539( .i (n12538), .o (n12539) );
  buffer buf_n12540( .i (n12539), .o (n12540) );
  buffer buf_n12541( .i (n12540), .o (n12541) );
  buffer buf_n12542( .i (n12541), .o (n12542) );
  buffer buf_n12543( .i (n12542), .o (n12543) );
  buffer buf_n12544( .i (n12543), .o (n12544) );
  buffer buf_n12545( .i (n12544), .o (n12545) );
  buffer buf_n12546( .i (n12545), .o (n12546) );
  buffer buf_n12547( .i (n12546), .o (n12547) );
  buffer buf_n12548( .i (n12547), .o (n12548) );
  buffer buf_n12549( .i (n12548), .o (n12549) );
  buffer buf_n12550( .i (n12549), .o (n12550) );
  buffer buf_n12551( .i (n12550), .o (n12551) );
  buffer buf_n12552( .i (n12551), .o (n12552) );
  buffer buf_n12553( .i (n12552), .o (n12553) );
  buffer buf_n12554( .i (n12553), .o (n12554) );
  buffer buf_n12555( .i (n12554), .o (n12555) );
  buffer buf_n12556( .i (n12555), .o (n12556) );
  buffer buf_n12557( .i (n12556), .o (n12557) );
  buffer buf_n12558( .i (n12557), .o (n12558) );
  buffer buf_n12559( .i (n12558), .o (n12559) );
  buffer buf_n12560( .i (n12559), .o (n12560) );
  buffer buf_n12561( .i (n12560), .o (n12561) );
  buffer buf_n12562( .i (n12561), .o (n12562) );
  buffer buf_n12563( .i (n12562), .o (n12563) );
  buffer buf_n12564( .i (n12563), .o (n12564) );
  buffer buf_n12565( .i (n12564), .o (n12565) );
  buffer buf_n12566( .i (n12565), .o (n12566) );
  buffer buf_n12567( .i (n12566), .o (n12567) );
  buffer buf_n12568( .i (n12567), .o (n12568) );
  buffer buf_n12569( .i (n12568), .o (n12569) );
  buffer buf_n12570( .i (n12569), .o (n12570) );
  buffer buf_n12571( .i (n12570), .o (n12571) );
  buffer buf_n12572( .i (n12571), .o (n12572) );
  buffer buf_n12573( .i (n12572), .o (n12573) );
  assign n12574 = n8854 & ~n12573 ;
  buffer buf_n4009( .i (n4008), .o (n4009) );
  buffer buf_n4010( .i (n4009), .o (n4010) );
  buffer buf_n4011( .i (n4010), .o (n4011) );
  assign n12575 = n4011 & n5746 ;
  buffer buf_n12576( .i (n12575), .o (n12576) );
  assign n12577 = n8939 | n12576 ;
  assign n12578 = ~n8942 & n12576 ;
  assign n12579 = n12577 & ~n12578 ;
  buffer buf_n12580( .i (n12579), .o (n12580) );
  buffer buf_n12581( .i (n12580), .o (n12581) );
  buffer buf_n12582( .i (n12581), .o (n12582) );
  buffer buf_n12583( .i (n12582), .o (n12583) );
  buffer buf_n12584( .i (n12583), .o (n12584) );
  buffer buf_n12585( .i (n12584), .o (n12585) );
  buffer buf_n12586( .i (n12585), .o (n12586) );
  buffer buf_n12587( .i (n12586), .o (n12587) );
  buffer buf_n12588( .i (n12587), .o (n12588) );
  buffer buf_n12589( .i (n12588), .o (n12589) );
  buffer buf_n12590( .i (n12589), .o (n12590) );
  buffer buf_n12591( .i (n12590), .o (n12591) );
  buffer buf_n12592( .i (n12591), .o (n12592) );
  buffer buf_n12593( .i (n12592), .o (n12593) );
  buffer buf_n12594( .i (n12593), .o (n12594) );
  buffer buf_n12595( .i (n12594), .o (n12595) );
  buffer buf_n12596( .i (n12595), .o (n12596) );
  buffer buf_n12597( .i (n12596), .o (n12597) );
  buffer buf_n12598( .i (n12597), .o (n12598) );
  buffer buf_n12599( .i (n12598), .o (n12599) );
  buffer buf_n12600( .i (n12599), .o (n12600) );
  buffer buf_n12601( .i (n12600), .o (n12601) );
  buffer buf_n12602( .i (n12601), .o (n12602) );
  buffer buf_n12603( .i (n12602), .o (n12603) );
  buffer buf_n12604( .i (n12603), .o (n12604) );
  buffer buf_n12605( .i (n12604), .o (n12605) );
  buffer buf_n12606( .i (n12605), .o (n12606) );
  buffer buf_n12607( .i (n12606), .o (n12607) );
  buffer buf_n12608( .i (n12607), .o (n12608) );
  buffer buf_n12609( .i (n12608), .o (n12609) );
  buffer buf_n12610( .i (n12609), .o (n12610) );
  buffer buf_n12611( .i (n12610), .o (n12611) );
  buffer buf_n12612( .i (n12611), .o (n12612) );
  buffer buf_n12613( .i (n12612), .o (n12613) );
  buffer buf_n12614( .i (n12613), .o (n12614) );
  buffer buf_n12615( .i (n12614), .o (n12615) );
  buffer buf_n12616( .i (n12615), .o (n12616) );
  buffer buf_n12617( .i (n12616), .o (n12617) );
  buffer buf_n12618( .i (n12617), .o (n12618) );
  buffer buf_n12619( .i (n12618), .o (n12619) );
  buffer buf_n12620( .i (n12619), .o (n12620) );
  buffer buf_n12621( .i (n12620), .o (n12621) );
  buffer buf_n12622( .i (n12621), .o (n12622) );
  buffer buf_n12623( .i (n12622), .o (n12623) );
  buffer buf_n12624( .i (n12623), .o (n12624) );
  buffer buf_n12625( .i (n12624), .o (n12625) );
  buffer buf_n12626( .i (n12625), .o (n12626) );
  buffer buf_n12627( .i (n12626), .o (n12627) );
  buffer buf_n12628( .i (n12627), .o (n12628) );
  buffer buf_n12629( .i (n12628), .o (n12629) );
  buffer buf_n12630( .i (n12629), .o (n12630) );
  buffer buf_n12631( .i (n12630), .o (n12631) );
  buffer buf_n12632( .i (n12631), .o (n12632) );
  buffer buf_n12633( .i (n12632), .o (n12633) );
  buffer buf_n12634( .i (n12633), .o (n12634) );
  buffer buf_n12635( .i (n12634), .o (n12635) );
  buffer buf_n12636( .i (n12635), .o (n12636) );
  buffer buf_n12637( .i (n12636), .o (n12637) );
  buffer buf_n12638( .i (n12637), .o (n12638) );
  buffer buf_n12639( .i (n12638), .o (n12639) );
  buffer buf_n12640( .i (n12639), .o (n12640) );
  buffer buf_n12641( .i (n12640), .o (n12641) );
  buffer buf_n12642( .i (n12641), .o (n12642) );
  buffer buf_n12643( .i (n12642), .o (n12643) );
  buffer buf_n12644( .i (n12643), .o (n12644) );
  buffer buf_n12645( .i (n12644), .o (n12645) );
  buffer buf_n12646( .i (n12645), .o (n12646) );
  buffer buf_n12647( .i (n12646), .o (n12647) );
  buffer buf_n12648( .i (n12647), .o (n12648) );
  buffer buf_n12649( .i (n12648), .o (n12649) );
  buffer buf_n12650( .i (n12649), .o (n12650) );
  buffer buf_n12651( .i (n12650), .o (n12651) );
  buffer buf_n12652( .i (n12651), .o (n12652) );
  buffer buf_n12653( .i (n12652), .o (n12653) );
  buffer buf_n12654( .i (n12653), .o (n12654) );
  buffer buf_n12655( .i (n12654), .o (n12655) );
  buffer buf_n12656( .i (n12655), .o (n12656) );
  buffer buf_n12657( .i (n12656), .o (n12657) );
  buffer buf_n12658( .i (n12657), .o (n12658) );
  buffer buf_n12659( .i (n12658), .o (n12659) );
  buffer buf_n12660( .i (n12659), .o (n12660) );
  buffer buf_n12661( .i (n12660), .o (n12661) );
  buffer buf_n12662( .i (n12661), .o (n12662) );
  buffer buf_n12663( .i (n12662), .o (n12663) );
  buffer buf_n12664( .i (n12663), .o (n12664) );
  buffer buf_n12665( .i (n12664), .o (n12665) );
  buffer buf_n12666( .i (n12665), .o (n12666) );
  buffer buf_n12667( .i (n12666), .o (n12667) );
  buffer buf_n12668( .i (n12667), .o (n12668) );
  buffer buf_n12669( .i (n12668), .o (n12669) );
  buffer buf_n12670( .i (n12669), .o (n12670) );
  buffer buf_n12671( .i (n12670), .o (n12671) );
  buffer buf_n12672( .i (n12671), .o (n12672) );
  buffer buf_n12673( .i (n12672), .o (n12673) );
  buffer buf_n12674( .i (n12673), .o (n12674) );
  buffer buf_n12675( .i (n12674), .o (n12675) );
  buffer buf_n12676( .i (n12675), .o (n12676) );
  buffer buf_n12677( .i (n12676), .o (n12677) );
  buffer buf_n12678( .i (n12677), .o (n12678) );
  buffer buf_n12679( .i (n12678), .o (n12679) );
  buffer buf_n12680( .i (n12679), .o (n12680) );
  buffer buf_n12681( .i (n12680), .o (n12681) );
  buffer buf_n12682( .i (n12681), .o (n12682) );
  buffer buf_n12683( .i (n12682), .o (n12683) );
  buffer buf_n12684( .i (n12683), .o (n12684) );
  buffer buf_n12685( .i (n12684), .o (n12685) );
  buffer buf_n12686( .i (n12685), .o (n12686) );
  buffer buf_n12687( .i (n12686), .o (n12687) );
  buffer buf_n12688( .i (n12687), .o (n12688) );
  buffer buf_n12689( .i (n12688), .o (n12689) );
  buffer buf_n12690( .i (n12689), .o (n12690) );
  buffer buf_n12691( .i (n12690), .o (n12691) );
  buffer buf_n12692( .i (n12691), .o (n12692) );
  buffer buf_n12693( .i (n12692), .o (n12693) );
  buffer buf_n12694( .i (n12693), .o (n12694) );
  buffer buf_n12695( .i (n12694), .o (n12695) );
  buffer buf_n12696( .i (n12695), .o (n12696) );
  buffer buf_n12697( .i (n12696), .o (n12697) );
  buffer buf_n12698( .i (n12697), .o (n12698) );
  buffer buf_n12699( .i (n12698), .o (n12699) );
  buffer buf_n12700( .i (n12699), .o (n12700) );
  buffer buf_n12701( .i (n12700), .o (n12701) );
  buffer buf_n12702( .i (n12701), .o (n12702) );
  assign n12703 = n12574 | n12702 ;
  assign n12704 = n5874 & n12703 ;
  assign n12705 = n12449 & ~n12704 ;
  assign n12706 = n12311 & ~n12705 ;
  assign n12707 = n10239 & ~n10752 ;
  assign n12708 = n10270 | n12707 ;
  buffer buf_n12709( .i (n12708), .o (n12709) );
  buffer buf_n12710( .i (n131), .o (n12710) );
  buffer buf_n12711( .i (n12710), .o (n12711) );
  buffer buf_n12712( .i (n12711), .o (n12712) );
  assign n12713 = n12709 & ~n12712 ;
  buffer buf_n12714( .i (n5949), .o (n12714) );
  assign n12715 = n12713 | n12714 ;
  buffer buf_n12716( .i (n12715), .o (n12716) );
  buffer buf_n12717( .i (n6100), .o (n12717) );
  assign n12718 = n12716 & n12717 ;
  assign n12719 = n121 & n4049 ;
  buffer buf_n12720( .i (n12719), .o (n12720) );
  buffer buf_n12721( .i (n10915), .o (n12721) );
  assign n12722 = n12720 & n12721 ;
  buffer buf_n4050( .i (n4049), .o (n4050) );
  buffer buf_n4051( .i (n4050), .o (n4051) );
  buffer buf_n12723( .i (n10204), .o (n12723) );
  assign n12724 = n122 & n12723 ;
  assign n12725 = n4051 | n12724 ;
  assign n12726 = ~n12722 & n12725 ;
  assign n12727 = n11523 | n12726 ;
  assign n12728 = n11198 & ~n12720 ;
  buffer buf_n12729( .i (n12728), .o (n12729) );
  assign n12730 = n12176 | n12729 ;
  assign n12731 = n12727 & ~n12730 ;
  buffer buf_n12732( .i (n12731), .o (n12732) );
  buffer buf_n12733( .i (n12732), .o (n12733) );
  assign n12734 = n11670 | n12733 ;
  buffer buf_n12735( .i (n12734), .o (n12735) );
  buffer buf_n12736( .i (n12735), .o (n12736) );
  buffer buf_n12737( .i (n12736), .o (n12737) );
  buffer buf_n12738( .i (n12737), .o (n12738) );
  buffer buf_n12739( .i (n12738), .o (n12739) );
  buffer buf_n12740( .i (n12739), .o (n12740) );
  buffer buf_n12741( .i (n12740), .o (n12741) );
  buffer buf_n12742( .i (n12741), .o (n12742) );
  assign n12743 = n12718 | n12742 ;
  assign n12744 = n10260 | n10752 ;
  buffer buf_n12745( .i (n10240), .o (n12745) );
  assign n12746 = ~n10268 & n12745 ;
  assign n12747 = n12744 & ~n12746 ;
  buffer buf_n12748( .i (n12747), .o (n12748) );
  assign n12749 = n12712 & ~n12748 ;
  buffer buf_n12750( .i (n12745), .o (n12750) );
  assign n12751 = n10254 & n12750 ;
  assign n12752 = n8927 & ~n11683 ;
  buffer buf_n8877( .i (n8876), .o (n8877) );
  assign n12753 = n8877 & n11683 ;
  assign n12754 = n12752 | n12753 ;
  assign n12755 = ~n12750 & n12754 ;
  assign n12756 = n12751 | n12755 ;
  assign n12757 = n12712 | n12756 ;
  assign n12758 = ~n12749 & n12757 ;
  buffer buf_n12759( .i (n12758), .o (n12759) );
  assign n12760 = n11509 & ~n12759 ;
  assign n12761 = n11511 & ~n12760 ;
  assign n12762 = n12743 & n12761 ;
  buffer buf_n4882( .i (n4881), .o (n4882) );
  buffer buf_n4883( .i (n4882), .o (n4883) );
  assign n12763 = n4874 & ~n4885 ;
  buffer buf_n12764( .i (n12763), .o (n12764) );
  assign n12765 = n4883 & n12764 ;
  assign n12766 = n4883 | n12764 ;
  assign n12767 = ~n12765 & n12766 ;
  buffer buf_n12768( .i (n12767), .o (n12768) );
  buffer buf_n12769( .i (n12768), .o (n12769) );
  buffer buf_n12770( .i (n12769), .o (n12770) );
  buffer buf_n12771( .i (n12770), .o (n12771) );
  buffer buf_n12772( .i (n12771), .o (n12772) );
  buffer buf_n12773( .i (n12772), .o (n12773) );
  buffer buf_n12774( .i (n12773), .o (n12774) );
  buffer buf_n12775( .i (n12774), .o (n12775) );
  buffer buf_n12776( .i (n12775), .o (n12776) );
  buffer buf_n12777( .i (n12776), .o (n12777) );
  buffer buf_n12778( .i (n12777), .o (n12778) );
  buffer buf_n12779( .i (n12778), .o (n12779) );
  buffer buf_n12780( .i (n12779), .o (n12780) );
  buffer buf_n12781( .i (n12780), .o (n12781) );
  buffer buf_n12782( .i (n12781), .o (n12782) );
  buffer buf_n12783( .i (n12782), .o (n12783) );
  buffer buf_n12784( .i (n12783), .o (n12784) );
  buffer buf_n12785( .i (n12784), .o (n12785) );
  buffer buf_n12786( .i (n12785), .o (n12786) );
  buffer buf_n12787( .i (n12786), .o (n12787) );
  buffer buf_n12788( .i (n12787), .o (n12788) );
  buffer buf_n12789( .i (n12788), .o (n12789) );
  buffer buf_n12790( .i (n12789), .o (n12790) );
  buffer buf_n12791( .i (n12790), .o (n12791) );
  buffer buf_n12792( .i (n12791), .o (n12792) );
  buffer buf_n12793( .i (n12792), .o (n12793) );
  buffer buf_n12794( .i (n12793), .o (n12794) );
  buffer buf_n12795( .i (n12794), .o (n12795) );
  assign n12910 = ~n5631 & n12795 ;
  assign n12911 = n12762 | n12910 ;
  buffer buf_n12912( .i (n12911), .o (n12912) );
  buffer buf_n12913( .i (n12912), .o (n12913) );
  buffer buf_n12914( .i (n12913), .o (n12914) );
  buffer buf_n12915( .i (n12914), .o (n12915) );
  buffer buf_n12916( .i (n12915), .o (n12916) );
  buffer buf_n12917( .i (n12916), .o (n12917) );
  buffer buf_n12918( .i (n12917), .o (n12918) );
  buffer buf_n12919( .i (n12918), .o (n12919) );
  buffer buf_n12920( .i (n12919), .o (n12920) );
  buffer buf_n12921( .i (n12920), .o (n12921) );
  buffer buf_n12922( .i (n12921), .o (n12922) );
  buffer buf_n12923( .i (n12922), .o (n12923) );
  buffer buf_n12924( .i (n12923), .o (n12924) );
  buffer buf_n12925( .i (n12924), .o (n12925) );
  buffer buf_n12926( .i (n12925), .o (n12926) );
  buffer buf_n12927( .i (n12926), .o (n12927) );
  buffer buf_n12928( .i (n12927), .o (n12928) );
  buffer buf_n12929( .i (n12928), .o (n12929) );
  buffer buf_n12930( .i (n12929), .o (n12930) );
  buffer buf_n12931( .i (n12930), .o (n12931) );
  buffer buf_n12932( .i (n12931), .o (n12932) );
  buffer buf_n12933( .i (n12932), .o (n12933) );
  buffer buf_n12934( .i (n12933), .o (n12934) );
  buffer buf_n12935( .i (n12934), .o (n12935) );
  buffer buf_n12936( .i (n12935), .o (n12936) );
  buffer buf_n12937( .i (n12936), .o (n12937) );
  buffer buf_n12938( .i (n12937), .o (n12938) );
  buffer buf_n12939( .i (n12938), .o (n12939) );
  buffer buf_n12940( .i (n12939), .o (n12940) );
  buffer buf_n12941( .i (n12940), .o (n12941) );
  buffer buf_n12942( .i (n12941), .o (n12942) );
  buffer buf_n12943( .i (n12942), .o (n12943) );
  buffer buf_n12944( .i (n12943), .o (n12944) );
  buffer buf_n12945( .i (n12944), .o (n12945) );
  buffer buf_n12946( .i (n12945), .o (n12946) );
  buffer buf_n12947( .i (n12946), .o (n12947) );
  buffer buf_n12948( .i (n12947), .o (n12948) );
  buffer buf_n12949( .i (n12948), .o (n12949) );
  buffer buf_n12950( .i (n12949), .o (n12950) );
  buffer buf_n12951( .i (n12950), .o (n12951) );
  buffer buf_n12952( .i (n12951), .o (n12952) );
  buffer buf_n12953( .i (n12952), .o (n12953) );
  buffer buf_n12954( .i (n12953), .o (n12954) );
  buffer buf_n12955( .i (n12954), .o (n12955) );
  buffer buf_n12956( .i (n12955), .o (n12956) );
  buffer buf_n12957( .i (n12956), .o (n12957) );
  buffer buf_n12958( .i (n12957), .o (n12958) );
  buffer buf_n12959( .i (n12958), .o (n12959) );
  buffer buf_n12960( .i (n12959), .o (n12960) );
  buffer buf_n12961( .i (n12960), .o (n12961) );
  buffer buf_n12962( .i (n12961), .o (n12962) );
  buffer buf_n12963( .i (n12962), .o (n12963) );
  buffer buf_n12964( .i (n12963), .o (n12964) );
  buffer buf_n12965( .i (n12964), .o (n12965) );
  buffer buf_n12966( .i (n12965), .o (n12966) );
  buffer buf_n12967( .i (n12966), .o (n12967) );
  buffer buf_n12968( .i (n12967), .o (n12968) );
  buffer buf_n12969( .i (n12968), .o (n12969) );
  buffer buf_n12970( .i (n12969), .o (n12970) );
  buffer buf_n12971( .i (n12970), .o (n12971) );
  buffer buf_n12972( .i (n12971), .o (n12972) );
  buffer buf_n12973( .i (n12972), .o (n12973) );
  buffer buf_n12974( .i (n12973), .o (n12974) );
  buffer buf_n12975( .i (n12974), .o (n12975) );
  buffer buf_n12976( .i (n12975), .o (n12976) );
  buffer buf_n12977( .i (n12976), .o (n12977) );
  buffer buf_n12978( .i (n12977), .o (n12978) );
  buffer buf_n12979( .i (n12978), .o (n12979) );
  buffer buf_n12980( .i (n12979), .o (n12980) );
  buffer buf_n12981( .i (n12980), .o (n12981) );
  buffer buf_n12982( .i (n12981), .o (n12982) );
  buffer buf_n12983( .i (n12982), .o (n12983) );
  buffer buf_n12984( .i (n12983), .o (n12984) );
  buffer buf_n12985( .i (n12984), .o (n12985) );
  buffer buf_n12986( .i (n12985), .o (n12986) );
  buffer buf_n12987( .i (n12986), .o (n12987) );
  buffer buf_n12988( .i (n12987), .o (n12988) );
  buffer buf_n12989( .i (n12988), .o (n12989) );
  buffer buf_n12990( .i (n12989), .o (n12990) );
  buffer buf_n12991( .i (n12990), .o (n12991) );
  buffer buf_n12992( .i (n12991), .o (n12992) );
  buffer buf_n12993( .i (n12992), .o (n12993) );
  buffer buf_n12994( .i (n12993), .o (n12994) );
  buffer buf_n12995( .i (n12994), .o (n12995) );
  buffer buf_n12996( .i (n12995), .o (n12996) );
  buffer buf_n12997( .i (n12996), .o (n12997) );
  buffer buf_n12998( .i (n12997), .o (n12998) );
  buffer buf_n12999( .i (n12998), .o (n12999) );
  buffer buf_n13000( .i (n12999), .o (n13000) );
  buffer buf_n13001( .i (n13000), .o (n13001) );
  buffer buf_n13002( .i (n13001), .o (n13002) );
  buffer buf_n13003( .i (n13002), .o (n13003) );
  buffer buf_n13004( .i (n13003), .o (n13004) );
  buffer buf_n13005( .i (n13004), .o (n13005) );
  buffer buf_n13006( .i (n13005), .o (n13006) );
  buffer buf_n13007( .i (n13006), .o (n13007) );
  buffer buf_n13008( .i (n13007), .o (n13008) );
  buffer buf_n13009( .i (n13008), .o (n13009) );
  buffer buf_n13010( .i (n13009), .o (n13010) );
  buffer buf_n13011( .i (n13010), .o (n13011) );
  buffer buf_n13012( .i (n13011), .o (n13012) );
  buffer buf_n13013( .i (n13012), .o (n13013) );
  buffer buf_n13014( .i (n13013), .o (n13014) );
  buffer buf_n13015( .i (n13014), .o (n13015) );
  buffer buf_n13016( .i (n13015), .o (n13016) );
  buffer buf_n13017( .i (n13016), .o (n13017) );
  buffer buf_n13018( .i (n13017), .o (n13018) );
  buffer buf_n13019( .i (n13018), .o (n13019) );
  buffer buf_n13020( .i (n13019), .o (n13020) );
  buffer buf_n13021( .i (n13020), .o (n13021) );
  buffer buf_n13022( .i (n13021), .o (n13022) );
  buffer buf_n13023( .i (n13022), .o (n13023) );
  buffer buf_n13024( .i (n5926), .o (n13024) );
  assign n13025 = ~n10248 & n13024 ;
  assign n13026 = n11511 & ~n13025 ;
  assign n13027 = n1680 & n3472 ;
  buffer buf_n13028( .i (n13027), .o (n13028) );
  buffer buf_n13029( .i (n13028), .o (n13029) );
  assign n13030 = n11658 & ~n13029 ;
  assign n13031 = n12176 | n13030 ;
  assign n13032 = n12721 & n13028 ;
  assign n13033 = n3473 & n12723 ;
  assign n13034 = n1682 | n13033 ;
  assign n13035 = ~n13032 & n13034 ;
  buffer buf_n13036( .i (n11198), .o (n13036) );
  buffer buf_n13037( .i (n13036), .o (n13037) );
  assign n13038 = n13035 | n13037 ;
  assign n13039 = ~n13031 & n13038 ;
  buffer buf_n13040( .i (n13039), .o (n13040) );
  buffer buf_n13041( .i (n13040), .o (n13041) );
  buffer buf_n13042( .i (n11669), .o (n13042) );
  assign n13043 = n13041 | n13042 ;
  buffer buf_n13044( .i (n13043), .o (n13044) );
  buffer buf_n13045( .i (n13044), .o (n13045) );
  buffer buf_n13046( .i (n13045), .o (n13046) );
  buffer buf_n13047( .i (n13046), .o (n13047) );
  buffer buf_n13048( .i (n13047), .o (n13048) );
  buffer buf_n13049( .i (n13048), .o (n13049) );
  buffer buf_n13050( .i (n13049), .o (n13050) );
  buffer buf_n13051( .i (n13050), .o (n13051) );
  assign n13052 = n10275 & n12717 ;
  assign n13053 = n13051 | n13052 ;
  assign n13054 = n13026 & n13053 ;
  buffer buf_n13055( .i (n13054), .o (n13055) );
  buffer buf_n13056( .i (n13055), .o (n13056) );
  buffer buf_n13057( .i (n13056), .o (n13057) );
  buffer buf_n13058( .i (n13057), .o (n13058) );
  buffer buf_n13059( .i (n13058), .o (n13059) );
  buffer buf_n13060( .i (n13059), .o (n13060) );
  buffer buf_n13061( .i (n13060), .o (n13061) );
  buffer buf_n13062( .i (n13061), .o (n13062) );
  buffer buf_n13063( .i (n13062), .o (n13063) );
  buffer buf_n13064( .i (n13063), .o (n13064) );
  buffer buf_n13065( .i (n13064), .o (n13065) );
  buffer buf_n13066( .i (n13065), .o (n13066) );
  buffer buf_n13067( .i (n13066), .o (n13067) );
  buffer buf_n13068( .i (n13067), .o (n13068) );
  buffer buf_n13069( .i (n13068), .o (n13069) );
  buffer buf_n13070( .i (n13069), .o (n13070) );
  buffer buf_n13071( .i (n13070), .o (n13071) );
  buffer buf_n13072( .i (n13071), .o (n13072) );
  buffer buf_n13073( .i (n13072), .o (n13073) );
  buffer buf_n13074( .i (n13073), .o (n13074) );
  buffer buf_n13075( .i (n13074), .o (n13075) );
  buffer buf_n13076( .i (n13075), .o (n13076) );
  buffer buf_n13077( .i (n13076), .o (n13077) );
  buffer buf_n13078( .i (n13077), .o (n13078) );
  buffer buf_n13079( .i (n13078), .o (n13079) );
  buffer buf_n13080( .i (n13079), .o (n13080) );
  buffer buf_n13081( .i (n13080), .o (n13081) );
  buffer buf_n13082( .i (n13081), .o (n13082) );
  buffer buf_n13083( .i (n13082), .o (n13083) );
  buffer buf_n13084( .i (n13083), .o (n13084) );
  buffer buf_n13085( .i (n13084), .o (n13085) );
  buffer buf_n13086( .i (n13085), .o (n13086) );
  buffer buf_n13087( .i (n13086), .o (n13087) );
  buffer buf_n13088( .i (n13087), .o (n13088) );
  buffer buf_n13089( .i (n13088), .o (n13089) );
  buffer buf_n13090( .i (n13089), .o (n13090) );
  buffer buf_n13091( .i (n13090), .o (n13091) );
  buffer buf_n13092( .i (n13091), .o (n13092) );
  buffer buf_n13093( .i (n13092), .o (n13093) );
  buffer buf_n13094( .i (n13093), .o (n13094) );
  buffer buf_n13095( .i (n13094), .o (n13095) );
  buffer buf_n13096( .i (n13095), .o (n13096) );
  buffer buf_n13097( .i (n13096), .o (n13097) );
  buffer buf_n13098( .i (n13097), .o (n13098) );
  buffer buf_n13099( .i (n13098), .o (n13099) );
  buffer buf_n13100( .i (n13099), .o (n13100) );
  buffer buf_n13101( .i (n13100), .o (n13101) );
  buffer buf_n13102( .i (n13101), .o (n13102) );
  buffer buf_n13103( .i (n13102), .o (n13103) );
  buffer buf_n13104( .i (n13103), .o (n13104) );
  buffer buf_n4709( .i (n4708), .o (n4709) );
  buffer buf_n4710( .i (n4709), .o (n4710) );
  assign n13105 = ~n5446 & n5449 ;
  buffer buf_n13106( .i (n13105), .o (n13106) );
  assign n13107 = n4710 & ~n13106 ;
  assign n13108 = ~n4710 & n13106 ;
  assign n13109 = n13107 | n13108 ;
  buffer buf_n13110( .i (n13109), .o (n13110) );
  assign n13175 = ~n5681 & n13110 ;
  assign n13176 = n13104 | n13175 ;
  buffer buf_n13177( .i (n13176), .o (n13177) );
  buffer buf_n13178( .i (n13177), .o (n13178) );
  buffer buf_n13179( .i (n13178), .o (n13179) );
  buffer buf_n13180( .i (n13179), .o (n13180) );
  buffer buf_n13181( .i (n13180), .o (n13181) );
  buffer buf_n13182( .i (n13181), .o (n13182) );
  buffer buf_n13183( .i (n13182), .o (n13183) );
  buffer buf_n13184( .i (n13183), .o (n13184) );
  buffer buf_n13185( .i (n13184), .o (n13185) );
  buffer buf_n13186( .i (n13185), .o (n13186) );
  buffer buf_n13187( .i (n13186), .o (n13187) );
  buffer buf_n13188( .i (n13187), .o (n13188) );
  buffer buf_n13189( .i (n13188), .o (n13189) );
  buffer buf_n13190( .i (n13189), .o (n13190) );
  buffer buf_n13191( .i (n13190), .o (n13191) );
  buffer buf_n13192( .i (n13191), .o (n13192) );
  buffer buf_n13193( .i (n13192), .o (n13193) );
  buffer buf_n13194( .i (n13193), .o (n13194) );
  buffer buf_n13195( .i (n13194), .o (n13195) );
  buffer buf_n13196( .i (n13195), .o (n13196) );
  buffer buf_n13197( .i (n13196), .o (n13197) );
  buffer buf_n13198( .i (n13197), .o (n13198) );
  buffer buf_n13199( .i (n13198), .o (n13199) );
  buffer buf_n13200( .i (n13199), .o (n13200) );
  buffer buf_n13201( .i (n13200), .o (n13201) );
  buffer buf_n13202( .i (n13201), .o (n13202) );
  buffer buf_n13203( .i (n13202), .o (n13203) );
  buffer buf_n13204( .i (n13203), .o (n13204) );
  buffer buf_n13205( .i (n13204), .o (n13205) );
  buffer buf_n13206( .i (n13205), .o (n13206) );
  buffer buf_n13207( .i (n13206), .o (n13207) );
  buffer buf_n13208( .i (n13207), .o (n13208) );
  buffer buf_n13209( .i (n13208), .o (n13209) );
  buffer buf_n13210( .i (n13209), .o (n13210) );
  buffer buf_n13211( .i (n13210), .o (n13211) );
  buffer buf_n13212( .i (n13211), .o (n13212) );
  buffer buf_n13213( .i (n13212), .o (n13213) );
  buffer buf_n13214( .i (n13213), .o (n13214) );
  buffer buf_n13215( .i (n13214), .o (n13215) );
  buffer buf_n13216( .i (n13215), .o (n13216) );
  buffer buf_n13217( .i (n13216), .o (n13217) );
  buffer buf_n13218( .i (n13217), .o (n13218) );
  buffer buf_n13219( .i (n13218), .o (n13219) );
  buffer buf_n13220( .i (n13219), .o (n13220) );
  buffer buf_n13221( .i (n13220), .o (n13221) );
  buffer buf_n13222( .i (n13221), .o (n13222) );
  buffer buf_n13223( .i (n13222), .o (n13223) );
  buffer buf_n13224( .i (n13223), .o (n13224) );
  buffer buf_n13225( .i (n13224), .o (n13225) );
  buffer buf_n13226( .i (n13225), .o (n13226) );
  buffer buf_n13227( .i (n13226), .o (n13227) );
  buffer buf_n13228( .i (n13227), .o (n13228) );
  buffer buf_n13229( .i (n13228), .o (n13229) );
  buffer buf_n13230( .i (n13229), .o (n13230) );
  buffer buf_n13231( .i (n13230), .o (n13231) );
  buffer buf_n13232( .i (n13231), .o (n13232) );
  buffer buf_n13233( .i (n13232), .o (n13233) );
  buffer buf_n13234( .i (n13233), .o (n13234) );
  buffer buf_n13235( .i (n13234), .o (n13235) );
  buffer buf_n13236( .i (n13235), .o (n13236) );
  buffer buf_n13237( .i (n13236), .o (n13237) );
  buffer buf_n13238( .i (n13237), .o (n13238) );
  buffer buf_n13111( .i (n13110), .o (n13111) );
  buffer buf_n13112( .i (n13111), .o (n13112) );
  buffer buf_n13113( .i (n13112), .o (n13113) );
  buffer buf_n13114( .i (n13113), .o (n13114) );
  buffer buf_n13115( .i (n13114), .o (n13115) );
  buffer buf_n13116( .i (n13115), .o (n13116) );
  buffer buf_n13117( .i (n13116), .o (n13117) );
  buffer buf_n13118( .i (n13117), .o (n13118) );
  buffer buf_n13119( .i (n13118), .o (n13119) );
  buffer buf_n13120( .i (n13119), .o (n13120) );
  buffer buf_n13121( .i (n13120), .o (n13121) );
  buffer buf_n13122( .i (n13121), .o (n13122) );
  buffer buf_n13123( .i (n13122), .o (n13123) );
  buffer buf_n13124( .i (n13123), .o (n13124) );
  buffer buf_n13125( .i (n13124), .o (n13125) );
  buffer buf_n13126( .i (n13125), .o (n13126) );
  buffer buf_n13127( .i (n13126), .o (n13127) );
  buffer buf_n13128( .i (n13127), .o (n13128) );
  buffer buf_n13129( .i (n13128), .o (n13129) );
  buffer buf_n13130( .i (n13129), .o (n13130) );
  buffer buf_n13131( .i (n13130), .o (n13131) );
  buffer buf_n13132( .i (n13131), .o (n13132) );
  buffer buf_n13133( .i (n13132), .o (n13133) );
  buffer buf_n13134( .i (n13133), .o (n13134) );
  buffer buf_n13135( .i (n13134), .o (n13135) );
  buffer buf_n13136( .i (n13135), .o (n13136) );
  buffer buf_n13137( .i (n13136), .o (n13137) );
  buffer buf_n13138( .i (n13137), .o (n13138) );
  buffer buf_n13139( .i (n13138), .o (n13139) );
  buffer buf_n13140( .i (n13139), .o (n13140) );
  buffer buf_n13141( .i (n13140), .o (n13141) );
  buffer buf_n13142( .i (n13141), .o (n13142) );
  buffer buf_n13143( .i (n13142), .o (n13143) );
  buffer buf_n13144( .i (n13143), .o (n13144) );
  buffer buf_n13145( .i (n13144), .o (n13145) );
  buffer buf_n13146( .i (n13145), .o (n13146) );
  buffer buf_n13147( .i (n13146), .o (n13147) );
  buffer buf_n13148( .i (n13147), .o (n13148) );
  buffer buf_n13149( .i (n13148), .o (n13149) );
  buffer buf_n13150( .i (n13149), .o (n13150) );
  buffer buf_n13151( .i (n13150), .o (n13151) );
  buffer buf_n13152( .i (n13151), .o (n13152) );
  buffer buf_n13153( .i (n13152), .o (n13153) );
  buffer buf_n13154( .i (n13153), .o (n13154) );
  buffer buf_n13155( .i (n13154), .o (n13155) );
  buffer buf_n13156( .i (n13155), .o (n13156) );
  buffer buf_n13157( .i (n13156), .o (n13157) );
  buffer buf_n13158( .i (n13157), .o (n13158) );
  buffer buf_n13159( .i (n13158), .o (n13159) );
  buffer buf_n13160( .i (n13159), .o (n13160) );
  buffer buf_n13161( .i (n13160), .o (n13161) );
  buffer buf_n13162( .i (n13161), .o (n13162) );
  buffer buf_n13163( .i (n13162), .o (n13163) );
  buffer buf_n13164( .i (n13163), .o (n13164) );
  buffer buf_n13165( .i (n13164), .o (n13165) );
  buffer buf_n13166( .i (n13165), .o (n13166) );
  buffer buf_n13167( .i (n13166), .o (n13167) );
  buffer buf_n13168( .i (n13167), .o (n13168) );
  buffer buf_n13169( .i (n13168), .o (n13169) );
  buffer buf_n13170( .i (n13169), .o (n13170) );
  buffer buf_n13171( .i (n13170), .o (n13171) );
  buffer buf_n13172( .i (n13171), .o (n13172) );
  buffer buf_n13173( .i (n13172), .o (n13173) );
  buffer buf_n13174( .i (n13173), .o (n13174) );
  assign n13239 = ~n5701 & n8024 ;
  assign n13240 = n6573 & ~n12712 ;
  assign n13241 = n12714 | n13240 ;
  buffer buf_n13242( .i (n13241), .o (n13242) );
  assign n13243 = n13024 & ~n13242 ;
  buffer buf_n13244( .i (n5883), .o (n13244) );
  assign n13245 = ~n13243 & n13244 ;
  buffer buf_n13246( .i (n12711), .o (n13246) );
  assign n13247 = n6640 & n13246 ;
  assign n13248 = n8896 | n12750 ;
  buffer buf_n8676( .i (n8675), .o (n8676) );
  assign n13249 = ~n8676 & n12750 ;
  assign n13250 = n13248 & ~n13249 ;
  assign n13251 = ~n13246 & n13250 ;
  assign n13252 = n13247 | n13251 ;
  buffer buf_n13253( .i (n13252), .o (n13253) );
  assign n13254 = n12717 & n13253 ;
  assign n13255 = n1628 & n1971 ;
  buffer buf_n13256( .i (n13255), .o (n13256) );
  buffer buf_n13257( .i (n13256), .o (n13257) );
  assign n13258 = n13036 & ~n13257 ;
  assign n13259 = n12176 | n13258 ;
  assign n13260 = n12721 & n13256 ;
  assign n13261 = n1629 & n12723 ;
  assign n13262 = n1973 | n13261 ;
  assign n13263 = ~n13260 & n13262 ;
  assign n13264 = n13037 | n13263 ;
  assign n13265 = ~n13259 & n13264 ;
  buffer buf_n13266( .i (n13265), .o (n13266) );
  buffer buf_n13267( .i (n13266), .o (n13267) );
  assign n13268 = n13042 | n13267 ;
  buffer buf_n13269( .i (n13268), .o (n13269) );
  buffer buf_n13270( .i (n13269), .o (n13270) );
  buffer buf_n13271( .i (n13270), .o (n13271) );
  buffer buf_n13272( .i (n13271), .o (n13272) );
  buffer buf_n13273( .i (n13272), .o (n13273) );
  buffer buf_n13274( .i (n13273), .o (n13274) );
  buffer buf_n13275( .i (n13274), .o (n13275) );
  buffer buf_n13276( .i (n13275), .o (n13276) );
  assign n13277 = n13254 | n13276 ;
  assign n13278 = n13245 & n13277 ;
  buffer buf_n13279( .i (n13278), .o (n13279) );
  buffer buf_n13280( .i (n13279), .o (n13280) );
  buffer buf_n13281( .i (n13280), .o (n13281) );
  buffer buf_n13282( .i (n13281), .o (n13282) );
  buffer buf_n13283( .i (n13282), .o (n13283) );
  buffer buf_n13284( .i (n13283), .o (n13284) );
  buffer buf_n13285( .i (n13284), .o (n13285) );
  buffer buf_n13286( .i (n13285), .o (n13286) );
  buffer buf_n13287( .i (n13286), .o (n13287) );
  buffer buf_n13288( .i (n13287), .o (n13288) );
  buffer buf_n13289( .i (n13288), .o (n13289) );
  buffer buf_n13290( .i (n13289), .o (n13290) );
  buffer buf_n13291( .i (n13290), .o (n13291) );
  buffer buf_n13292( .i (n13291), .o (n13292) );
  buffer buf_n13293( .i (n13292), .o (n13293) );
  buffer buf_n13294( .i (n13293), .o (n13294) );
  buffer buf_n13295( .i (n13294), .o (n13295) );
  buffer buf_n13296( .i (n13295), .o (n13296) );
  buffer buf_n13297( .i (n13296), .o (n13297) );
  buffer buf_n13298( .i (n13297), .o (n13298) );
  buffer buf_n13299( .i (n13298), .o (n13299) );
  buffer buf_n13300( .i (n13299), .o (n13300) );
  buffer buf_n13301( .i (n13300), .o (n13301) );
  buffer buf_n13302( .i (n13301), .o (n13302) );
  buffer buf_n13303( .i (n13302), .o (n13303) );
  buffer buf_n13304( .i (n13303), .o (n13304) );
  buffer buf_n13305( .i (n13304), .o (n13305) );
  buffer buf_n13306( .i (n13305), .o (n13306) );
  buffer buf_n13307( .i (n13306), .o (n13307) );
  buffer buf_n13308( .i (n13307), .o (n13308) );
  buffer buf_n13309( .i (n13308), .o (n13309) );
  buffer buf_n13310( .i (n13309), .o (n13310) );
  buffer buf_n13311( .i (n13310), .o (n13311) );
  buffer buf_n13312( .i (n13311), .o (n13312) );
  buffer buf_n13313( .i (n13312), .o (n13313) );
  buffer buf_n13314( .i (n13313), .o (n13314) );
  buffer buf_n13315( .i (n13314), .o (n13315) );
  buffer buf_n13316( .i (n13315), .o (n13316) );
  buffer buf_n13317( .i (n13316), .o (n13317) );
  buffer buf_n13318( .i (n13317), .o (n13318) );
  buffer buf_n13319( .i (n13318), .o (n13319) );
  buffer buf_n13320( .i (n13319), .o (n13320) );
  buffer buf_n13321( .i (n13320), .o (n13321) );
  buffer buf_n13322( .i (n13321), .o (n13322) );
  buffer buf_n13323( .i (n13322), .o (n13323) );
  buffer buf_n13324( .i (n13323), .o (n13324) );
  buffer buf_n13325( .i (n13324), .o (n13325) );
  buffer buf_n13326( .i (n13325), .o (n13326) );
  buffer buf_n13327( .i (n13326), .o (n13327) );
  buffer buf_n13328( .i (n13327), .o (n13328) );
  buffer buf_n13329( .i (n13328), .o (n13329) );
  buffer buf_n13330( .i (n13329), .o (n13330) );
  buffer buf_n13331( .i (n13330), .o (n13331) );
  buffer buf_n13332( .i (n13331), .o (n13332) );
  buffer buf_n13333( .i (n13332), .o (n13333) );
  buffer buf_n13334( .i (n13333), .o (n13334) );
  buffer buf_n13335( .i (n13334), .o (n13335) );
  buffer buf_n13336( .i (n13335), .o (n13336) );
  buffer buf_n13337( .i (n13336), .o (n13337) );
  buffer buf_n13338( .i (n13337), .o (n13338) );
  buffer buf_n13339( .i (n13338), .o (n13339) );
  buffer buf_n13340( .i (n13339), .o (n13340) );
  buffer buf_n13341( .i (n13340), .o (n13341) );
  buffer buf_n13342( .i (n13341), .o (n13342) );
  buffer buf_n13343( .i (n13342), .o (n13343) );
  buffer buf_n13344( .i (n13343), .o (n13344) );
  buffer buf_n13345( .i (n13344), .o (n13345) );
  buffer buf_n13346( .i (n13345), .o (n13346) );
  buffer buf_n13347( .i (n13346), .o (n13347) );
  buffer buf_n13348( .i (n13347), .o (n13348) );
  assign n13349 = n13239 | n13348 ;
  buffer buf_n13350( .i (n13349), .o (n13350) );
  buffer buf_n13351( .i (n13350), .o (n13351) );
  buffer buf_n13352( .i (n13351), .o (n13352) );
  buffer buf_n13353( .i (n13352), .o (n13353) );
  buffer buf_n13354( .i (n13353), .o (n13354) );
  buffer buf_n13355( .i (n13354), .o (n13355) );
  buffer buf_n13356( .i (n13355), .o (n13356) );
  buffer buf_n13357( .i (n13356), .o (n13357) );
  buffer buf_n13358( .i (n13357), .o (n13358) );
  buffer buf_n13359( .i (n13358), .o (n13359) );
  buffer buf_n13360( .i (n13359), .o (n13360) );
  buffer buf_n13361( .i (n13360), .o (n13361) );
  buffer buf_n13362( .i (n13361), .o (n13362) );
  buffer buf_n13363( .i (n13362), .o (n13363) );
  buffer buf_n13364( .i (n13363), .o (n13364) );
  buffer buf_n13365( .i (n13364), .o (n13365) );
  buffer buf_n13366( .i (n13365), .o (n13366) );
  buffer buf_n13367( .i (n13366), .o (n13367) );
  buffer buf_n13368( .i (n13367), .o (n13368) );
  buffer buf_n13369( .i (n13368), .o (n13369) );
  buffer buf_n13370( .i (n13369), .o (n13370) );
  buffer buf_n13371( .i (n13370), .o (n13371) );
  buffer buf_n13372( .i (n13371), .o (n13372) );
  buffer buf_n13373( .i (n13372), .o (n13373) );
  buffer buf_n13374( .i (n13373), .o (n13374) );
  buffer buf_n13375( .i (n13374), .o (n13375) );
  buffer buf_n13376( .i (n13375), .o (n13376) );
  buffer buf_n13377( .i (n13376), .o (n13377) );
  buffer buf_n13378( .i (n13377), .o (n13378) );
  buffer buf_n13379( .i (n13378), .o (n13379) );
  buffer buf_n13380( .i (n13379), .o (n13380) );
  buffer buf_n13381( .i (n13380), .o (n13381) );
  buffer buf_n13382( .i (n13381), .o (n13382) );
  buffer buf_n13383( .i (n13382), .o (n13383) );
  buffer buf_n13384( .i (n13383), .o (n13384) );
  buffer buf_n13385( .i (n13384), .o (n13385) );
  buffer buf_n13386( .i (n13385), .o (n13386) );
  buffer buf_n13387( .i (n13386), .o (n13387) );
  buffer buf_n13388( .i (n13387), .o (n13388) );
  buffer buf_n13389( .i (n13388), .o (n13389) );
  buffer buf_n13390( .i (n13389), .o (n13390) );
  buffer buf_n13391( .i (n13390), .o (n13391) );
  buffer buf_n13392( .i (n5630), .o (n13392) );
  assign n13393 = n8299 & ~n13392 ;
  assign n13394 = n13024 & ~n13253 ;
  assign n13395 = n13244 & ~n13394 ;
  buffer buf_n13396( .i (n6054), .o (n13396) );
  assign n13397 = n1477 & ~n13396 ;
  buffer buf_n13398( .i (n13397), .o (n13398) );
  buffer buf_n2440( .i (n2439), .o (n2440) );
  buffer buf_n2441( .i (n2440), .o (n2441) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  buffer buf_n2443( .i (n2442), .o (n2443) );
  buffer buf_n2444( .i (n2443), .o (n2444) );
  buffer buf_n2445( .i (n2444), .o (n2445) );
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n2448( .i (n2447), .o (n2448) );
  buffer buf_n2449( .i (n2448), .o (n2449) );
  buffer buf_n2450( .i (n2449), .o (n2450) );
  buffer buf_n2451( .i (n2450), .o (n2451) );
  buffer buf_n2452( .i (n2451), .o (n2452) );
  buffer buf_n2453( .i (n2452), .o (n2453) );
  buffer buf_n2454( .i (n2453), .o (n2454) );
  buffer buf_n2455( .i (n2454), .o (n2455) );
  buffer buf_n13399( .i (n6065), .o (n13399) );
  assign n13400 = n1477 | n13399 ;
  assign n13401 = n2455 & n13400 ;
  assign n13402 = n13398 | n13401 ;
  buffer buf_n13403( .i (n13402), .o (n13403) );
  buffer buf_n13404( .i (n13403), .o (n13404) );
  assign n13405 = n2455 & n10915 ;
  assign n13406 = n13398 & n13405 ;
  buffer buf_n13407( .i (n13406), .o (n13407) );
  buffer buf_n13408( .i (n10767), .o (n13408) );
  assign n13409 = n13407 | n13408 ;
  assign n13410 = n13404 & ~n13409 ;
  buffer buf_n13411( .i (n13410), .o (n13411) );
  buffer buf_n13412( .i (n13411), .o (n13412) );
  assign n13413 = n13042 | n13412 ;
  buffer buf_n13414( .i (n13413), .o (n13414) );
  buffer buf_n13415( .i (n13414), .o (n13415) );
  buffer buf_n13416( .i (n13415), .o (n13416) );
  buffer buf_n13417( .i (n13416), .o (n13417) );
  buffer buf_n13418( .i (n13417), .o (n13418) );
  buffer buf_n13419( .i (n13418), .o (n13419) );
  buffer buf_n13420( .i (n13419), .o (n13420) );
  buffer buf_n13421( .i (n13420), .o (n13421) );
  assign n13422 = n12717 & n13242 ;
  assign n13423 = n13421 | n13422 ;
  assign n13424 = n13395 & n13423 ;
  assign n13425 = n13393 | n13424 ;
  buffer buf_n13426( .i (n13425), .o (n13426) );
  buffer buf_n13427( .i (n13426), .o (n13427) );
  buffer buf_n13428( .i (n13427), .o (n13428) );
  buffer buf_n13429( .i (n13428), .o (n13429) );
  buffer buf_n13430( .i (n13429), .o (n13430) );
  buffer buf_n13431( .i (n13430), .o (n13431) );
  buffer buf_n13432( .i (n13431), .o (n13432) );
  buffer buf_n13433( .i (n13432), .o (n13433) );
  buffer buf_n13434( .i (n13433), .o (n13434) );
  buffer buf_n13435( .i (n13434), .o (n13435) );
  buffer buf_n13436( .i (n13435), .o (n13436) );
  buffer buf_n13437( .i (n13436), .o (n13437) );
  buffer buf_n13438( .i (n13437), .o (n13438) );
  buffer buf_n13439( .i (n13438), .o (n13439) );
  buffer buf_n13440( .i (n13439), .o (n13440) );
  buffer buf_n13441( .i (n13440), .o (n13441) );
  buffer buf_n13442( .i (n13441), .o (n13442) );
  buffer buf_n13443( .i (n13442), .o (n13443) );
  buffer buf_n13444( .i (n13443), .o (n13444) );
  buffer buf_n13445( .i (n13444), .o (n13445) );
  buffer buf_n13446( .i (n13445), .o (n13446) );
  buffer buf_n13447( .i (n13446), .o (n13447) );
  buffer buf_n13448( .i (n13447), .o (n13448) );
  buffer buf_n13449( .i (n13448), .o (n13449) );
  buffer buf_n13450( .i (n13449), .o (n13450) );
  buffer buf_n13451( .i (n13450), .o (n13451) );
  buffer buf_n13452( .i (n13451), .o (n13452) );
  buffer buf_n13453( .i (n13452), .o (n13453) );
  buffer buf_n13454( .i (n13453), .o (n13454) );
  buffer buf_n13455( .i (n13454), .o (n13455) );
  buffer buf_n13456( .i (n13455), .o (n13456) );
  buffer buf_n13457( .i (n13456), .o (n13457) );
  buffer buf_n13458( .i (n13457), .o (n13458) );
  buffer buf_n13459( .i (n13458), .o (n13459) );
  buffer buf_n13460( .i (n13459), .o (n13460) );
  buffer buf_n13461( .i (n13460), .o (n13461) );
  buffer buf_n13462( .i (n13461), .o (n13462) );
  buffer buf_n13463( .i (n13462), .o (n13463) );
  buffer buf_n13464( .i (n13463), .o (n13464) );
  buffer buf_n13465( .i (n13464), .o (n13465) );
  buffer buf_n13466( .i (n13465), .o (n13466) );
  buffer buf_n13467( .i (n13466), .o (n13467) );
  buffer buf_n13468( .i (n13467), .o (n13468) );
  buffer buf_n13469( .i (n13468), .o (n13469) );
  buffer buf_n13470( .i (n13469), .o (n13470) );
  buffer buf_n13471( .i (n13470), .o (n13471) );
  buffer buf_n13472( .i (n13471), .o (n13472) );
  buffer buf_n13473( .i (n13472), .o (n13473) );
  buffer buf_n13474( .i (n13473), .o (n13474) );
  buffer buf_n13475( .i (n13474), .o (n13475) );
  buffer buf_n13476( .i (n13475), .o (n13476) );
  buffer buf_n13477( .i (n13476), .o (n13477) );
  buffer buf_n13478( .i (n13477), .o (n13478) );
  buffer buf_n13479( .i (n13478), .o (n13479) );
  buffer buf_n13480( .i (n13479), .o (n13480) );
  buffer buf_n13481( .i (n13480), .o (n13481) );
  buffer buf_n13482( .i (n13481), .o (n13482) );
  buffer buf_n13483( .i (n13482), .o (n13483) );
  buffer buf_n13484( .i (n13483), .o (n13484) );
  buffer buf_n13485( .i (n13484), .o (n13485) );
  buffer buf_n13486( .i (n13485), .o (n13486) );
  buffer buf_n13487( .i (n13486), .o (n13487) );
  buffer buf_n13488( .i (n13487), .o (n13488) );
  buffer buf_n13489( .i (n13488), .o (n13489) );
  buffer buf_n13490( .i (n13489), .o (n13490) );
  buffer buf_n13491( .i (n13490), .o (n13491) );
  buffer buf_n13492( .i (n13491), .o (n13492) );
  buffer buf_n13493( .i (n13492), .o (n13493) );
  buffer buf_n13494( .i (n13493), .o (n13494) );
  buffer buf_n13495( .i (n13494), .o (n13495) );
  buffer buf_n13496( .i (n13495), .o (n13496) );
  buffer buf_n13497( .i (n13496), .o (n13497) );
  buffer buf_n13498( .i (n13497), .o (n13498) );
  buffer buf_n13499( .i (n13498), .o (n13499) );
  buffer buf_n13500( .i (n13499), .o (n13500) );
  buffer buf_n13501( .i (n13500), .o (n13501) );
  buffer buf_n13502( .i (n13501), .o (n13502) );
  buffer buf_n13503( .i (n13502), .o (n13503) );
  buffer buf_n13504( .i (n13503), .o (n13504) );
  buffer buf_n13505( .i (n13504), .o (n13505) );
  buffer buf_n13506( .i (n13505), .o (n13506) );
  buffer buf_n13507( .i (n13506), .o (n13507) );
  buffer buf_n13508( .i (n13507), .o (n13508) );
  buffer buf_n13509( .i (n13508), .o (n13509) );
  buffer buf_n13510( .i (n13509), .o (n13510) );
  buffer buf_n13511( .i (n13510), .o (n13511) );
  buffer buf_n13512( .i (n13511), .o (n13512) );
  buffer buf_n13513( .i (n13512), .o (n13513) );
  buffer buf_n13514( .i (n13513), .o (n13514) );
  buffer buf_n13515( .i (n13514), .o (n13515) );
  buffer buf_n13516( .i (n13515), .o (n13516) );
  buffer buf_n13517( .i (n13516), .o (n13517) );
  buffer buf_n13518( .i (n13517), .o (n13518) );
  buffer buf_n13519( .i (n13518), .o (n13519) );
  buffer buf_n13520( .i (n13519), .o (n13520) );
  buffer buf_n13521( .i (n13520), .o (n13521) );
  buffer buf_n13522( .i (n13521), .o (n13522) );
  buffer buf_n13523( .i (n13522), .o (n13523) );
  buffer buf_n13524( .i (n13523), .o (n13524) );
  buffer buf_n13525( .i (n13524), .o (n13525) );
  buffer buf_n13526( .i (n13525), .o (n13526) );
  buffer buf_n13527( .i (n13526), .o (n13527) );
  buffer buf_n13528( .i (n13527), .o (n13528) );
  buffer buf_n13529( .i (n13528), .o (n13529) );
  buffer buf_n13530( .i (n13529), .o (n13530) );
  buffer buf_n13531( .i (n13530), .o (n13531) );
  buffer buf_n13532( .i (n13531), .o (n13532) );
  buffer buf_n13533( .i (n13532), .o (n13533) );
  buffer buf_n13534( .i (n13533), .o (n13534) );
  buffer buf_n13535( .i (n13534), .o (n13535) );
  buffer buf_n13536( .i (n13535), .o (n13536) );
  buffer buf_n13537( .i (n13536), .o (n13537) );
  buffer buf_n4647( .i (n4646), .o (n4647) );
  buffer buf_n4648( .i (n4647), .o (n4648) );
  assign n13538 = ~n5454 & n5457 ;
  buffer buf_n13539( .i (n13538), .o (n13539) );
  assign n13540 = n4648 & n13539 ;
  assign n13541 = n4648 | n13539 ;
  assign n13542 = ~n13540 & n13541 ;
  buffer buf_n13543( .i (n13542), .o (n13543) );
  buffer buf_n13544( .i (n13543), .o (n13544) );
  buffer buf_n13545( .i (n13544), .o (n13545) );
  buffer buf_n13546( .i (n13545), .o (n13546) );
  buffer buf_n13547( .i (n13546), .o (n13547) );
  buffer buf_n13548( .i (n13547), .o (n13548) );
  buffer buf_n13549( .i (n13548), .o (n13549) );
  buffer buf_n13550( .i (n13549), .o (n13550) );
  buffer buf_n13551( .i (n13550), .o (n13551) );
  buffer buf_n13552( .i (n13551), .o (n13552) );
  buffer buf_n13553( .i (n13552), .o (n13553) );
  buffer buf_n13554( .i (n13553), .o (n13554) );
  buffer buf_n13555( .i (n13554), .o (n13555) );
  buffer buf_n13556( .i (n13555), .o (n13556) );
  buffer buf_n13557( .i (n13556), .o (n13557) );
  buffer buf_n13558( .i (n13557), .o (n13558) );
  buffer buf_n13559( .i (n13558), .o (n13559) );
  buffer buf_n13560( .i (n13559), .o (n13560) );
  buffer buf_n13561( .i (n13560), .o (n13561) );
  buffer buf_n13562( .i (n13561), .o (n13562) );
  buffer buf_n13563( .i (n13562), .o (n13563) );
  buffer buf_n13564( .i (n13563), .o (n13564) );
  buffer buf_n13565( .i (n13564), .o (n13565) );
  buffer buf_n13566( .i (n13565), .o (n13566) );
  buffer buf_n13567( .i (n13566), .o (n13567) );
  buffer buf_n13568( .i (n13567), .o (n13568) );
  buffer buf_n13569( .i (n13568), .o (n13569) );
  buffer buf_n13570( .i (n13569), .o (n13570) );
  buffer buf_n13571( .i (n13570), .o (n13571) );
  buffer buf_n13572( .i (n13571), .o (n13572) );
  buffer buf_n13573( .i (n13572), .o (n13573) );
  buffer buf_n13574( .i (n13573), .o (n13574) );
  buffer buf_n13575( .i (n13574), .o (n13575) );
  buffer buf_n13576( .i (n13575), .o (n13576) );
  buffer buf_n13577( .i (n13576), .o (n13577) );
  buffer buf_n13578( .i (n13577), .o (n13578) );
  buffer buf_n13579( .i (n13578), .o (n13579) );
  buffer buf_n13580( .i (n13579), .o (n13580) );
  buffer buf_n13581( .i (n13580), .o (n13581) );
  buffer buf_n13582( .i (n13581), .o (n13582) );
  buffer buf_n13583( .i (n13582), .o (n13583) );
  buffer buf_n13584( .i (n13583), .o (n13584) );
  buffer buf_n13585( .i (n13584), .o (n13585) );
  buffer buf_n13586( .i (n13585), .o (n13586) );
  buffer buf_n13587( .i (n13586), .o (n13587) );
  buffer buf_n13588( .i (n13587), .o (n13588) );
  buffer buf_n13589( .i (n13588), .o (n13589) );
  buffer buf_n13590( .i (n13589), .o (n13590) );
  buffer buf_n13591( .i (n13590), .o (n13591) );
  buffer buf_n13592( .i (n13591), .o (n13592) );
  buffer buf_n13593( .i (n13592), .o (n13593) );
  buffer buf_n13594( .i (n13593), .o (n13594) );
  buffer buf_n13595( .i (n13594), .o (n13595) );
  buffer buf_n13596( .i (n13595), .o (n13596) );
  buffer buf_n13597( .i (n13596), .o (n13597) );
  buffer buf_n13598( .i (n13597), .o (n13598) );
  buffer buf_n13599( .i (n13598), .o (n13599) );
  buffer buf_n13600( .i (n13599), .o (n13600) );
  buffer buf_n13601( .i (n13600), .o (n13601) );
  buffer buf_n13602( .i (n13601), .o (n13602) );
  assign n13603 = n12748 & ~n13246 ;
  assign n13604 = n12714 | n13603 ;
  buffer buf_n13605( .i (n13604), .o (n13605) );
  assign n13606 = n13024 & ~n13605 ;
  assign n13607 = n13244 & ~n13606 ;
  assign n13608 = ~n12709 & n13246 ;
  assign n13609 = n6599 & ~n10735 ;
  assign n13610 = n6607 & n10735 ;
  assign n13611 = n13609 | n13610 ;
  buffer buf_n13612( .i (n13611), .o (n13612) );
  buffer buf_n13613( .i (n12745), .o (n13613) );
  assign n13614 = n13612 & ~n13613 ;
  assign n13615 = n10232 & n12745 ;
  assign n13616 = n12710 | n13615 ;
  assign n13617 = n13614 | n13616 ;
  buffer buf_n13618( .i (n13617), .o (n13618) );
  assign n13619 = ~n13608 & n13618 ;
  buffer buf_n13620( .i (n13619), .o (n13620) );
  buffer buf_n13621( .i (n6099), .o (n13621) );
  buffer buf_n13622( .i (n13621), .o (n13622) );
  assign n13623 = n13620 & n13622 ;
  assign n13624 = n2610 & n12723 ;
  assign n13625 = n616 | n13624 ;
  assign n13626 = n614 & n2609 ;
  buffer buf_n13627( .i (n13626), .o (n13627) );
  assign n13629 = n12721 & n13627 ;
  assign n13630 = n13625 & ~n13629 ;
  assign n13631 = n13037 | n13630 ;
  buffer buf_n13628( .i (n13627), .o (n13628) );
  assign n13632 = n13036 & ~n13628 ;
  assign n13633 = n13408 | n13632 ;
  assign n13634 = n13631 & ~n13633 ;
  buffer buf_n13635( .i (n13634), .o (n13635) );
  buffer buf_n13636( .i (n13635), .o (n13636) );
  assign n13637 = n13042 | n13636 ;
  buffer buf_n13638( .i (n13637), .o (n13638) );
  buffer buf_n13639( .i (n13638), .o (n13639) );
  buffer buf_n13640( .i (n13639), .o (n13640) );
  buffer buf_n13641( .i (n13640), .o (n13641) );
  buffer buf_n13642( .i (n13641), .o (n13642) );
  buffer buf_n13643( .i (n13642), .o (n13643) );
  buffer buf_n13644( .i (n13643), .o (n13644) );
  buffer buf_n13645( .i (n13644), .o (n13645) );
  assign n13646 = n13623 | n13645 ;
  assign n13647 = n13607 & n13646 ;
  buffer buf_n13648( .i (n13647), .o (n13648) );
  buffer buf_n13649( .i (n13648), .o (n13649) );
  buffer buf_n13650( .i (n13649), .o (n13650) );
  buffer buf_n13651( .i (n13650), .o (n13651) );
  buffer buf_n13652( .i (n13651), .o (n13652) );
  buffer buf_n13653( .i (n13652), .o (n13653) );
  buffer buf_n13654( .i (n13653), .o (n13654) );
  buffer buf_n13655( .i (n13654), .o (n13655) );
  buffer buf_n13656( .i (n13655), .o (n13656) );
  buffer buf_n13657( .i (n13656), .o (n13657) );
  buffer buf_n13658( .i (n13657), .o (n13658) );
  buffer buf_n13659( .i (n13658), .o (n13659) );
  buffer buf_n13660( .i (n13659), .o (n13660) );
  buffer buf_n13661( .i (n13660), .o (n13661) );
  buffer buf_n13662( .i (n13661), .o (n13662) );
  buffer buf_n13663( .i (n13662), .o (n13663) );
  buffer buf_n13664( .i (n13663), .o (n13664) );
  buffer buf_n13665( .i (n13664), .o (n13665) );
  buffer buf_n13666( .i (n13665), .o (n13666) );
  buffer buf_n13667( .i (n13666), .o (n13667) );
  buffer buf_n13668( .i (n13667), .o (n13668) );
  buffer buf_n13669( .i (n13668), .o (n13669) );
  buffer buf_n13670( .i (n13669), .o (n13670) );
  buffer buf_n13671( .i (n13670), .o (n13671) );
  buffer buf_n13672( .i (n13671), .o (n13672) );
  buffer buf_n13673( .i (n13672), .o (n13673) );
  buffer buf_n13674( .i (n13673), .o (n13674) );
  buffer buf_n13675( .i (n13674), .o (n13675) );
  buffer buf_n13676( .i (n13675), .o (n13676) );
  buffer buf_n13677( .i (n13676), .o (n13677) );
  buffer buf_n13678( .i (n13677), .o (n13678) );
  buffer buf_n13679( .i (n13678), .o (n13679) );
  buffer buf_n13680( .i (n13679), .o (n13680) );
  buffer buf_n13681( .i (n13680), .o (n13681) );
  buffer buf_n13682( .i (n13681), .o (n13682) );
  buffer buf_n13683( .i (n13682), .o (n13683) );
  buffer buf_n13684( .i (n13683), .o (n13684) );
  buffer buf_n13685( .i (n13684), .o (n13685) );
  buffer buf_n13686( .i (n13685), .o (n13686) );
  buffer buf_n13687( .i (n13686), .o (n13687) );
  buffer buf_n13688( .i (n13687), .o (n13688) );
  buffer buf_n13689( .i (n13688), .o (n13689) );
  buffer buf_n13690( .i (n13689), .o (n13690) );
  buffer buf_n13691( .i (n13690), .o (n13691) );
  buffer buf_n13692( .i (n13691), .o (n13692) );
  buffer buf_n13693( .i (n13692), .o (n13693) );
  buffer buf_n13694( .i (n13693), .o (n13694) );
  buffer buf_n13695( .i (n13694), .o (n13695) );
  buffer buf_n13696( .i (n13695), .o (n13696) );
  buffer buf_n13697( .i (n13696), .o (n13697) );
  buffer buf_n13698( .i (n13697), .o (n13698) );
  buffer buf_n13699( .i (n13698), .o (n13699) );
  buffer buf_n13700( .i (n13699), .o (n13700) );
  buffer buf_n13701( .i (n13700), .o (n13701) );
  buffer buf_n13702( .i (n13701), .o (n13702) );
  assign n13703 = ~n5686 & n13543 ;
  assign n13704 = n13702 | n13703 ;
  buffer buf_n13705( .i (n13704), .o (n13705) );
  buffer buf_n13706( .i (n13705), .o (n13706) );
  buffer buf_n13707( .i (n13706), .o (n13707) );
  buffer buf_n13708( .i (n13707), .o (n13708) );
  buffer buf_n13709( .i (n13708), .o (n13709) );
  buffer buf_n13710( .i (n13709), .o (n13710) );
  buffer buf_n13711( .i (n13710), .o (n13711) );
  buffer buf_n13712( .i (n13711), .o (n13712) );
  buffer buf_n13713( .i (n13712), .o (n13713) );
  buffer buf_n13714( .i (n13713), .o (n13714) );
  buffer buf_n13715( .i (n13714), .o (n13715) );
  buffer buf_n13716( .i (n13715), .o (n13716) );
  buffer buf_n13717( .i (n13716), .o (n13717) );
  buffer buf_n13718( .i (n13717), .o (n13718) );
  buffer buf_n13719( .i (n13718), .o (n13719) );
  buffer buf_n13720( .i (n13719), .o (n13720) );
  buffer buf_n13721( .i (n13720), .o (n13721) );
  buffer buf_n13722( .i (n13721), .o (n13722) );
  buffer buf_n13723( .i (n13722), .o (n13723) );
  buffer buf_n13724( .i (n13723), .o (n13724) );
  buffer buf_n13725( .i (n13724), .o (n13725) );
  buffer buf_n13726( .i (n13725), .o (n13726) );
  buffer buf_n13727( .i (n13726), .o (n13727) );
  buffer buf_n13728( .i (n13727), .o (n13728) );
  buffer buf_n13729( .i (n13728), .o (n13729) );
  buffer buf_n13730( .i (n13729), .o (n13730) );
  buffer buf_n13731( .i (n13730), .o (n13731) );
  buffer buf_n13732( .i (n13731), .o (n13732) );
  buffer buf_n13733( .i (n13732), .o (n13733) );
  buffer buf_n13734( .i (n13733), .o (n13734) );
  buffer buf_n13735( .i (n13734), .o (n13735) );
  buffer buf_n13736( .i (n13735), .o (n13736) );
  buffer buf_n13737( .i (n13736), .o (n13737) );
  buffer buf_n13738( .i (n13737), .o (n13738) );
  buffer buf_n13739( .i (n13738), .o (n13739) );
  buffer buf_n13740( .i (n13739), .o (n13740) );
  buffer buf_n13741( .i (n13740), .o (n13741) );
  buffer buf_n13742( .i (n13741), .o (n13742) );
  buffer buf_n13743( .i (n13742), .o (n13743) );
  buffer buf_n13744( .i (n13743), .o (n13744) );
  buffer buf_n13745( .i (n13744), .o (n13745) );
  buffer buf_n13746( .i (n13745), .o (n13746) );
  buffer buf_n13747( .i (n13746), .o (n13747) );
  buffer buf_n13748( .i (n13747), .o (n13748) );
  buffer buf_n13749( .i (n13748), .o (n13749) );
  buffer buf_n13750( .i (n13749), .o (n13750) );
  buffer buf_n13751( .i (n13750), .o (n13751) );
  buffer buf_n13752( .i (n13751), .o (n13752) );
  buffer buf_n13753( .i (n13752), .o (n13753) );
  buffer buf_n13754( .i (n13753), .o (n13754) );
  buffer buf_n13755( .i (n13754), .o (n13755) );
  buffer buf_n13756( .i (n13755), .o (n13756) );
  buffer buf_n13757( .i (n13756), .o (n13757) );
  buffer buf_n13758( .i (n13757), .o (n13758) );
  buffer buf_n13759( .i (n13758), .o (n13759) );
  buffer buf_n13760( .i (n13759), .o (n13760) );
  buffer buf_n13761( .i (n13760), .o (n13761) );
  buffer buf_n9366( .i (n9365), .o (n9366) );
  buffer buf_n9367( .i (n9366), .o (n9367) );
  buffer buf_n9368( .i (n9367), .o (n9368) );
  buffer buf_n9369( .i (n9368), .o (n9369) );
  buffer buf_n9370( .i (n9369), .o (n9370) );
  buffer buf_n9371( .i (n9370), .o (n9371) );
  buffer buf_n9372( .i (n9371), .o (n9372) );
  buffer buf_n9373( .i (n9372), .o (n9373) );
  buffer buf_n9374( .i (n9373), .o (n9374) );
  buffer buf_n9375( .i (n9374), .o (n9375) );
  buffer buf_n9376( .i (n9375), .o (n9376) );
  buffer buf_n9377( .i (n9376), .o (n9377) );
  buffer buf_n9378( .i (n9377), .o (n9378) );
  buffer buf_n9379( .i (n9378), .o (n9379) );
  buffer buf_n9380( .i (n9379), .o (n9380) );
  buffer buf_n9381( .i (n9380), .o (n9381) );
  buffer buf_n9382( .i (n9381), .o (n9382) );
  buffer buf_n9383( .i (n9382), .o (n9383) );
  buffer buf_n9384( .i (n9383), .o (n9384) );
  buffer buf_n9385( .i (n9384), .o (n9385) );
  buffer buf_n9386( .i (n9385), .o (n9386) );
  buffer buf_n9387( .i (n9386), .o (n9387) );
  buffer buf_n9388( .i (n9387), .o (n9388) );
  buffer buf_n9389( .i (n9388), .o (n9389) );
  buffer buf_n9390( .i (n9389), .o (n9390) );
  buffer buf_n9391( .i (n9390), .o (n9391) );
  buffer buf_n9392( .i (n9391), .o (n9392) );
  buffer buf_n9393( .i (n9392), .o (n9393) );
  buffer buf_n9394( .i (n9393), .o (n9394) );
  buffer buf_n9395( .i (n9394), .o (n9395) );
  buffer buf_n9396( .i (n9395), .o (n9396) );
  buffer buf_n9397( .i (n9396), .o (n9397) );
  buffer buf_n9398( .i (n9397), .o (n9398) );
  buffer buf_n9399( .i (n9398), .o (n9399) );
  buffer buf_n7534( .i (n7533), .o (n7534) );
  buffer buf_n7535( .i (n7534), .o (n7535) );
  assign n13762 = ~n7445 & n7538 ;
  buffer buf_n13763( .i (n13762), .o (n13763) );
  assign n13764 = ~n7535 & n13763 ;
  assign n13765 = n7535 & ~n13763 ;
  assign n13766 = n13764 | n13765 ;
  buffer buf_n13767( .i (n13766), .o (n13767) );
  buffer buf_n13768( .i (n13767), .o (n13768) );
  buffer buf_n13769( .i (n13768), .o (n13769) );
  buffer buf_n13770( .i (n13769), .o (n13770) );
  buffer buf_n13771( .i (n13770), .o (n13771) );
  buffer buf_n13772( .i (n13771), .o (n13772) );
  buffer buf_n13773( .i (n13772), .o (n13773) );
  buffer buf_n13774( .i (n13773), .o (n13774) );
  buffer buf_n13775( .i (n13774), .o (n13775) );
  buffer buf_n13776( .i (n13775), .o (n13776) );
  buffer buf_n13777( .i (n13776), .o (n13777) );
  buffer buf_n13778( .i (n13777), .o (n13778) );
  buffer buf_n13779( .i (n13778), .o (n13779) );
  buffer buf_n8557( .i (n8556), .o (n8557) );
  buffer buf_n8558( .i (n8557), .o (n8558) );
  buffer buf_n8559( .i (n8558), .o (n8559) );
  buffer buf_n8560( .i (n8559), .o (n8560) );
  buffer buf_n8561( .i (n8560), .o (n8561) );
  buffer buf_n8562( .i (n8561), .o (n8562) );
  buffer buf_n8563( .i (n8562), .o (n8563) );
  buffer buf_n8564( .i (n8563), .o (n8564) );
  buffer buf_n8565( .i (n8564), .o (n8565) );
  buffer buf_n8566( .i (n8565), .o (n8566) );
  buffer buf_n8567( .i (n8566), .o (n8567) );
  buffer buf_n8568( .i (n8567), .o (n8568) );
  buffer buf_n8569( .i (n8568), .o (n8569) );
  buffer buf_n8570( .i (n8569), .o (n8570) );
  buffer buf_n8571( .i (n8570), .o (n8571) );
  buffer buf_n8572( .i (n8571), .o (n8572) );
  buffer buf_n8573( .i (n8572), .o (n8573) );
  buffer buf_n8574( .i (n8573), .o (n8574) );
  buffer buf_n8575( .i (n8574), .o (n8575) );
  buffer buf_n8576( .i (n8575), .o (n8576) );
  buffer buf_n8577( .i (n8576), .o (n8577) );
  buffer buf_n8578( .i (n8577), .o (n8578) );
  buffer buf_n8579( .i (n8578), .o (n8579) );
  buffer buf_n8580( .i (n8579), .o (n8580) );
  buffer buf_n8581( .i (n8580), .o (n8581) );
  buffer buf_n8582( .i (n8581), .o (n8582) );
  buffer buf_n8583( .i (n8582), .o (n8583) );
  buffer buf_n8584( .i (n8583), .o (n8584) );
  buffer buf_n8585( .i (n8584), .o (n8585) );
  buffer buf_n8586( .i (n8585), .o (n8586) );
  buffer buf_n8587( .i (n8586), .o (n8587) );
  buffer buf_n8588( .i (n8587), .o (n8588) );
  buffer buf_n8589( .i (n8588), .o (n8589) );
  buffer buf_n8590( .i (n8589), .o (n8590) );
  buffer buf_n8591( .i (n8590), .o (n8591) );
  buffer buf_n8592( .i (n8591), .o (n8592) );
  buffer buf_n8593( .i (n8592), .o (n8593) );
  buffer buf_n8594( .i (n8593), .o (n8594) );
  buffer buf_n8595( .i (n8594), .o (n8595) );
  buffer buf_n8596( .i (n8595), .o (n8596) );
  buffer buf_n8597( .i (n8596), .o (n8597) );
  buffer buf_n8598( .i (n8597), .o (n8598) );
  buffer buf_n8599( .i (n8598), .o (n8599) );
  buffer buf_n8600( .i (n8599), .o (n8600) );
  buffer buf_n8601( .i (n8600), .o (n8601) );
  buffer buf_n8602( .i (n8601), .o (n8602) );
  buffer buf_n8603( .i (n8602), .o (n8603) );
  buffer buf_n8604( .i (n8603), .o (n8604) );
  buffer buf_n8605( .i (n8604), .o (n8605) );
  buffer buf_n8606( .i (n8605), .o (n8606) );
  buffer buf_n8607( .i (n8606), .o (n8607) );
  buffer buf_n8608( .i (n8607), .o (n8608) );
  buffer buf_n8609( .i (n8608), .o (n8609) );
  buffer buf_n8610( .i (n8609), .o (n8610) );
  buffer buf_n8611( .i (n8610), .o (n8611) );
  buffer buf_n8612( .i (n8611), .o (n8612) );
  buffer buf_n8613( .i (n8612), .o (n8613) );
  buffer buf_n8614( .i (n8613), .o (n8614) );
  buffer buf_n8615( .i (n8614), .o (n8615) );
  buffer buf_n8616( .i (n8615), .o (n8616) );
  buffer buf_n8617( .i (n8616), .o (n8617) );
  buffer buf_n8618( .i (n8617), .o (n8618) );
  buffer buf_n8619( .i (n8618), .o (n8619) );
  buffer buf_n8620( .i (n8619), .o (n8620) );
  buffer buf_n8621( .i (n8620), .o (n8621) );
  buffer buf_n8622( .i (n8621), .o (n8622) );
  buffer buf_n8623( .i (n8622), .o (n8623) );
  buffer buf_n8624( .i (n8623), .o (n8624) );
  buffer buf_n8625( .i (n8624), .o (n8625) );
  buffer buf_n8626( .i (n8625), .o (n8626) );
  buffer buf_n8627( .i (n8626), .o (n8627) );
  buffer buf_n8628( .i (n8627), .o (n8628) );
  buffer buf_n8629( .i (n8628), .o (n8629) );
  buffer buf_n8630( .i (n8629), .o (n8630) );
  buffer buf_n8631( .i (n8630), .o (n8631) );
  buffer buf_n8632( .i (n8631), .o (n8632) );
  buffer buf_n8633( .i (n8632), .o (n8633) );
  buffer buf_n8634( .i (n8633), .o (n8634) );
  buffer buf_n8635( .i (n8634), .o (n8635) );
  buffer buf_n8636( .i (n8635), .o (n8636) );
  buffer buf_n8637( .i (n8636), .o (n8637) );
  buffer buf_n8638( .i (n8637), .o (n8638) );
  buffer buf_n8639( .i (n8638), .o (n8639) );
  buffer buf_n8640( .i (n8639), .o (n8640) );
  buffer buf_n4866( .i (n4865), .o (n4866) );
  buffer buf_n4867( .i (n4866), .o (n4867) );
  assign n13780 = n4858 & ~n4869 ;
  buffer buf_n13781( .i (n13780), .o (n13781) );
  assign n13782 = n4867 & ~n13781 ;
  assign n13783 = ~n4867 & n13781 ;
  assign n13784 = n13782 | n13783 ;
  buffer buf_n13785( .i (n13784), .o (n13785) );
  buffer buf_n13786( .i (n13785), .o (n13786) );
  buffer buf_n13787( .i (n13786), .o (n13787) );
  buffer buf_n13788( .i (n13787), .o (n13788) );
  buffer buf_n13789( .i (n13788), .o (n13789) );
  buffer buf_n13790( .i (n13789), .o (n13790) );
  buffer buf_n13791( .i (n13790), .o (n13791) );
  buffer buf_n13792( .i (n13791), .o (n13792) );
  buffer buf_n13793( .i (n13792), .o (n13793) );
  buffer buf_n13794( .i (n13793), .o (n13794) );
  buffer buf_n13795( .i (n13794), .o (n13795) );
  buffer buf_n13796( .i (n13795), .o (n13796) );
  buffer buf_n13797( .i (n13796), .o (n13797) );
  buffer buf_n13798( .i (n13797), .o (n13798) );
  buffer buf_n13799( .i (n13798), .o (n13799) );
  buffer buf_n13800( .i (n13799), .o (n13800) );
  buffer buf_n13801( .i (n13800), .o (n13801) );
  buffer buf_n13802( .i (n13801), .o (n13802) );
  buffer buf_n13803( .i (n13802), .o (n13803) );
  buffer buf_n13804( .i (n13803), .o (n13804) );
  buffer buf_n13805( .i (n13804), .o (n13805) );
  buffer buf_n13806( .i (n13805), .o (n13806) );
  buffer buf_n13807( .i (n13806), .o (n13807) );
  buffer buf_n13808( .i (n13807), .o (n13808) );
  buffer buf_n13809( .i (n13808), .o (n13809) );
  buffer buf_n13810( .i (n13809), .o (n13810) );
  buffer buf_n13811( .i (n13810), .o (n13811) );
  buffer buf_n13812( .i (n13811), .o (n13812) );
  buffer buf_n13813( .i (n13812), .o (n13813) );
  buffer buf_n13814( .i (n13813), .o (n13814) );
  buffer buf_n13815( .i (n13814), .o (n13815) );
  buffer buf_n13816( .i (n13815), .o (n13816) );
  buffer buf_n13817( .i (n13816), .o (n13817) );
  assign n13932 = ~n13392 & n13817 ;
  assign n13933 = n6593 & n11683 ;
  assign n13934 = n8118 & n9261 ;
  buffer buf_n13935( .i (n13934), .o (n13935) );
  assign n13936 = ~n45 & n8101 ;
  assign n13937 = n13935 | n13936 ;
  buffer buf_n13938( .i (n11494), .o (n13938) );
  buffer buf_n13939( .i (n13938), .o (n13939) );
  assign n13940 = n13937 & ~n13939 ;
  assign n13941 = n13933 | n13940 ;
  assign n13942 = ~n13613 & n13941 ;
  assign n13943 = n13612 & n13613 ;
  assign n13944 = n13942 | n13943 ;
  buffer buf_n13945( .i (n12711), .o (n13945) );
  assign n13946 = n13944 & ~n13945 ;
  assign n13947 = n10244 & n13945 ;
  assign n13948 = n13946 | n13947 ;
  buffer buf_n13949( .i (n13948), .o (n13949) );
  buffer buf_n13950( .i (n5925), .o (n13950) );
  buffer buf_n13951( .i (n13950), .o (n13951) );
  assign n13952 = ~n13949 & n13951 ;
  assign n13953 = n13244 & ~n13952 ;
  assign n13954 = n10272 & ~n13945 ;
  assign n13955 = n12714 | n13954 ;
  buffer buf_n13956( .i (n13955), .o (n13956) );
  assign n13957 = n13622 & n13956 ;
  assign n13958 = n483 & n1851 ;
  buffer buf_n13959( .i (n13958), .o (n13959) );
  buffer buf_n13960( .i (n13959), .o (n13960) );
  buffer buf_n13961( .i (n13960), .o (n13961) );
  assign n13962 = n6056 & n13961 ;
  buffer buf_n13963( .i (n6064), .o (n13963) );
  assign n13964 = n1853 & n13963 ;
  assign n13965 = n486 | n13964 ;
  assign n13966 = n6077 & n13959 ;
  assign n13967 = n13396 | n13966 ;
  assign n13968 = n13965 & ~n13967 ;
  assign n13969 = n13962 | n13968 ;
  buffer buf_n13970( .i (n13969), .o (n13970) );
  buffer buf_n13971( .i (n13970), .o (n13971) );
  assign n13972 = ~n6090 & n13971 ;
  buffer buf_n13973( .i (n13972), .o (n13973) );
  buffer buf_n13974( .i (n13973), .o (n13974) );
  buffer buf_n13975( .i (n11669), .o (n13975) );
  assign n13976 = n13974 | n13975 ;
  buffer buf_n13977( .i (n13976), .o (n13977) );
  buffer buf_n13978( .i (n13977), .o (n13978) );
  buffer buf_n13979( .i (n13978), .o (n13979) );
  buffer buf_n13980( .i (n13979), .o (n13980) );
  buffer buf_n13981( .i (n13980), .o (n13981) );
  buffer buf_n13982( .i (n13981), .o (n13982) );
  buffer buf_n13983( .i (n13982), .o (n13983) );
  buffer buf_n13984( .i (n13983), .o (n13984) );
  assign n13985 = n13957 | n13984 ;
  assign n13986 = n13953 & n13985 ;
  assign n13987 = n13932 | n13986 ;
  buffer buf_n13988( .i (n13987), .o (n13988) );
  buffer buf_n13989( .i (n13988), .o (n13989) );
  buffer buf_n13990( .i (n13989), .o (n13990) );
  buffer buf_n13991( .i (n13990), .o (n13991) );
  buffer buf_n13992( .i (n13991), .o (n13992) );
  buffer buf_n13993( .i (n13992), .o (n13993) );
  buffer buf_n13994( .i (n13993), .o (n13994) );
  buffer buf_n13995( .i (n13994), .o (n13995) );
  buffer buf_n13996( .i (n13995), .o (n13996) );
  buffer buf_n13997( .i (n13996), .o (n13997) );
  buffer buf_n13998( .i (n13997), .o (n13998) );
  buffer buf_n13999( .i (n13998), .o (n13999) );
  buffer buf_n14000( .i (n13999), .o (n14000) );
  buffer buf_n14001( .i (n14000), .o (n14001) );
  buffer buf_n14002( .i (n14001), .o (n14002) );
  buffer buf_n14003( .i (n14002), .o (n14003) );
  buffer buf_n14004( .i (n14003), .o (n14004) );
  buffer buf_n14005( .i (n14004), .o (n14005) );
  buffer buf_n14006( .i (n14005), .o (n14006) );
  buffer buf_n14007( .i (n14006), .o (n14007) );
  buffer buf_n14008( .i (n14007), .o (n14008) );
  buffer buf_n14009( .i (n14008), .o (n14009) );
  buffer buf_n14010( .i (n14009), .o (n14010) );
  buffer buf_n14011( .i (n14010), .o (n14011) );
  buffer buf_n14012( .i (n14011), .o (n14012) );
  buffer buf_n14013( .i (n14012), .o (n14013) );
  buffer buf_n14014( .i (n14013), .o (n14014) );
  buffer buf_n14015( .i (n14014), .o (n14015) );
  buffer buf_n14016( .i (n14015), .o (n14016) );
  buffer buf_n14017( .i (n14016), .o (n14017) );
  buffer buf_n14018( .i (n14017), .o (n14018) );
  buffer buf_n14019( .i (n14018), .o (n14019) );
  buffer buf_n14020( .i (n14019), .o (n14020) );
  buffer buf_n14021( .i (n14020), .o (n14021) );
  buffer buf_n14022( .i (n14021), .o (n14022) );
  buffer buf_n14023( .i (n14022), .o (n14023) );
  buffer buf_n14024( .i (n14023), .o (n14024) );
  buffer buf_n14025( .i (n14024), .o (n14025) );
  buffer buf_n14026( .i (n14025), .o (n14026) );
  buffer buf_n14027( .i (n14026), .o (n14027) );
  buffer buf_n14028( .i (n14027), .o (n14028) );
  buffer buf_n14029( .i (n14028), .o (n14029) );
  buffer buf_n14030( .i (n14029), .o (n14030) );
  buffer buf_n14031( .i (n14030), .o (n14031) );
  buffer buf_n14032( .i (n14031), .o (n14032) );
  buffer buf_n14033( .i (n14032), .o (n14033) );
  buffer buf_n14034( .i (n14033), .o (n14034) );
  buffer buf_n14035( .i (n14034), .o (n14035) );
  buffer buf_n14036( .i (n14035), .o (n14036) );
  buffer buf_n14037( .i (n14036), .o (n14037) );
  buffer buf_n14038( .i (n14037), .o (n14038) );
  buffer buf_n14039( .i (n14038), .o (n14039) );
  buffer buf_n14040( .i (n14039), .o (n14040) );
  buffer buf_n14041( .i (n14040), .o (n14041) );
  buffer buf_n14042( .i (n14041), .o (n14042) );
  buffer buf_n14043( .i (n14042), .o (n14043) );
  buffer buf_n14044( .i (n14043), .o (n14044) );
  buffer buf_n14045( .i (n14044), .o (n14045) );
  buffer buf_n14046( .i (n14045), .o (n14046) );
  buffer buf_n14047( .i (n14046), .o (n14047) );
  buffer buf_n14048( .i (n14047), .o (n14048) );
  buffer buf_n14049( .i (n14048), .o (n14049) );
  buffer buf_n14050( .i (n14049), .o (n14050) );
  buffer buf_n14051( .i (n14050), .o (n14051) );
  buffer buf_n14052( .i (n14051), .o (n14052) );
  buffer buf_n14053( .i (n14052), .o (n14053) );
  buffer buf_n14054( .i (n14053), .o (n14054) );
  buffer buf_n14055( .i (n14054), .o (n14055) );
  buffer buf_n14056( .i (n14055), .o (n14056) );
  buffer buf_n14057( .i (n14056), .o (n14057) );
  buffer buf_n14058( .i (n14057), .o (n14058) );
  buffer buf_n14059( .i (n14058), .o (n14059) );
  buffer buf_n14060( .i (n14059), .o (n14060) );
  buffer buf_n14061( .i (n14060), .o (n14061) );
  buffer buf_n14062( .i (n14061), .o (n14062) );
  buffer buf_n14063( .i (n14062), .o (n14063) );
  buffer buf_n14064( .i (n14063), .o (n14064) );
  buffer buf_n14065( .i (n14064), .o (n14065) );
  buffer buf_n14066( .i (n14065), .o (n14066) );
  buffer buf_n14067( .i (n14066), .o (n14067) );
  buffer buf_n14068( .i (n14067), .o (n14068) );
  buffer buf_n14069( .i (n14068), .o (n14069) );
  buffer buf_n14070( .i (n14069), .o (n14070) );
  buffer buf_n14071( .i (n14070), .o (n14071) );
  buffer buf_n14072( .i (n14071), .o (n14072) );
  buffer buf_n14073( .i (n14072), .o (n14073) );
  buffer buf_n14074( .i (n14073), .o (n14074) );
  buffer buf_n14075( .i (n14074), .o (n14075) );
  buffer buf_n14076( .i (n14075), .o (n14076) );
  buffer buf_n14077( .i (n14076), .o (n14077) );
  buffer buf_n14078( .i (n14077), .o (n14078) );
  buffer buf_n14079( .i (n14078), .o (n14079) );
  buffer buf_n14080( .i (n14079), .o (n14080) );
  buffer buf_n14081( .i (n14080), .o (n14081) );
  buffer buf_n14082( .i (n14081), .o (n14082) );
  buffer buf_n14083( .i (n14082), .o (n14083) );
  buffer buf_n14084( .i (n14083), .o (n14084) );
  buffer buf_n14085( .i (n14084), .o (n14085) );
  buffer buf_n14086( .i (n14085), .o (n14086) );
  buffer buf_n14087( .i (n14086), .o (n14087) );
  buffer buf_n14088( .i (n14087), .o (n14088) );
  buffer buf_n14089( .i (n14088), .o (n14089) );
  buffer buf_n14090( .i (n14089), .o (n14090) );
  buffer buf_n14091( .i (n14090), .o (n14091) );
  buffer buf_n14092( .i (n14091), .o (n14092) );
  buffer buf_n14093( .i (n14092), .o (n14093) );
  buffer buf_n14094( .i (n14093), .o (n14094) );
  buffer buf_n14095( .i (n14094), .o (n14095) );
  buffer buf_n14096( .i (n14095), .o (n14096) );
  buffer buf_n14097( .i (n14096), .o (n14097) );
  buffer buf_n14098( .i (n14097), .o (n14098) );
  buffer buf_n14099( .i (n14098), .o (n14099) );
  assign n14100 = n13951 & ~n13956 ;
  buffer buf_n14101( .i (n5882), .o (n14101) );
  buffer buf_n14102( .i (n14101), .o (n14102) );
  assign n14103 = ~n14100 & n14102 ;
  buffer buf_n14104( .i (n13399), .o (n14104) );
  assign n14105 = n949 & n14104 ;
  assign n14106 = n2311 | n14105 ;
  assign n14107 = n948 & n2309 ;
  buffer buf_n14108( .i (n14107), .o (n14108) );
  buffer buf_n14110( .i (n10915), .o (n14110) );
  assign n14111 = n14108 & n14110 ;
  assign n14112 = n14106 & ~n14111 ;
  assign n14113 = n13037 | n14112 ;
  buffer buf_n14109( .i (n14108), .o (n14109) );
  assign n14114 = n13036 & ~n14109 ;
  assign n14115 = n13408 | n14114 ;
  assign n14116 = n14113 & ~n14115 ;
  buffer buf_n14117( .i (n14116), .o (n14117) );
  buffer buf_n14118( .i (n14117), .o (n14118) );
  assign n14119 = n13975 | n14118 ;
  buffer buf_n14120( .i (n14119), .o (n14120) );
  buffer buf_n14121( .i (n14120), .o (n14121) );
  buffer buf_n14122( .i (n14121), .o (n14122) );
  buffer buf_n14123( .i (n14122), .o (n14123) );
  buffer buf_n14124( .i (n14123), .o (n14124) );
  buffer buf_n14125( .i (n14124), .o (n14125) );
  buffer buf_n14126( .i (n14125), .o (n14126) );
  buffer buf_n14127( .i (n14126), .o (n14127) );
  assign n14128 = n13622 & n13949 ;
  assign n14129 = n14127 | n14128 ;
  assign n14130 = n14103 & n14129 ;
  buffer buf_n14131( .i (n14130), .o (n14131) );
  buffer buf_n14132( .i (n14131), .o (n14132) );
  buffer buf_n14133( .i (n14132), .o (n14133) );
  buffer buf_n14134( .i (n14133), .o (n14134) );
  buffer buf_n14135( .i (n14134), .o (n14135) );
  buffer buf_n14136( .i (n14135), .o (n14136) );
  buffer buf_n14137( .i (n14136), .o (n14137) );
  buffer buf_n14138( .i (n14137), .o (n14138) );
  buffer buf_n14139( .i (n14138), .o (n14139) );
  buffer buf_n14140( .i (n14139), .o (n14140) );
  buffer buf_n14141( .i (n14140), .o (n14141) );
  buffer buf_n14142( .i (n14141), .o (n14142) );
  buffer buf_n14143( .i (n14142), .o (n14143) );
  buffer buf_n14144( .i (n14143), .o (n14144) );
  buffer buf_n14145( .i (n14144), .o (n14145) );
  buffer buf_n14146( .i (n14145), .o (n14146) );
  buffer buf_n14147( .i (n14146), .o (n14147) );
  buffer buf_n14148( .i (n14147), .o (n14148) );
  buffer buf_n14149( .i (n14148), .o (n14149) );
  buffer buf_n14150( .i (n14149), .o (n14150) );
  buffer buf_n14151( .i (n14150), .o (n14151) );
  buffer buf_n14152( .i (n14151), .o (n14152) );
  buffer buf_n14153( .i (n14152), .o (n14153) );
  buffer buf_n14154( .i (n14153), .o (n14154) );
  buffer buf_n14155( .i (n14154), .o (n14155) );
  buffer buf_n14156( .i (n14155), .o (n14156) );
  buffer buf_n14157( .i (n14156), .o (n14157) );
  buffer buf_n14158( .i (n14157), .o (n14158) );
  buffer buf_n14159( .i (n14158), .o (n14159) );
  buffer buf_n14160( .i (n14159), .o (n14160) );
  buffer buf_n14161( .i (n14160), .o (n14161) );
  buffer buf_n14162( .i (n14161), .o (n14162) );
  buffer buf_n14163( .i (n14162), .o (n14163) );
  buffer buf_n14164( .i (n14163), .o (n14164) );
  buffer buf_n14165( .i (n14164), .o (n14165) );
  buffer buf_n14166( .i (n14165), .o (n14166) );
  buffer buf_n14167( .i (n14166), .o (n14167) );
  buffer buf_n14168( .i (n14167), .o (n14168) );
  buffer buf_n14169( .i (n14168), .o (n14169) );
  buffer buf_n14170( .i (n14169), .o (n14170) );
  buffer buf_n14171( .i (n14170), .o (n14171) );
  buffer buf_n14172( .i (n14171), .o (n14172) );
  buffer buf_n14173( .i (n14172), .o (n14173) );
  buffer buf_n14174( .i (n14173), .o (n14174) );
  buffer buf_n14175( .i (n14174), .o (n14175) );
  buffer buf_n14176( .i (n14175), .o (n14176) );
  buffer buf_n14177( .i (n14176), .o (n14177) );
  buffer buf_n14178( .i (n14177), .o (n14178) );
  buffer buf_n14179( .i (n14178), .o (n14179) );
  buffer buf_n14180( .i (n14179), .o (n14180) );
  buffer buf_n14181( .i (n14180), .o (n14181) );
  buffer buf_n14182( .i (n14181), .o (n14182) );
  buffer buf_n14183( .i (n14182), .o (n14183) );
  buffer buf_n14184( .i (n14183), .o (n14184) );
  buffer buf_n14185( .i (n14184), .o (n14185) );
  buffer buf_n14186( .i (n14185), .o (n14186) );
  buffer buf_n14187( .i (n14186), .o (n14187) );
  buffer buf_n14188( .i (n14187), .o (n14188) );
  buffer buf_n14189( .i (n14188), .o (n14189) );
  buffer buf_n14190( .i (n14189), .o (n14190) );
  buffer buf_n14191( .i (n14190), .o (n14191) );
  buffer buf_n14192( .i (n14191), .o (n14192) );
  buffer buf_n14193( .i (n14192), .o (n14193) );
  buffer buf_n14194( .i (n14193), .o (n14194) );
  buffer buf_n14195( .i (n14194), .o (n14195) );
  buffer buf_n14196( .i (n14195), .o (n14196) );
  buffer buf_n14197( .i (n14196), .o (n14197) );
  buffer buf_n14198( .i (n14197), .o (n14198) );
  buffer buf_n14199( .i (n14198), .o (n14199) );
  buffer buf_n14200( .i (n14199), .o (n14200) );
  buffer buf_n14201( .i (n14200), .o (n14201) );
  buffer buf_n14202( .i (n14201), .o (n14202) );
  buffer buf_n14203( .i (n14202), .o (n14203) );
  buffer buf_n14204( .i (n14203), .o (n14204) );
  buffer buf_n14205( .i (n14204), .o (n14205) );
  buffer buf_n14206( .i (n14205), .o (n14206) );
  buffer buf_n14207( .i (n14206), .o (n14207) );
  buffer buf_n14208( .i (n14207), .o (n14208) );
  buffer buf_n14209( .i (n14208), .o (n14209) );
  buffer buf_n14210( .i (n14209), .o (n14210) );
  buffer buf_n14211( .i (n14210), .o (n14211) );
  buffer buf_n14212( .i (n14211), .o (n14212) );
  buffer buf_n14213( .i (n14212), .o (n14213) );
  buffer buf_n14214( .i (n14213), .o (n14214) );
  buffer buf_n14215( .i (n14214), .o (n14215) );
  buffer buf_n14216( .i (n14215), .o (n14216) );
  buffer buf_n14217( .i (n14216), .o (n14217) );
  buffer buf_n14218( .i (n14217), .o (n14218) );
  buffer buf_n14219( .i (n14218), .o (n14219) );
  buffer buf_n14220( .i (n14219), .o (n14220) );
  buffer buf_n14221( .i (n14220), .o (n14221) );
  buffer buf_n14222( .i (n14221), .o (n14222) );
  buffer buf_n14223( .i (n14222), .o (n14223) );
  buffer buf_n14224( .i (n14223), .o (n14224) );
  buffer buf_n14225( .i (n14224), .o (n14225) );
  buffer buf_n14226( .i (n14225), .o (n14226) );
  assign n14227 = n7437 & ~n7441 ;
  buffer buf_n6985( .i (n6984), .o (n6985) );
  buffer buf_n6986( .i (n6985), .o (n6986) );
  buffer buf_n7435( .i (n7434), .o (n7435) );
  assign n14228 = n7435 & ~n7440 ;
  assign n14229 = n6986 | n14228 ;
  assign n14230 = ~n14227 & n14229 ;
  buffer buf_n14231( .i (n14230), .o (n14231) );
  assign n14250 = ~n5727 & n14231 ;
  assign n14251 = n14226 | n14250 ;
  buffer buf_n14252( .i (n14251), .o (n14252) );
  buffer buf_n14253( .i (n14252), .o (n14253) );
  buffer buf_n14254( .i (n14253), .o (n14254) );
  buffer buf_n14255( .i (n14254), .o (n14255) );
  buffer buf_n14256( .i (n14255), .o (n14256) );
  buffer buf_n14257( .i (n14256), .o (n14257) );
  buffer buf_n14258( .i (n14257), .o (n14258) );
  buffer buf_n14259( .i (n14258), .o (n14259) );
  buffer buf_n14260( .i (n14259), .o (n14260) );
  buffer buf_n14261( .i (n14260), .o (n14261) );
  buffer buf_n14262( .i (n14261), .o (n14262) );
  buffer buf_n14263( .i (n14262), .o (n14263) );
  buffer buf_n14264( .i (n14263), .o (n14264) );
  buffer buf_n14265( .i (n14264), .o (n14265) );
  buffer buf_n14266( .i (n14265), .o (n14266) );
  buffer buf_n14267( .i (n14266), .o (n14267) );
  buffer buf_n7427( .i (n7426), .o (n7427) );
  buffer buf_n7428( .i (n7427), .o (n7428) );
  buffer buf_n7342( .i (n7341), .o (n7342) );
  assign n14268 = n7338 & ~n7342 ;
  assign n14269 = n7428 & ~n14268 ;
  assign n14270 = n7339 & ~n7430 ;
  assign n14271 = n14269 | n14270 ;
  buffer buf_n14272( .i (n14271), .o (n14272) );
  assign n14297 = ~n5721 & n14272 ;
  assign n14298 = n889 & n14104 ;
  assign n14299 = n3604 | n14298 ;
  assign n14300 = n888 & n3602 ;
  buffer buf_n14301( .i (n14300), .o (n14301) );
  assign n14303 = n14110 & n14301 ;
  assign n14304 = n14299 & ~n14303 ;
  buffer buf_n14305( .i (n13396), .o (n14305) );
  buffer buf_n14306( .i (n14305), .o (n14306) );
  buffer buf_n14307( .i (n14306), .o (n14307) );
  buffer buf_n14308( .i (n14307), .o (n14308) );
  assign n14309 = n14304 | n14308 ;
  buffer buf_n14302( .i (n14301), .o (n14302) );
  assign n14310 = ~n14302 & n14307 ;
  assign n14311 = n13408 | n14310 ;
  assign n14312 = n14309 & ~n14311 ;
  buffer buf_n14313( .i (n14312), .o (n14313) );
  buffer buf_n14314( .i (n14313), .o (n14314) );
  assign n14315 = n13975 | n14314 ;
  buffer buf_n14316( .i (n14315), .o (n14316) );
  buffer buf_n14317( .i (n14316), .o (n14317) );
  buffer buf_n14318( .i (n14317), .o (n14318) );
  buffer buf_n14319( .i (n14318), .o (n14319) );
  buffer buf_n14320( .i (n14319), .o (n14320) );
  buffer buf_n14321( .i (n14320), .o (n14321) );
  buffer buf_n14322( .i (n14321), .o (n14322) );
  buffer buf_n14323( .i (n14322), .o (n14323) );
  assign n14324 = n12759 & n13622 ;
  assign n14325 = n14323 | n14324 ;
  assign n14326 = ~n12716 & n13951 ;
  assign n14327 = n14102 & ~n14326 ;
  assign n14328 = n14325 & n14327 ;
  buffer buf_n14329( .i (n14328), .o (n14329) );
  buffer buf_n14330( .i (n14329), .o (n14330) );
  buffer buf_n14331( .i (n14330), .o (n14331) );
  buffer buf_n14332( .i (n14331), .o (n14332) );
  buffer buf_n14333( .i (n14332), .o (n14333) );
  buffer buf_n14334( .i (n14333), .o (n14334) );
  buffer buf_n14335( .i (n14334), .o (n14335) );
  buffer buf_n14336( .i (n14335), .o (n14336) );
  buffer buf_n14337( .i (n14336), .o (n14337) );
  buffer buf_n14338( .i (n14337), .o (n14338) );
  buffer buf_n14339( .i (n14338), .o (n14339) );
  buffer buf_n14340( .i (n14339), .o (n14340) );
  buffer buf_n14341( .i (n14340), .o (n14341) );
  buffer buf_n14342( .i (n14341), .o (n14342) );
  buffer buf_n14343( .i (n14342), .o (n14343) );
  buffer buf_n14344( .i (n14343), .o (n14344) );
  buffer buf_n14345( .i (n14344), .o (n14345) );
  buffer buf_n14346( .i (n14345), .o (n14346) );
  buffer buf_n14347( .i (n14346), .o (n14347) );
  buffer buf_n14348( .i (n14347), .o (n14348) );
  buffer buf_n14349( .i (n14348), .o (n14349) );
  buffer buf_n14350( .i (n14349), .o (n14350) );
  buffer buf_n14351( .i (n14350), .o (n14351) );
  buffer buf_n14352( .i (n14351), .o (n14352) );
  buffer buf_n14353( .i (n14352), .o (n14353) );
  buffer buf_n14354( .i (n14353), .o (n14354) );
  buffer buf_n14355( .i (n14354), .o (n14355) );
  buffer buf_n14356( .i (n14355), .o (n14356) );
  buffer buf_n14357( .i (n14356), .o (n14357) );
  buffer buf_n14358( .i (n14357), .o (n14358) );
  buffer buf_n14359( .i (n14358), .o (n14359) );
  buffer buf_n14360( .i (n14359), .o (n14360) );
  buffer buf_n14361( .i (n14360), .o (n14361) );
  buffer buf_n14362( .i (n14361), .o (n14362) );
  buffer buf_n14363( .i (n14362), .o (n14363) );
  buffer buf_n14364( .i (n14363), .o (n14364) );
  buffer buf_n14365( .i (n14364), .o (n14365) );
  buffer buf_n14366( .i (n14365), .o (n14366) );
  buffer buf_n14367( .i (n14366), .o (n14367) );
  buffer buf_n14368( .i (n14367), .o (n14368) );
  buffer buf_n14369( .i (n14368), .o (n14369) );
  buffer buf_n14370( .i (n14369), .o (n14370) );
  buffer buf_n14371( .i (n14370), .o (n14371) );
  buffer buf_n14372( .i (n14371), .o (n14372) );
  buffer buf_n14373( .i (n14372), .o (n14373) );
  buffer buf_n14374( .i (n14373), .o (n14374) );
  buffer buf_n14375( .i (n14374), .o (n14375) );
  buffer buf_n14376( .i (n14375), .o (n14376) );
  buffer buf_n14377( .i (n14376), .o (n14377) );
  buffer buf_n14378( .i (n14377), .o (n14378) );
  buffer buf_n14379( .i (n14378), .o (n14379) );
  buffer buf_n14380( .i (n14379), .o (n14380) );
  buffer buf_n14381( .i (n14380), .o (n14381) );
  buffer buf_n14382( .i (n14381), .o (n14382) );
  buffer buf_n14383( .i (n14382), .o (n14383) );
  buffer buf_n14384( .i (n14383), .o (n14384) );
  buffer buf_n14385( .i (n14384), .o (n14385) );
  buffer buf_n14386( .i (n14385), .o (n14386) );
  buffer buf_n14387( .i (n14386), .o (n14387) );
  buffer buf_n14388( .i (n14387), .o (n14388) );
  buffer buf_n14389( .i (n14388), .o (n14389) );
  buffer buf_n14390( .i (n14389), .o (n14390) );
  buffer buf_n14391( .i (n14390), .o (n14391) );
  buffer buf_n14392( .i (n14391), .o (n14392) );
  buffer buf_n14393( .i (n14392), .o (n14393) );
  buffer buf_n14394( .i (n14393), .o (n14394) );
  buffer buf_n14395( .i (n14394), .o (n14395) );
  buffer buf_n14396( .i (n14395), .o (n14396) );
  buffer buf_n14397( .i (n14396), .o (n14397) );
  buffer buf_n14398( .i (n14397), .o (n14398) );
  buffer buf_n14399( .i (n14398), .o (n14399) );
  buffer buf_n14400( .i (n14399), .o (n14400) );
  buffer buf_n14401( .i (n14400), .o (n14401) );
  buffer buf_n14402( .i (n14401), .o (n14402) );
  buffer buf_n14403( .i (n14402), .o (n14403) );
  buffer buf_n14404( .i (n14403), .o (n14404) );
  buffer buf_n14405( .i (n14404), .o (n14405) );
  buffer buf_n14406( .i (n14405), .o (n14406) );
  buffer buf_n14407( .i (n14406), .o (n14407) );
  buffer buf_n14408( .i (n14407), .o (n14408) );
  buffer buf_n14409( .i (n14408), .o (n14409) );
  buffer buf_n14410( .i (n14409), .o (n14410) );
  buffer buf_n14411( .i (n14410), .o (n14411) );
  buffer buf_n14412( .i (n14411), .o (n14412) );
  buffer buf_n14413( .i (n14412), .o (n14413) );
  buffer buf_n14414( .i (n14413), .o (n14414) );
  buffer buf_n14415( .i (n14414), .o (n14415) );
  buffer buf_n14416( .i (n14415), .o (n14416) );
  buffer buf_n14417( .i (n14416), .o (n14417) );
  buffer buf_n14418( .i (n14417), .o (n14418) );
  assign n14419 = n14297 | n14418 ;
  buffer buf_n14420( .i (n14419), .o (n14420) );
  buffer buf_n14421( .i (n14420), .o (n14421) );
  buffer buf_n14422( .i (n14421), .o (n14422) );
  buffer buf_n14423( .i (n14422), .o (n14423) );
  buffer buf_n14424( .i (n14423), .o (n14424) );
  buffer buf_n14425( .i (n14424), .o (n14425) );
  buffer buf_n14426( .i (n14425), .o (n14426) );
  buffer buf_n14427( .i (n14426), .o (n14427) );
  buffer buf_n14428( .i (n14427), .o (n14428) );
  buffer buf_n14429( .i (n14428), .o (n14429) );
  buffer buf_n14430( .i (n14429), .o (n14430) );
  buffer buf_n14431( .i (n14430), .o (n14431) );
  buffer buf_n14432( .i (n14431), .o (n14432) );
  buffer buf_n14433( .i (n14432), .o (n14433) );
  buffer buf_n14434( .i (n14433), .o (n14434) );
  buffer buf_n14435( .i (n14434), .o (n14435) );
  buffer buf_n14436( .i (n14435), .o (n14436) );
  buffer buf_n14437( .i (n14436), .o (n14437) );
  buffer buf_n14438( .i (n14437), .o (n14438) );
  buffer buf_n14439( .i (n14438), .o (n14439) );
  buffer buf_n14440( .i (n14439), .o (n14440) );
  buffer buf_n14441( .i (n14440), .o (n14441) );
  buffer buf_n5079( .i (n5078), .o (n5079) );
  buffer buf_n5080( .i (n5079), .o (n5080) );
  buffer buf_n5045( .i (n5044), .o (n5045) );
  assign n14442 = ~n5045 & n5085 ;
  assign n14443 = n5080 & ~n14442 ;
  assign n14444 = ~n5082 & n5086 ;
  assign n14445 = n14443 | n14444 ;
  buffer buf_n14446( .i (n14445), .o (n14446) );
  buffer buf_n14447( .i (n14446), .o (n14447) );
  buffer buf_n14448( .i (n14447), .o (n14448) );
  buffer buf_n14449( .i (n14448), .o (n14449) );
  buffer buf_n14450( .i (n14449), .o (n14450) );
  buffer buf_n14451( .i (n14450), .o (n14451) );
  buffer buf_n14452( .i (n14451), .o (n14452) );
  buffer buf_n14453( .i (n14452), .o (n14453) );
  buffer buf_n14454( .i (n14453), .o (n14454) );
  buffer buf_n14455( .i (n14454), .o (n14455) );
  buffer buf_n14456( .i (n14455), .o (n14456) );
  buffer buf_n14457( .i (n14456), .o (n14457) );
  buffer buf_n14458( .i (n14457), .o (n14458) );
  buffer buf_n14459( .i (n14458), .o (n14459) );
  buffer buf_n14460( .i (n14459), .o (n14460) );
  buffer buf_n14461( .i (n14460), .o (n14461) );
  buffer buf_n14462( .i (n14461), .o (n14462) );
  buffer buf_n14463( .i (n14462), .o (n14463) );
  buffer buf_n14464( .i (n14463), .o (n14464) );
  buffer buf_n14465( .i (n14464), .o (n14465) );
  buffer buf_n14466( .i (n14465), .o (n14466) );
  buffer buf_n14467( .i (n14466), .o (n14467) );
  buffer buf_n14468( .i (n14467), .o (n14468) );
  buffer buf_n14469( .i (n14468), .o (n14469) );
  buffer buf_n14470( .i (n14469), .o (n14470) );
  buffer buf_n14471( .i (n14470), .o (n14471) );
  buffer buf_n14472( .i (n14471), .o (n14472) );
  buffer buf_n14473( .i (n14472), .o (n14473) );
  buffer buf_n14474( .i (n14473), .o (n14474) );
  buffer buf_n14475( .i (n14474), .o (n14475) );
  buffer buf_n14476( .i (n14475), .o (n14476) );
  buffer buf_n14477( .i (n14476), .o (n14477) );
  buffer buf_n14478( .i (n14477), .o (n14478) );
  buffer buf_n14479( .i (n14478), .o (n14479) );
  buffer buf_n14480( .i (n14479), .o (n14480) );
  buffer buf_n14481( .i (n14480), .o (n14481) );
  buffer buf_n14482( .i (n14481), .o (n14482) );
  buffer buf_n14483( .i (n14482), .o (n14483) );
  buffer buf_n14484( .i (n14483), .o (n14484) );
  buffer buf_n14485( .i (n14484), .o (n14485) );
  buffer buf_n14486( .i (n14485), .o (n14486) );
  buffer buf_n14487( .i (n14486), .o (n14487) );
  buffer buf_n14488( .i (n14487), .o (n14488) );
  buffer buf_n14489( .i (n14488), .o (n14489) );
  buffer buf_n14490( .i (n14489), .o (n14490) );
  buffer buf_n14491( .i (n14490), .o (n14491) );
  buffer buf_n14492( .i (n14491), .o (n14492) );
  buffer buf_n14493( .i (n14492), .o (n14493) );
  buffer buf_n14494( .i (n14493), .o (n14494) );
  buffer buf_n14495( .i (n14494), .o (n14495) );
  buffer buf_n14496( .i (n14495), .o (n14496) );
  buffer buf_n14497( .i (n14496), .o (n14497) );
  buffer buf_n14498( .i (n14497), .o (n14498) );
  buffer buf_n14499( .i (n14498), .o (n14499) );
  buffer buf_n14500( .i (n14499), .o (n14500) );
  buffer buf_n14501( .i (n14500), .o (n14501) );
  buffer buf_n14502( .i (n14501), .o (n14502) );
  buffer buf_n14503( .i (n14502), .o (n14503) );
  buffer buf_n14504( .i (n14503), .o (n14504) );
  buffer buf_n14505( .i (n14504), .o (n14505) );
  buffer buf_n14506( .i (n14505), .o (n14506) );
  buffer buf_n14507( .i (n14506), .o (n14507) );
  buffer buf_n14508( .i (n14507), .o (n14508) );
  buffer buf_n14509( .i (n14508), .o (n14509) );
  buffer buf_n14510( .i (n14509), .o (n14510) );
  buffer buf_n14511( .i (n14510), .o (n14511) );
  buffer buf_n14512( .i (n14511), .o (n14512) );
  buffer buf_n14513( .i (n14512), .o (n14513) );
  buffer buf_n14514( .i (n14513), .o (n14514) );
  buffer buf_n14515( .i (n14514), .o (n14515) );
  buffer buf_n14516( .i (n14515), .o (n14516) );
  buffer buf_n14517( .i (n14516), .o (n14517) );
  buffer buf_n14518( .i (n14517), .o (n14518) );
  buffer buf_n14519( .i (n14518), .o (n14519) );
  buffer buf_n14520( .i (n14519), .o (n14520) );
  buffer buf_n14521( .i (n14520), .o (n14521) );
  buffer buf_n14522( .i (n14521), .o (n14522) );
  buffer buf_n14523( .i (n14522), .o (n14523) );
  buffer buf_n14524( .i (n14523), .o (n14524) );
  buffer buf_n14525( .i (n14524), .o (n14525) );
  buffer buf_n14526( .i (n14525), .o (n14526) );
  buffer buf_n14527( .i (n14526), .o (n14527) );
  buffer buf_n14528( .i (n14527), .o (n14528) );
  buffer buf_n14529( .i (n14528), .o (n14529) );
  buffer buf_n14530( .i (n14529), .o (n14530) );
  buffer buf_n14531( .i (n14530), .o (n14531) );
  buffer buf_n14532( .i (n14531), .o (n14532) );
  buffer buf_n14533( .i (n14532), .o (n14533) );
  buffer buf_n14534( .i (n14533), .o (n14534) );
  buffer buf_n14535( .i (n14534), .o (n14535) );
  buffer buf_n14536( .i (n14535), .o (n14536) );
  buffer buf_n14537( .i (n14536), .o (n14537) );
  buffer buf_n14538( .i (n14537), .o (n14538) );
  buffer buf_n14539( .i (n14538), .o (n14539) );
  buffer buf_n14540( .i (n14539), .o (n14540) );
  buffer buf_n14541( .i (n14540), .o (n14541) );
  buffer buf_n14542( .i (n14541), .o (n14542) );
  buffer buf_n14543( .i (n14542), .o (n14543) );
  buffer buf_n14544( .i (n14543), .o (n14544) );
  buffer buf_n14545( .i (n14544), .o (n14545) );
  buffer buf_n14546( .i (n14545), .o (n14546) );
  buffer buf_n14547( .i (n14546), .o (n14547) );
  buffer buf_n14548( .i (n14547), .o (n14548) );
  buffer buf_n14549( .i (n14548), .o (n14549) );
  buffer buf_n14550( .i (n14549), .o (n14550) );
  buffer buf_n14551( .i (n14550), .o (n14551) );
  buffer buf_n14552( .i (n14551), .o (n14552) );
  assign n14553 = ~n5632 & n10090 ;
  buffer buf_n14554( .i (n13621), .o (n14554) );
  assign n14555 = n11697 & n14554 ;
  assign n14556 = n754 & ~n6053 ;
  buffer buf_n14557( .i (n14556), .o (n14557) );
  buffer buf_n2644( .i (n2643), .o (n2644) );
  buffer buf_n2645( .i (n2644), .o (n2645) );
  buffer buf_n2646( .i (n2645), .o (n2646) );
  buffer buf_n2647( .i (n2646), .o (n2647) );
  buffer buf_n2648( .i (n2647), .o (n2648) );
  buffer buf_n2649( .i (n2648), .o (n2649) );
  buffer buf_n2650( .i (n2649), .o (n2650) );
  buffer buf_n2651( .i (n2650), .o (n2651) );
  buffer buf_n2652( .i (n2651), .o (n2652) );
  buffer buf_n2653( .i (n2652), .o (n2653) );
  buffer buf_n2654( .i (n2653), .o (n2654) );
  assign n14558 = n2654 & n6077 ;
  assign n14559 = n14557 & ~n14558 ;
  buffer buf_n2655( .i (n2654), .o (n2655) );
  assign n14560 = n2655 & ~n14557 ;
  assign n14561 = n14559 | n14560 ;
  assign n14562 = n756 | n13399 ;
  assign n14563 = ~n6086 & n14562 ;
  assign n14564 = n14561 & n14563 ;
  buffer buf_n14565( .i (n14564), .o (n14565) );
  buffer buf_n14566( .i (n14565), .o (n14566) );
  buffer buf_n14567( .i (n14566), .o (n14567) );
  buffer buf_n14568( .i (n14567), .o (n14568) );
  buffer buf_n14569( .i (n14568), .o (n14569) );
  assign n14570 = n13975 | n14569 ;
  buffer buf_n14571( .i (n14570), .o (n14571) );
  buffer buf_n14572( .i (n14571), .o (n14572) );
  buffer buf_n14573( .i (n14572), .o (n14573) );
  buffer buf_n14574( .i (n14573), .o (n14574) );
  buffer buf_n14575( .i (n14574), .o (n14575) );
  buffer buf_n14576( .i (n14575), .o (n14576) );
  buffer buf_n14577( .i (n14576), .o (n14577) );
  buffer buf_n14578( .i (n14577), .o (n14578) );
  assign n14579 = n14555 | n14578 ;
  buffer buf_n14580( .i (n14579), .o (n14580) );
  assign n14581 = ~n11692 & n12168 ;
  assign n14582 = n12170 & ~n14581 ;
  assign n14583 = n14580 & n14582 ;
  assign n14584 = n14553 | n14583 ;
  buffer buf_n14585( .i (n14584), .o (n14585) );
  buffer buf_n14586( .i (n14585), .o (n14586) );
  buffer buf_n14587( .i (n14586), .o (n14587) );
  buffer buf_n14588( .i (n14587), .o (n14588) );
  buffer buf_n14589( .i (n14588), .o (n14589) );
  buffer buf_n14590( .i (n14589), .o (n14590) );
  buffer buf_n14591( .i (n14590), .o (n14591) );
  buffer buf_n14592( .i (n14591), .o (n14592) );
  buffer buf_n14593( .i (n14592), .o (n14593) );
  buffer buf_n14594( .i (n14593), .o (n14594) );
  buffer buf_n14595( .i (n14594), .o (n14595) );
  buffer buf_n14596( .i (n14595), .o (n14596) );
  buffer buf_n14597( .i (n14596), .o (n14597) );
  buffer buf_n14598( .i (n14597), .o (n14598) );
  buffer buf_n14599( .i (n14598), .o (n14599) );
  buffer buf_n14600( .i (n14599), .o (n14600) );
  buffer buf_n14601( .i (n14600), .o (n14601) );
  buffer buf_n14602( .i (n14601), .o (n14602) );
  buffer buf_n14603( .i (n14602), .o (n14603) );
  buffer buf_n14604( .i (n14603), .o (n14604) );
  buffer buf_n14605( .i (n14604), .o (n14605) );
  buffer buf_n14606( .i (n14605), .o (n14606) );
  buffer buf_n14607( .i (n14606), .o (n14607) );
  buffer buf_n14608( .i (n14607), .o (n14608) );
  buffer buf_n14609( .i (n14608), .o (n14609) );
  buffer buf_n14610( .i (n14609), .o (n14610) );
  buffer buf_n14611( .i (n14610), .o (n14611) );
  buffer buf_n14612( .i (n14611), .o (n14612) );
  buffer buf_n14613( .i (n14612), .o (n14613) );
  buffer buf_n14614( .i (n14613), .o (n14614) );
  buffer buf_n14615( .i (n14614), .o (n14615) );
  buffer buf_n14616( .i (n14615), .o (n14616) );
  buffer buf_n14617( .i (n14616), .o (n14617) );
  buffer buf_n14618( .i (n14617), .o (n14618) );
  buffer buf_n14619( .i (n14618), .o (n14619) );
  buffer buf_n14620( .i (n14619), .o (n14620) );
  buffer buf_n14621( .i (n14620), .o (n14621) );
  buffer buf_n14622( .i (n14621), .o (n14622) );
  buffer buf_n14623( .i (n14622), .o (n14623) );
  buffer buf_n14624( .i (n14623), .o (n14624) );
  buffer buf_n14625( .i (n14624), .o (n14625) );
  buffer buf_n14626( .i (n14625), .o (n14626) );
  buffer buf_n14627( .i (n14626), .o (n14627) );
  buffer buf_n14628( .i (n14627), .o (n14628) );
  buffer buf_n14629( .i (n14628), .o (n14629) );
  buffer buf_n14630( .i (n14629), .o (n14630) );
  buffer buf_n14631( .i (n14630), .o (n14631) );
  buffer buf_n14632( .i (n14631), .o (n14632) );
  buffer buf_n14633( .i (n14632), .o (n14633) );
  buffer buf_n14634( .i (n14633), .o (n14634) );
  buffer buf_n14635( .i (n14634), .o (n14635) );
  buffer buf_n14636( .i (n14635), .o (n14636) );
  buffer buf_n14637( .i (n14636), .o (n14637) );
  buffer buf_n14638( .i (n14637), .o (n14638) );
  buffer buf_n14639( .i (n14638), .o (n14639) );
  buffer buf_n14640( .i (n14639), .o (n14640) );
  buffer buf_n14641( .i (n14640), .o (n14641) );
  buffer buf_n14642( .i (n14641), .o (n14642) );
  buffer buf_n14643( .i (n14642), .o (n14643) );
  buffer buf_n14644( .i (n14643), .o (n14644) );
  buffer buf_n14645( .i (n14644), .o (n14645) );
  buffer buf_n14646( .i (n14645), .o (n14646) );
  buffer buf_n14647( .i (n14646), .o (n14647) );
  buffer buf_n14648( .i (n14647), .o (n14648) );
  buffer buf_n14649( .i (n14648), .o (n14649) );
  buffer buf_n14650( .i (n14649), .o (n14650) );
  buffer buf_n14651( .i (n14650), .o (n14651) );
  buffer buf_n14652( .i (n14651), .o (n14652) );
  buffer buf_n14653( .i (n14652), .o (n14653) );
  buffer buf_n14654( .i (n14653), .o (n14654) );
  buffer buf_n14655( .i (n14654), .o (n14655) );
  buffer buf_n14656( .i (n14655), .o (n14656) );
  buffer buf_n14657( .i (n14656), .o (n14657) );
  buffer buf_n14658( .i (n14657), .o (n14658) );
  buffer buf_n14659( .i (n14658), .o (n14659) );
  buffer buf_n14660( .i (n14659), .o (n14660) );
  buffer buf_n14661( .i (n14660), .o (n14661) );
  buffer buf_n14662( .i (n14661), .o (n14662) );
  buffer buf_n14663( .i (n14662), .o (n14663) );
  buffer buf_n14664( .i (n14663), .o (n14664) );
  buffer buf_n14665( .i (n14664), .o (n14665) );
  buffer buf_n14666( .i (n14665), .o (n14666) );
  buffer buf_n14667( .i (n14666), .o (n14667) );
  buffer buf_n14668( .i (n14667), .o (n14668) );
  buffer buf_n14669( .i (n14668), .o (n14669) );
  buffer buf_n14670( .i (n14669), .o (n14670) );
  buffer buf_n14671( .i (n14670), .o (n14671) );
  buffer buf_n14672( .i (n14671), .o (n14672) );
  buffer buf_n14673( .i (n14672), .o (n14673) );
  buffer buf_n14674( .i (n14673), .o (n14674) );
  buffer buf_n14675( .i (n14674), .o (n14675) );
  buffer buf_n14676( .i (n14675), .o (n14676) );
  buffer buf_n14677( .i (n14676), .o (n14677) );
  buffer buf_n14678( .i (n14677), .o (n14678) );
  buffer buf_n14679( .i (n14678), .o (n14679) );
  buffer buf_n14680( .i (n14679), .o (n14680) );
  buffer buf_n14681( .i (n14680), .o (n14681) );
  buffer buf_n14682( .i (n14681), .o (n14682) );
  buffer buf_n14683( .i (n14682), .o (n14683) );
  buffer buf_n14684( .i (n14683), .o (n14684) );
  buffer buf_n14685( .i (n14684), .o (n14685) );
  buffer buf_n14686( .i (n14685), .o (n14686) );
  buffer buf_n14687( .i (n14686), .o (n14687) );
  buffer buf_n14688( .i (n14687), .o (n14688) );
  buffer buf_n14689( .i (n14688), .o (n14689) );
  buffer buf_n14690( .i (n14689), .o (n14690) );
  buffer buf_n14691( .i (n14690), .o (n14691) );
  buffer buf_n14692( .i (n14691), .o (n14692) );
  buffer buf_n14693( .i (n14692), .o (n14693) );
  buffer buf_n14694( .i (n14693), .o (n14694) );
  buffer buf_n14695( .i (n14694), .o (n14695) );
  buffer buf_n12796( .i (n12795), .o (n12796) );
  buffer buf_n12797( .i (n12796), .o (n12797) );
  buffer buf_n12798( .i (n12797), .o (n12798) );
  buffer buf_n12799( .i (n12798), .o (n12799) );
  buffer buf_n12800( .i (n12799), .o (n12800) );
  buffer buf_n12801( .i (n12800), .o (n12801) );
  buffer buf_n12802( .i (n12801), .o (n12802) );
  buffer buf_n12803( .i (n12802), .o (n12803) );
  buffer buf_n12804( .i (n12803), .o (n12804) );
  buffer buf_n12805( .i (n12804), .o (n12805) );
  buffer buf_n12806( .i (n12805), .o (n12806) );
  buffer buf_n12807( .i (n12806), .o (n12807) );
  buffer buf_n12808( .i (n12807), .o (n12808) );
  buffer buf_n12809( .i (n12808), .o (n12809) );
  buffer buf_n12810( .i (n12809), .o (n12810) );
  buffer buf_n12811( .i (n12810), .o (n12811) );
  buffer buf_n12812( .i (n12811), .o (n12812) );
  buffer buf_n12813( .i (n12812), .o (n12813) );
  buffer buf_n12814( .i (n12813), .o (n12814) );
  buffer buf_n12815( .i (n12814), .o (n12815) );
  buffer buf_n12816( .i (n12815), .o (n12816) );
  buffer buf_n12817( .i (n12816), .o (n12817) );
  buffer buf_n12818( .i (n12817), .o (n12818) );
  buffer buf_n12819( .i (n12818), .o (n12819) );
  buffer buf_n12820( .i (n12819), .o (n12820) );
  buffer buf_n12821( .i (n12820), .o (n12821) );
  buffer buf_n12822( .i (n12821), .o (n12822) );
  buffer buf_n12823( .i (n12822), .o (n12823) );
  buffer buf_n12824( .i (n12823), .o (n12824) );
  buffer buf_n12825( .i (n12824), .o (n12825) );
  buffer buf_n12826( .i (n12825), .o (n12826) );
  buffer buf_n12827( .i (n12826), .o (n12827) );
  buffer buf_n12828( .i (n12827), .o (n12828) );
  buffer buf_n12829( .i (n12828), .o (n12829) );
  buffer buf_n12830( .i (n12829), .o (n12830) );
  buffer buf_n12831( .i (n12830), .o (n12831) );
  buffer buf_n12832( .i (n12831), .o (n12832) );
  buffer buf_n12833( .i (n12832), .o (n12833) );
  buffer buf_n12834( .i (n12833), .o (n12834) );
  buffer buf_n12835( .i (n12834), .o (n12835) );
  buffer buf_n12836( .i (n12835), .o (n12836) );
  buffer buf_n12837( .i (n12836), .o (n12837) );
  buffer buf_n12838( .i (n12837), .o (n12838) );
  buffer buf_n12839( .i (n12838), .o (n12839) );
  buffer buf_n12840( .i (n12839), .o (n12840) );
  buffer buf_n12841( .i (n12840), .o (n12841) );
  buffer buf_n12842( .i (n12841), .o (n12842) );
  buffer buf_n12843( .i (n12842), .o (n12843) );
  buffer buf_n12844( .i (n12843), .o (n12844) );
  buffer buf_n12845( .i (n12844), .o (n12845) );
  buffer buf_n12846( .i (n12845), .o (n12846) );
  buffer buf_n12847( .i (n12846), .o (n12847) );
  buffer buf_n12848( .i (n12847), .o (n12848) );
  buffer buf_n12849( .i (n12848), .o (n12849) );
  buffer buf_n12850( .i (n12849), .o (n12850) );
  buffer buf_n12851( .i (n12850), .o (n12851) );
  buffer buf_n12852( .i (n12851), .o (n12852) );
  buffer buf_n12853( .i (n12852), .o (n12853) );
  buffer buf_n12854( .i (n12853), .o (n12854) );
  buffer buf_n12855( .i (n12854), .o (n12855) );
  buffer buf_n12856( .i (n12855), .o (n12856) );
  buffer buf_n12857( .i (n12856), .o (n12857) );
  buffer buf_n12858( .i (n12857), .o (n12858) );
  buffer buf_n12859( .i (n12858), .o (n12859) );
  buffer buf_n12860( .i (n12859), .o (n12860) );
  buffer buf_n12861( .i (n12860), .o (n12861) );
  buffer buf_n12862( .i (n12861), .o (n12862) );
  buffer buf_n12863( .i (n12862), .o (n12863) );
  buffer buf_n12864( .i (n12863), .o (n12864) );
  buffer buf_n12865( .i (n12864), .o (n12865) );
  buffer buf_n12866( .i (n12865), .o (n12866) );
  buffer buf_n12867( .i (n12866), .o (n12867) );
  buffer buf_n12868( .i (n12867), .o (n12868) );
  buffer buf_n12869( .i (n12868), .o (n12869) );
  buffer buf_n12870( .i (n12869), .o (n12870) );
  buffer buf_n12871( .i (n12870), .o (n12871) );
  buffer buf_n12872( .i (n12871), .o (n12872) );
  buffer buf_n12873( .i (n12872), .o (n12873) );
  buffer buf_n12874( .i (n12873), .o (n12874) );
  buffer buf_n12875( .i (n12874), .o (n12875) );
  buffer buf_n12876( .i (n12875), .o (n12876) );
  buffer buf_n12877( .i (n12876), .o (n12877) );
  buffer buf_n12878( .i (n12877), .o (n12878) );
  buffer buf_n12879( .i (n12878), .o (n12879) );
  buffer buf_n12880( .i (n12879), .o (n12880) );
  buffer buf_n12881( .i (n12880), .o (n12881) );
  buffer buf_n12882( .i (n12881), .o (n12882) );
  buffer buf_n12883( .i (n12882), .o (n12883) );
  buffer buf_n12884( .i (n12883), .o (n12884) );
  buffer buf_n12885( .i (n12884), .o (n12885) );
  buffer buf_n12886( .i (n12885), .o (n12886) );
  buffer buf_n12887( .i (n12886), .o (n12887) );
  buffer buf_n12888( .i (n12887), .o (n12888) );
  buffer buf_n12889( .i (n12888), .o (n12889) );
  buffer buf_n12890( .i (n12889), .o (n12890) );
  buffer buf_n12891( .i (n12890), .o (n12891) );
  buffer buf_n12892( .i (n12891), .o (n12892) );
  buffer buf_n12893( .i (n12892), .o (n12893) );
  buffer buf_n12894( .i (n12893), .o (n12894) );
  buffer buf_n12895( .i (n12894), .o (n12895) );
  buffer buf_n12896( .i (n12895), .o (n12896) );
  buffer buf_n12897( .i (n12896), .o (n12897) );
  buffer buf_n12898( .i (n12897), .o (n12898) );
  buffer buf_n12899( .i (n12898), .o (n12899) );
  buffer buf_n12900( .i (n12899), .o (n12900) );
  buffer buf_n12901( .i (n12900), .o (n12901) );
  buffer buf_n12902( .i (n12901), .o (n12902) );
  buffer buf_n12903( .i (n12902), .o (n12903) );
  buffer buf_n12904( .i (n12903), .o (n12904) );
  buffer buf_n12905( .i (n12904), .o (n12905) );
  buffer buf_n12906( .i (n12905), .o (n12906) );
  buffer buf_n12907( .i (n12906), .o (n12907) );
  buffer buf_n12908( .i (n12907), .o (n12908) );
  buffer buf_n12909( .i (n12908), .o (n12909) );
  buffer buf_n14696( .i (n13392), .o (n14696) );
  assign n14697 = n10507 & ~n14696 ;
  assign n14698 = ~n6292 & n12168 ;
  assign n14699 = n12170 & ~n14698 ;
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  buffer buf_n1813( .i (n1812), .o (n1813) );
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  assign n14700 = n1816 & n10914 ;
  buffer buf_n14701( .i (n6052), .o (n14701) );
  assign n14702 = n3267 & ~n14701 ;
  buffer buf_n14703( .i (n14702), .o (n14703) );
  buffer buf_n14704( .i (n14703), .o (n14704) );
  assign n14705 = ~n14700 & n14704 ;
  assign n14706 = n3269 | n13399 ;
  assign n14707 = n1816 & ~n14703 ;
  assign n14708 = n14706 & n14707 ;
  assign n14709 = n14705 | n14708 ;
  buffer buf_n14710( .i (n14709), .o (n14710) );
  buffer buf_n14711( .i (n14710), .o (n14711) );
  buffer buf_n14712( .i (n10767), .o (n14712) );
  buffer buf_n14713( .i (n14712), .o (n14713) );
  assign n14714 = n14711 & ~n14713 ;
  buffer buf_n14715( .i (n14714), .o (n14715) );
  buffer buf_n14716( .i (n14715), .o (n14716) );
  buffer buf_n14717( .i (n11669), .o (n14717) );
  assign n14718 = n14716 | n14717 ;
  buffer buf_n14719( .i (n14718), .o (n14719) );
  buffer buf_n14720( .i (n14719), .o (n14720) );
  buffer buf_n14721( .i (n14720), .o (n14721) );
  buffer buf_n14722( .i (n14721), .o (n14722) );
  buffer buf_n14723( .i (n14722), .o (n14723) );
  buffer buf_n14724( .i (n14723), .o (n14724) );
  buffer buf_n14725( .i (n14724), .o (n14725) );
  buffer buf_n14726( .i (n14725), .o (n14726) );
  assign n14727 = n6047 & n14554 ;
  assign n14728 = n14726 | n14727 ;
  buffer buf_n14729( .i (n14728), .o (n14729) );
  assign n14730 = n14699 & n14729 ;
  assign n14731 = n14697 | n14730 ;
  buffer buf_n14732( .i (n14731), .o (n14732) );
  buffer buf_n14733( .i (n14732), .o (n14733) );
  buffer buf_n14734( .i (n14733), .o (n14734) );
  buffer buf_n14735( .i (n14734), .o (n14735) );
  buffer buf_n14736( .i (n14735), .o (n14736) );
  buffer buf_n14737( .i (n14736), .o (n14737) );
  buffer buf_n14738( .i (n14737), .o (n14738) );
  buffer buf_n14739( .i (n14738), .o (n14739) );
  buffer buf_n14740( .i (n14739), .o (n14740) );
  buffer buf_n14741( .i (n14740), .o (n14741) );
  buffer buf_n14742( .i (n14741), .o (n14742) );
  buffer buf_n14743( .i (n14742), .o (n14743) );
  buffer buf_n14744( .i (n14743), .o (n14744) );
  buffer buf_n14745( .i (n14744), .o (n14745) );
  buffer buf_n14746( .i (n14745), .o (n14746) );
  buffer buf_n14747( .i (n14746), .o (n14747) );
  buffer buf_n14748( .i (n14747), .o (n14748) );
  buffer buf_n14749( .i (n14748), .o (n14749) );
  buffer buf_n14750( .i (n14749), .o (n14750) );
  buffer buf_n14751( .i (n14750), .o (n14751) );
  buffer buf_n14752( .i (n14751), .o (n14752) );
  buffer buf_n14753( .i (n14752), .o (n14753) );
  buffer buf_n14754( .i (n14753), .o (n14754) );
  buffer buf_n14755( .i (n14754), .o (n14755) );
  buffer buf_n14756( .i (n14755), .o (n14756) );
  buffer buf_n14757( .i (n14756), .o (n14757) );
  buffer buf_n14758( .i (n14757), .o (n14758) );
  buffer buf_n14759( .i (n14758), .o (n14759) );
  buffer buf_n14760( .i (n14759), .o (n14760) );
  buffer buf_n14761( .i (n14760), .o (n14761) );
  buffer buf_n14762( .i (n14761), .o (n14762) );
  buffer buf_n14763( .i (n14762), .o (n14763) );
  buffer buf_n14764( .i (n14763), .o (n14764) );
  buffer buf_n14765( .i (n14764), .o (n14765) );
  buffer buf_n14766( .i (n14765), .o (n14766) );
  buffer buf_n14767( .i (n14766), .o (n14767) );
  buffer buf_n14768( .i (n14767), .o (n14768) );
  buffer buf_n14769( .i (n14768), .o (n14769) );
  buffer buf_n14770( .i (n14769), .o (n14770) );
  buffer buf_n14771( .i (n14770), .o (n14771) );
  buffer buf_n14772( .i (n14771), .o (n14772) );
  buffer buf_n14773( .i (n14772), .o (n14773) );
  buffer buf_n14774( .i (n14773), .o (n14774) );
  buffer buf_n14775( .i (n14774), .o (n14775) );
  buffer buf_n14776( .i (n14775), .o (n14776) );
  buffer buf_n14777( .i (n14776), .o (n14777) );
  buffer buf_n14778( .i (n14777), .o (n14778) );
  buffer buf_n14779( .i (n14778), .o (n14779) );
  buffer buf_n14780( .i (n14779), .o (n14780) );
  buffer buf_n14781( .i (n14780), .o (n14781) );
  buffer buf_n14782( .i (n14781), .o (n14782) );
  buffer buf_n14783( .i (n14782), .o (n14783) );
  buffer buf_n14784( .i (n14783), .o (n14784) );
  buffer buf_n14785( .i (n14784), .o (n14785) );
  buffer buf_n14786( .i (n14785), .o (n14786) );
  buffer buf_n14787( .i (n14786), .o (n14787) );
  buffer buf_n14788( .i (n14787), .o (n14788) );
  buffer buf_n14789( .i (n14788), .o (n14789) );
  buffer buf_n14790( .i (n14789), .o (n14790) );
  buffer buf_n14791( .i (n14790), .o (n14791) );
  buffer buf_n14792( .i (n14791), .o (n14792) );
  buffer buf_n14793( .i (n14792), .o (n14793) );
  buffer buf_n14794( .i (n14793), .o (n14794) );
  buffer buf_n14795( .i (n14794), .o (n14795) );
  buffer buf_n14796( .i (n14795), .o (n14796) );
  buffer buf_n14797( .i (n14796), .o (n14797) );
  buffer buf_n14798( .i (n14797), .o (n14798) );
  buffer buf_n14799( .i (n14798), .o (n14799) );
  buffer buf_n14800( .i (n14799), .o (n14800) );
  buffer buf_n14801( .i (n14800), .o (n14801) );
  buffer buf_n14802( .i (n14801), .o (n14802) );
  buffer buf_n14803( .i (n14802), .o (n14803) );
  buffer buf_n14804( .i (n14803), .o (n14804) );
  buffer buf_n14805( .i (n14804), .o (n14805) );
  buffer buf_n14806( .i (n14805), .o (n14806) );
  buffer buf_n14807( .i (n14806), .o (n14807) );
  buffer buf_n14808( .i (n14807), .o (n14808) );
  buffer buf_n14809( .i (n14808), .o (n14809) );
  buffer buf_n14810( .i (n14809), .o (n14810) );
  buffer buf_n14811( .i (n14810), .o (n14811) );
  buffer buf_n14812( .i (n14811), .o (n14812) );
  buffer buf_n14813( .i (n14812), .o (n14813) );
  buffer buf_n14814( .i (n14813), .o (n14814) );
  buffer buf_n14815( .i (n14814), .o (n14815) );
  buffer buf_n14816( .i (n14815), .o (n14816) );
  buffer buf_n14817( .i (n14816), .o (n14817) );
  buffer buf_n14818( .i (n14817), .o (n14818) );
  buffer buf_n14819( .i (n14818), .o (n14819) );
  buffer buf_n14820( .i (n14819), .o (n14820) );
  buffer buf_n14821( .i (n14820), .o (n14821) );
  buffer buf_n14822( .i (n14821), .o (n14822) );
  buffer buf_n14823( .i (n14822), .o (n14823) );
  buffer buf_n14824( .i (n14823), .o (n14824) );
  buffer buf_n14825( .i (n14824), .o (n14825) );
  buffer buf_n14826( .i (n14825), .o (n14826) );
  buffer buf_n14827( .i (n14826), .o (n14827) );
  buffer buf_n14828( .i (n14827), .o (n14828) );
  buffer buf_n14829( .i (n14828), .o (n14829) );
  buffer buf_n14830( .i (n14829), .o (n14830) );
  buffer buf_n14831( .i (n14830), .o (n14831) );
  buffer buf_n14832( .i (n14831), .o (n14832) );
  buffer buf_n14833( .i (n14832), .o (n14833) );
  buffer buf_n14834( .i (n14833), .o (n14834) );
  buffer buf_n14835( .i (n14834), .o (n14835) );
  buffer buf_n14836( .i (n14835), .o (n14836) );
  buffer buf_n14837( .i (n14836), .o (n14837) );
  buffer buf_n14838( .i (n14837), .o (n14838) );
  buffer buf_n14839( .i (n14838), .o (n14839) );
  buffer buf_n14840( .i (n14839), .o (n14840) );
  buffer buf_n14841( .i (n14840), .o (n14841) );
  buffer buf_n14842( .i (n14841), .o (n14842) );
  buffer buf_n14232( .i (n14231), .o (n14232) );
  buffer buf_n14233( .i (n14232), .o (n14233) );
  buffer buf_n14234( .i (n14233), .o (n14234) );
  buffer buf_n14235( .i (n14234), .o (n14235) );
  buffer buf_n14236( .i (n14235), .o (n14236) );
  buffer buf_n14237( .i (n14236), .o (n14237) );
  buffer buf_n14238( .i (n14237), .o (n14238) );
  buffer buf_n14239( .i (n14238), .o (n14239) );
  buffer buf_n14240( .i (n14239), .o (n14240) );
  buffer buf_n14241( .i (n14240), .o (n14241) );
  buffer buf_n14242( .i (n14241), .o (n14242) );
  buffer buf_n14243( .i (n14242), .o (n14243) );
  buffer buf_n14244( .i (n14243), .o (n14244) );
  buffer buf_n14245( .i (n14244), .o (n14245) );
  buffer buf_n14246( .i (n14245), .o (n14246) );
  buffer buf_n14247( .i (n14246), .o (n14247) );
  buffer buf_n14248( .i (n14247), .o (n14248) );
  buffer buf_n14249( .i (n14248), .o (n14249) );
  buffer buf_n11002( .i (n11001), .o (n11002) );
  buffer buf_n11003( .i (n11002), .o (n11003) );
  buffer buf_n11004( .i (n11003), .o (n11004) );
  buffer buf_n11005( .i (n11004), .o (n11005) );
  buffer buf_n11006( .i (n11005), .o (n11006) );
  buffer buf_n11007( .i (n11006), .o (n11007) );
  buffer buf_n11008( .i (n11007), .o (n11008) );
  buffer buf_n11009( .i (n11008), .o (n11009) );
  buffer buf_n11010( .i (n11009), .o (n11010) );
  buffer buf_n11011( .i (n11010), .o (n11011) );
  buffer buf_n11012( .i (n11011), .o (n11012) );
  buffer buf_n11013( .i (n11012), .o (n11013) );
  buffer buf_n11014( .i (n11013), .o (n11014) );
  buffer buf_n11015( .i (n11014), .o (n11015) );
  buffer buf_n11016( .i (n11015), .o (n11016) );
  buffer buf_n11017( .i (n11016), .o (n11017) );
  buffer buf_n11018( .i (n11017), .o (n11018) );
  buffer buf_n11019( .i (n11018), .o (n11019) );
  buffer buf_n11020( .i (n11019), .o (n11020) );
  buffer buf_n11021( .i (n11020), .o (n11021) );
  buffer buf_n11022( .i (n11021), .o (n11022) );
  buffer buf_n11023( .i (n11022), .o (n11023) );
  buffer buf_n11024( .i (n11023), .o (n11024) );
  buffer buf_n11025( .i (n11024), .o (n11025) );
  buffer buf_n11026( .i (n11025), .o (n11026) );
  buffer buf_n11027( .i (n11026), .o (n11027) );
  buffer buf_n11028( .i (n11027), .o (n11028) );
  buffer buf_n11029( .i (n11028), .o (n11029) );
  buffer buf_n11030( .i (n11029), .o (n11030) );
  buffer buf_n11031( .i (n11030), .o (n11031) );
  buffer buf_n11032( .i (n11031), .o (n11032) );
  buffer buf_n11033( .i (n11032), .o (n11033) );
  buffer buf_n11034( .i (n11033), .o (n11034) );
  buffer buf_n11035( .i (n11034), .o (n11035) );
  buffer buf_n11036( .i (n11035), .o (n11036) );
  buffer buf_n11037( .i (n11036), .o (n11037) );
  buffer buf_n11038( .i (n11037), .o (n11038) );
  buffer buf_n11039( .i (n11038), .o (n11039) );
  buffer buf_n11040( .i (n11039), .o (n11040) );
  buffer buf_n11041( .i (n11040), .o (n11041) );
  buffer buf_n11042( .i (n11041), .o (n11042) );
  buffer buf_n11043( .i (n11042), .o (n11043) );
  buffer buf_n11044( .i (n11043), .o (n11044) );
  buffer buf_n11045( .i (n11044), .o (n11045) );
  buffer buf_n11046( .i (n11045), .o (n11046) );
  buffer buf_n11047( .i (n11046), .o (n11047) );
  buffer buf_n11048( .i (n11047), .o (n11048) );
  buffer buf_n11049( .i (n11048), .o (n11049) );
  buffer buf_n11050( .i (n11049), .o (n11050) );
  buffer buf_n11051( .i (n11050), .o (n11051) );
  buffer buf_n11052( .i (n11051), .o (n11052) );
  buffer buf_n11053( .i (n11052), .o (n11053) );
  buffer buf_n11054( .i (n11053), .o (n11054) );
  buffer buf_n11055( .i (n11054), .o (n11055) );
  buffer buf_n9984( .i (n9983), .o (n9984) );
  buffer buf_n9985( .i (n9984), .o (n9985) );
  buffer buf_n9986( .i (n9985), .o (n9986) );
  buffer buf_n9987( .i (n9986), .o (n9987) );
  buffer buf_n9988( .i (n9987), .o (n9988) );
  buffer buf_n9989( .i (n9988), .o (n9989) );
  buffer buf_n9990( .i (n9989), .o (n9990) );
  buffer buf_n9991( .i (n9990), .o (n9991) );
  buffer buf_n9992( .i (n9991), .o (n9992) );
  buffer buf_n9993( .i (n9992), .o (n9993) );
  buffer buf_n9994( .i (n9993), .o (n9994) );
  buffer buf_n9995( .i (n9994), .o (n9995) );
  buffer buf_n9996( .i (n9995), .o (n9996) );
  buffer buf_n9997( .i (n9996), .o (n9997) );
  buffer buf_n9998( .i (n9997), .o (n9998) );
  buffer buf_n9999( .i (n9998), .o (n9999) );
  buffer buf_n10000( .i (n9999), .o (n10000) );
  buffer buf_n10001( .i (n10000), .o (n10001) );
  buffer buf_n10002( .i (n10001), .o (n10002) );
  buffer buf_n10003( .i (n10002), .o (n10003) );
  buffer buf_n10004( .i (n10003), .o (n10004) );
  buffer buf_n10005( .i (n10004), .o (n10005) );
  buffer buf_n10006( .i (n10005), .o (n10006) );
  buffer buf_n10007( .i (n10006), .o (n10007) );
  buffer buf_n10008( .i (n10007), .o (n10008) );
  buffer buf_n10009( .i (n10008), .o (n10009) );
  buffer buf_n10010( .i (n10009), .o (n10010) );
  buffer buf_n10011( .i (n10010), .o (n10011) );
  buffer buf_n10012( .i (n10011), .o (n10012) );
  buffer buf_n10013( .i (n10012), .o (n10013) );
  buffer buf_n10014( .i (n10013), .o (n10014) );
  buffer buf_n10015( .i (n10014), .o (n10015) );
  buffer buf_n10016( .i (n10015), .o (n10016) );
  buffer buf_n10017( .i (n10016), .o (n10017) );
  buffer buf_n10018( .i (n10017), .o (n10018) );
  buffer buf_n10019( .i (n10018), .o (n10019) );
  buffer buf_n10020( .i (n10019), .o (n10020) );
  buffer buf_n10021( .i (n10020), .o (n10021) );
  buffer buf_n10022( .i (n10021), .o (n10022) );
  assign n14843 = ~n5733 & n13767 ;
  assign n14844 = n11508 & n14554 ;
  assign n14845 = n2693 & n2995 ;
  buffer buf_n14846( .i (n14845), .o (n14846) );
  buffer buf_n14847( .i (n14846), .o (n14847) );
  assign n14848 = n14307 & ~n14847 ;
  assign n14849 = n14712 | n14848 ;
  assign n14850 = n2694 & n14104 ;
  assign n14851 = n2997 | n14850 ;
  assign n14852 = n14110 & n14846 ;
  assign n14853 = n14851 & ~n14852 ;
  assign n14854 = n14308 | n14853 ;
  assign n14855 = ~n14849 & n14854 ;
  buffer buf_n14856( .i (n14855), .o (n14856) );
  buffer buf_n14857( .i (n14856), .o (n14857) );
  assign n14858 = n14717 | n14857 ;
  buffer buf_n14859( .i (n14858), .o (n14859) );
  buffer buf_n14860( .i (n14859), .o (n14860) );
  buffer buf_n14861( .i (n14860), .o (n14861) );
  buffer buf_n14862( .i (n14861), .o (n14862) );
  buffer buf_n14863( .i (n14862), .o (n14863) );
  buffer buf_n14864( .i (n14863), .o (n14864) );
  buffer buf_n14865( .i (n14864), .o (n14865) );
  buffer buf_n14866( .i (n14865), .o (n14866) );
  assign n14867 = n14844 | n14866 ;
  buffer buf_n14868( .i (n14867), .o (n14868) );
  assign n14869 = ~n11540 & n12168 ;
  assign n14870 = n12170 & ~n14869 ;
  assign n14871 = n14868 & n14870 ;
  buffer buf_n14872( .i (n14871), .o (n14872) );
  buffer buf_n14873( .i (n14872), .o (n14873) );
  buffer buf_n14874( .i (n14873), .o (n14874) );
  buffer buf_n14875( .i (n14874), .o (n14875) );
  buffer buf_n14876( .i (n14875), .o (n14876) );
  buffer buf_n14877( .i (n14876), .o (n14877) );
  buffer buf_n14878( .i (n14877), .o (n14878) );
  buffer buf_n14879( .i (n14878), .o (n14879) );
  buffer buf_n14880( .i (n14879), .o (n14880) );
  buffer buf_n14881( .i (n14880), .o (n14881) );
  buffer buf_n14882( .i (n14881), .o (n14882) );
  buffer buf_n14883( .i (n14882), .o (n14883) );
  buffer buf_n14884( .i (n14883), .o (n14884) );
  buffer buf_n14885( .i (n14884), .o (n14885) );
  buffer buf_n14886( .i (n14885), .o (n14886) );
  buffer buf_n14887( .i (n14886), .o (n14887) );
  buffer buf_n14888( .i (n14887), .o (n14888) );
  buffer buf_n14889( .i (n14888), .o (n14889) );
  buffer buf_n14890( .i (n14889), .o (n14890) );
  buffer buf_n14891( .i (n14890), .o (n14891) );
  buffer buf_n14892( .i (n14891), .o (n14892) );
  buffer buf_n14893( .i (n14892), .o (n14893) );
  buffer buf_n14894( .i (n14893), .o (n14894) );
  buffer buf_n14895( .i (n14894), .o (n14895) );
  buffer buf_n14896( .i (n14895), .o (n14896) );
  buffer buf_n14897( .i (n14896), .o (n14897) );
  buffer buf_n14898( .i (n14897), .o (n14898) );
  buffer buf_n14899( .i (n14898), .o (n14899) );
  buffer buf_n14900( .i (n14899), .o (n14900) );
  buffer buf_n14901( .i (n14900), .o (n14901) );
  buffer buf_n14902( .i (n14901), .o (n14902) );
  buffer buf_n14903( .i (n14902), .o (n14903) );
  buffer buf_n14904( .i (n14903), .o (n14904) );
  buffer buf_n14905( .i (n14904), .o (n14905) );
  buffer buf_n14906( .i (n14905), .o (n14906) );
  buffer buf_n14907( .i (n14906), .o (n14907) );
  buffer buf_n14908( .i (n14907), .o (n14908) );
  buffer buf_n14909( .i (n14908), .o (n14909) );
  buffer buf_n14910( .i (n14909), .o (n14910) );
  buffer buf_n14911( .i (n14910), .o (n14911) );
  buffer buf_n14912( .i (n14911), .o (n14912) );
  buffer buf_n14913( .i (n14912), .o (n14913) );
  buffer buf_n14914( .i (n14913), .o (n14914) );
  buffer buf_n14915( .i (n14914), .o (n14915) );
  buffer buf_n14916( .i (n14915), .o (n14916) );
  buffer buf_n14917( .i (n14916), .o (n14917) );
  buffer buf_n14918( .i (n14917), .o (n14918) );
  buffer buf_n14919( .i (n14918), .o (n14919) );
  buffer buf_n14920( .i (n14919), .o (n14920) );
  buffer buf_n14921( .i (n14920), .o (n14921) );
  buffer buf_n14922( .i (n14921), .o (n14922) );
  buffer buf_n14923( .i (n14922), .o (n14923) );
  buffer buf_n14924( .i (n14923), .o (n14924) );
  buffer buf_n14925( .i (n14924), .o (n14925) );
  buffer buf_n14926( .i (n14925), .o (n14926) );
  buffer buf_n14927( .i (n14926), .o (n14927) );
  buffer buf_n14928( .i (n14927), .o (n14928) );
  buffer buf_n14929( .i (n14928), .o (n14929) );
  buffer buf_n14930( .i (n14929), .o (n14930) );
  buffer buf_n14931( .i (n14930), .o (n14931) );
  buffer buf_n14932( .i (n14931), .o (n14932) );
  buffer buf_n14933( .i (n14932), .o (n14933) );
  buffer buf_n14934( .i (n14933), .o (n14934) );
  buffer buf_n14935( .i (n14934), .o (n14935) );
  buffer buf_n14936( .i (n14935), .o (n14936) );
  buffer buf_n14937( .i (n14936), .o (n14937) );
  buffer buf_n14938( .i (n14937), .o (n14938) );
  buffer buf_n14939( .i (n14938), .o (n14939) );
  buffer buf_n14940( .i (n14939), .o (n14940) );
  buffer buf_n14941( .i (n14940), .o (n14941) );
  buffer buf_n14942( .i (n14941), .o (n14942) );
  buffer buf_n14943( .i (n14942), .o (n14943) );
  buffer buf_n14944( .i (n14943), .o (n14944) );
  buffer buf_n14945( .i (n14944), .o (n14945) );
  buffer buf_n14946( .i (n14945), .o (n14946) );
  buffer buf_n14947( .i (n14946), .o (n14947) );
  buffer buf_n14948( .i (n14947), .o (n14948) );
  buffer buf_n14949( .i (n14948), .o (n14949) );
  buffer buf_n14950( .i (n14949), .o (n14950) );
  buffer buf_n14951( .i (n14950), .o (n14951) );
  buffer buf_n14952( .i (n14951), .o (n14952) );
  buffer buf_n14953( .i (n14952), .o (n14953) );
  buffer buf_n14954( .i (n14953), .o (n14954) );
  buffer buf_n14955( .i (n14954), .o (n14955) );
  buffer buf_n14956( .i (n14955), .o (n14956) );
  buffer buf_n14957( .i (n14956), .o (n14957) );
  buffer buf_n14958( .i (n14957), .o (n14958) );
  buffer buf_n14959( .i (n14958), .o (n14959) );
  buffer buf_n14960( .i (n14959), .o (n14960) );
  buffer buf_n14961( .i (n14960), .o (n14961) );
  buffer buf_n14962( .i (n14961), .o (n14962) );
  buffer buf_n14963( .i (n14962), .o (n14963) );
  buffer buf_n14964( .i (n14963), .o (n14964) );
  buffer buf_n14965( .i (n14964), .o (n14965) );
  buffer buf_n14966( .i (n14965), .o (n14966) );
  buffer buf_n14967( .i (n14966), .o (n14967) );
  buffer buf_n14968( .i (n14967), .o (n14968) );
  buffer buf_n14969( .i (n14968), .o (n14969) );
  buffer buf_n14970( .i (n14969), .o (n14970) );
  buffer buf_n14971( .i (n14970), .o (n14971) );
  buffer buf_n14972( .i (n14971), .o (n14972) );
  assign n14973 = n14843 | n14972 ;
  buffer buf_n14974( .i (n14973), .o (n14974) );
  buffer buf_n14975( .i (n14974), .o (n14975) );
  buffer buf_n14976( .i (n14975), .o (n14976) );
  buffer buf_n14977( .i (n14976), .o (n14977) );
  buffer buf_n14978( .i (n14977), .o (n14978) );
  buffer buf_n14979( .i (n14978), .o (n14979) );
  buffer buf_n14980( .i (n14979), .o (n14980) );
  buffer buf_n14981( .i (n14980), .o (n14981) );
  buffer buf_n14982( .i (n14981), .o (n14982) );
  buffer buf_n14983( .i (n14982), .o (n14983) );
  buffer buf_n14273( .i (n14272), .o (n14273) );
  buffer buf_n14274( .i (n14273), .o (n14274) );
  buffer buf_n14275( .i (n14274), .o (n14275) );
  buffer buf_n14276( .i (n14275), .o (n14276) );
  buffer buf_n14277( .i (n14276), .o (n14277) );
  buffer buf_n14278( .i (n14277), .o (n14278) );
  buffer buf_n14279( .i (n14278), .o (n14279) );
  buffer buf_n14280( .i (n14279), .o (n14280) );
  buffer buf_n14281( .i (n14280), .o (n14281) );
  buffer buf_n14282( .i (n14281), .o (n14282) );
  buffer buf_n14283( .i (n14282), .o (n14283) );
  buffer buf_n14284( .i (n14283), .o (n14284) );
  buffer buf_n14285( .i (n14284), .o (n14285) );
  buffer buf_n14286( .i (n14285), .o (n14286) );
  buffer buf_n14287( .i (n14286), .o (n14287) );
  buffer buf_n14288( .i (n14287), .o (n14288) );
  buffer buf_n14289( .i (n14288), .o (n14289) );
  buffer buf_n14290( .i (n14289), .o (n14290) );
  buffer buf_n14291( .i (n14290), .o (n14291) );
  buffer buf_n14292( .i (n14291), .o (n14292) );
  buffer buf_n14293( .i (n14292), .o (n14293) );
  buffer buf_n14294( .i (n14293), .o (n14294) );
  buffer buf_n14295( .i (n14294), .o (n14295) );
  buffer buf_n14296( .i (n14295), .o (n14296) );
  assign n14984 = ~n5666 & n11115 ;
  assign n14985 = ~n8683 & n13951 ;
  assign n14986 = n14102 & ~n14985 ;
  assign n14987 = n173 & n2871 ;
  buffer buf_n14988( .i (n14987), .o (n14988) );
  buffer buf_n14989( .i (n14988), .o (n14989) );
  assign n14990 = n14307 & ~n14989 ;
  assign n14991 = n14712 | n14990 ;
  assign n14992 = n14110 & n14988 ;
  assign n14993 = n174 & n14104 ;
  assign n14994 = n2873 | n14993 ;
  assign n14995 = ~n14992 & n14994 ;
  assign n14996 = n14308 | n14995 ;
  assign n14997 = ~n14991 & n14996 ;
  buffer buf_n14998( .i (n14997), .o (n14998) );
  buffer buf_n14999( .i (n14998), .o (n14999) );
  assign n15000 = n14717 | n14999 ;
  buffer buf_n15001( .i (n15000), .o (n15001) );
  buffer buf_n15002( .i (n15001), .o (n15002) );
  buffer buf_n15003( .i (n15002), .o (n15003) );
  buffer buf_n15004( .i (n15003), .o (n15004) );
  buffer buf_n15005( .i (n15004), .o (n15005) );
  buffer buf_n15006( .i (n15005), .o (n15006) );
  buffer buf_n15007( .i (n15006), .o (n15007) );
  buffer buf_n15008( .i (n15007), .o (n15008) );
  assign n15009 = n8732 & n14554 ;
  assign n15010 = n15008 | n15009 ;
  assign n15011 = n14986 & n15010 ;
  buffer buf_n15012( .i (n15011), .o (n15012) );
  buffer buf_n15013( .i (n15012), .o (n15013) );
  buffer buf_n15014( .i (n15013), .o (n15014) );
  buffer buf_n15015( .i (n15014), .o (n15015) );
  buffer buf_n15016( .i (n15015), .o (n15016) );
  buffer buf_n15017( .i (n15016), .o (n15017) );
  buffer buf_n15018( .i (n15017), .o (n15018) );
  buffer buf_n15019( .i (n15018), .o (n15019) );
  buffer buf_n15020( .i (n15019), .o (n15020) );
  buffer buf_n15021( .i (n15020), .o (n15021) );
  buffer buf_n15022( .i (n15021), .o (n15022) );
  buffer buf_n15023( .i (n15022), .o (n15023) );
  buffer buf_n15024( .i (n15023), .o (n15024) );
  buffer buf_n15025( .i (n15024), .o (n15025) );
  buffer buf_n15026( .i (n15025), .o (n15026) );
  buffer buf_n15027( .i (n15026), .o (n15027) );
  buffer buf_n15028( .i (n15027), .o (n15028) );
  buffer buf_n15029( .i (n15028), .o (n15029) );
  buffer buf_n15030( .i (n15029), .o (n15030) );
  buffer buf_n15031( .i (n15030), .o (n15031) );
  buffer buf_n15032( .i (n15031), .o (n15032) );
  buffer buf_n15033( .i (n15032), .o (n15033) );
  buffer buf_n15034( .i (n15033), .o (n15034) );
  buffer buf_n15035( .i (n15034), .o (n15035) );
  buffer buf_n15036( .i (n15035), .o (n15036) );
  buffer buf_n15037( .i (n15036), .o (n15037) );
  buffer buf_n15038( .i (n15037), .o (n15038) );
  buffer buf_n15039( .i (n15038), .o (n15039) );
  buffer buf_n15040( .i (n15039), .o (n15040) );
  buffer buf_n15041( .i (n15040), .o (n15041) );
  buffer buf_n15042( .i (n15041), .o (n15042) );
  buffer buf_n15043( .i (n15042), .o (n15043) );
  buffer buf_n15044( .i (n15043), .o (n15044) );
  buffer buf_n15045( .i (n15044), .o (n15045) );
  buffer buf_n15046( .i (n15045), .o (n15046) );
  assign n15047 = n14984 | n15046 ;
  buffer buf_n15048( .i (n15047), .o (n15048) );
  buffer buf_n15049( .i (n15048), .o (n15049) );
  buffer buf_n15050( .i (n15049), .o (n15050) );
  buffer buf_n15051( .i (n15050), .o (n15051) );
  buffer buf_n15052( .i (n15051), .o (n15052) );
  buffer buf_n15053( .i (n15052), .o (n15053) );
  buffer buf_n15054( .i (n15053), .o (n15054) );
  buffer buf_n15055( .i (n15054), .o (n15055) );
  buffer buf_n15056( .i (n15055), .o (n15056) );
  buffer buf_n15057( .i (n15056), .o (n15057) );
  buffer buf_n15058( .i (n15057), .o (n15058) );
  buffer buf_n15059( .i (n15058), .o (n15059) );
  buffer buf_n15060( .i (n15059), .o (n15060) );
  buffer buf_n15061( .i (n15060), .o (n15061) );
  buffer buf_n15062( .i (n15061), .o (n15062) );
  buffer buf_n15063( .i (n15062), .o (n15063) );
  buffer buf_n15064( .i (n15063), .o (n15064) );
  buffer buf_n15065( .i (n15064), .o (n15065) );
  buffer buf_n15066( .i (n15065), .o (n15066) );
  buffer buf_n15067( .i (n15066), .o (n15067) );
  buffer buf_n15068( .i (n15067), .o (n15068) );
  buffer buf_n15069( .i (n15068), .o (n15069) );
  buffer buf_n15070( .i (n15069), .o (n15070) );
  buffer buf_n15071( .i (n15070), .o (n15071) );
  buffer buf_n15072( .i (n15071), .o (n15072) );
  buffer buf_n15073( .i (n15072), .o (n15073) );
  buffer buf_n15074( .i (n15073), .o (n15074) );
  buffer buf_n15075( .i (n15074), .o (n15075) );
  buffer buf_n15076( .i (n15075), .o (n15076) );
  buffer buf_n15077( .i (n15076), .o (n15077) );
  buffer buf_n15078( .i (n15077), .o (n15078) );
  buffer buf_n15079( .i (n15078), .o (n15079) );
  buffer buf_n15080( .i (n15079), .o (n15080) );
  buffer buf_n15081( .i (n15080), .o (n15081) );
  buffer buf_n15082( .i (n15081), .o (n15082) );
  buffer buf_n15083( .i (n15082), .o (n15083) );
  buffer buf_n15084( .i (n15083), .o (n15084) );
  buffer buf_n15085( .i (n15084), .o (n15085) );
  buffer buf_n15086( .i (n15085), .o (n15086) );
  buffer buf_n15087( .i (n15086), .o (n15087) );
  buffer buf_n15088( .i (n15087), .o (n15088) );
  buffer buf_n15089( .i (n15088), .o (n15089) );
  buffer buf_n15090( .i (n15089), .o (n15090) );
  buffer buf_n15091( .i (n15090), .o (n15091) );
  buffer buf_n15092( .i (n15091), .o (n15092) );
  buffer buf_n15093( .i (n15092), .o (n15093) );
  buffer buf_n15094( .i (n15093), .o (n15094) );
  buffer buf_n15095( .i (n15094), .o (n15095) );
  buffer buf_n15096( .i (n15095), .o (n15096) );
  buffer buf_n15097( .i (n15096), .o (n15097) );
  buffer buf_n15098( .i (n15097), .o (n15098) );
  buffer buf_n15099( .i (n15098), .o (n15099) );
  buffer buf_n15100( .i (n15099), .o (n15100) );
  buffer buf_n15101( .i (n15100), .o (n15101) );
  buffer buf_n15102( .i (n15101), .o (n15102) );
  buffer buf_n15103( .i (n15102), .o (n15103) );
  buffer buf_n15104( .i (n15103), .o (n15104) );
  buffer buf_n15105( .i (n15104), .o (n15105) );
  buffer buf_n15106( .i (n15105), .o (n15106) );
  buffer buf_n15107( .i (n15106), .o (n15107) );
  buffer buf_n15108( .i (n15107), .o (n15108) );
  buffer buf_n15109( .i (n15108), .o (n15109) );
  buffer buf_n15110( .i (n15109), .o (n15110) );
  buffer buf_n15111( .i (n15110), .o (n15111) );
  buffer buf_n15112( .i (n15111), .o (n15112) );
  buffer buf_n15113( .i (n15112), .o (n15113) );
  buffer buf_n15114( .i (n15113), .o (n15114) );
  buffer buf_n15115( .i (n15114), .o (n15115) );
  buffer buf_n15116( .i (n15115), .o (n15116) );
  buffer buf_n15117( .i (n15116), .o (n15117) );
  buffer buf_n15118( .i (n15117), .o (n15118) );
  buffer buf_n15119( .i (n15118), .o (n15119) );
  buffer buf_n15120( .i (n15119), .o (n15120) );
  buffer buf_n15121( .i (n15120), .o (n15121) );
  buffer buf_n15122( .i (n15121), .o (n15122) );
  buffer buf_n15123( .i (n15122), .o (n15123) );
  buffer buf_n15124( .i (n15123), .o (n15124) );
  assign n15125 = ~n5639 & n14446 ;
  buffer buf_n15126( .i (n13950), .o (n15126) );
  assign n15127 = ~n13620 & n15126 ;
  assign n15128 = n14102 & ~n15127 ;
  assign n15129 = n212 & ~n13396 ;
  buffer buf_n15130( .i (n15129), .o (n15130) );
  buffer buf_n3733( .i (n3732), .o (n3733) );
  buffer buf_n3734( .i (n3733), .o (n3734) );
  buffer buf_n3735( .i (n3734), .o (n3735) );
  buffer buf_n3736( .i (n3735), .o (n3736) );
  buffer buf_n3737( .i (n3736), .o (n3737) );
  buffer buf_n3738( .i (n3737), .o (n3738) );
  buffer buf_n3739( .i (n3738), .o (n3739) );
  buffer buf_n3740( .i (n3739), .o (n3740) );
  buffer buf_n3741( .i (n3740), .o (n3741) );
  buffer buf_n3742( .i (n3741), .o (n3742) );
  buffer buf_n15131( .i (n13963), .o (n15131) );
  assign n15132 = n212 | n15131 ;
  assign n15133 = n3742 & n15132 ;
  assign n15134 = n15130 | n15133 ;
  buffer buf_n15135( .i (n15134), .o (n15135) );
  buffer buf_n15136( .i (n15135), .o (n15136) );
  buffer buf_n15137( .i (n10914), .o (n15137) );
  assign n15138 = n3742 & n15137 ;
  assign n15139 = n15130 & n15138 ;
  buffer buf_n15140( .i (n15139), .o (n15140) );
  assign n15141 = n14712 | n15140 ;
  assign n15142 = n15136 & ~n15141 ;
  buffer buf_n15143( .i (n15142), .o (n15143) );
  buffer buf_n15144( .i (n15143), .o (n15144) );
  assign n15145 = n14717 | n15144 ;
  buffer buf_n15146( .i (n15145), .o (n15146) );
  buffer buf_n15147( .i (n15146), .o (n15147) );
  buffer buf_n15148( .i (n15147), .o (n15148) );
  buffer buf_n15149( .i (n15148), .o (n15149) );
  buffer buf_n15150( .i (n15149), .o (n15150) );
  buffer buf_n15151( .i (n15150), .o (n15151) );
  buffer buf_n15152( .i (n15151), .o (n15152) );
  buffer buf_n15153( .i (n15152), .o (n15153) );
  buffer buf_n15154( .i (n13621), .o (n15154) );
  assign n15155 = n13605 & n15154 ;
  assign n15156 = n15153 | n15155 ;
  assign n15157 = n15128 & n15156 ;
  buffer buf_n15158( .i (n15157), .o (n15158) );
  buffer buf_n15159( .i (n15158), .o (n15159) );
  buffer buf_n15160( .i (n15159), .o (n15160) );
  buffer buf_n15161( .i (n15160), .o (n15161) );
  buffer buf_n15162( .i (n15161), .o (n15162) );
  buffer buf_n15163( .i (n15162), .o (n15163) );
  buffer buf_n15164( .i (n15163), .o (n15164) );
  buffer buf_n15165( .i (n15164), .o (n15165) );
  assign n15166 = n15125 | n15165 ;
  buffer buf_n15167( .i (n15166), .o (n15167) );
  buffer buf_n15168( .i (n15167), .o (n15168) );
  buffer buf_n15169( .i (n15168), .o (n15169) );
  buffer buf_n15170( .i (n15169), .o (n15170) );
  buffer buf_n15171( .i (n15170), .o (n15171) );
  buffer buf_n15172( .i (n15171), .o (n15172) );
  buffer buf_n15173( .i (n15172), .o (n15173) );
  buffer buf_n15174( .i (n15173), .o (n15174) );
  buffer buf_n15175( .i (n15174), .o (n15175) );
  buffer buf_n15176( .i (n15175), .o (n15176) );
  buffer buf_n15177( .i (n15176), .o (n15177) );
  buffer buf_n15178( .i (n15177), .o (n15178) );
  buffer buf_n15179( .i (n15178), .o (n15179) );
  buffer buf_n15180( .i (n15179), .o (n15180) );
  buffer buf_n15181( .i (n15180), .o (n15181) );
  buffer buf_n15182( .i (n15181), .o (n15182) );
  buffer buf_n15183( .i (n15182), .o (n15183) );
  buffer buf_n15184( .i (n15183), .o (n15184) );
  buffer buf_n15185( .i (n15184), .o (n15185) );
  buffer buf_n15186( .i (n15185), .o (n15186) );
  buffer buf_n15187( .i (n15186), .o (n15187) );
  buffer buf_n15188( .i (n15187), .o (n15188) );
  buffer buf_n15189( .i (n15188), .o (n15189) );
  buffer buf_n15190( .i (n15189), .o (n15190) );
  buffer buf_n15191( .i (n15190), .o (n15191) );
  buffer buf_n15192( .i (n15191), .o (n15192) );
  buffer buf_n15193( .i (n15192), .o (n15193) );
  buffer buf_n15194( .i (n15193), .o (n15194) );
  buffer buf_n15195( .i (n15194), .o (n15195) );
  buffer buf_n15196( .i (n15195), .o (n15196) );
  buffer buf_n15197( .i (n15196), .o (n15197) );
  buffer buf_n15198( .i (n15197), .o (n15198) );
  buffer buf_n15199( .i (n15198), .o (n15199) );
  buffer buf_n15200( .i (n15199), .o (n15200) );
  buffer buf_n15201( .i (n15200), .o (n15201) );
  buffer buf_n15202( .i (n15201), .o (n15202) );
  buffer buf_n15203( .i (n15202), .o (n15203) );
  buffer buf_n15204( .i (n15203), .o (n15204) );
  buffer buf_n15205( .i (n15204), .o (n15205) );
  buffer buf_n15206( .i (n15205), .o (n15206) );
  buffer buf_n15207( .i (n15206), .o (n15207) );
  buffer buf_n15208( .i (n15207), .o (n15208) );
  buffer buf_n15209( .i (n15208), .o (n15209) );
  buffer buf_n15210( .i (n15209), .o (n15210) );
  buffer buf_n15211( .i (n15210), .o (n15211) );
  buffer buf_n15212( .i (n15211), .o (n15212) );
  buffer buf_n15213( .i (n15212), .o (n15213) );
  buffer buf_n15214( .i (n15213), .o (n15214) );
  buffer buf_n15215( .i (n15214), .o (n15215) );
  buffer buf_n15216( .i (n15215), .o (n15216) );
  buffer buf_n15217( .i (n15216), .o (n15217) );
  buffer buf_n15218( .i (n15217), .o (n15218) );
  buffer buf_n15219( .i (n15218), .o (n15219) );
  buffer buf_n15220( .i (n15219), .o (n15220) );
  buffer buf_n15221( .i (n15220), .o (n15221) );
  buffer buf_n15222( .i (n15221), .o (n15222) );
  buffer buf_n15223( .i (n15222), .o (n15223) );
  buffer buf_n15224( .i (n15223), .o (n15224) );
  buffer buf_n15225( .i (n15224), .o (n15225) );
  buffer buf_n15226( .i (n15225), .o (n15226) );
  buffer buf_n15227( .i (n15226), .o (n15227) );
  buffer buf_n15228( .i (n15227), .o (n15228) );
  buffer buf_n15229( .i (n15228), .o (n15229) );
  buffer buf_n15230( .i (n15229), .o (n15230) );
  buffer buf_n15231( .i (n15230), .o (n15231) );
  buffer buf_n15232( .i (n15231), .o (n15232) );
  buffer buf_n15233( .i (n15232), .o (n15233) );
  buffer buf_n15234( .i (n15233), .o (n15234) );
  buffer buf_n15235( .i (n15234), .o (n15235) );
  buffer buf_n15236( .i (n15235), .o (n15236) );
  buffer buf_n15237( .i (n15236), .o (n15237) );
  buffer buf_n15238( .i (n15237), .o (n15238) );
  buffer buf_n15239( .i (n15238), .o (n15239) );
  buffer buf_n15240( .i (n15239), .o (n15240) );
  buffer buf_n15241( .i (n15240), .o (n15241) );
  buffer buf_n15242( .i (n15241), .o (n15242) );
  buffer buf_n15243( .i (n15242), .o (n15243) );
  buffer buf_n15244( .i (n15243), .o (n15244) );
  buffer buf_n15245( .i (n15244), .o (n15245) );
  buffer buf_n15246( .i (n15245), .o (n15246) );
  buffer buf_n15247( .i (n15246), .o (n15247) );
  buffer buf_n15248( .i (n15247), .o (n15248) );
  buffer buf_n15249( .i (n15248), .o (n15249) );
  buffer buf_n15250( .i (n15249), .o (n15250) );
  buffer buf_n15251( .i (n15250), .o (n15251) );
  buffer buf_n15252( .i (n15251), .o (n15252) );
  buffer buf_n15253( .i (n15252), .o (n15253) );
  buffer buf_n15254( .i (n15253), .o (n15254) );
  buffer buf_n15255( .i (n15254), .o (n15255) );
  buffer buf_n15256( .i (n15255), .o (n15256) );
  buffer buf_n15257( .i (n15256), .o (n15257) );
  buffer buf_n15258( .i (n15257), .o (n15258) );
  buffer buf_n15259( .i (n15258), .o (n15259) );
  buffer buf_n15260( .i (n15259), .o (n15260) );
  buffer buf_n15261( .i (n15260), .o (n15261) );
  buffer buf_n15262( .i (n15261), .o (n15262) );
  buffer buf_n15263( .i (n15262), .o (n15263) );
  buffer buf_n15264( .i (n15263), .o (n15264) );
  buffer buf_n15265( .i (n15264), .o (n15265) );
  buffer buf_n15266( .i (n15265), .o (n15266) );
  buffer buf_n15267( .i (n15266), .o (n15267) );
  buffer buf_n15268( .i (n15267), .o (n15268) );
  buffer buf_n15269( .i (n15268), .o (n15269) );
  buffer buf_n15270( .i (n15269), .o (n15270) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  assign n15271 = n716 & n1777 ;
  buffer buf_n15272( .i (n15271), .o (n15272) );
  buffer buf_n15273( .i (n15272), .o (n15273) );
  assign n15274 = n14305 & ~n15273 ;
  assign n15275 = n6087 | n15274 ;
  buffer buf_n1778( .i (n1777), .o (n1778) );
  assign n15276 = n1778 & n13963 ;
  assign n15277 = n718 | n15276 ;
  assign n15278 = n10914 & n15272 ;
  assign n15279 = n15277 & ~n15278 ;
  assign n15280 = n14306 | n15279 ;
  assign n15281 = ~n15275 & n15280 ;
  buffer buf_n15282( .i (n15281), .o (n15282) );
  buffer buf_n15283( .i (n15282), .o (n15283) );
  buffer buf_n15284( .i (n15283), .o (n15284) );
  buffer buf_n15285( .i (n15284), .o (n15285) );
  buffer buf_n15286( .i (n5917), .o (n15286) );
  buffer buf_n15287( .i (n15286), .o (n15287) );
  assign n15288 = n15285 | n15287 ;
  buffer buf_n15289( .i (n15288), .o (n15289) );
  buffer buf_n15290( .i (n15289), .o (n15290) );
  buffer buf_n15291( .i (n15290), .o (n15291) );
  buffer buf_n15292( .i (n15291), .o (n15292) );
  buffer buf_n15293( .i (n15292), .o (n15293) );
  buffer buf_n15294( .i (n15293), .o (n15294) );
  buffer buf_n15295( .i (n15294), .o (n15295) );
  buffer buf_n15296( .i (n15295), .o (n15296) );
  buffer buf_n15297( .i (n15296), .o (n15297) );
  assign n15298 = n9277 & n11541 ;
  assign n15299 = n15297 | n15298 ;
  assign n15300 = ~n9271 & n15126 ;
  buffer buf_n15301( .i (n14101), .o (n15301) );
  assign n15302 = ~n15300 & n15301 ;
  buffer buf_n15303( .i (n15302), .o (n15303) );
  assign n15304 = n15299 & n15303 ;
  assign n15305 = n11978 & ~n14696 ;
  assign n15306 = n15304 | n15305 ;
  buffer buf_n15307( .i (n15306), .o (n15307) );
  buffer buf_n15308( .i (n15307), .o (n15308) );
  buffer buf_n15309( .i (n15308), .o (n15309) );
  buffer buf_n15310( .i (n15309), .o (n15310) );
  buffer buf_n15311( .i (n15310), .o (n15311) );
  buffer buf_n15312( .i (n15311), .o (n15312) );
  buffer buf_n15313( .i (n15312), .o (n15313) );
  buffer buf_n15314( .i (n15313), .o (n15314) );
  buffer buf_n15315( .i (n15314), .o (n15315) );
  buffer buf_n15316( .i (n15315), .o (n15316) );
  buffer buf_n15317( .i (n15316), .o (n15317) );
  buffer buf_n15318( .i (n15317), .o (n15318) );
  buffer buf_n15319( .i (n15318), .o (n15319) );
  buffer buf_n15320( .i (n15319), .o (n15320) );
  buffer buf_n15321( .i (n15320), .o (n15321) );
  buffer buf_n15322( .i (n15321), .o (n15322) );
  buffer buf_n15323( .i (n15322), .o (n15323) );
  buffer buf_n15324( .i (n15323), .o (n15324) );
  buffer buf_n15325( .i (n15324), .o (n15325) );
  buffer buf_n15326( .i (n15325), .o (n15326) );
  buffer buf_n15327( .i (n15326), .o (n15327) );
  buffer buf_n15328( .i (n15327), .o (n15328) );
  buffer buf_n15329( .i (n15328), .o (n15329) );
  buffer buf_n15330( .i (n15329), .o (n15330) );
  buffer buf_n15331( .i (n15330), .o (n15331) );
  buffer buf_n15332( .i (n15331), .o (n15332) );
  buffer buf_n15333( .i (n15332), .o (n15333) );
  buffer buf_n15334( .i (n15333), .o (n15334) );
  buffer buf_n15335( .i (n15334), .o (n15335) );
  buffer buf_n15336( .i (n15335), .o (n15336) );
  buffer buf_n15337( .i (n15336), .o (n15337) );
  buffer buf_n15338( .i (n15337), .o (n15338) );
  buffer buf_n15339( .i (n15338), .o (n15339) );
  buffer buf_n15340( .i (n15339), .o (n15340) );
  buffer buf_n15341( .i (n15340), .o (n15341) );
  buffer buf_n15342( .i (n15341), .o (n15342) );
  buffer buf_n15343( .i (n15342), .o (n15343) );
  buffer buf_n15344( .i (n15343), .o (n15344) );
  buffer buf_n15345( .i (n15344), .o (n15345) );
  buffer buf_n15346( .i (n15345), .o (n15346) );
  buffer buf_n15347( .i (n15346), .o (n15347) );
  buffer buf_n15348( .i (n15347), .o (n15348) );
  buffer buf_n15349( .i (n15348), .o (n15349) );
  buffer buf_n15350( .i (n15349), .o (n15350) );
  buffer buf_n15351( .i (n15350), .o (n15351) );
  buffer buf_n15352( .i (n15351), .o (n15352) );
  buffer buf_n15353( .i (n15352), .o (n15353) );
  buffer buf_n15354( .i (n15353), .o (n15354) );
  buffer buf_n15355( .i (n15354), .o (n15355) );
  buffer buf_n15356( .i (n15355), .o (n15356) );
  buffer buf_n15357( .i (n15356), .o (n15357) );
  buffer buf_n15358( .i (n15357), .o (n15358) );
  buffer buf_n15359( .i (n15358), .o (n15359) );
  buffer buf_n15360( .i (n15359), .o (n15360) );
  buffer buf_n15361( .i (n15360), .o (n15361) );
  buffer buf_n15362( .i (n15361), .o (n15362) );
  buffer buf_n15363( .i (n15362), .o (n15363) );
  buffer buf_n15364( .i (n15363), .o (n15364) );
  buffer buf_n15365( .i (n15364), .o (n15365) );
  buffer buf_n15366( .i (n15365), .o (n15366) );
  buffer buf_n15367( .i (n15366), .o (n15367) );
  buffer buf_n15368( .i (n15367), .o (n15368) );
  buffer buf_n15369( .i (n15368), .o (n15369) );
  buffer buf_n15370( .i (n15369), .o (n15370) );
  buffer buf_n15371( .i (n15370), .o (n15371) );
  buffer buf_n15372( .i (n15371), .o (n15372) );
  buffer buf_n15373( .i (n15372), .o (n15373) );
  buffer buf_n15374( .i (n15373), .o (n15374) );
  buffer buf_n15375( .i (n15374), .o (n15375) );
  buffer buf_n15376( .i (n15375), .o (n15376) );
  buffer buf_n15377( .i (n15376), .o (n15377) );
  buffer buf_n15378( .i (n15377), .o (n15378) );
  buffer buf_n15379( .i (n15378), .o (n15379) );
  buffer buf_n15380( .i (n15379), .o (n15380) );
  buffer buf_n15381( .i (n15380), .o (n15381) );
  buffer buf_n15382( .i (n15381), .o (n15382) );
  buffer buf_n15383( .i (n15382), .o (n15383) );
  buffer buf_n15384( .i (n15383), .o (n15384) );
  buffer buf_n15385( .i (n15384), .o (n15385) );
  buffer buf_n15386( .i (n15385), .o (n15386) );
  buffer buf_n15387( .i (n15386), .o (n15387) );
  buffer buf_n15388( .i (n15387), .o (n15388) );
  buffer buf_n15389( .i (n15388), .o (n15389) );
  buffer buf_n15390( .i (n15389), .o (n15390) );
  buffer buf_n15391( .i (n15390), .o (n15391) );
  buffer buf_n15392( .i (n15391), .o (n15392) );
  buffer buf_n15393( .i (n15392), .o (n15393) );
  buffer buf_n15394( .i (n15393), .o (n15394) );
  buffer buf_n15395( .i (n15394), .o (n15395) );
  buffer buf_n15396( .i (n15395), .o (n15396) );
  buffer buf_n15397( .i (n15396), .o (n15397) );
  buffer buf_n15398( .i (n15397), .o (n15398) );
  buffer buf_n15399( .i (n15398), .o (n15399) );
  buffer buf_n15400( .i (n15399), .o (n15400) );
  buffer buf_n15401( .i (n15400), .o (n15401) );
  buffer buf_n15402( .i (n15401), .o (n15402) );
  buffer buf_n15403( .i (n15402), .o (n15403) );
  buffer buf_n15404( .i (n15403), .o (n15404) );
  buffer buf_n15405( .i (n15404), .o (n15405) );
  buffer buf_n15406( .i (n15405), .o (n15406) );
  buffer buf_n15407( .i (n15406), .o (n15407) );
  buffer buf_n15408( .i (n15407), .o (n15408) );
  buffer buf_n15409( .i (n15408), .o (n15409) );
  buffer buf_n15410( .i (n15409), .o (n15410) );
  buffer buf_n15411( .i (n15410), .o (n15411) );
  buffer buf_n15412( .i (n15411), .o (n15412) );
  buffer buf_n15413( .i (n15412), .o (n15413) );
  buffer buf_n15414( .i (n15413), .o (n15414) );
  buffer buf_n15415( .i (n15414), .o (n15415) );
  buffer buf_n15416( .i (n15415), .o (n15416) );
  buffer buf_n15417( .i (n15416), .o (n15417) );
  buffer buf_n13818( .i (n13817), .o (n13818) );
  buffer buf_n13819( .i (n13818), .o (n13819) );
  buffer buf_n13820( .i (n13819), .o (n13820) );
  buffer buf_n13821( .i (n13820), .o (n13821) );
  buffer buf_n13822( .i (n13821), .o (n13822) );
  buffer buf_n13823( .i (n13822), .o (n13823) );
  buffer buf_n13824( .i (n13823), .o (n13824) );
  buffer buf_n13825( .i (n13824), .o (n13825) );
  buffer buf_n13826( .i (n13825), .o (n13826) );
  buffer buf_n13827( .i (n13826), .o (n13827) );
  buffer buf_n13828( .i (n13827), .o (n13828) );
  buffer buf_n13829( .i (n13828), .o (n13829) );
  buffer buf_n13830( .i (n13829), .o (n13830) );
  buffer buf_n13831( .i (n13830), .o (n13831) );
  buffer buf_n13832( .i (n13831), .o (n13832) );
  buffer buf_n13833( .i (n13832), .o (n13833) );
  buffer buf_n13834( .i (n13833), .o (n13834) );
  buffer buf_n13835( .i (n13834), .o (n13835) );
  buffer buf_n13836( .i (n13835), .o (n13836) );
  buffer buf_n13837( .i (n13836), .o (n13837) );
  buffer buf_n13838( .i (n13837), .o (n13838) );
  buffer buf_n13839( .i (n13838), .o (n13839) );
  buffer buf_n13840( .i (n13839), .o (n13840) );
  buffer buf_n13841( .i (n13840), .o (n13841) );
  buffer buf_n13842( .i (n13841), .o (n13842) );
  buffer buf_n13843( .i (n13842), .o (n13843) );
  buffer buf_n13844( .i (n13843), .o (n13844) );
  buffer buf_n13845( .i (n13844), .o (n13845) );
  buffer buf_n13846( .i (n13845), .o (n13846) );
  buffer buf_n13847( .i (n13846), .o (n13847) );
  buffer buf_n13848( .i (n13847), .o (n13848) );
  buffer buf_n13849( .i (n13848), .o (n13849) );
  buffer buf_n13850( .i (n13849), .o (n13850) );
  buffer buf_n13851( .i (n13850), .o (n13851) );
  buffer buf_n13852( .i (n13851), .o (n13852) );
  buffer buf_n13853( .i (n13852), .o (n13853) );
  buffer buf_n13854( .i (n13853), .o (n13854) );
  buffer buf_n13855( .i (n13854), .o (n13855) );
  buffer buf_n13856( .i (n13855), .o (n13856) );
  buffer buf_n13857( .i (n13856), .o (n13857) );
  buffer buf_n13858( .i (n13857), .o (n13858) );
  buffer buf_n13859( .i (n13858), .o (n13859) );
  buffer buf_n13860( .i (n13859), .o (n13860) );
  buffer buf_n13861( .i (n13860), .o (n13861) );
  buffer buf_n13862( .i (n13861), .o (n13862) );
  buffer buf_n13863( .i (n13862), .o (n13863) );
  buffer buf_n13864( .i (n13863), .o (n13864) );
  buffer buf_n13865( .i (n13864), .o (n13865) );
  buffer buf_n13866( .i (n13865), .o (n13866) );
  buffer buf_n13867( .i (n13866), .o (n13867) );
  buffer buf_n13868( .i (n13867), .o (n13868) );
  buffer buf_n13869( .i (n13868), .o (n13869) );
  buffer buf_n13870( .i (n13869), .o (n13870) );
  buffer buf_n13871( .i (n13870), .o (n13871) );
  buffer buf_n13872( .i (n13871), .o (n13872) );
  buffer buf_n13873( .i (n13872), .o (n13873) );
  buffer buf_n13874( .i (n13873), .o (n13874) );
  buffer buf_n13875( .i (n13874), .o (n13875) );
  buffer buf_n13876( .i (n13875), .o (n13876) );
  buffer buf_n13877( .i (n13876), .o (n13877) );
  buffer buf_n13878( .i (n13877), .o (n13878) );
  buffer buf_n13879( .i (n13878), .o (n13879) );
  buffer buf_n13880( .i (n13879), .o (n13880) );
  buffer buf_n13881( .i (n13880), .o (n13881) );
  buffer buf_n13882( .i (n13881), .o (n13882) );
  buffer buf_n13883( .i (n13882), .o (n13883) );
  buffer buf_n13884( .i (n13883), .o (n13884) );
  buffer buf_n13885( .i (n13884), .o (n13885) );
  buffer buf_n13886( .i (n13885), .o (n13886) );
  buffer buf_n13887( .i (n13886), .o (n13887) );
  buffer buf_n13888( .i (n13887), .o (n13888) );
  buffer buf_n13889( .i (n13888), .o (n13889) );
  buffer buf_n13890( .i (n13889), .o (n13890) );
  buffer buf_n13891( .i (n13890), .o (n13891) );
  buffer buf_n13892( .i (n13891), .o (n13892) );
  buffer buf_n13893( .i (n13892), .o (n13893) );
  buffer buf_n13894( .i (n13893), .o (n13894) );
  buffer buf_n13895( .i (n13894), .o (n13895) );
  buffer buf_n13896( .i (n13895), .o (n13896) );
  buffer buf_n13897( .i (n13896), .o (n13897) );
  buffer buf_n13898( .i (n13897), .o (n13898) );
  buffer buf_n13899( .i (n13898), .o (n13899) );
  buffer buf_n13900( .i (n13899), .o (n13900) );
  buffer buf_n13901( .i (n13900), .o (n13901) );
  buffer buf_n13902( .i (n13901), .o (n13902) );
  buffer buf_n13903( .i (n13902), .o (n13903) );
  buffer buf_n13904( .i (n13903), .o (n13904) );
  buffer buf_n13905( .i (n13904), .o (n13905) );
  buffer buf_n13906( .i (n13905), .o (n13906) );
  buffer buf_n13907( .i (n13906), .o (n13907) );
  buffer buf_n13908( .i (n13907), .o (n13908) );
  buffer buf_n13909( .i (n13908), .o (n13909) );
  buffer buf_n13910( .i (n13909), .o (n13910) );
  buffer buf_n13911( .i (n13910), .o (n13911) );
  buffer buf_n13912( .i (n13911), .o (n13912) );
  buffer buf_n13913( .i (n13912), .o (n13913) );
  buffer buf_n13914( .i (n13913), .o (n13914) );
  buffer buf_n13915( .i (n13914), .o (n13915) );
  buffer buf_n13916( .i (n13915), .o (n13916) );
  buffer buf_n13917( .i (n13916), .o (n13917) );
  buffer buf_n13918( .i (n13917), .o (n13918) );
  buffer buf_n13919( .i (n13918), .o (n13919) );
  buffer buf_n13920( .i (n13919), .o (n13920) );
  buffer buf_n13921( .i (n13920), .o (n13921) );
  buffer buf_n13922( .i (n13921), .o (n13922) );
  buffer buf_n13923( .i (n13922), .o (n13923) );
  buffer buf_n13924( .i (n13923), .o (n13924) );
  buffer buf_n13925( .i (n13924), .o (n13925) );
  buffer buf_n13926( .i (n13925), .o (n13926) );
  buffer buf_n13927( .i (n13926), .o (n13927) );
  buffer buf_n13928( .i (n13927), .o (n13928) );
  buffer buf_n13929( .i (n13928), .o (n13929) );
  buffer buf_n13930( .i (n13929), .o (n13930) );
  buffer buf_n13931( .i (n13930), .o (n13931) );
  buffer buf_n12098( .i (n12097), .o (n12098) );
  buffer buf_n12099( .i (n12098), .o (n12099) );
  buffer buf_n12100( .i (n12099), .o (n12100) );
  buffer buf_n12101( .i (n12100), .o (n12101) );
  buffer buf_n12102( .i (n12101), .o (n12102) );
  buffer buf_n12103( .i (n12102), .o (n12103) );
  buffer buf_n12104( .i (n12103), .o (n12104) );
  buffer buf_n12105( .i (n12104), .o (n12105) );
  buffer buf_n12106( .i (n12105), .o (n12106) );
  buffer buf_n12107( .i (n12106), .o (n12107) );
  buffer buf_n12108( .i (n12107), .o (n12108) );
  buffer buf_n12109( .i (n12108), .o (n12109) );
  buffer buf_n12110( .i (n12109), .o (n12110) );
  buffer buf_n12111( .i (n12110), .o (n12111) );
  buffer buf_n12112( .i (n12111), .o (n12112) );
  buffer buf_n12113( .i (n12112), .o (n12113) );
  buffer buf_n12114( .i (n12113), .o (n12114) );
  buffer buf_n12115( .i (n12114), .o (n12115) );
  buffer buf_n12116( .i (n12115), .o (n12116) );
  buffer buf_n12117( .i (n12116), .o (n12117) );
  buffer buf_n12118( .i (n12117), .o (n12118) );
  buffer buf_n12119( .i (n12118), .o (n12119) );
  buffer buf_n12120( .i (n12119), .o (n12120) );
  buffer buf_n12121( .i (n12120), .o (n12121) );
  buffer buf_n12122( .i (n12121), .o (n12122) );
  buffer buf_n12123( .i (n12122), .o (n12123) );
  buffer buf_n12124( .i (n12123), .o (n12124) );
  buffer buf_n12125( .i (n12124), .o (n12125) );
  buffer buf_n12126( .i (n12125), .o (n12126) );
  buffer buf_n12127( .i (n12126), .o (n12127) );
  buffer buf_n12128( .i (n12127), .o (n12128) );
  buffer buf_n12129( .i (n12128), .o (n12129) );
  buffer buf_n12130( .i (n12129), .o (n12130) );
  buffer buf_n12131( .i (n12130), .o (n12131) );
  buffer buf_n12132( .i (n12131), .o (n12132) );
  buffer buf_n12133( .i (n12132), .o (n12133) );
  buffer buf_n12134( .i (n12133), .o (n12134) );
  buffer buf_n12135( .i (n12134), .o (n12135) );
  buffer buf_n12136( .i (n12135), .o (n12136) );
  buffer buf_n12137( .i (n12136), .o (n12137) );
  buffer buf_n12138( .i (n12137), .o (n12138) );
  buffer buf_n12139( .i (n12138), .o (n12139) );
  buffer buf_n12140( .i (n12139), .o (n12140) );
  buffer buf_n12141( .i (n12140), .o (n12141) );
  buffer buf_n12142( .i (n12141), .o (n12142) );
  buffer buf_n12143( .i (n12142), .o (n12143) );
  buffer buf_n12144( .i (n12143), .o (n12144) );
  buffer buf_n12145( .i (n12144), .o (n12145) );
  buffer buf_n12146( .i (n12145), .o (n12146) );
  buffer buf_n12147( .i (n12146), .o (n12147) );
  buffer buf_n12148( .i (n12147), .o (n12148) );
  buffer buf_n12149( .i (n12148), .o (n12149) );
  buffer buf_n12150( .i (n12149), .o (n12150) );
  buffer buf_n12151( .i (n12150), .o (n12151) );
  buffer buf_n12152( .i (n12151), .o (n12152) );
  buffer buf_n12153( .i (n12152), .o (n12153) );
  buffer buf_n12154( .i (n12153), .o (n12154) );
  buffer buf_n12155( .i (n12154), .o (n12155) );
  buffer buf_n12156( .i (n12155), .o (n12156) );
  buffer buf_n12157( .i (n12156), .o (n12157) );
  buffer buf_n12158( .i (n12157), .o (n12158) );
  buffer buf_n12159( .i (n12158), .o (n12159) );
  buffer buf_n12160( .i (n12159), .o (n12160) );
  buffer buf_n12161( .i (n12160), .o (n12161) );
  buffer buf_n12162( .i (n12161), .o (n12162) );
  buffer buf_n12163( .i (n12162), .o (n12163) );
  buffer buf_n12164( .i (n12163), .o (n12164) );
  buffer buf_n12165( .i (n12164), .o (n12165) );
  buffer buf_n12166( .i (n12165), .o (n12166) );
  assign y0 = n6407 ;
  assign y1 = n5601 ;
  assign y2 = n6782 ;
  assign y3 = n7741 ;
  assign y4 = n7821 ;
  assign y5 = n7856 ;
  assign y6 = n8018 ;
  assign y7 = n8068 ;
  assign y8 = n8286 ;
  assign y9 = n8413 ;
  assign y10 = n8550 ;
  assign y11 = n6539 ;
  assign y12 = n8848 ;
  assign y13 = n9095 ;
  assign y14 = n9212 ;
  assign y15 = n9433 ;
  assign y16 = n9621 ;
  assign y17 = n9873 ;
  assign y18 = n10061 ;
  assign y19 = n10203 ;
  assign y20 = n10498 ;
  assign y21 = n10620 ;
  assign y22 = n10632 ;
  assign y23 = n10398 ;
  assign y24 = n10732 ;
  assign y25 = n10902 ;
  assign y26 = n11109 ;
  assign y27 = n11194 ;
  assign y28 = n11333 ;
  assign y29 = n11490 ;
  assign y30 = n11656 ;
  assign y31 = n8859 ;
  assign y32 = n9784 ;
  assign y33 = n11813 ;
  assign y34 = n11954 ;
  assign y35 = n12091 ;
  assign y36 = n12310 ;
  assign y37 = n12706 ;
  assign y38 = n13023 ;
  assign y39 = n13238 ;
  assign y40 = n13174 ;
  assign y41 = n13391 ;
  assign y42 = n13537 ;
  assign y43 = n13602 ;
  assign y44 = n13761 ;
  assign y45 = n9399 ;
  assign y46 = n13779 ;
  assign y47 = n8640 ;
  assign y48 = n14099 ;
  assign y49 = n14267 ;
  assign y50 = n14441 ;
  assign y51 = n14552 ;
  assign y52 = n14695 ;
  assign y53 = n12909 ;
  assign y54 = n14842 ;
  assign y55 = n14249 ;
  assign y56 = n11055 ;
  assign y57 = n10022 ;
  assign y58 = n14983 ;
  assign y59 = n14296 ;
  assign y60 = n15124 ;
  assign y61 = n15270 ;
  assign y62 = n15417 ;
  assign y63 = n13931 ;
  assign y64 = n12166 ;
endmodule
