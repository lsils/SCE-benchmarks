module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G158 , G159 , G16 , G160 , G161 , G162 , G163 , G164 , G165 , G166 , G167 , G168 , G169 , G17 , G170 , G171 , G172 , G173 , G174 , G175 , G176 , G177 , G178 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 , G5193 , G5194 , G5195 , G5196 , G5197 , G5198 , G5199 , G5200 , G5201 , G5202 , G5203 , G5204 , G5205 , G5206 , G5207 , G5208 , G5209 , G5210 , G5211 , G5212 , G5213 , G5214 , G5215 , G5216 , G5217 , G5218 , G5219 , G5220 , G5221 , G5222 , G5223 , G5224 , G5225 , G5226 , G5227 , G5228 , G5229 , G5230 , G5231 , G5232 , G5233 , G5234 , G5235 , G5236 , G5237 , G5238 , G5239 , G5240 , G5241 , G5242 , G5243 , G5244 , G5245 , G5246 , G5247 , G5248 , G5249 , G5250 , G5251 , G5252 , G5253 , G5254 , G5255 , G5256 , G5257 , G5258 , G5259 , G5260 , G5261 , G5262 , G5263 , G5264 , G5265 , G5266 , G5267 , G5268 , G5269 , G5270 , G5271 , G5272 , G5273 , G5274 , G5275 , G5276 , G5277 , G5278 , G5279 , G5280 , G5281 , G5282 , G5283 , G5284 , G5285 , G5286 , G5287 , G5288 , G5289 , G5290 , G5291 , G5292 , G5293 , G5294 , G5295 , G5296 , G5297 , G5298 , G5299 , G5300 , G5301 , G5302 , G5303 , G5304 , G5305 , G5306 , G5307 , G5308 , G5309 , G5310 , G5311 , G5312 , G5313 , G5314 , G5315 );
  input G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G158 , G159 , G16 , G160 , G161 , G162 , G163 , G164 , G165 , G166 , G167 , G168 , G169 , G17 , G170 , G171 , G172 , G173 , G174 , G175 , G176 , G177 , G178 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 ;
  output G5193 , G5194 , G5195 , G5196 , G5197 , G5198 , G5199 , G5200 , G5201 , G5202 , G5203 , G5204 , G5205 , G5206 , G5207 , G5208 , G5209 , G5210 , G5211 , G5212 , G5213 , G5214 , G5215 , G5216 , G5217 , G5218 , G5219 , G5220 , G5221 , G5222 , G5223 , G5224 , G5225 , G5226 , G5227 , G5228 , G5229 , G5230 , G5231 , G5232 , G5233 , G5234 , G5235 , G5236 , G5237 , G5238 , G5239 , G5240 , G5241 , G5242 , G5243 , G5244 , G5245 , G5246 , G5247 , G5248 , G5249 , G5250 , G5251 , G5252 , G5253 , G5254 , G5255 , G5256 , G5257 , G5258 , G5259 , G5260 , G5261 , G5262 , G5263 , G5264 , G5265 , G5266 , G5267 , G5268 , G5269 , G5270 , G5271 , G5272 , G5273 , G5274 , G5275 , G5276 , G5277 , G5278 , G5279 , G5280 , G5281 , G5282 , G5283 , G5284 , G5285 , G5286 , G5287 , G5288 , G5289 , G5290 , G5291 , G5292 , G5293 , G5294 , G5295 , G5296 , G5297 , G5298 , G5299 , G5300 , G5301 , G5302 , G5303 , G5304 , G5305 , G5306 , G5307 , G5308 , G5309 , G5310 , G5311 , G5312 , G5313 , G5314 , G5315 ;
  wire n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 ;
  assign n179 = G153 & G156 ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = G66 & G67 ;
  assign n182 = G1 & G134 ;
  assign n183 = ~G165 & G63 ;
  assign n184 = ~G11 | G164 ;
  assign n185 = G136 & G154 ;
  buffer buf_n186( .i (n185), .o (n186) );
  inverter inv_n2980( .i (n186), .o (n2980) );
  assign n187 = G11 & G12 ;
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  assign n192 = ~G65 | ~n191 ;
  inverter inv_n2981( .i (n188), .o (n2981) );
  assign n193 = G163 & G34 ;
  assign n194 = ~G163 & G33 ;
  assign n195 = n193 | n194 ;
  assign n196 = ~n191 | ~n195 ;
  assign n197 = G13 & G163 ;
  assign n198 = ~G163 & G35 ;
  assign n199 = n197 | n198 ;
  assign n200 = n190 & n199 ;
  inverter inv_n201( .i (n200), .o (n201) );
  assign n202 = ~G32 | ~n191 ;
  assign n203 = ~G163 & G9 ;
  assign n204 = G163 & G8 ;
  assign n205 = n189 & ~n204 ;
  assign n206 = ~n203 & n205 ;
  assign n207 = G66 & ~n206 ;
  assign n208 = ~G163 & G30 ;
  assign n209 = G10 & G163 ;
  assign n210 = n189 & ~n209 ;
  assign n211 = ~n208 & n210 ;
  assign n212 = G66 & ~n211 ;
  assign n213 = ~G163 & G7 ;
  assign n214 = G163 & G28 ;
  assign n215 = n189 & ~n214 ;
  assign n216 = ~n213 & n215 ;
  assign n217 = G66 & ~n216 ;
  assign n218 = ~G163 & G29 ;
  assign n219 = G163 & G31 ;
  buffer buf_n220( .i (n188), .o (n220) );
  assign n221 = ~n219 & n220 ;
  assign n222 = ~n218 & n221 ;
  assign n223 = G66 & ~n222 ;
  assign n224 = G100 | G117 ;
  assign n225 = ~G101 & G117 ;
  assign n226 = n224 & ~n225 ;
  assign n227 = G145 & ~n226 ;
  assign n228 = G102 & G117 ;
  assign n229 = ~G117 & G98 ;
  assign n230 = n228 | n229 ;
  assign n231 = ~G145 & n230 ;
  assign n232 = n227 | n231 ;
  buffer buf_n233( .i (n232), .o (n233) );
  assign n243 = G100 | G119 ;
  assign n244 = ~G101 & G119 ;
  assign n245 = n243 & ~n244 ;
  assign n246 = G146 & ~n245 ;
  assign n247 = G102 & G119 ;
  assign n248 = ~G119 & G98 ;
  assign n249 = n247 | n248 ;
  assign n250 = ~G146 & n249 ;
  assign n251 = n246 | n250 ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n262 = n233 & n252 ;
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  assign n274 = G128 | G169 ;
  assign n275 = G128 & ~G168 ;
  assign n276 = n274 & ~n275 ;
  assign n277 = G150 & ~n276 ;
  assign n278 = G128 & G167 ;
  assign n279 = ~G128 & G166 ;
  assign n280 = n278 | n279 ;
  assign n281 = ~G150 & n280 ;
  assign n282 = n277 | n281 ;
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  assign n285 = G113 | G98 ;
  assign n286 = ~G102 & G113 ;
  assign n287 = n285 & ~n286 ;
  buffer buf_n288( .i (n287), .o (n288) );
  assign n304 = G100 | G115 ;
  assign n305 = ~G101 & G115 ;
  assign n306 = n304 & ~n305 ;
  buffer buf_n307( .i (n306), .o (n307) );
  assign n318 = n288 & ~n307 ;
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  assign n327 = G100 | G130 ;
  assign n328 = ~G101 & G130 ;
  assign n329 = n327 & ~n328 ;
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  assign n343 = ~G148 & G166 ;
  assign n344 = G148 & ~G169 ;
  assign n345 = n343 | n344 ;
  buffer buf_n346( .i (n345), .o (n346) );
  assign n347 = ~n340 & n346 ;
  assign n348 = n326 & n347 ;
  assign n349 = n284 & n348 ;
  assign n350 = G121 | G169 ;
  assign n351 = G121 & ~G168 ;
  assign n352 = n350 & ~n351 ;
  assign n353 = G147 & ~n352 ;
  assign n354 = G121 & G167 ;
  assign n355 = ~G121 & G166 ;
  assign n356 = n354 | n355 ;
  assign n357 = ~G147 & n356 ;
  assign n358 = n353 | n357 ;
  buffer buf_n359( .i (n358), .o (n359) );
  assign n360 = G126 | G169 ;
  assign n361 = G126 & ~G168 ;
  assign n362 = n360 & ~n361 ;
  assign n363 = G149 & ~n362 ;
  assign n364 = G126 & G167 ;
  assign n365 = ~G126 & G166 ;
  assign n366 = n364 | n365 ;
  assign n367 = ~G149 & n366 ;
  assign n368 = n363 | n367 ;
  buffer buf_n369( .i (n368), .o (n369) );
  assign n370 = n359 & n369 ;
  assign n371 = n349 & n370 ;
  assign n372 = n273 & n371 ;
  assign n373 = G169 | G94 ;
  assign n374 = ~G168 & G94 ;
  assign n375 = n373 & ~n374 ;
  assign n376 = G140 & ~n375 ;
  assign n377 = G167 & G94 ;
  assign n378 = G166 & ~G94 ;
  assign n379 = n377 | n378 ;
  assign n380 = ~G140 & n379 ;
  assign n381 = n376 | n380 ;
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  assign n385 = G169 | G90 ;
  assign n386 = ~G168 & G90 ;
  assign n387 = n385 & ~n386 ;
  assign n388 = G143 & ~n387 ;
  assign n389 = G167 & G90 ;
  assign n390 = G166 & ~G90 ;
  assign n391 = n389 | n390 ;
  assign n392 = ~G143 & n391 ;
  assign n393 = n388 | n392 ;
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  assign n396 = G169 | G92 ;
  assign n397 = ~G168 & G92 ;
  assign n398 = n396 & ~n397 ;
  assign n399 = G144 & ~n398 ;
  assign n400 = G167 & G92 ;
  assign n401 = G166 & ~G92 ;
  assign n402 = n400 | n401 ;
  assign n403 = ~G144 & n402 ;
  assign n404 = n399 | n403 ;
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  assign n407 = n395 & n406 ;
  assign n408 = n384 & n407 ;
  assign n409 = G109 | G169 ;
  assign n410 = G109 & ~G168 ;
  assign n411 = n409 & ~n410 ;
  assign n412 = G135 & ~n411 ;
  assign n413 = G109 & G167 ;
  assign n414 = ~G109 & G166 ;
  assign n415 = n413 | n414 ;
  assign n416 = ~G135 & n415 ;
  assign n417 = n412 | n416 ;
  buffer buf_n418( .i (n417), .o (n418) );
  assign n419 = G169 | G96 ;
  assign n420 = ~G168 & G96 ;
  assign n421 = n419 & ~n420 ;
  assign n422 = G141 & ~n421 ;
  assign n423 = G167 & G96 ;
  assign n424 = G166 & ~G96 ;
  assign n425 = n423 | n424 ;
  assign n426 = ~G141 & n425 ;
  assign n427 = n422 | n426 ;
  buffer buf_n428( .i (n427), .o (n428) );
  assign n429 = n418 & n428 ;
  assign n430 = G107 | G169 ;
  assign n431 = G107 & ~G168 ;
  assign n432 = n430 & ~n431 ;
  assign n433 = G139 & ~n432 ;
  assign n434 = G107 & G167 ;
  assign n435 = ~G107 & G166 ;
  assign n436 = n434 | n435 ;
  assign n437 = ~G139 & n436 ;
  assign n438 = n433 | n437 ;
  buffer buf_n439( .i (n438), .o (n439) );
  assign n440 = G101 | G88 ;
  assign n441 = ~G100 & G88 ;
  assign n442 = n440 & ~n441 ;
  assign n443 = G142 & ~n442 ;
  assign n444 = G88 & G98 ;
  assign n445 = G102 & ~G88 ;
  assign n446 = n444 | n445 ;
  assign n447 = ~G142 & n446 ;
  assign n448 = n443 | n447 ;
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  assign n459 = n439 & n456 ;
  assign n460 = G103 | G169 ;
  assign n461 = G103 & ~G168 ;
  assign n462 = n460 & ~n461 ;
  assign n463 = G137 & ~n462 ;
  assign n464 = G103 & G167 ;
  assign n465 = ~G103 & G166 ;
  assign n466 = n464 | n465 ;
  assign n467 = ~G137 & n466 ;
  assign n468 = n463 | n467 ;
  buffer buf_n469( .i (n468), .o (n469) );
  assign n470 = G105 | G169 ;
  assign n471 = G105 & ~G168 ;
  assign n472 = n470 & ~n471 ;
  assign n473 = G138 & ~n472 ;
  assign n474 = G105 & G167 ;
  assign n475 = ~G105 & G166 ;
  assign n476 = n474 | n475 ;
  assign n477 = ~G138 & n476 ;
  assign n478 = n473 | n477 ;
  buffer buf_n479( .i (n478), .o (n479) );
  assign n480 = n469 & n479 ;
  assign n481 = n459 & n480 ;
  assign n482 = n429 & n481 ;
  assign n483 = n408 & n482 ;
  assign n484 = G124 & G96 ;
  assign n485 = ~G124 & G97 ;
  assign n486 = n484 | n485 ;
  buffer buf_n487( .i (n486), .o (n487) );
  assign n505 = G141 & n487 ;
  buffer buf_n506( .i (n505), .o (n506) );
  assign n510 = G141 | n487 ;
  buffer buf_n511( .i (n510), .o (n511) );
  assign n514 = ~n506 & n511 ;
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  assign n523 = G109 & G124 ;
  assign n524 = G110 & ~G124 ;
  assign n525 = n523 | n524 ;
  buffer buf_n526( .i (n525), .o (n526) );
  assign n549 = G135 & n526 ;
  buffer buf_n550( .i (n549), .o (n550) );
  assign n562 = G135 | n526 ;
  buffer buf_n563( .i (n562), .o (n563) );
  assign n572 = ~n550 & n563 ;
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  assign n590 = G107 & G124 ;
  assign n591 = G108 & ~G124 ;
  assign n592 = n590 | n591 ;
  buffer buf_n593( .i (n592), .o (n593) );
  assign n616 = G139 | n593 ;
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  assign n626 = G139 & n593 ;
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  assign n643 = n618 & ~n628 ;
  buffer buf_n644( .i (n643), .o (n644) );
  assign n659 = n574 & n644 ;
  buffer buf_n660( .i (n659), .o (n660) );
  assign n664 = G105 & G124 ;
  assign n665 = G106 & ~G124 ;
  assign n666 = n664 | n665 ;
  buffer buf_n667( .i (n666), .o (n667) );
  assign n689 = G138 & n667 ;
  buffer buf_n690( .i (n689), .o (n690) );
  assign n691 = G138 | n667 ;
  buffer buf_n692( .i (n691), .o (n692) );
  assign n695 = ~n690 & n692 ;
  buffer buf_n696( .i (n695), .o (n696) );
  assign n711 = G103 & G124 ;
  assign n712 = G104 & ~G124 ;
  assign n713 = n711 | n712 ;
  buffer buf_n714( .i (n713), .o (n714) );
  assign n736 = G137 | n714 ;
  buffer buf_n737( .i (n736), .o (n737) );
  assign n743 = G137 & n714 ;
  buffer buf_n744( .i (n743), .o (n744) );
  assign n751 = n737 & ~n744 ;
  buffer buf_n752( .i (n751), .o (n752) );
  assign n767 = n696 & n752 ;
  buffer buf_n768( .i (n767), .o (n768) );
  assign n778 = n660 & n768 ;
  buffer buf_n779( .i (n778), .o (n779) );
  assign n790 = n518 & n779 ;
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  assign n801 = G124 & G88 ;
  assign n802 = ~G124 & G89 ;
  assign n803 = n801 | n802 ;
  buffer buf_n804( .i (n803), .o (n804) );
  assign n825 = G142 & n804 ;
  buffer buf_n826( .i (n825), .o (n826) );
  assign n846 = G142 | n804 ;
  buffer buf_n847( .i (n846), .o (n847) );
  assign n866 = ~n826 & n847 ;
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  assign n886 = G124 & G90 ;
  assign n887 = ~G124 & G91 ;
  assign n888 = n886 | n887 ;
  buffer buf_n889( .i (n888), .o (n889) );
  assign n913 = G143 & n889 ;
  buffer buf_n914( .i (n913), .o (n914) );
  assign n931 = G143 | n889 ;
  buffer buf_n932( .i (n931), .o (n932) );
  assign n941 = ~n914 & n932 ;
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  assign n959 = G124 & G92 ;
  assign n960 = ~G124 & G93 ;
  assign n961 = n959 | n960 ;
  buffer buf_n962( .i (n961), .o (n962) );
  assign n988 = G144 & n962 ;
  buffer buf_n989( .i (n988), .o (n989) );
  assign n992 = G144 | n962 ;
  buffer buf_n993( .i (n992), .o (n993) );
  assign n994 = ~n989 & n993 ;
  buffer buf_n995( .i (n994), .o (n995) );
  assign n1014 = G124 & G94 ;
  assign n1015 = ~G124 & G95 ;
  assign n1016 = n1014 | n1015 ;
  buffer buf_n1017( .i (n1016), .o (n1017) );
  assign n1040 = G140 & n1017 ;
  buffer buf_n1041( .i (n1040), .o (n1041) );
  assign n1059 = G140 | n1017 ;
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1078 = ~n1041 & n1060 ;
  buffer buf_n1079( .i (n1078), .o (n1079) );
  assign n1098 = n995 & n1079 ;
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  assign n1113 = n955 & n1112 ;
  buffer buf_n1114( .i (n1113), .o (n1114) );
  assign n1115 = n882 & n1114 ;
  buffer buf_n1116( .i (n1115), .o (n1116) );
  assign n1117 = n800 & n1116 ;
  buffer buf_n1118( .i (n1117), .o (n1118) );
  assign n1119 = G123 | G125 ;
  buffer buf_n1120( .i (n1119), .o (n1120) );
  assign n1135 = G148 & n1120 ;
  buffer buf_n1136( .i (n1135), .o (n1136) );
  assign n1145 = G148 | n1120 ;
  buffer buf_n1146( .i (n1145), .o (n1146) );
  assign n1155 = ~n1136 & n1146 ;
  buffer buf_n1156( .i (n1155), .o (n1156) );
  assign n1167 = G123 & G128 ;
  assign n1168 = ~G123 & G129 ;
  assign n1169 = n1167 | n1168 ;
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  assign n1189 = G150 | n1172 ;
  buffer buf_n1190( .i (n1189), .o (n1190) );
  assign n1205 = G123 & G130 ;
  assign n1206 = ~G123 & G131 ;
  assign n1207 = n1205 | n1206 ;
  buffer buf_n1208( .i (n1207), .o (n1208) );
  assign n1228 = G150 & n1170 ;
  buffer buf_n1229( .i (n1228), .o (n1229) );
  assign n1246 = n1208 | n1229 ;
  buffer buf_n1247( .i (n1246), .o (n1247) );
  assign n1252 = n1190 & ~n1247 ;
  buffer buf_n1253( .i (n1252), .o (n1253) );
  assign n1268 = G123 & G126 ;
  assign n1269 = ~G123 & G127 ;
  assign n1270 = n1268 | n1269 ;
  buffer buf_n1271( .i (n1270), .o (n1271) );
  assign n1288 = G149 & n1271 ;
  buffer buf_n1289( .i (n1288), .o (n1289) );
  assign n1292 = G149 | n1271 ;
  buffer buf_n1293( .i (n1292), .o (n1293) );
  assign n1295 = ~n1289 & n1293 ;
  buffer buf_n1296( .i (n1295), .o (n1296) );
  assign n1311 = n1253 & n1296 ;
  buffer buf_n1312( .i (n1311), .o (n1312) );
  assign n1317 = n1156 & n1312 ;
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  assign n1332 = G117 & G123 ;
  assign n1333 = G118 & ~G123 ;
  assign n1334 = n1332 | n1333 ;
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  assign n1339 = G145 & n1336 ;
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  assign n1346 = G145 | n1337 ;
  buffer buf_n1347( .i (n1346), .o (n1347) );
  assign n1351 = ~n1341 & n1347 ;
  buffer buf_n1352( .i (n1351), .o (n1352) );
  assign n1357 = G119 & G123 ;
  assign n1358 = G120 & ~G123 ;
  assign n1359 = n1357 | n1358 ;
  buffer buf_n1360( .i (n1359), .o (n1360) );
  assign n1375 = G146 & n1360 ;
  buffer buf_n1376( .i (n1375), .o (n1376) );
  assign n1384 = G146 | n1360 ;
  buffer buf_n1385( .i (n1384), .o (n1385) );
  assign n1393 = ~n1376 & n1385 ;
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  assign n1403 = n1352 & n1398 ;
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  buffer buf_n1409( .i (n1408), .o (n1409) );
  assign n1410 = G113 & G123 ;
  assign n1411 = G114 & ~G123 ;
  assign n1412 = n1410 | n1411 ;
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  assign n1428 = G115 & G123 ;
  assign n1429 = G116 & ~G123 ;
  assign n1430 = n1428 | n1429 ;
  buffer buf_n1431( .i (n1430), .o (n1431) );
  assign n1434 = n1421 | n1431 ;
  buffer buf_n1435( .i (n1434), .o (n1435) );
  assign n1436 = G122 | G123 ;
  buffer buf_n1437( .i (n1436), .o (n1437) );
  assign n1454 = ~G121 & G123 ;
  assign n1455 = n1437 & ~n1454 ;
  buffer buf_n1456( .i (n1455), .o (n1456) );
  assign n1471 = G147 & n1456 ;
  buffer buf_n1472( .i (n1471), .o (n1472) );
  assign n1480 = G147 | n1456 ;
  buffer buf_n1481( .i (n1480), .o (n1481) );
  assign n1488 = ~n1472 & n1481 ;
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  assign n1503 = ~n1435 & n1502 ;
  assign n1504 = n1409 & n1503 ;
  assign n1505 = n1331 & n1504 ;
  buffer buf_n1506( .i (n1505), .o (n1506) );
  assign n1507 = G113 | G115 ;
  assign n1508 = G113 & G115 ;
  assign n1509 = n1507 & ~n1508 ;
  buffer buf_n1510( .i (n1509), .o (n1510) );
  assign n1511 = G117 & ~G119 ;
  assign n1512 = ~G117 & G119 ;
  assign n1513 = n1511 | n1512 ;
  buffer buf_n1514( .i (n1513), .o (n1514) );
  assign n1515 = ~n1510 & n1514 ;
  assign n1516 = n1510 & ~n1514 ;
  assign n1517 = n1515 | n1516 ;
  buffer buf_n1518( .i (n1517), .o (n1518) );
  assign n1519 = G130 & ~G132 ;
  assign n1520 = ~G130 & G132 ;
  assign n1521 = n1519 | n1520 ;
  buffer buf_n1522( .i (n1521), .o (n1522) );
  assign n1523 = G121 & ~n1522 ;
  assign n1524 = ~G121 & n1522 ;
  assign n1525 = n1523 | n1524 ;
  buffer buf_n1526( .i (n1525), .o (n1526) );
  assign n1527 = G126 & ~G128 ;
  assign n1528 = ~G126 & G128 ;
  assign n1529 = n1527 | n1528 ;
  buffer buf_n1530( .i (n1529), .o (n1530) );
  assign n1531 = n1526 & ~n1530 ;
  assign n1532 = ~n1526 & n1530 ;
  assign n1533 = n1531 | n1532 ;
  buffer buf_n1534( .i (n1533), .o (n1534) );
  assign n1535 = n1518 | n1534 ;
  assign n1536 = n1518 & n1534 ;
  assign n1537 = n1535 & ~n1536 ;
  buffer buf_n1538( .i (n1537), .o (n1538) );
  inverter inv_n2982( .i (n1538), .o (n2982) );
  assign n1539 = G88 | G90 ;
  assign n1540 = G88 & G90 ;
  assign n1541 = n1539 & ~n1540 ;
  buffer buf_n1542( .i (n1541), .o (n1542) );
  assign n1543 = G92 & ~G94 ;
  assign n1544 = ~G92 & G94 ;
  assign n1545 = n1543 | n1544 ;
  buffer buf_n1546( .i (n1545), .o (n1546) );
  assign n1547 = ~n1542 & n1546 ;
  assign n1548 = n1542 & ~n1546 ;
  assign n1549 = n1547 | n1548 ;
  buffer buf_n1550( .i (n1549), .o (n1550) );
  assign n1551 = G103 | G96 ;
  assign n1552 = G103 & G96 ;
  assign n1553 = n1551 & ~n1552 ;
  buffer buf_n1554( .i (n1553), .o (n1554) );
  assign n1555 = G109 & ~G111 ;
  assign n1556 = ~G109 & G111 ;
  assign n1557 = n1555 | n1556 ;
  buffer buf_n1558( .i (n1557), .o (n1558) );
  assign n1559 = n1554 | n1558 ;
  assign n1560 = n1554 & n1558 ;
  assign n1561 = n1559 & ~n1560 ;
  buffer buf_n1562( .i (n1561), .o (n1562) );
  assign n1563 = G105 & ~G107 ;
  assign n1564 = ~G105 & G107 ;
  assign n1565 = n1563 | n1564 ;
  buffer buf_n1566( .i (n1565), .o (n1566) );
  assign n1567 = n1562 & ~n1566 ;
  assign n1568 = ~n1562 & n1566 ;
  assign n1569 = n1567 | n1568 ;
  buffer buf_n1570( .i (n1569), .o (n1570) );
  assign n1571 = n1550 & n1570 ;
  assign n1572 = n1550 | n1570 ;
  assign n1573 = ~n1571 & n1572 ;
  buffer buf_n1574( .i (n1573), .o (n1574) );
  inverter inv_n2983( .i (n1574), .o (n2983) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  assign n1575 = n550 & n617 ;
  buffer buf_n1576( .i (n1575), .o (n1576) );
  assign n1582 = n628 | n690 ;
  assign n1583 = n1576 | n1582 ;
  assign n1584 = n694 & n1583 ;
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n753( .i (n752), .o (n753) );
  assign n1595 = n515 & n753 ;
  assign n1596 = n1585 & n1595 ;
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  assign n1597 = n513 & n747 ;
  assign n1598 = n509 | n1597 ;
  assign n1599 = n1596 | n1598 ;
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  assign n1611 = n1116 & n1610 ;
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  assign n1612 = n993 & n1041 ;
  buffer buf_n1613( .i (n1612), .o (n1613) );
  assign n1619 = n991 | n1613 ;
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  assign n1635 = n936 & n1622 ;
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n1637( .i (n1636), .o (n1637) );
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  assign n1647 = n930 | n1646 ;
  buffer buf_n1648( .i (n1647), .o (n1648) );
  assign n1649 = n865 & n1648 ;
  assign n1650 = n845 | n1649 ;
  assign n1651 = n1611 | n1650 ;
  buffer buf_n1652( .i (n1651), .o (n1652) );
  assign n1653 = ~n1421 & n1431 ;
  inverter inv_n1654( .i (n1653), .o (n1654) );
  assign n1655 = G176 & ~G177 ;
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  buffer buf_n1658( .i (n1657), .o (n1658) );
  assign n1665 = G60 & n1658 ;
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  assign n1666 = ~G21 & n1226 ;
  assign n1667 = G21 & ~n1226 ;
  assign n1668 = n1666 | n1667 ;
  buffer buf_n1669( .i (n1668), .o (n1669) );
  assign n1670 = ~G176 & n1669 ;
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  assign n1671 = G176 & ~n342 ;
  assign n1672 = G177 & ~n1671 ;
  assign n1673 = ~n1670 & n1672 ;
  assign n1674 = n1665 | n1673 ;
  buffer buf_n1675( .i (n1674), .o (n1675) );
  inverter inv_n2984( .i (n1675), .o (n2984) );
  assign n1677 = G58 & n1657 ;
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  assign n1678 = n1204 & ~n1245 ;
  assign n1679 = n1225 & ~n1678 ;
  assign n1680 = n1267 | n1679 ;
  buffer buf_n1681( .i (n1680), .o (n1681) );
  assign n1684 = G176 | n1681 ;
  assign n1685 = G176 & n283 ;
  assign n1686 = G177 & ~n1685 ;
  assign n1687 = n1684 & n1686 ;
  assign n1688 = n1677 | n1687 ;
  buffer buf_n1689( .i (n1688), .o (n1689) );
  inverter inv_n2985( .i (n1689), .o (n2985) );
  assign n1692 = G48 & n1658 ;
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  assign n1693 = G2 & n580 ;
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  assign n1703 = G2 | n589 ;
  assign n1704 = ~n1702 & n1703 ;
  buffer buf_n1705( .i (n1704), .o (n1705) );
  assign n1706 = G176 | n1705 ;
  assign n1707 = G176 & n418 ;
  assign n1708 = G177 & ~n1707 ;
  assign n1709 = n1706 & n1708 ;
  assign n1710 = n1692 | n1709 ;
  buffer buf_n1711( .i (n1710), .o (n1711) );
  inverter inv_n2986( .i (n1711), .o (n2986) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  assign n1714 = n1422 & n1432 ;
  assign n1715 = n1435 & ~n1714 ;
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  assign n1724 = G173 | n1713 ;
  buffer buf_n1676( .i (n1675), .o (n1676) );
  assign n1725 = G173 & ~n1676 ;
  assign n1726 = G172 & ~n1725 ;
  assign n1727 = n1724 & n1726 ;
  assign n1728 = ~G172 & G173 ;
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  assign n1731 = G3 & n1730 ;
  assign n1732 = G172 | G173 ;
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  assign n1735 = G22 & ~n1734 ;
  assign n1736 = n1731 | n1735 ;
  assign n1737 = n1727 | n1736 ;
  assign n1738 = G19 & n1658 ;
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  assign n1739 = n1232 & n1294 ;
  assign n1740 = n1291 | n1739 ;
  buffer buf_n1741( .i (n1740), .o (n1741) );
  assign n1746 = n1138 | n1741 ;
  assign n1747 = n1149 & n1746 ;
  assign n1748 = n1318 | n1747 ;
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  assign n1758 = n1501 | n1757 ;
  assign n1759 = n1501 & n1757 ;
  assign n1760 = n1758 & ~n1759 ;
  buffer buf_n1761( .i (n1760), .o (n1761) );
  assign n1766 = ~G176 & n1761 ;
  assign n1767 = G176 & n359 ;
  assign n1768 = G177 & ~n1767 ;
  assign n1769 = ~n1766 & n1768 ;
  assign n1770 = n1738 | n1769 ;
  buffer buf_n1771( .i (n1770), .o (n1771) );
  inverter inv_n2987( .i (n1771), .o (n2987) );
  assign n1773 = G59 & n1656 ;
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  assign n1774 = n1316 | n1745 ;
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  assign n1780 = ~n1166 & n1779 ;
  assign n1781 = n1166 & ~n1779 ;
  assign n1782 = n1780 | n1781 ;
  buffer buf_n1783( .i (n1782), .o (n1783) );
  assign n1789 = ~G176 & n1783 ;
  assign n1790 = G176 & n346 ;
  assign n1791 = G177 & ~n1790 ;
  assign n1792 = ~n1789 & n1791 ;
  assign n1793 = n1773 | n1792 ;
  buffer buf_n1794( .i (n1793), .o (n1794) );
  inverter inv_n2988( .i (n1794), .o (n2988) );
  buffer buf_n1798( .i (n1657), .o (n1798) );
  assign n1799 = G50 & n1798 ;
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  assign n1800 = n1245 | n1265 ;
  buffer buf_n1801( .i (n1800), .o (n1801) );
  assign n1802 = n1310 | n1801 ;
  assign n1803 = n1310 & n1801 ;
  assign n1804 = n1802 & ~n1803 ;
  buffer buf_n1805( .i (n1804), .o (n1805) );
  assign n1808 = ~G176 & n1805 ;
  assign n1809 = G176 & n369 ;
  assign n1810 = G177 & ~n1809 ;
  assign n1811 = ~n1808 & n1810 ;
  assign n1812 = n1799 | n1811 ;
  buffer buf_n1813( .i (n1812), .o (n1813) );
  inverter inv_n2989( .i (n1813), .o (n2989) );
  assign n1815 = G174 | n1713 ;
  assign n1816 = G174 & ~n1676 ;
  assign n1817 = G175 & ~n1816 ;
  assign n1818 = n1815 & n1817 ;
  assign n1819 = G174 & ~G175 ;
  buffer buf_n1820( .i (n1819), .o (n1820) );
  buffer buf_n1821( .i (n1820), .o (n1821) );
  assign n1822 = G3 & n1821 ;
  assign n1823 = G174 | G175 ;
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1825( .i (n1824), .o (n1825) );
  assign n1826 = G22 & ~n1825 ;
  assign n1827 = n1822 | n1826 ;
  assign n1828 = n1818 | n1827 ;
  assign n1829 = G53 & n1798 ;
  assign n1830 = G2 & n791 ;
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  assign n1840 = G2 & n789 ;
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  assign n1841 = n742 & n1586 ;
  assign n1842 = n750 | n1841 ;
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  assign n1846 = ~n522 & n1845 ;
  assign n1847 = n522 & ~n1845 ;
  assign n1848 = n1846 | n1847 ;
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  assign n1854 = n1840 | n1853 ;
  assign n1855 = ~n1839 & n1854 ;
  buffer buf_n1856( .i (n1855), .o (n1856) );
  assign n1860 = ~G176 & n1856 ;
  assign n1861 = G176 & n428 ;
  assign n1862 = G177 & ~n1861 ;
  assign n1863 = ~n1860 & n1862 ;
  assign n1864 = n1829 | n1863 ;
  buffer buf_n1865( .i (n1864), .o (n1865) );
  inverter inv_n2990( .i (n1865), .o (n2990) );
  assign n1868 = G57 & n1657 ;
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  assign n1869 = n663 & n701 ;
  assign n1870 = n1589 | n1869 ;
  buffer buf_n1871( .i (n1870), .o (n1871) );
  buffer buf_n1872( .i (n1871), .o (n1872) );
  buffer buf_n1873( .i (n1872), .o (n1873) );
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  assign n1876 = G2 | n1594 ;
  assign n1877 = n1875 & n1876 ;
  buffer buf_n1878( .i (n1877), .o (n1878) );
  assign n1879 = ~n766 & n1878 ;
  assign n1880 = n766 & ~n1878 ;
  assign n1881 = n1879 | n1880 ;
  buffer buf_n1882( .i (n1881), .o (n1882) );
  assign n1885 = ~G176 & n1882 ;
  assign n1886 = G176 & n469 ;
  assign n1887 = G177 & ~n1886 ;
  assign n1888 = ~n1885 & n1887 ;
  assign n1889 = n1868 | n1888 ;
  buffer buf_n1890( .i (n1889), .o (n1890) );
  inverter inv_n2991( .i (n1890), .o (n2991) );
  buffer buf_n1894( .i (n1656), .o (n1894) );
  assign n1895 = G56 & n1894 ;
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  assign n1896 = n561 | n1694 ;
  buffer buf_n1897( .i (n1896), .o (n1897) );
  assign n1902 = n654 & n1897 ;
  buffer buf_n1903( .i (n1902), .o (n1903) );
  assign n1907 = n642 | n1903 ;
  buffer buf_n1908( .i (n1907), .o (n1908) );
  assign n1909 = n710 | n1908 ;
  assign n1910 = n710 & n1908 ;
  assign n1911 = n1909 & ~n1910 ;
  buffer buf_n1912( .i (n1911), .o (n1912) );
  assign n1916 = ~G176 & n1912 ;
  assign n1917 = G176 & n479 ;
  assign n1918 = G177 & ~n1917 ;
  assign n1919 = ~n1916 & n1918 ;
  assign n1920 = n1895 | n1919 ;
  buffer buf_n1921( .i (n1920), .o (n1921) );
  inverter inv_n2992( .i (n1921), .o (n2992) );
  assign n1925 = G55 & n1894 ;
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  assign n1926 = n658 | n1901 ;
  assign n1927 = ~n1906 & n1926 ;
  buffer buf_n1928( .i (n1927), .o (n1928) );
  assign n1930 = ~G176 & n1928 ;
  assign n1931 = G176 & n439 ;
  assign n1932 = G177 & ~n1931 ;
  assign n1933 = ~n1930 & n1932 ;
  assign n1934 = n1925 | n1933 ;
  buffer buf_n1935( .i (n1934), .o (n1935) );
  inverter inv_n2993( .i (n1935), .o (n2993) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  assign n1939 = n1338 & n1414 ;
  assign n1940 = n1338 | n1414 ;
  assign n1941 = ~n1939 & n1940 ;
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  assign n1952 = n1374 & n1433 ;
  assign n1953 = n1374 | n1433 ;
  assign n1954 = ~n1952 & n1953 ;
  buffer buf_n1955( .i (n1954), .o (n1955) );
  assign n1956 = ~n1951 & n1955 ;
  assign n1957 = n1951 & ~n1955 ;
  assign n1958 = n1956 | n1957 ;
  buffer buf_n1959( .i (n1958), .o (n1959) );
  assign n1960 = G123 & G132 ;
  assign n1961 = ~G123 & G133 ;
  assign n1962 = n1960 | n1961 ;
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  assign n1964 = n1188 | n1287 ;
  assign n1965 = n1188 & n1287 ;
  assign n1966 = n1964 & ~n1965 ;
  buffer buf_n1967( .i (n1966), .o (n1967) );
  assign n1968 = n1963 | n1967 ;
  assign n1969 = n1963 & n1967 ;
  assign n1970 = n1968 & ~n1969 ;
  buffer buf_n1971( .i (n1970), .o (n1971) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  assign n1972 = n1134 & n1470 ;
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  assign n1973 = G125 | n1453 ;
  assign n1974 = ~n1972 & n1973 ;
  buffer buf_n1975( .i (n1974), .o (n1975) );
  assign n1976 = ~n1227 & n1975 ;
  assign n1977 = n1227 & ~n1975 ;
  assign n1978 = n1976 | n1977 ;
  buffer buf_n1979( .i (n1978), .o (n1979) );
  assign n1980 = n1971 & ~n1979 ;
  assign n1981 = ~n1971 & n1979 ;
  assign n1982 = n1980 | n1981 ;
  buffer buf_n1983( .i (n1982), .o (n1983) );
  assign n1984 = ~n1959 & n1983 ;
  assign n1985 = n1959 & ~n1983 ;
  assign n1986 = n1984 | n1985 ;
  buffer buf_n1987( .i (n1986), .o (n1987) );
  inverter inv_n2994( .i (n1987), .o (n2994) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  assign n1988 = n688 & n735 ;
  assign n1989 = n688 | n735 ;
  assign n1990 = ~n1988 & n1989 ;
  buffer buf_n1991( .i (n1990), .o (n1991) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  assign n1992 = ~n548 & n615 ;
  assign n1993 = n548 & ~n615 ;
  assign n1994 = n1992 | n1993 ;
  buffer buf_n1995( .i (n1994), .o (n1995) );
  assign n1996 = n1991 | n1995 ;
  assign n1997 = n1991 & n1995 ;
  assign n1998 = n1996 & ~n1997 ;
  buffer buf_n1999( .i (n1998), .o (n1999) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  assign n2000 = n912 & n987 ;
  assign n2001 = n912 | n987 ;
  assign n2002 = ~n2000 & n2001 ;
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  assign n2004 = G111 & G124 ;
  assign n2005 = G112 & ~G124 ;
  assign n2006 = n2004 | n2005 ;
  buffer buf_n2007( .i (n2006), .o (n2007) );
  assign n2008 = n1039 & ~n2007 ;
  assign n2009 = ~n1039 & n2007 ;
  assign n2010 = n2008 | n2009 ;
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  assign n2012 = ~n504 & n824 ;
  assign n2013 = n504 & ~n824 ;
  assign n2014 = n2012 | n2013 ;
  buffer buf_n2015( .i (n2014), .o (n2015) );
  assign n2016 = ~n2011 & n2015 ;
  assign n2017 = n2011 & ~n2015 ;
  assign n2018 = n2016 | n2017 ;
  buffer buf_n2019( .i (n2018), .o (n2019) );
  assign n2020 = ~n2003 & n2019 ;
  assign n2021 = n2003 & ~n2019 ;
  assign n2022 = n2020 | n2021 ;
  buffer buf_n2023( .i (n2022), .o (n2023) );
  assign n2024 = ~n1999 & n2023 ;
  assign n2025 = n1999 & ~n2023 ;
  assign n2026 = n2024 | n2025 ;
  buffer buf_n2027( .i (n2026), .o (n2027) );
  inverter inv_n2995( .i (n2027), .o (n2995) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  assign n2028 = n1603 | n1831 ;
  buffer buf_n2029( .i (n2028), .o (n2029) );
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n2031( .i (n2030), .o (n2031) );
  buffer buf_n2032( .i (n2031), .o (n2032) );
  assign n2034 = n1114 & n2032 ;
  assign n2035 = n1648 | n2034 ;
  buffer buf_n2036( .i (n2035), .o (n2036) );
  assign n2037 = n885 | n2036 ;
  assign n2038 = n885 & n2036 ;
  assign n2039 = n2037 & ~n2038 ;
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n2033( .i (n2032), .o (n2033) );
  assign n2045 = n1097 | n2033 ;
  assign n2046 = n1097 & n2033 ;
  assign n2047 = n2045 & ~n2046 ;
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n1915( .i (n1914), .o (n1915) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  assign n2054 = ~n1705 & n1929 ;
  assign n2055 = n1884 & n2054 ;
  assign n2056 = n1915 & n2055 ;
  assign n2057 = n1859 & n2056 ;
  assign n2058 = ~n2053 & n2057 ;
  assign n2059 = n2044 & n2058 ;
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n1633( .i (n1632), .o (n1633) );
  buffer buf_n1634( .i (n1633), .o (n1634) );
  assign n2060 = n1112 & n2030 ;
  assign n2061 = n1634 | n2060 ;
  buffer buf_n2062( .i (n2061), .o (n2062) );
  assign n2063 = ~n958 & n2062 ;
  assign n2064 = n958 & ~n2062 ;
  assign n2065 = n2063 | n2064 ;
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  assign n2073 = n1077 & n2030 ;
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  assign n2074 = n1058 | n2030 ;
  assign n2075 = ~n2073 & n2074 ;
  buffer buf_n2076( .i (n2075), .o (n2076) );
  assign n2077 = n1013 | n2076 ;
  assign n2078 = n1013 & n2076 ;
  assign n2079 = n2077 & ~n2078 ;
  buffer buf_n2080( .i (n2079), .o (n2080) );
  buffer buf_n2081( .i (n2080), .o (n2081) );
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  assign n2087 = n2072 & ~n2086 ;
  assign n2088 = n2059 & n2087 ;
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  assign n2089 = n1487 & n1749 ;
  assign n2090 = n1479 | n2089 ;
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  assign n2096 = n1392 & n2092 ;
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  assign n2097 = n1383 | n2092 ;
  assign n2098 = ~n2096 & n2097 ;
  buffer buf_n2099( .i (n2098), .o (n2099) );
  assign n2100 = n1356 & n2099 ;
  assign n2101 = n1356 | n2099 ;
  assign n2102 = ~n2100 & n2101 ;
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n2111( .i (n2110), .o (n2111) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  assign n2112 = n1350 & n1383 ;
  assign n2113 = n1345 | n2112 ;
  buffer buf_n2093( .i (n2092), .o (n2093) );
  assign n2114 = n1404 & n2093 ;
  assign n2115 = n2113 | n2114 ;
  buffer buf_n2116( .i (n2115), .o (n2116) );
  assign n2117 = n1432 | n2116 ;
  assign n2118 = n1432 & n2116 ;
  assign n2119 = n2117 & ~n2118 ;
  buffer buf_n2120( .i (n2119), .o (n2120) );
  buffer buf_n2121( .i (n2120), .o (n2121) );
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  assign n2127 = n1402 & n2095 ;
  assign n2128 = n1402 | n2095 ;
  assign n2129 = ~n2127 & n2128 ;
  buffer buf_n2130( .i (n2129), .o (n2130) );
  buffer buf_n2131( .i (n2130), .o (n2131) );
  buffer buf_n2132( .i (n2131), .o (n2132) );
  buffer buf_n2133( .i (n2132), .o (n2133) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  assign n2137 = n1669 & n1716 ;
  assign n2138 = ~n1683 & n2137 ;
  assign n2139 = n1807 & n2138 ;
  assign n2140 = n1788 & n2139 ;
  assign n2141 = n1765 & n2140 ;
  assign n2142 = ~n2136 & n2141 ;
  assign n2143 = ~n2126 & n2142 ;
  assign n2144 = ~n2111 & n2143 ;
  assign n2145 = G158 | n1712 ;
  assign n2146 = G158 & ~n1675 ;
  assign n2147 = G159 & ~n2146 ;
  assign n2148 = n2145 & n2147 ;
  assign n2149 = G158 | G159 ;
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  assign n2152 = G81 & ~n2151 ;
  assign n2153 = G158 & ~G159 ;
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n2155( .i (n2154), .o (n2155) );
  assign n2156 = G80 & n2155 ;
  assign n2157 = n2152 | n2156 ;
  assign n2158 = n2148 | n2157 ;
  assign n2159 = G64 & n2158 ;
  assign n2160 = G160 | n1712 ;
  assign n2161 = G160 & ~n1675 ;
  assign n2162 = G161 & ~n2161 ;
  assign n2163 = n2160 & n2162 ;
  assign n2164 = G160 | G161 ;
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n2166( .i (n2165), .o (n2166) );
  assign n2167 = G81 & ~n2166 ;
  assign n2168 = G160 & ~G161 ;
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  assign n2171 = G80 & n2170 ;
  assign n2172 = n2167 | n2171 ;
  assign n2173 = n2163 | n2172 ;
  assign n2174 = G64 & n2173 ;
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  assign n2175 = G173 | n1867 ;
  buffer buf_n1772( .i (n1771), .o (n1772) );
  assign n2176 = G173 & ~n1772 ;
  assign n2177 = G172 & ~n2176 ;
  assign n2178 = n2175 & n2177 ;
  assign n2179 = G16 & n1730 ;
  assign n2180 = G14 & ~n1734 ;
  assign n2181 = n2179 | n2180 ;
  assign n2182 = n2178 | n2181 ;
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  assign n2183 = G173 | n1893 ;
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  assign n2184 = G173 & ~n1797 ;
  assign n2185 = G172 & ~n2184 ;
  assign n2186 = n2183 & n2185 ;
  assign n2187 = G6 & ~n1734 ;
  assign n2188 = G27 & n1730 ;
  assign n2189 = n2187 | n2188 ;
  assign n2190 = n2186 | n2189 ;
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  assign n2191 = G173 | n1924 ;
  buffer buf_n1814( .i (n1813), .o (n1814) );
  assign n2192 = G173 & ~n1814 ;
  assign n2193 = G172 & ~n2192 ;
  assign n2194 = n2191 & n2193 ;
  assign n2195 = G26 & n1730 ;
  assign n2196 = G5 & ~n1734 ;
  assign n2197 = n2195 | n2196 ;
  assign n2198 = n2194 | n2197 ;
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  assign n2199 = G173 | n1938 ;
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  assign n2200 = G173 & ~n1691 ;
  assign n2201 = G172 & ~n2200 ;
  assign n2202 = n2199 & n2201 ;
  buffer buf_n2203( .i (n1729), .o (n2203) );
  assign n2204 = G24 & n2203 ;
  buffer buf_n2205( .i (n1733), .o (n2205) );
  assign n2206 = G25 & ~n2205 ;
  assign n2207 = n2204 | n2206 ;
  assign n2208 = n2202 | n2207 ;
  assign n2209 = G174 | n1867 ;
  assign n2210 = G174 & ~n1772 ;
  assign n2211 = G175 & ~n2210 ;
  assign n2212 = n2209 & n2211 ;
  assign n2213 = G14 & ~n1825 ;
  assign n2214 = G16 & n1821 ;
  assign n2215 = n2213 | n2214 ;
  assign n2216 = n2212 | n2215 ;
  assign n2217 = G174 | n1893 ;
  assign n2218 = G174 & ~n1797 ;
  assign n2219 = G175 & ~n2218 ;
  assign n2220 = n2217 & n2219 ;
  assign n2221 = G27 & n1821 ;
  assign n2222 = G6 & ~n1825 ;
  assign n2223 = n2221 | n2222 ;
  assign n2224 = n2220 | n2223 ;
  assign n2225 = G174 | n1924 ;
  assign n2226 = G174 & ~n1814 ;
  assign n2227 = G175 & ~n2226 ;
  assign n2228 = n2225 & n2227 ;
  assign n2229 = G5 & ~n1825 ;
  assign n2230 = G26 & n1821 ;
  assign n2231 = n2229 | n2230 ;
  assign n2232 = n2228 | n2231 ;
  assign n2233 = G174 | n1938 ;
  assign n2234 = G174 & ~n1691 ;
  assign n2235 = G175 & ~n2234 ;
  assign n2236 = n2233 & n2235 ;
  buffer buf_n2237( .i (n1820), .o (n2237) );
  assign n2238 = G24 & n2237 ;
  buffer buf_n2239( .i (n1824), .o (n2239) );
  assign n2240 = G25 & ~n2239 ;
  assign n2241 = n2238 | n2240 ;
  assign n2242 = n2236 | n2241 ;
  assign n2243 = G158 | n1866 ;
  assign n2244 = G158 & ~n1771 ;
  assign n2245 = G159 & ~n2244 ;
  assign n2246 = n2243 & n2245 ;
  assign n2247 = G76 & ~n2151 ;
  assign n2248 = G86 & n2155 ;
  assign n2249 = n2247 | n2248 ;
  assign n2250 = n2246 | n2249 ;
  assign n2251 = G64 & n2250 ;
  assign n2252 = G158 | n1937 ;
  assign n2253 = G158 & ~n1690 ;
  assign n2254 = G159 & ~n2253 ;
  assign n2255 = n2252 & n2254 ;
  assign n2256 = G72 & ~n2151 ;
  assign n2257 = G82 & n2155 ;
  assign n2258 = n2256 | n2257 ;
  assign n2259 = n2255 | n2258 ;
  assign n2260 = G64 & n2259 ;
  assign n2261 = G158 | n1923 ;
  assign n2262 = G158 & ~n1813 ;
  assign n2263 = G159 & ~n2262 ;
  assign n2264 = n2261 & n2263 ;
  assign n2265 = G70 & ~n2151 ;
  assign n2266 = G71 & n2155 ;
  assign n2267 = n2265 | n2266 ;
  assign n2268 = n2264 | n2267 ;
  assign n2269 = G64 & n2268 ;
  assign n2270 = G158 | n1892 ;
  assign n2271 = G158 & ~n1796 ;
  assign n2272 = G159 & ~n2271 ;
  assign n2273 = n2270 & n2272 ;
  buffer buf_n2274( .i (n2150), .o (n2274) );
  assign n2275 = G68 & ~n2274 ;
  buffer buf_n2276( .i (n2154), .o (n2276) );
  assign n2277 = G69 & n2276 ;
  assign n2278 = n2275 | n2277 ;
  assign n2279 = n2273 | n2278 ;
  assign n2280 = G64 & n2279 ;
  assign n2281 = G160 | n1866 ;
  assign n2282 = G160 & ~n1771 ;
  assign n2283 = G161 & ~n2282 ;
  assign n2284 = n2281 & n2283 ;
  assign n2285 = G76 & ~n2166 ;
  assign n2286 = G86 & n2170 ;
  assign n2287 = n2285 | n2286 ;
  assign n2288 = n2284 | n2287 ;
  assign n2289 = G64 & n2288 ;
  assign n2290 = G160 | n1937 ;
  assign n2291 = G160 & ~n1690 ;
  assign n2292 = G161 & ~n2291 ;
  assign n2293 = n2290 & n2292 ;
  assign n2294 = G72 & ~n2166 ;
  assign n2295 = G82 & n2170 ;
  assign n2296 = n2294 | n2295 ;
  assign n2297 = n2293 | n2296 ;
  assign n2298 = G64 & n2297 ;
  assign n2299 = G160 | n1923 ;
  assign n2300 = G160 & ~n1813 ;
  assign n2301 = G161 & ~n2300 ;
  assign n2302 = n2299 & n2301 ;
  assign n2303 = G70 & ~n2166 ;
  assign n2304 = G71 & n2170 ;
  assign n2305 = n2303 | n2304 ;
  assign n2306 = n2302 | n2305 ;
  assign n2307 = G64 & n2306 ;
  assign n2308 = G160 | n1892 ;
  assign n2309 = G160 & ~n1796 ;
  assign n2310 = G161 & ~n2309 ;
  assign n2311 = n2308 & n2310 ;
  buffer buf_n2312( .i (n2165), .o (n2312) );
  assign n2313 = G68 & ~n2312 ;
  buffer buf_n2314( .i (n2169), .o (n2314) );
  assign n2315 = G69 & n2314 ;
  assign n2316 = n2313 | n2315 ;
  assign n2317 = n2311 | n2316 ;
  assign n2318 = G64 & n2317 ;
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  assign n2319 = G170 & n1721 ;
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  assign n2320 = ~G61 & n1427 ;
  assign n2321 = G61 & ~n1427 ;
  assign n2322 = n2320 | n2321 ;
  buffer buf_n2323( .i (n2322), .o (n2323) );
  assign n2326 = G170 | n2323 ;
  assign n2327 = ~n2319 & n2326 ;
  assign n2328 = G171 & ~n2327 ;
  assign n2329 = G178 & G62 ;
  assign n2330 = G170 & ~G54 ;
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  assign n2331 = G170 | n303 ;
  assign n2332 = ~n2330 & n2331 ;
  assign n2333 = G171 | n2332 ;
  assign n2334 = ~n2329 & n2333 ;
  assign n2335 = ~n2328 & n2334 ;
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2325( .i (n2324), .o (n2325) );
  assign n2336 = n1723 & n2325 ;
  assign n2337 = n1723 | n2325 ;
  assign n2338 = n2336 | ~n2337 ;
  assign n2339 = G54 & n1798 ;
  assign n2340 = ~G176 & n1716 ;
  assign n2341 = G176 & ~n298 ;
  assign n2342 = G177 & ~n2341 ;
  assign n2343 = ~n2340 & n2342 ;
  assign n2344 = n2339 | n2343 ;
  buffer buf_n2345( .i (n2344), .o (n2345) );
  inverter inv_n2996( .i (n2345), .o (n2996) );
  assign n2347 = G52 & n1798 ;
  assign n2348 = G176 | n2120 ;
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  assign n2349 = G176 & ~n317 ;
  assign n2350 = G177 & ~n2349 ;
  assign n2351 = n2348 & n2350 ;
  assign n2352 = n2347 | n2351 ;
  buffer buf_n2353( .i (n2352), .o (n2353) );
  inverter inv_n2997( .i (n2353), .o (n2997) );
  assign n2356 = G47 & n1894 ;
  assign n2357 = G176 | n2103 ;
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  assign n2358 = G176 & n242 ;
  assign n2359 = G177 & ~n2358 ;
  assign n2360 = n2357 & n2359 ;
  assign n2361 = n2356 | n2360 ;
  buffer buf_n2362( .i (n2361), .o (n2362) );
  inverter inv_n2998( .i (n2362), .o (n2998) );
  assign n2366 = G43 & n1894 ;
  assign n2367 = G176 | n2130 ;
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  assign n2368 = G176 & n261 ;
  assign n2369 = G177 & ~n2368 ;
  assign n2370 = n2367 & n2369 ;
  assign n2371 = n2366 | n2370 ;
  buffer buf_n2372( .i (n2371), .o (n2372) );
  inverter inv_n2999( .i (n2372), .o (n2999) );
  assign n2376 = G155 & G99 ;
  assign n2377 = n186 & n2376 ;
  assign n2378 = n180 & n2377 ;
  assign n2379 = ~n1538 & n2378 ;
  assign n2380 = ~n1574 & n2379 ;
  assign n2381 = ~n1987 & n2380 ;
  assign n2382 = ~n2027 & n2381 ;
  buffer buf_n1659( .i (n1658), .o (n1659) );
  assign n2383 = G46 & n1659 ;
  assign n2384 = ~G176 & n2040 ;
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  assign n2385 = G176 & n458 ;
  assign n2386 = G177 & ~n2385 ;
  assign n2387 = ~n2384 & n2386 ;
  assign n2388 = n2383 | n2387 ;
  buffer buf_n2389( .i (n2388), .o (n2389) );
  inverter inv_n3000( .i (n2389), .o (n3000) );
  buffer buf_n2391( .i (n1656), .o (n2391) );
  assign n2392 = G45 & n2391 ;
  assign n2393 = ~G176 & n2066 ;
  assign n2394 = G176 & n394 ;
  assign n2395 = G177 & ~n2394 ;
  assign n2396 = ~n2393 & n2395 ;
  assign n2397 = n2392 | n2396 ;
  buffer buf_n2398( .i (n2397), .o (n2398) );
  inverter inv_n3001( .i (n2398), .o (n3001) );
  assign n2402 = G20 & n2391 ;
  assign n2403 = G176 | n2080 ;
  assign n2404 = G176 & n405 ;
  assign n2405 = G177 & ~n2404 ;
  assign n2406 = n2403 & n2405 ;
  assign n2407 = n2402 | n2406 ;
  buffer buf_n2408( .i (n2407), .o (n2408) );
  inverter inv_n3002( .i (n2408), .o (n3002) );
  assign n2412 = G44 & n2391 ;
  assign n2413 = G176 | n2048 ;
  assign n2414 = G176 & n382 ;
  assign n2415 = G177 & ~n2414 ;
  assign n2416 = n2413 & n2415 ;
  assign n2417 = n2412 | n2416 ;
  buffer buf_n2418( .i (n2417), .o (n2418) );
  inverter inv_n3003( .i (n2418), .o (n3003) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  assign n2422 = G174 | n2390 ;
  buffer buf_n2346( .i (n2345), .o (n2346) );
  assign n2423 = G174 & ~n2346 ;
  assign n2424 = G175 & ~n2423 ;
  assign n2425 = n2422 & n2424 ;
  assign n2426 = G41 & ~n2239 ;
  assign n2427 = G42 & n2237 ;
  assign n2428 = n2426 | n2427 ;
  assign n2429 = n2425 | n2428 ;
  assign n2430 = G173 | n2390 ;
  assign n2431 = G173 & ~n2346 ;
  assign n2432 = G172 & ~n2431 ;
  assign n2433 = n2430 & n2432 ;
  assign n2434 = G41 & ~n2205 ;
  assign n2435 = G42 & n2203 ;
  assign n2436 = n2434 | n2435 ;
  assign n2437 = n2433 | n2436 ;
  buffer buf_n2354( .i (n2353), .o (n2354) );
  buffer buf_n2355( .i (n2354), .o (n2355) );
  assign n2438 = G173 & ~n2355 ;
  buffer buf_n2399( .i (n2398), .o (n2399) );
  buffer buf_n2400( .i (n2399), .o (n2400) );
  assign n2439 = G173 | n2400 ;
  assign n2440 = G172 & n2439 ;
  assign n2441 = ~n2438 & n2440 ;
  assign n2442 = G17 & n2203 ;
  assign n2443 = G18 & ~n2205 ;
  assign n2444 = n2442 | n2443 ;
  assign n2445 = n2441 | n2444 ;
  buffer buf_n2363( .i (n2362), .o (n2363) );
  buffer buf_n2364( .i (n2363), .o (n2364) );
  buffer buf_n2365( .i (n2364), .o (n2365) );
  assign n2446 = G173 & ~n2365 ;
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  assign n2447 = G173 | n2410 ;
  assign n2448 = G172 & n2447 ;
  assign n2449 = ~n2446 & n2448 ;
  assign n2450 = G39 & n2203 ;
  assign n2451 = G40 & ~n2205 ;
  assign n2452 = n2450 | n2451 ;
  assign n2453 = n2449 | n2452 ;
  buffer buf_n2373( .i (n2372), .o (n2373) );
  buffer buf_n2374( .i (n2373), .o (n2374) );
  buffer buf_n2375( .i (n2374), .o (n2375) );
  assign n2454 = G173 & ~n2375 ;
  buffer buf_n2419( .i (n2418), .o (n2419) );
  buffer buf_n2420( .i (n2419), .o (n2420) );
  assign n2455 = G173 | n2420 ;
  assign n2456 = G172 & n2455 ;
  assign n2457 = ~n2454 & n2456 ;
  buffer buf_n2458( .i (n1729), .o (n2458) );
  assign n2459 = G36 & n2458 ;
  buffer buf_n2460( .i (n1733), .o (n2460) );
  assign n2461 = G15 & ~n2460 ;
  assign n2462 = n2459 | n2461 ;
  assign n2463 = n2457 | n2462 ;
  buffer buf_n2401( .i (n2400), .o (n2401) );
  assign n2464 = G174 | n2401 ;
  assign n2465 = G174 & ~n2354 ;
  assign n2466 = G175 & ~n2465 ;
  assign n2467 = n2464 & n2466 ;
  assign n2468 = G17 & n2237 ;
  assign n2469 = G18 & ~n2239 ;
  assign n2470 = n2468 | n2469 ;
  assign n2471 = n2467 | n2470 ;
  buffer buf_n2411( .i (n2410), .o (n2411) );
  assign n2472 = G174 | n2411 ;
  assign n2473 = G174 & ~n2364 ;
  assign n2474 = G175 & ~n2473 ;
  assign n2475 = n2472 & n2474 ;
  assign n2476 = G39 & n2237 ;
  assign n2477 = G40 & ~n2239 ;
  assign n2478 = n2476 | n2477 ;
  assign n2479 = n2475 | n2478 ;
  buffer buf_n2421( .i (n2420), .o (n2421) );
  assign n2480 = G174 | n2421 ;
  assign n2481 = G174 & ~n2374 ;
  assign n2482 = G175 & ~n2481 ;
  assign n2483 = n2480 & n2482 ;
  buffer buf_n2484( .i (n1820), .o (n2484) );
  assign n2485 = G36 & n2484 ;
  buffer buf_n2486( .i (n1824), .o (n2486) );
  assign n2487 = G15 & ~n2486 ;
  assign n2488 = n2485 | n2487 ;
  assign n2489 = n2483 | n2488 ;
  assign n2490 = G158 & ~n2374 ;
  assign n2491 = G158 | n2419 ;
  assign n2492 = G159 & n2491 ;
  assign n2493 = ~n2490 & n2492 ;
  assign n2494 = G77 & ~n2274 ;
  assign n2495 = G87 & n2276 ;
  assign n2496 = n2494 | n2495 ;
  assign n2497 = n2493 | n2496 ;
  assign n2498 = G64 & n2497 ;
  assign n2499 = G158 & ~n2364 ;
  assign n2500 = G158 | n2409 ;
  assign n2501 = G159 & n2500 ;
  assign n2502 = ~n2499 & n2501 ;
  assign n2503 = G75 & ~n2274 ;
  assign n2504 = G85 & n2276 ;
  assign n2505 = n2503 | n2504 ;
  assign n2506 = n2502 | n2505 ;
  assign n2507 = G64 & n2506 ;
  assign n2508 = G158 & ~n2354 ;
  assign n2509 = G158 | n2399 ;
  assign n2510 = G159 & n2509 ;
  assign n2511 = ~n2508 & n2510 ;
  assign n2512 = G84 & n2276 ;
  assign n2513 = G74 & ~n2274 ;
  assign n2514 = n2512 | n2513 ;
  assign n2515 = n2511 | n2514 ;
  assign n2516 = G64 & n2515 ;
  assign n2517 = G158 | n2389 ;
  assign n2518 = G158 & ~n2345 ;
  assign n2519 = G159 & ~n2518 ;
  assign n2520 = n2517 & n2519 ;
  buffer buf_n2521( .i (n2150), .o (n2521) );
  assign n2522 = G73 & ~n2521 ;
  buffer buf_n2523( .i (n2154), .o (n2523) );
  assign n2524 = G83 & n2523 ;
  assign n2525 = n2522 | n2524 ;
  assign n2526 = n2520 | n2525 ;
  assign n2527 = G64 & n2526 ;
  assign n2528 = G160 | n2420 ;
  assign n2529 = G160 & ~n2373 ;
  assign n2530 = G161 & ~n2529 ;
  assign n2531 = n2528 & n2530 ;
  assign n2532 = G77 & ~n2312 ;
  assign n2533 = G87 & n2314 ;
  assign n2534 = n2532 | n2533 ;
  assign n2535 = n2531 | n2534 ;
  assign n2536 = G64 & n2535 ;
  assign n2537 = G160 | n2410 ;
  assign n2538 = G160 & ~n2363 ;
  assign n2539 = G161 & ~n2538 ;
  assign n2540 = n2537 & n2539 ;
  assign n2541 = G85 & n2314 ;
  assign n2542 = G75 & ~n2312 ;
  assign n2543 = n2541 | n2542 ;
  assign n2544 = n2540 | n2543 ;
  assign n2545 = G64 & n2544 ;
  assign n2546 = G160 & ~n2354 ;
  assign n2547 = G160 | n2399 ;
  assign n2548 = G161 & n2547 ;
  assign n2549 = ~n2546 & n2548 ;
  assign n2550 = G74 & ~n2312 ;
  assign n2551 = G84 & n2314 ;
  assign n2552 = n2550 | n2551 ;
  assign n2553 = n2549 | n2552 ;
  assign n2554 = G64 & n2553 ;
  assign n2555 = G160 | n2389 ;
  assign n2556 = G160 & ~n2345 ;
  assign n2557 = G161 & ~n2556 ;
  assign n2558 = n2555 & n2557 ;
  buffer buf_n2559( .i (n2165), .o (n2559) );
  assign n2560 = G73 & ~n2559 ;
  buffer buf_n2561( .i (n2169), .o (n2561) );
  assign n2562 = G83 & n2561 ;
  assign n2563 = n2560 | n2562 ;
  assign n2564 = n2558 | n2563 ;
  assign n2565 = G64 & n2564 ;
  assign n2566 = ~G145 & n1335 ;
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n2568( .i (n2567), .o (n2568) );
  assign n2569 = n1379 & ~n2568 ;
  assign n2570 = G145 & ~n1386 ;
  assign n2571 = n2567 | n2570 ;
  assign n2572 = n1337 & ~n1394 ;
  assign n2573 = n2571 & ~n2572 ;
  assign n2574 = n2569 | n2573 ;
  buffer buf_n2575( .i (n2574), .o (n2575) );
  assign n2576 = n1942 & n2575 ;
  assign n2577 = n1942 | n2575 ;
  assign n2578 = ~n2576 & n2577 ;
  assign n2579 = n2093 & ~n2578 ;
  assign n2580 = ~n1340 & n1379 ;
  assign n2581 = n1347 & ~n2580 ;
  buffer buf_n2582( .i (n2581), .o (n2582) );
  assign n2583 = ~n1388 & n1414 ;
  buffer buf_n2584( .i (n1413), .o (n2584) );
  assign n2585 = n1388 & ~n2584 ;
  assign n2586 = n2583 | n2585 ;
  buffer buf_n2587( .i (n2586), .o (n2587) );
  assign n2588 = n2582 & n2587 ;
  assign n2589 = n2582 | n2587 ;
  assign n2590 = ~n2588 & n2589 ;
  assign n2591 = n2093 | n2590 ;
  assign n2592 = ~n2579 & n2591 ;
  buffer buf_n2593( .i (n2592), .o (n2593) );
  buffer buf_n2594( .i (n2593), .o (n2594) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  assign n2595 = n1144 & ~n1775 ;
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  assign n2596 = ~n1154 & n1775 ;
  assign n2597 = n2595 | n2596 ;
  buffer buf_n2598( .i (n2597), .o (n2598) );
  assign n2599 = G162 & n1213 ;
  assign n2600 = n1194 & n2599 ;
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  assign n2601 = G162 | n1193 ;
  assign n2602 = n1251 & n2601 ;
  assign n2603 = ~n2600 & n2602 ;
  buffer buf_n2604( .i (n2603), .o (n2604) );
  assign n2605 = ~n1156 & n1489 ;
  assign n2606 = n1156 & ~n1489 ;
  assign n2607 = n2605 | n2606 ;
  buffer buf_n2608( .i (n2607), .o (n2608) );
  assign n2609 = n2604 & n2608 ;
  assign n2610 = n2604 | n2608 ;
  assign n2611 = ~n2609 & n2610 ;
  buffer buf_n2612( .i (n2611), .o (n2612) );
  assign n2613 = ~n1304 & n2612 ;
  assign n2614 = n1304 & ~n2612 ;
  assign n2615 = n2613 | n2614 ;
  buffer buf_n2616( .i (n2615), .o (n2616) );
  assign n2617 = n2598 & ~n2616 ;
  assign n2618 = ~n2598 & n2616 ;
  assign n2619 = n2617 | n2618 ;
  buffer buf_n2620( .i (n2619), .o (n2620) );
  buffer buf_n2621( .i (n2620), .o (n2621) );
  assign n2622 = n2594 | n2621 ;
  assign n2623 = n2593 & n2620 ;
  assign n2624 = G176 | n2623 ;
  assign n2625 = n2622 & ~n2624 ;
  assign n2626 = ~G148 & G98 ;
  assign n2627 = ~G100 & G148 ;
  assign n2628 = n2626 | n2627 ;
  buffer buf_n2629( .i (n2628), .o (n2629) );
  assign n2630 = ~n330 & n2629 ;
  assign n2631 = n330 & ~n2629 ;
  assign n2632 = n2630 | n2631 ;
  buffer buf_n2633( .i (n2632), .o (n2633) );
  assign n2634 = G100 | G121 ;
  assign n2635 = ~G101 & G121 ;
  assign n2636 = n2634 & ~n2635 ;
  assign n2637 = G147 & ~n2636 ;
  assign n2638 = G102 & G121 ;
  assign n2639 = ~G121 & G98 ;
  assign n2640 = n2638 | n2639 ;
  assign n2641 = ~G147 & n2640 ;
  assign n2642 = n2637 | n2641 ;
  buffer buf_n2643( .i (n2642), .o (n2643) );
  assign n2644 = n2633 | n2643 ;
  assign n2645 = n2633 & n2643 ;
  assign n2646 = n2644 & ~n2645 ;
  buffer buf_n2647( .i (n2646), .o (n2647) );
  assign n2648 = G100 | G128 ;
  assign n2649 = ~G101 & G128 ;
  assign n2650 = n2648 & ~n2649 ;
  assign n2651 = G150 & ~n2650 ;
  assign n2652 = G102 & G128 ;
  assign n2653 = ~G128 & G98 ;
  assign n2654 = n2652 | n2653 ;
  assign n2655 = ~G150 & n2654 ;
  assign n2656 = n2651 | n2655 ;
  buffer buf_n2657( .i (n2656), .o (n2657) );
  assign n2658 = G100 | G126 ;
  assign n2659 = ~G101 & G126 ;
  assign n2660 = n2658 & ~n2659 ;
  assign n2661 = G149 & ~n2660 ;
  assign n2662 = G102 & G126 ;
  assign n2663 = ~G126 & G98 ;
  assign n2664 = n2662 | n2663 ;
  assign n2665 = ~G149 & n2664 ;
  assign n2666 = n2661 | n2665 ;
  buffer buf_n2667( .i (n2666), .o (n2667) );
  assign n2668 = n2657 | n2667 ;
  assign n2669 = n2657 & n2667 ;
  assign n2670 = n2668 & ~n2669 ;
  buffer buf_n2671( .i (n2670), .o (n2671) );
  assign n2672 = n2647 | n2671 ;
  assign n2673 = n2647 & n2671 ;
  assign n2674 = n2672 & ~n2673 ;
  buffer buf_n2675( .i (n2674), .o (n2675) );
  buffer buf_n2676( .i (n2675), .o (n2676) );
  assign n2677 = n234 | n253 ;
  assign n2678 = ~n263 & n2677 ;
  buffer buf_n2679( .i (n2678), .o (n2679) );
  assign n2680 = ~n289 & n308 ;
  assign n2681 = n319 | n2680 ;
  buffer buf_n2682( .i (n2681), .o (n2682) );
  assign n2683 = n2679 | n2682 ;
  assign n2684 = n2679 & n2682 ;
  assign n2685 = n2683 & ~n2684 ;
  buffer buf_n2686( .i (n2685), .o (n2686) );
  buffer buf_n2687( .i (n2686), .o (n2687) );
  assign n2688 = n2676 | n2687 ;
  assign n2689 = n2675 & n2686 ;
  assign n2690 = G176 & ~n2689 ;
  assign n2691 = n2688 & n2690 ;
  assign n2692 = G177 & ~n2691 ;
  assign n2693 = ~n2625 & n2692 ;
  buffer buf_n2694( .i (n2693), .o (n2694) );
  buffer buf_n2695( .i (n2694), .o (n2695) );
  buffer buf_n2696( .i (n2695), .o (n2696) );
  buffer buf_n2697( .i (n2696), .o (n2697) );
  buffer buf_n2698( .i (n2697), .o (n2698) );
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n2700( .i (n2699), .o (n2700) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  assign n2701 = ~G51 & n1664 ;
  assign n2702 = ~n2700 & ~n2701 ;
  assign n2703 = n579 & n635 ;
  assign n2704 = n576 | n646 ;
  assign n2705 = ~n661 & n2704 ;
  buffer buf_n2706( .i (n2705), .o (n2706) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  assign n2707 = n556 | n633 ;
  assign n2708 = ~n1581 & n2707 ;
  assign n2709 = n2706 | n2708 ;
  assign n2710 = ~n2703 & n2709 ;
  buffer buf_n2711( .i (n2710), .o (n2711) );
  assign n2712 = n1591 & ~n2711 ;
  assign n2713 = ~n1591 & n2711 ;
  assign n2714 = n2712 | n2713 ;
  buffer buf_n2715( .i (n2714), .o (n2715) );
  buffer buf_n2716( .i (n2715), .o (n2716) );
  assign n2717 = n1850 | n2716 ;
  assign n2718 = n1849 & n2715 ;
  assign n2719 = G157 | n2718 ;
  assign n2720 = n2717 & ~n2719 ;
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  assign n2721 = n571 & n625 ;
  assign n2722 = n571 | n635 ;
  assign n2723 = ~n2721 & n2722 ;
  buffer buf_n2724( .i (n2723), .o (n2724) );
  assign n2725 = n1871 & ~n2724 ;
  assign n2726 = ~n1871 & n2724 ;
  assign n2727 = n2725 | n2726 ;
  buffer buf_n2728( .i (n2727), .o (n2728) );
  buffer buf_n2729( .i (n2728), .o (n2729) );
  assign n2730 = n519 | n2706 ;
  assign n2731 = n519 & n2706 ;
  assign n2732 = n2730 & ~n2731 ;
  buffer buf_n2733( .i (n2732), .o (n2733) );
  assign n2734 = n781 | n1843 ;
  buffer buf_n2735( .i (n2734), .o (n2735) );
  assign n2736 = n2733 & ~n2735 ;
  assign n2737 = ~n2733 & n2735 ;
  assign n2738 = n2736 | n2737 ;
  buffer buf_n2739( .i (n2738), .o (n2739) );
  buffer buf_n2740( .i (n2739), .o (n2740) );
  assign n2741 = n2729 & n2740 ;
  assign n2742 = n2728 | n2739 ;
  assign n2743 = G157 & n2742 ;
  assign n2744 = ~n2741 & n2743 ;
  assign n2745 = n2720 | n2744 ;
  buffer buf_n2746( .i (n2745), .o (n2746) );
  buffer buf_n2747( .i (n2746), .o (n2747) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  assign n2748 = n1099 | n1620 ;
  buffer buf_n2749( .i (n2748), .o (n2749) );
  buffer buf_n2750( .i (n2749), .o (n2750) );
  buffer buf_n2751( .i (n2750), .o (n2751) );
  buffer buf_n2752( .i (n2751), .o (n2752) );
  assign n2753 = ~n921 & n2752 ;
  assign n2754 = n940 & ~n2753 ;
  buffer buf_n2755( .i (n2754), .o (n2755) );
  assign n2756 = n867 | n997 ;
  assign n2757 = n867 & n997 ;
  assign n2758 = n2756 & ~n2757 ;
  buffer buf_n2759( .i (n2758), .o (n2759) );
  buffer buf_n2760( .i (n2759), .o (n2760) );
  buffer buf_n2761( .i (n2760), .o (n2761) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  assign n2762 = n1047 | n2749 ;
  assign n2763 = ~n1618 & n2762 ;
  buffer buf_n2764( .i (n2763), .o (n2764) );
  assign n2765 = n2761 & n2764 ;
  assign n2766 = n2761 | n2764 ;
  assign n2767 = ~n2765 & n2766 ;
  buffer buf_n2768( .i (n2767), .o (n2768) );
  assign n2769 = n2755 & n2768 ;
  assign n2770 = n2755 | n2768 ;
  assign n2771 = ~n2769 & n2770 ;
  buffer buf_n2772( .i (n2771), .o (n2772) );
  assign n2773 = n1604 & n2772 ;
  assign n2774 = n919 | n1623 ;
  assign n2775 = ~n1636 & n2774 ;
  buffer buf_n2776( .i (n2775), .o (n2776) );
  buffer buf_n2777( .i (n2776), .o (n2777) );
  assign n2778 = ~n942 & n1064 ;
  assign n2779 = n942 & ~n1064 ;
  assign n2780 = n2778 | n2779 ;
  buffer buf_n2781( .i (n2780), .o (n2781) );
  assign n2782 = n2759 & ~n2781 ;
  assign n2783 = ~n2759 & n2781 ;
  assign n2784 = n2782 | n2783 ;
  buffer buf_n2785( .i (n2784), .o (n2785) );
  buffer buf_n2786( .i (n2785), .o (n2786) );
  assign n2787 = n2777 | n2786 ;
  assign n2788 = n2776 & n2785 ;
  assign n2789 = n1600 | n2788 ;
  assign n2790 = n2787 & ~n2789 ;
  buffer buf_n2791( .i (n2790), .o (n2791) );
  buffer buf_n2792( .i (n2791), .o (n2792) );
  assign n2793 = G157 | n2792 ;
  assign n2794 = n2773 | n2793 ;
  assign n2795 = n793 | n1603 ;
  assign n2796 = n2772 & n2795 ;
  assign n2797 = ~n793 & n2791 ;
  assign n2798 = G157 & ~n2797 ;
  assign n2799 = ~n2796 & n2798 ;
  assign n2800 = n2794 & ~n2799 ;
  buffer buf_n2801( .i (n2800), .o (n2801) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  assign n2802 = n706 | n762 ;
  assign n2803 = ~n777 & n2802 ;
  buffer buf_n2804( .i (n2803), .o (n2804) );
  assign n2805 = n2801 & ~n2804 ;
  assign n2806 = ~n2801 & n2804 ;
  assign n2807 = n2805 | n2806 ;
  buffer buf_n2808( .i (n2807), .o (n2808) );
  buffer buf_n2809( .i (n2808), .o (n2809) );
  assign n2810 = ~n2747 & n2809 ;
  assign n2811 = n2746 & ~n2808 ;
  assign n2812 = G176 | n2811 ;
  assign n2813 = n2810 | n2812 ;
  assign n2814 = G100 | G90 ;
  assign n2815 = ~G101 & G90 ;
  assign n2816 = n2814 & ~n2815 ;
  assign n2817 = G143 & ~n2816 ;
  assign n2818 = G102 & G90 ;
  assign n2819 = ~G90 & G98 ;
  assign n2820 = n2818 | n2819 ;
  assign n2821 = ~G143 & n2820 ;
  assign n2822 = n2817 | n2821 ;
  buffer buf_n2823( .i (n2822), .o (n2823) );
  assign n2824 = G100 | G92 ;
  assign n2825 = ~G101 & G92 ;
  assign n2826 = n2824 & ~n2825 ;
  assign n2827 = G144 & ~n2826 ;
  assign n2828 = G102 & G92 ;
  assign n2829 = ~G92 & G98 ;
  assign n2830 = n2828 | n2829 ;
  assign n2831 = ~G144 & n2830 ;
  assign n2832 = n2827 | n2831 ;
  buffer buf_n2833( .i (n2832), .o (n2833) );
  assign n2834 = n2823 & ~n2833 ;
  assign n2835 = ~n2823 & n2833 ;
  assign n2836 = n2834 | n2835 ;
  buffer buf_n2837( .i (n2836), .o (n2837) );
  assign n2838 = G100 | G94 ;
  assign n2839 = ~G101 & G94 ;
  assign n2840 = n2838 & ~n2839 ;
  assign n2841 = G140 & ~n2840 ;
  assign n2842 = G102 & G94 ;
  assign n2843 = ~G94 & G98 ;
  assign n2844 = n2842 | n2843 ;
  assign n2845 = ~G140 & n2844 ;
  assign n2846 = n2841 | n2845 ;
  buffer buf_n2847( .i (n2846), .o (n2847) );
  assign n2848 = n449 & n2847 ;
  assign n2849 = n449 | n2847 ;
  assign n2850 = ~n2848 & n2849 ;
  buffer buf_n2851( .i (n2850), .o (n2851) );
  assign n2852 = ~n2837 & n2851 ;
  assign n2853 = n2837 & ~n2851 ;
  assign n2854 = n2852 | n2853 ;
  buffer buf_n2855( .i (n2854), .o (n2855) );
  buffer buf_n2856( .i (n2855), .o (n2856) );
  assign n2857 = G100 | G107 ;
  assign n2858 = ~G101 & G107 ;
  assign n2859 = n2857 & ~n2858 ;
  assign n2860 = G139 & ~n2859 ;
  assign n2861 = G102 & G107 ;
  assign n2862 = ~G107 & G98 ;
  assign n2863 = n2861 | n2862 ;
  assign n2864 = ~G139 & n2863 ;
  assign n2865 = n2860 | n2864 ;
  buffer buf_n2866( .i (n2865), .o (n2866) );
  assign n2867 = G100 | G105 ;
  assign n2868 = ~G101 & G105 ;
  assign n2869 = n2867 & ~n2868 ;
  assign n2870 = G138 & ~n2869 ;
  assign n2871 = G102 & G105 ;
  assign n2872 = ~G105 & G98 ;
  assign n2873 = n2871 | n2872 ;
  assign n2874 = ~G138 & n2873 ;
  assign n2875 = n2870 | n2874 ;
  buffer buf_n2876( .i (n2875), .o (n2876) );
  assign n2877 = n2866 & n2876 ;
  assign n2878 = n2866 | n2876 ;
  assign n2879 = ~n2877 & n2878 ;
  buffer buf_n2880( .i (n2879), .o (n2880) );
  assign n2881 = G100 | G96 ;
  assign n2882 = ~G101 & G96 ;
  assign n2883 = n2881 & ~n2882 ;
  assign n2884 = G141 & ~n2883 ;
  assign n2885 = G102 & G96 ;
  assign n2886 = ~G96 & G98 ;
  assign n2887 = n2885 | n2886 ;
  assign n2888 = ~G141 & n2887 ;
  assign n2889 = n2884 | n2888 ;
  buffer buf_n2890( .i (n2889), .o (n2890) );
  assign n2891 = G100 | G109 ;
  assign n2892 = ~G101 & G109 ;
  assign n2893 = n2891 & ~n2892 ;
  assign n2894 = G135 & ~n2893 ;
  assign n2895 = G102 & G109 ;
  assign n2896 = ~G109 & G98 ;
  assign n2897 = n2895 | n2896 ;
  assign n2898 = ~G135 & n2897 ;
  assign n2899 = n2894 | n2898 ;
  buffer buf_n2900( .i (n2899), .o (n2900) );
  assign n2901 = G100 | G103 ;
  assign n2902 = ~G101 & G103 ;
  assign n2903 = n2901 & ~n2902 ;
  assign n2904 = G137 & ~n2903 ;
  assign n2905 = G102 & G103 ;
  assign n2906 = ~G103 & G98 ;
  assign n2907 = n2905 | n2906 ;
  assign n2908 = ~G137 & n2907 ;
  assign n2909 = n2904 | n2908 ;
  buffer buf_n2910( .i (n2909), .o (n2910) );
  assign n2911 = n2900 & n2910 ;
  assign n2912 = n2900 | n2910 ;
  assign n2913 = ~n2911 & n2912 ;
  buffer buf_n2914( .i (n2913), .o (n2914) );
  assign n2915 = n2890 & ~n2914 ;
  assign n2916 = ~n2890 & n2914 ;
  assign n2917 = n2915 | n2916 ;
  buffer buf_n2918( .i (n2917), .o (n2918) );
  assign n2919 = ~n2880 & n2918 ;
  assign n2920 = n2880 & ~n2918 ;
  assign n2921 = n2919 | n2920 ;
  buffer buf_n2922( .i (n2921), .o (n2922) );
  buffer buf_n2923( .i (n2922), .o (n2923) );
  assign n2924 = ~n2856 & n2923 ;
  assign n2925 = n2855 & ~n2922 ;
  assign n2926 = G176 & ~n2925 ;
  assign n2927 = ~n2924 & n2926 ;
  assign n2928 = G177 & ~n2927 ;
  assign n2929 = n2813 & n2928 ;
  buffer buf_n2930( .i (n2929), .o (n2930) );
  buffer buf_n2931( .i (n2930), .o (n2931) );
  buffer buf_n2932( .i (n2931), .o (n2932) );
  buffer buf_n2933( .i (n2932), .o (n2933) );
  buffer buf_n2934( .i (n2933), .o (n2934) );
  buffer buf_n2935( .i (n2934), .o (n2935) );
  assign n2936 = ~G49 & n1664 ;
  assign n2937 = ~n2935 & ~n2936 ;
  assign n2938 = ~G177 & G38 ;
  assign n2939 = n2930 | n2938 ;
  buffer buf_n2940( .i (n2939), .o (n2940) );
  buffer buf_n2941( .i (n2940), .o (n2941) );
  assign n2942 = G173 | n2941 ;
  assign n2943 = ~G177 & G37 ;
  assign n2944 = n2694 | n2943 ;
  buffer buf_n2945( .i (n2944), .o (n2945) );
  buffer buf_n2946( .i (n2945), .o (n2946) );
  assign n2947 = G173 & ~n2946 ;
  assign n2948 = G172 & ~n2947 ;
  assign n2949 = n2942 & n2948 ;
  assign n2950 = G23 & ~n2460 ;
  assign n2951 = G4 & n2458 ;
  assign n2952 = n2950 | n2951 ;
  assign n2953 = n2949 | n2952 ;
  assign n2954 = G174 | n2941 ;
  assign n2955 = G174 & ~n2946 ;
  assign n2956 = G175 & ~n2955 ;
  assign n2957 = n2954 & n2956 ;
  assign n2958 = G23 & ~n2486 ;
  assign n2959 = G4 & n2484 ;
  assign n2960 = n2958 | n2959 ;
  assign n2961 = n2957 | n2960 ;
  assign n2962 = G158 | n2940 ;
  assign n2963 = G158 & ~n2945 ;
  assign n2964 = G159 & ~n2963 ;
  assign n2965 = n2962 & n2964 ;
  assign n2966 = G79 & ~n2521 ;
  assign n2967 = G78 & n2523 ;
  assign n2968 = n2966 | n2967 ;
  assign n2969 = n2965 | n2968 ;
  assign n2970 = ~G64 | ~n2969 ;
  assign n2971 = G160 | n2940 ;
  assign n2972 = G160 & ~n2945 ;
  assign n2973 = G161 & ~n2972 ;
  assign n2974 = n2971 & n2973 ;
  assign n2975 = G79 & ~n2559 ;
  assign n2976 = G78 & n2561 ;
  assign n2977 = n2975 | n2976 ;
  assign n2978 = n2974 | n2977 ;
  assign n2979 = ~G64 | ~n2978 ;
  assign G5193 = ~G66 ;
  assign G5194 = ~G113 ;
  assign G5195 = ~G165 ;
  assign G5196 = ~G151 ;
  assign G5197 = ~G127 ;
  assign G5198 = ~G131 ;
  assign G5199 = n180 ;
  assign G5200 = ~G152 ;
  assign G5201 = ~G151 ;
  assign G5202 = ~G151 ;
  assign G5203 = ~G125 ;
  assign G5204 = ~G129 ;
  assign G5205 = n181 ;
  assign G5206 = ~G99 ;
  assign G5207 = ~G153 ;
  assign G5208 = ~G156 ;
  assign G5209 = ~G155 ;
  assign G5210 = n182 ;
  assign G5211 = n183 ;
  assign G5212 = n184 ;
  assign G5213 = n2980 ;
  assign G5214 = G64 ;
  assign G5215 = G66 ;
  assign G5216 = G1 ;
  assign G5217 = G152 ;
  assign G5218 = G114 ;
  assign G5219 = G152 ;
  assign G5220 = n192 ;
  assign G5221 = n2981 ;
  assign G5222 = ~G1 ;
  assign G5223 = ~G1 ;
  assign G5224 = ~G1 ;
  assign G5225 = ~G1 ;
  assign G5226 = ~G114 ;
  assign G5227 = ~G114 ;
  assign G5228 = n196 ;
  assign G5229 = n201 ;
  assign G5230 = n201 ;
  assign G5231 = n202 ;
  assign G5232 = n207 ;
  assign G5233 = n212 ;
  assign G5234 = n217 ;
  assign G5235 = n223 ;
  assign G5236 = n372 ;
  assign G5237 = n483 ;
  assign G5238 = n1118 ;
  assign G5239 = n1506 ;
  assign G5240 = n1506 ;
  assign G5241 = n1118 ;
  assign G5242 = n2982 ;
  assign G5243 = n2983 ;
  assign G5244 = n1652 ;
  assign G5245 = n1654 ;
  assign G5246 = n1652 ;
  assign G5247 = n1654 ;
  assign G5248 = n2984 ;
  assign G5249 = n2985 ;
  assign G5250 = n2986 ;
  assign G5251 = n1716 ;
  assign G5252 = n1737 ;
  assign G5253 = n2987 ;
  assign G5254 = n2988 ;
  assign G5255 = n2989 ;
  assign G5256 = n1828 ;
  assign G5257 = n2990 ;
  assign G5258 = n2991 ;
  assign G5259 = n2992 ;
  assign G5260 = n2993 ;
  assign G5261 = n2994 ;
  assign G5262 = n2995 ;
  assign G5263 = n2088 ;
  assign G5264 = n2144 ;
  assign G5265 = n2159 ;
  assign G5266 = n2174 ;
  assign G5267 = n2182 ;
  assign G5268 = n2190 ;
  assign G5269 = n2198 ;
  assign G5270 = n2208 ;
  assign G5271 = n2216 ;
  assign G5272 = n2224 ;
  assign G5273 = n2232 ;
  assign G5274 = n2242 ;
  assign G5275 = n2251 ;
  assign G5276 = n2260 ;
  assign G5277 = n2269 ;
  assign G5278 = n2280 ;
  assign G5279 = n2289 ;
  assign G5280 = n2298 ;
  assign G5281 = n2307 ;
  assign G5282 = n2318 ;
  assign G5283 = n2335 ;
  assign G5284 = n2338 ;
  assign G5285 = n2996 ;
  assign G5286 = n2997 ;
  assign G5287 = n2998 ;
  assign G5288 = n2999 ;
  assign G5289 = n2382 ;
  assign G5290 = n3000 ;
  assign G5291 = n3001 ;
  assign G5292 = n3002 ;
  assign G5293 = n3003 ;
  assign G5294 = n2429 ;
  assign G5295 = n2437 ;
  assign G5296 = n2445 ;
  assign G5297 = n2453 ;
  assign G5298 = n2463 ;
  assign G5299 = n2471 ;
  assign G5300 = n2479 ;
  assign G5301 = n2489 ;
  assign G5302 = n2498 ;
  assign G5303 = n2507 ;
  assign G5304 = n2516 ;
  assign G5305 = n2527 ;
  assign G5306 = n2536 ;
  assign G5307 = n2545 ;
  assign G5308 = n2554 ;
  assign G5309 = n2565 ;
  assign G5310 = n2702 ;
  assign G5311 = n2937 ;
  assign G5312 = n2953 ;
  assign G5313 = n2961 ;
  assign G5314 = n2970 ;
  assign G5315 = n2979 ;
endmodule
