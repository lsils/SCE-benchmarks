module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G6 , G7 , G8 , G9 , G3519 , G3520 , G3521 , G3522 , G3523 , G3524 , G3525 , G3526 , G3527 , G3528 , G3529 , G3530 , G3531 , G3532 , G3533 , G3534 , G3535 , G3536 , G3537 , G3538 , G3539 , G3540 );
  input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G6 , G7 , G8 , G9 ;
  output G3519 , G3520 , G3521 , G3522 , G3523 , G3524 , G3525 , G3526 , G3527 , G3528 , G3529 , G3530 , G3531 , G3532 , G3533 , G3534 , G3535 , G3536 , G3537 , G3538 , G3539 , G3540 ;
  wire n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 ;
  buffer buf_n440( .i (G8), .o (n440) );
  buffer buf_n452( .i (G9), .o (n452) );
  assign n465 = n440 | n452 ;
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n79( .i (G10), .o (n79) );
  buffer buf_n427( .i (G7), .o (n427) );
  assign n467 = n79 | n427 ;
  buffer buf_n468( .i (n467), .o (n468) );
  assign n471 = ~n466 & ~n468 ;
  buffer buf_n91( .i (G11), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n103( .i (G12), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n115( .i (G13), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  assign n472 = n104 | n116 ;
  buffer buf_n473( .i (n472), .o (n473) );
  assign n474 = ~n94 | ~n473 ;
  buffer buf_n51( .i (G1), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n243( .i (G3), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  assign n475 = n54 | n246 ;
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n263( .i (G32), .o (n263) );
  assign n477 = n263 & ~n452 ;
  buffer buf_n258( .i (G31), .o (n258) );
  assign n478 = n258 & ~n440 ;
  assign n479 = n477 | n478 ;
  buffer buf_n284( .i (G36), .o (n284) );
  assign n480 = ~n115 & n284 ;
  buffer buf_n128( .i (G14), .o (n128) );
  buffer buf_n289( .i (G37), .o (n289) );
  assign n481 = ~n128 & n289 ;
  assign n482 = n480 | n481 ;
  assign n483 = n479 | n482 ;
  buffer buf_n273( .i (G34), .o (n273) );
  assign n484 = ~n91 & n273 ;
  buffer buf_n279( .i (G35), .o (n279) );
  assign n485 = ~n103 & n279 ;
  assign n486 = n484 | n485 ;
  buffer buf_n268( .i (G33), .o (n268) );
  assign n487 = ~n79 & n268 ;
  buffer buf_n253( .i (G30), .o (n253) );
  assign n488 = n253 & ~n427 ;
  assign n489 = n487 | n488 ;
  assign n490 = n486 | n489 ;
  assign n491 = n483 | n490 ;
  assign n492 = n476 & n491 ;
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n154( .i (G2), .o (n154) );
  assign n496 = ~n52 & n154 ;
  buffer buf_n497( .i (n496), .o (n497) );
  assign n500 = ~n246 & n497 ;
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  assign n502 = ~n429 & n466 ;
  buffer buf_n503( .i (n502), .o (n503) );
  assign n508 = n501 & n503 ;
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  assign n511 = n158 | n476 ;
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  assign n513 = n283 | n288 ;
  assign n514 = n278 & n513 ;
  assign n515 = ~n512 & n514 ;
  assign n516 = n510 | n515 ;
  assign n517 = ~n495 & ~n516 ;
  assign n518 = n284 | n289 ;
  assign n519 = n284 & n289 ;
  assign n520 = n518 & ~n519 ;
  buffer buf_n521( .i (n520), .o (n521) );
  assign n522 = n273 & ~n279 ;
  assign n523 = ~n273 & n279 ;
  assign n524 = n522 | n523 ;
  buffer buf_n525( .i (n524), .o (n525) );
  assign n526 = n521 | n525 ;
  assign n527 = n521 & n525 ;
  assign n528 = n526 & ~n527 ;
  buffer buf_n529( .i (n528), .o (n529) );
  assign n530 = n253 & ~n258 ;
  assign n531 = ~n253 & n258 ;
  assign n532 = n530 | n531 ;
  buffer buf_n533( .i (n532), .o (n533) );
  assign n534 = n263 | n268 ;
  assign n535 = n263 & n268 ;
  assign n536 = n534 & ~n535 ;
  buffer buf_n537( .i (n536), .o (n537) );
  assign n538 = n533 | n537 ;
  assign n539 = n533 & n537 ;
  assign n540 = n538 & ~n539 ;
  buffer buf_n541( .i (n540), .o (n541) );
  assign n542 = n529 | n541 ;
  assign n543 = n529 & n541 ;
  assign n544 = n542 & ~n543 ;
  assign n545 = n440 & n452 ;
  buffer buf_n546( .i (n545), .o (n546) );
  assign n547 = n466 & ~n546 ;
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n80( .i (n79), .o (n80) );
  assign n549 = n80 & n428 ;
  assign n550 = n468 & ~n549 ;
  buffer buf_n551( .i (n550), .o (n551) );
  assign n552 = ~n548 & n551 ;
  assign n553 = n548 & ~n551 ;
  assign n554 = n552 | n553 ;
  buffer buf_n555( .i (n554), .o (n555) );
  assign n556 = ~n91 & n115 ;
  assign n557 = n91 & ~n115 ;
  assign n558 = n556 | n557 ;
  buffer buf_n559( .i (n558), .o (n559) );
  assign n560 = n103 | n128 ;
  assign n561 = n103 & n128 ;
  assign n562 = n560 & ~n561 ;
  buffer buf_n563( .i (n562), .o (n563) );
  assign n564 = n559 & ~n563 ;
  assign n565 = ~n559 & n563 ;
  assign n566 = n564 | n565 ;
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  assign n569 = n555 & n568 ;
  assign n570 = n555 | n568 ;
  assign n571 = ~n569 & n570 ;
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  assign n572 = n246 & n497 ;
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  assign n578 = n435 | n577 ;
  assign n579 = ~n53 & n245 ;
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  assign n584 = n52 & n154 ;
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n310( .i (G4), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  assign n588 = n53 & n245 ;
  assign n589 = n313 & n588 ;
  assign n590 = n586 | n589 ;
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  assign n594 = n583 | n592 ;
  buffer buf_n595( .i (n594), .o (n595) );
  assign n596 = n435 & n595 ;
  assign n597 = n578 & ~n596 ;
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n247( .i (n246), .o (n247) );
  assign n598 = n429 | n466 ;
  assign n599 = n247 & n598 ;
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n163( .i (G21), .o (n163) );
  buffer buf_n602( .i (n245), .o (n602) );
  assign n603 = n313 | n602 ;
  buffer buf_n604( .i (n603), .o (n604) );
  assign n605 = n163 & ~n604 ;
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n606( .i (n244), .o (n606) );
  assign n607 = n312 & ~n606 ;
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  assign n610 = ~n444 & n609 ;
  assign n611 = n605 | n610 ;
  assign n612 = n601 | n611 ;
  assign n613 = n593 & n612 ;
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  assign n616 = n597 | n615 ;
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n190( .i (G25), .o (n190) );
  buffer buf_n192( .i (G26), .o (n192) );
  assign n619 = n190 | n192 ;
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n403( .i (G5), .o (n403) );
  buffer buf_n418( .i (G6), .o (n418) );
  assign n631 = n403 | n418 ;
  assign n632 = ~n53 & n631 ;
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n294( .i (G38), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  assign n639 = n313 & n405 ;
  buffer buf_n640( .i (n639), .o (n640) );
  assign n644 = n587 & ~n640 ;
  buffer buf_n645( .i (n644), .o (n645) );
  assign n647 = n298 & ~n645 ;
  buffer buf_n648( .i (n647), .o (n648) );
  assign n649 = n638 & n648 ;
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  assign n651 = n257 & ~n634 ;
  assign n652 = G49 | n312 ;
  buffer buf_n653( .i (n652), .o (n653) );
  assign n655 = G28 & ~n653 ;
  assign n656 = n80 & ~n312 ;
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n240( .i (G29), .o (n240) );
  buffer buf_n658( .i (n311), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  assign n660 = n240 & n659 ;
  assign n661 = n657 | n660 ;
  assign n662 = n655 | n661 ;
  assign n663 = n651 | n662 ;
  assign n664 = ~n645 & n663 ;
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  assign n668 = n650 | n667 ;
  buffer buf_n669( .i (n668), .o (n669) );
  assign n670 = n630 & ~n669 ;
  assign n671 = n618 | n670 ;
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n180( .i (G23), .o (n180) );
  buffer buf_n181( .i (G24), .o (n181) );
  assign n673 = n180 | n181 ;
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  assign n684 = ~n669 & n683 ;
  assign n685 = n618 & n684 ;
  buffer buf_n686( .i (n685), .o (n686) );
  assign n688 = n672 & ~n686 ;
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  assign n690 = n448 & n595 ;
  assign n691 = n448 | n577 ;
  assign n692 = ~n690 & n691 ;
  buffer buf_n248( .i (n247), .o (n248) );
  assign n693 = n248 & n548 ;
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  assign n694 = ~n455 & n608 ;
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n171( .i (G22), .o (n171) );
  assign n695 = n171 & ~n606 ;
  buffer buf_n696( .i (n695), .o (n696) );
  assign n704 = ~n314 & n696 ;
  assign n705 = n694 | n704 ;
  assign n706 = n693 | n705 ;
  assign n707 = n592 & n706 ;
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  assign n711 = n692 | n710 ;
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  assign n714 = n262 & ~n634 ;
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n654( .i (n653), .o (n654) );
  assign n716 = n242 & ~n654 ;
  assign n717 = n92 | n658 ;
  buffer buf_n718( .i (n717), .o (n718) );
  assign n719 = ~n255 & n659 ;
  assign n720 = n718 & ~n719 ;
  buffer buf_n721( .i (n720), .o (n721) );
  assign n722 = n716 | n721 ;
  assign n723 = n715 | n722 ;
  assign n724 = ~n646 & n723 ;
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  assign n727 = n650 | n726 ;
  buffer buf_n728( .i (n727), .o (n728) );
  assign n729 = n630 & ~n728 ;
  assign n730 = n713 | n729 ;
  buffer buf_n731( .i (n730), .o (n731) );
  assign n732 = n683 & ~n728 ;
  assign n733 = n713 & n732 ;
  buffer buf_n734( .i (n733), .o (n734) );
  assign n735 = n731 & ~n734 ;
  buffer buf_n736( .i (n735), .o (n736) );
  assign n737 = n689 & n736 ;
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  assign n739 = n250 & n592 ;
  buffer buf_n740( .i (n739), .o (n740) );
  assign n741 = n595 & ~n740 ;
  assign n742 = n88 & ~n741 ;
  assign n743 = ~n85 & n575 ;
  assign n744 = n444 | n604 ;
  buffer buf_n95( .i (n94), .o (n95) );
  assign n745 = ~n95 & n609 ;
  assign n746 = n744 & ~n745 ;
  buffer buf_n747( .i (n591), .o (n747) );
  assign n748 = ~n746 & n747 ;
  assign n749 = n743 | n748 ;
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  assign n752 = n742 | n751 ;
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  assign n755 = n272 & ~n634 ;
  buffer buf_n756( .i (n755), .o (n756) );
  assign n757 = n262 & ~n654 ;
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  assign n758 = n118 | n314 ;
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  assign n759 = ~n266 & n314 ;
  assign n760 = n758 & ~n759 ;
  assign n761 = n757 | n760 ;
  assign n762 = n756 | n761 ;
  assign n763 = ~n646 & n762 ;
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  assign n766 = n650 | n765 ;
  buffer buf_n767( .i (n766), .o (n767) );
  assign n768 = n630 & ~n767 ;
  assign n769 = n754 | n768 ;
  buffer buf_n770( .i (n769), .o (n770) );
  assign n771 = n683 & ~n767 ;
  assign n772 = n754 & n771 ;
  buffer buf_n773( .i (n772), .o (n773) );
  assign n774 = n770 & ~n773 ;
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  assign n786 = n577 | n740 ;
  buffer buf_n787( .i (n786), .o (n787) );
  assign n788 = ~n462 & n787 ;
  assign n789 = n431 & ~n604 ;
  assign n790 = n83 & n609 ;
  assign n791 = n789 | n790 ;
  assign n792 = n747 & n791 ;
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  assign n795 = n460 & ~n595 ;
  assign n796 = n794 | n795 ;
  buffer buf_n797( .i (n796), .o (n797) );
  assign n798 = n788 | n797 ;
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n800( .i (n633), .o (n800) );
  assign n801 = n267 & ~n800 ;
  buffer buf_n802( .i (n801), .o (n802) );
  assign n803 = n257 & ~n654 ;
  assign n804 = n104 | n658 ;
  buffer buf_n805( .i (n804), .o (n805) );
  assign n806 = ~n260 & n659 ;
  assign n807 = n805 & ~n806 ;
  buffer buf_n808( .i (n807), .o (n808) );
  assign n809 = n803 | n808 ;
  assign n810 = n802 | n809 ;
  assign n811 = ~n646 & n810 ;
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  assign n814 = n650 | n813 ;
  buffer buf_n815( .i (n814), .o (n815) );
  assign n816 = n630 & ~n815 ;
  assign n817 = n799 | n816 ;
  buffer buf_n818( .i (n817), .o (n818) );
  assign n819 = n683 & ~n815 ;
  assign n820 = n799 & n819 ;
  buffer buf_n821( .i (n820), .o (n821) );
  assign n823 = n818 & ~n821 ;
  buffer buf_n824( .i (n823), .o (n824) );
  assign n825 = n775 & n824 ;
  buffer buf_n826( .i (n825), .o (n826) );
  assign n827 = n738 & n826 ;
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  assign n835 = n94 | n473 ;
  assign n836 = n248 & n835 ;
  buffer buf_n837( .i (n836), .o (n837) );
  assign n838 = n456 | n604 ;
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  assign n839 = ~n107 & n609 ;
  assign n840 = n838 & ~n839 ;
  assign n841 = ~n837 & n840 ;
  assign n842 = n593 & ~n841 ;
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n315( .i (n314), .o (n315) );
  assign n845 = ~n56 & n315 ;
  assign n846 = n574 | n845 ;
  assign n847 = n747 | n846 ;
  buffer buf_n848( .i (n847), .o (n848) );
  assign n849 = n99 & ~n848 ;
  assign n850 = ~n99 & n577 ;
  assign n851 = n849 | n850 ;
  assign n852 = n844 | n851 ;
  buffer buf_n853( .i (n852), .o (n853) );
  assign n854 = n267 & ~n654 ;
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n855( .i (n659), .o (n855) );
  assign n856 = n131 | n855 ;
  assign n857 = ~n271 & n855 ;
  assign n858 = n856 & ~n857 ;
  assign n859 = n854 | n858 ;
  assign n860 = n52 | n418 ;
  buffer buf_n861( .i (n860), .o (n861) );
  assign n863 = n294 | n861 ;
  assign n864 = ~n275 & n861 ;
  assign n865 = n863 & ~n864 ;
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  assign n868 = n859 | n867 ;
  assign n869 = ~n646 & n868 ;
  buffer buf_n870( .i (n869), .o (n870) );
  assign n871 = n680 & ~n870 ;
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  assign n874 = n853 & n873 ;
  buffer buf_n875( .i (n874), .o (n875) );
  assign n878 = n627 & ~n870 ;
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  assign n881 = n853 | n880 ;
  buffer buf_n882( .i (n881), .o (n882) );
  assign n884 = ~n875 & n882 ;
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n887( .i (n576), .o (n887) );
  assign n888 = n111 | n887 ;
  assign n889 = n111 & n848 ;
  assign n890 = n888 & ~n889 ;
  assign n891 = n105 & n117 ;
  assign n892 = n473 & ~n891 ;
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  assign n897 = n740 & n896 ;
  assign n898 = n585 & ~n602 ;
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n658), .o (n900) );
  assign n901 = n117 & n900 ;
  assign n902 = n657 | n901 ;
  assign n903 = n899 & n902 ;
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  assign n908 = n897 | n907 ;
  assign n909 = n890 | n908 ;
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  assign n912 = n405 | n861 ;
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  assign n918 = n648 & ~n917 ;
  buffer buf_n919( .i (n918), .o (n919) );
  assign n920 = n283 & n913 ;
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n653), .o (n922) );
  assign n923 = n272 & ~n922 ;
  buffer buf_n299( .i (G39), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  assign n924 = n300 | n855 ;
  assign n925 = ~n276 & n855 ;
  assign n926 = n924 & ~n925 ;
  assign n927 = n923 | n926 ;
  assign n928 = n921 | n927 ;
  buffer buf_n929( .i (n645), .o (n929) );
  assign n930 = n928 & ~n929 ;
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  assign n933 = n919 | n932 ;
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n682), .o (n935) );
  assign n936 = ~n934 & n935 ;
  assign n937 = n911 & n936 ;
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n629), .o (n939) );
  assign n940 = ~n934 & n939 ;
  assign n941 = n911 | n940 ;
  buffer buf_n942( .i (n941), .o (n942) );
  assign n943 = ~n938 & n942 ;
  buffer buf_n944( .i (n943), .o (n944) );
  assign n945 = n886 & n944 ;
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  assign n947 = ~n125 & n787 ;
  assign n948 = n123 & ~n848 ;
  assign n949 = n130 & n900 ;
  assign n950 = n718 & ~n949 ;
  assign n951 = n899 & ~n950 ;
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  assign n956 = n948 | n955 ;
  buffer buf_n957( .i (n956), .o (n957) );
  assign n958 = n947 | n957 ;
  buffer buf_n959( .i (n958), .o (n959) );
  assign n960 = n288 & n913 ;
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n900), .o (n962) );
  assign n963 = n282 & n962 ;
  buffer buf_n325( .i (G40), .o (n325) );
  assign n964 = n325 & ~n962 ;
  assign n965 = n963 | n964 ;
  assign n966 = n277 & ~n922 ;
  assign n967 = n965 | n966 ;
  assign n968 = n961 | n967 ;
  assign n969 = ~n929 & n968 ;
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  assign n972 = n919 | n971 ;
  buffer buf_n973( .i (n972), .o (n973) );
  assign n974 = n935 & ~n973 ;
  assign n975 = n959 & n974 ;
  buffer buf_n976( .i (n975), .o (n976) );
  assign n981 = n939 & ~n973 ;
  assign n982 = n959 | n981 ;
  buffer buf_n983( .i (n982), .o (n983) );
  assign n984 = ~n976 & n983 ;
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  assign n988 = n946 & n987 ;
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  assign n990 = ~n740 & n848 ;
  assign n991 = n137 & ~n990 ;
  assign n992 = ~n133 & n574 ;
  assign n993 = n299 & n900 ;
  assign n994 = n805 & ~n993 ;
  assign n995 = n899 & ~n994 ;
  buffer buf_n996( .i (n995), .o (n996) );
  assign n997 = n992 | n996 ;
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  assign n1001 = n991 | n1000 ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  assign n1004 = n293 & n913 ;
  buffer buf_n1005( .i (n1004), .o (n1005) );
  assign n1006 = n287 & n962 ;
  buffer buf_n333( .i (G41), .o (n333) );
  assign n1007 = n333 & ~n962 ;
  assign n1008 = n1006 | n1007 ;
  assign n1009 = n283 & ~n922 ;
  assign n1010 = n1008 | n1009 ;
  assign n1011 = n1005 | n1010 ;
  assign n1012 = ~n929 & n1011 ;
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  assign n1015 = n919 | n1014 ;
  buffer buf_n1016( .i (n1015), .o (n1016) );
  assign n1017 = n935 & ~n1016 ;
  assign n1018 = n1003 & n1017 ;
  buffer buf_n1019( .i (n1018), .o (n1019) );
  assign n1026 = n939 & ~n1016 ;
  assign n1027 = n1003 | n1026 ;
  buffer buf_n1028( .i (n1027), .o (n1028) );
  assign n1029 = ~n1019 & n1028 ;
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  assign n1035 = n989 & n1034 ;
  buffer buf_n1036( .i (n1035), .o (n1036) );
  assign n1037 = n830 & n1036 ;
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  assign n1038 = n989 & n1025 ;
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  assign n1039 = n946 & n980 ;
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n883( .i (n882), .o (n883) );
  assign n1040 = n883 & n938 ;
  assign n1041 = n877 | n1040 ;
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  assign n1045 = n1039 | n1044 ;
  buffer buf_n1046( .i (n1045), .o (n1046) );
  assign n1047 = n1038 | n1046 ;
  buffer buf_n1048( .i (n1047), .o (n1048) );
  assign n1049 = n831 & n1048 ;
  buffer buf_n822( .i (n821), .o (n822) );
  assign n1050 = n773 & n818 ;
  assign n1051 = n822 | n1050 ;
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  assign n1054 = n738 & n1053 ;
  buffer buf_n687( .i (n686), .o (n687) );
  assign n1055 = n672 & n734 ;
  assign n1056 = n687 | n1055 ;
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  assign n1060 = n1054 | n1059 ;
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  assign n1068 = n1049 | n1064 ;
  buffer buf_n196( .i (G27), .o (n196) );
  buffer buf_n361( .i (G48), .o (n361) );
  assign n1069 = n196 & n361 ;
  buffer buf_n1070( .i (n1069), .o (n1070) );
  assign n1113 = ~n512 & n1070 ;
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  assign n1131 = n959 & n1119 ;
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  assign n1135 = n985 | n1134 ;
  assign n1136 = n985 & n1134 ;
  assign n1137 = n1135 & ~n1136 ;
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n354( .i (G47), .o (n354) );
  assign n1140 = n1002 & n1118 ;
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  assign n1145 = n1030 | n1144 ;
  assign n1146 = n1030 & n1144 ;
  assign n1147 = n1145 & ~n1146 ;
  buffer buf_n1148( .i (n1147), .o (n1148) );
  assign n1149 = n354 & n1148 ;
  assign n1150 = ~n1139 & n1149 ;
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  assign n1157 = n409 & ~n512 ;
  buffer buf_n1158( .i (n1157), .o (n1158) );
  assign n1188 = n507 & ~n1158 ;
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n1207 = n1048 & ~n1130 ;
  buffer buf_n1208( .i (n1207), .o (n1208) );
  assign n1215 = ~n78 & n1208 ;
  assign n1216 = n1206 | n1215 ;
  buffer buf_n1217( .i (n608), .o (n1217) );
  assign n1218 = ~n158 & n1217 ;
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  assign n1234 = n1148 & n1233 ;
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  assign n1235 = ~n426 & n1158 ;
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  assign n1258 = ~n180 & n606 ;
  assign n1259 = n497 & ~n1258 ;
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n191( .i (n190), .o (n191) );
  assign n1273 = n191 & n606 ;
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n1277( .i (n244), .o (n1277) );
  assign n1278 = n181 & n1277 ;
  buffer buf_n1279( .i (n1278), .o (n1279) );
  assign n1280 = n195 & ~n1279 ;
  buffer buf_n1281( .i (n1280), .o (n1281) );
  assign n1282 = n1276 & n1281 ;
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n341( .i (G43), .o (n341) );
  assign n1286 = n299 | n341 ;
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  assign n1292 = ~n1284 & n1291 ;
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  assign n1293 = ~n251 & n337 ;
  assign n1294 = n319 & ~n1293 ;
  assign n1295 = ~n1292 & n1294 ;
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n182( .i (n181), .o (n182) );
  assign n1297 = n182 | n620 ;
  assign n1298 = n247 & n1297 ;
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  assign n1301 = n328 & n1300 ;
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n348( .i (G44), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  assign n1304 = n195 | n1279 ;
  buffer buf_n1305( .i (n1304), .o (n1305) );
  assign n1306 = n1276 | n1305 ;
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  assign n1310 = n353 & n1308 ;
  assign n1311 = n1303 | n1310 ;
  assign n1312 = ~n1276 & n1281 ;
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  assign n1316 = G45 | n333 ;
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  assign n1321 = ~n1314 & n1320 ;
  assign n1322 = n1276 & ~n1305 ;
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n339( .i (G42), .o (n339) );
  assign n1326 = G46 | n339 ;
  assign n1327 = ~n1324 & n1326 ;
  assign n1328 = n1321 | n1327 ;
  assign n1329 = n1311 | n1328 ;
  assign n1330 = n1296 & ~n1329 ;
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n252( .i (n251), .o (n252) );
  assign n1334 = n252 & n1314 ;
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  assign n1338 = n102 | n1336 ;
  buffer buf_n1339( .i (n1338), .o (n1339) );
  assign n1340 = n123 | n1284 ;
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  assign n1345 = n1339 & n1344 ;
  assign n1346 = n460 | n1284 ;
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  assign n1348 = n436 | n1315 ;
  assign n1349 = n1347 & n1348 ;
  buffer buf_n1325( .i (n1324), .o (n1325) );
  assign n1350 = n88 | n1325 ;
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  assign n1351 = ~n449 & n1309 ;
  assign n1352 = n1350 & ~n1351 ;
  assign n1353 = n1349 & n1352 ;
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  assign n1355 = n179 & ~n1325 ;
  assign n1356 = n321 | n1355 ;
  buffer buf_n1357( .i (n1356), .o (n1357) );
  assign n1358 = ~n109 & n1300 ;
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  assign n1364 = n1357 | n1363 ;
  assign n1365 = n1354 & ~n1364 ;
  assign n1366 = n1345 & n1365 ;
  assign n1367 = n1333 | n1366 ;
  assign n1368 = ~n1272 & n1367 ;
  assign n1369 = n1243 & ~n1368 ;
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  assign n1373 = ~n1234 & n1372 ;
  buffer buf_n1374( .i (n1373), .o (n1374) );
  assign n1375 = n354 & ~n1148 ;
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n1247( .i (n1246), .o (n1247) );
  assign n1379 = ~n354 & n1148 ;
  assign n1380 = n1247 | n1379 ;
  assign n1381 = n1376 | n1380 ;
  assign n1382 = ~n1374 & n1381 ;
  buffer buf_n1383( .i (n1382), .o (n1383) );
  inverter inv_n2496( .i (n1383), .o (n2496) );
  assign n1392 = n753 & n1118 ;
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  assign n1397 = n775 | n1396 ;
  assign n1398 = n775 & n1396 ;
  assign n1399 = n1397 & ~n1398 ;
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1409( .i (n311), .o (n1409) );
  assign n1410 = ~n155 & n1409 ;
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  assign n1429 = n1400 & n1428 ;
  buffer buf_n159( .i (G20), .o (n159) );
  assign n1430 = n159 & n1308 ;
  assign n1431 = ~n446 & n1300 ;
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n152( .i (G19), .o (n152) );
  assign n1433 = n152 & ~n1313 ;
  assign n1434 = n1432 | n1433 ;
  assign n1435 = n1430 | n1434 ;
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  assign n1440 = n439 | n1337 ;
  buffer buf_n143( .i (G18), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  assign n1441 = n150 & ~n1324 ;
  assign n1442 = ~n163 & n456 ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1283), .o (n1446) );
  assign n1447 = n1445 | n1446 ;
  assign n1448 = ~n1441 & n1447 ;
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  assign n1451 = ~n1357 & n1450 ;
  assign n1452 = n1440 & n1451 ;
  assign n1453 = ~n1439 & n1452 ;
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  assign n1454 = n330 & n1308 ;
  assign n1455 = n1360 | n1454 ;
  buffer buf_n338( .i (n337), .o (n338) );
  assign n1456 = n338 & ~n1314 ;
  assign n1457 = n93 & ~n299 ;
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  assign n1464 = n1446 | n1462 ;
  assign n1465 = ~n1456 & n1464 ;
  assign n1466 = ~n1455 & n1465 ;
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  assign n1470 = n127 | n1337 ;
  assign n1471 = n135 & ~n339 ;
  buffer buf_n1472( .i (n1471), .o (n1472) );
  assign n1473 = n1325 | n1472 ;
  assign n1474 = n321 & n1473 ;
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  assign n1477 = n1470 & n1476 ;
  assign n1478 = n1469 & n1477 ;
  assign n1479 = n1453 | n1478 ;
  assign n1480 = ~n1272 & n1479 ;
  assign n1481 = n1243 & ~n1480 ;
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  assign n1485 = ~n1429 & n1484 ;
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n1488( .i (n1487), .o (n1488) );
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  assign n1497 = n970 | n1013 ;
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  assign n1498 = n189 | n870 ;
  assign n1499 = n1497 | n1498 ;
  buffer buf_n1500( .i (n1499), .o (n1500) );
  assign n1501 = n934 | n1500 ;
  buffer buf_n1502( .i (n1501), .o (n1502) );
  assign n1503 = n973 & n1016 ;
  assign n1504 = n189 & n870 ;
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  assign n1507 = n934 & n1506 ;
  assign n1508 = n1503 & n1507 ;
  assign n1509 = n1502 & ~n1508 ;
  assign n1510 = n1121 | n1509 ;
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1518( .i (n1517), .o (n1518) );
  assign n1519 = n1036 & n1129 ;
  assign n1520 = n1518 & ~n1519 ;
  buffer buf_n1521( .i (n1520), .o (n1521) );
  assign n1522 = n360 & ~n1521 ;
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  assign n1526 = ~n1208 & n1406 ;
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  assign n1528 = ~n785 & n1209 ;
  assign n1529 = n1527 | n1528 ;
  buffer buf_n1530( .i (n1529), .o (n1530) );
  assign n1531 = n1525 | n1530 ;
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  assign n1533 = n1525 & n1530 ;
  assign n1534 = n1257 | n1533 ;
  assign n1535 = n1532 & ~n1534 ;
  assign n1536 = n1496 | n1535 ;
  buffer buf_n1537( .i (n1536), .o (n1537) );
  assign n1545 = n360 & n1521 ;
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  assign n1549 = n799 & n1119 ;
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  assign n1553 = n824 & ~n1552 ;
  assign n1554 = ~n824 & n1552 ;
  assign n1555 = n1553 | n1554 ;
  buffer buf_n1556( .i (n1555), .o (n1556) );
  assign n1566 = n1400 & n1556 ;
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  assign n1574 = n198 & ~n512 ;
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  assign n1583 = n712 & n1579 ;
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  assign n1588 = n736 | n1587 ;
  assign n1589 = n736 & n1587 ;
  assign n1590 = n1588 & ~n1589 ;
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  assign n1595 = n1567 & n1593 ;
  buffer buf_n1596( .i (n1595), .o (n1596) );
  assign n1602 = n831 & n1596 ;
  assign n1603 = n831 | n1596 ;
  assign n1604 = ~n1602 & n1603 ;
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  assign n1608 = n1547 & ~n1607 ;
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  assign n1612 = n834 | n1209 ;
  assign n1613 = ~n1067 & n1612 ;
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  assign n1615 = n821 & ~n1121 ;
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n1620( .i (n1619), .o (n1620) );
  assign n1621 = n773 & ~n1121 ;
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  assign n1634 = n1556 & ~n1625 ;
  assign n1635 = n1620 | n1634 ;
  buffer buf_n1636( .i (n1635), .o (n1636) );
  assign n1637 = n1594 & n1636 ;
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  assign n1639 = n734 & ~n1582 ;
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  assign n1649 = n1638 | n1648 ;
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  assign n1654 = n1614 & n1653 ;
  assign n1655 = n1614 | n1653 ;
  assign n1656 = ~n1654 & n1655 ;
  buffer buf_n1657( .i (n1656), .o (n1657) );
  assign n1658 = n1611 & n1657 ;
  assign n1659 = n1611 | n1657 ;
  assign n1660 = ~n1658 & n1659 ;
  buffer buf_n1661( .i (n51), .o (n1661) );
  assign n1662 = n154 | n1661 ;
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  assign n1668 = n476 & n1665 ;
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  assign n1699 = ~n1660 & n1698 ;
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  assign n1700 = n431 & ~n456 ;
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  assign n1701 = n470 | n548 ;
  assign n1702 = ~n1700 & n1701 ;
  assign n1703 = n1667 | n1702 ;
  assign n1704 = ~n132 & n501 ;
  assign n1705 = ~n893 & n1704 ;
  buffer buf_n1706( .i (n1705), .o (n1706) );
  assign n1707 = n1703 & ~n1706 ;
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  assign n1736 = n1699 | ~n1735 ;
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n862( .i (n861), .o (n862) );
  assign n1737 = ~n580 & n862 ;
  assign n1738 = ~n499 & n1737 ;
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1772( .i (n1120), .o (n1772) );
  assign n1773 = n1019 & ~n1772 ;
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  assign n1778 = n1138 | n1777 ;
  buffer buf_n1779( .i (n1778), .o (n1779) );
  assign n1780 = n985 & n1774 ;
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  assign n1785 = n1779 & ~n1784 ;
  buffer buf_n1786( .i (n1785), .o (n1786) );
  assign n1787 = n1378 | n1786 ;
  assign n1788 = n1378 & n1786 ;
  assign n1789 = n1787 & ~n1788 ;
  buffer buf_n1790( .i (n1789), .o (n1790) );
  assign n1791 = n1209 & n1790 ;
  assign n1792 = n1178 | n1791 ;
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  assign n1797 = n910 & n1118 ;
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  assign n1802 = n944 | n1801 ;
  assign n1803 = n944 & n1801 ;
  assign n1804 = n1802 & ~n1803 ;
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  assign n1810 = n976 & ~n1772 ;
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  buffer buf_n1813( .i (n1812), .o (n1813) );
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  assign n1817 = n1779 & ~n1816 ;
  buffer buf_n1818( .i (n1817), .o (n1818) );
  assign n1819 = n1809 | n1818 ;
  buffer buf_n1820( .i (n1819), .o (n1820) );
  assign n1821 = n1809 & n1818 ;
  buffer buf_n1822( .i (n1821), .o (n1822) );
  assign n1823 = n1820 & ~n1822 ;
  buffer buf_n1824( .i (n1823), .o (n1824) );
  assign n1825 = ~n1156 & n1824 ;
  buffer buf_n1826( .i (n1825), .o (n1826) );
  assign n1827 = n1156 & ~n1824 ;
  buffer buf_n1828( .i (n1827), .o (n1828) );
  assign n1830 = n1826 | n1828 ;
  buffer buf_n1831( .i (n1830), .o (n1831) );
  assign n1832 = n1214 & ~n1831 ;
  assign n1833 = n1796 | n1832 ;
  assign n1834 = ~n1767 & n1833 ;
  buffer buf_n1829( .i (n1828), .o (n1829) );
  assign n1835 = n938 & ~n1772 ;
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  assign n1846 = n1820 & ~n1845 ;
  buffer buf_n1847( .i (n1846), .o (n1847) );
  buffer buf_n1848( .i (n1117), .o (n1848) );
  assign n1849 = n853 & n1848 ;
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  assign n1853 = n885 | n1852 ;
  assign n1854 = n885 & n1852 ;
  assign n1855 = n1853 & ~n1854 ;
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  assign n1866 = n1847 & ~n1865 ;
  assign n1867 = ~n1847 & n1865 ;
  assign n1868 = n1866 | n1867 ;
  buffer buf_n1869( .i (n1868), .o (n1869) );
  assign n1870 = n1829 & ~n1869 ;
  assign n1871 = ~n1829 & n1869 ;
  assign n1872 = n1870 | n1871 ;
  buffer buf_n1873( .i (n1872), .o (n1873) );
  buffer buf_n1874( .i (n1873), .o (n1874) );
  assign n1875 = ~n1834 & n1874 ;
  assign n1876 = n1232 & n1856 ;
  assign n1877 = ~n152 & n434 ;
  buffer buf_n1878( .i (n1877), .o (n1878) );
  assign n1879 = n1325 | n1878 ;
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n1880( .i (n1307), .o (n1880) );
  assign n1881 = n167 & n1880 ;
  buffer buf_n1882( .i (n1313), .o (n1882) );
  assign n1883 = n159 & ~n1882 ;
  assign n1884 = n1881 | n1883 ;
  assign n1885 = n1879 & ~n1884 ;
  assign n1886 = n80 & ~n171 ;
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n1888( .i (n1887), .o (n1888) );
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  assign n1893 = n1446 | n1892 ;
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  assign n1896 = n1885 & n1895 ;
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  assign n1899 = ~n458 & n1300 ;
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  assign n1905 = n451 | n1336 ;
  assign n1906 = ~n1904 & n1905 ;
  assign n1907 = ~n324 & n1906 ;
  assign n1908 = n1898 & n1907 ;
  assign n1909 = n1291 & ~n1324 ;
  assign n1910 = n106 & ~n325 ;
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  assign n1916 = n1446 | n1914 ;
  assign n1917 = ~n1909 & n1916 ;
  buffer buf_n1918( .i (n1917), .o (n1918) );
  buffer buf_n1919( .i (n1918), .o (n1919) );
  buffer buf_n1920( .i (n1919), .o (n1920) );
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n340( .i (n339), .o (n340) );
  assign n1922 = n340 & ~n1882 ;
  assign n1923 = n338 & n1880 ;
  assign n1924 = n1922 | n1923 ;
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  assign n1928 = n139 | n1336 ;
  buffer buf_n1929( .i (n1299), .o (n1929) );
  assign n1930 = ~n121 & n1929 ;
  assign n1931 = n318 & ~n1930 ;
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n1934( .i (n1933), .o (n1934) );
  buffer buf_n1935( .i (n1934), .o (n1935) );
  assign n1936 = n1928 & n1935 ;
  assign n1937 = ~n1927 & n1936 ;
  assign n1938 = n1921 & n1937 ;
  assign n1939 = n1908 | n1938 ;
  assign n1940 = ~n1272 & n1939 ;
  assign n1941 = n1243 & ~n1940 ;
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  assign n1944 = ~n1876 & n1943 ;
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  buffer buf_n1954( .i (n1953), .o (n1954) );
  buffer buf_n1955( .i (n1954), .o (n1955) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  assign n1960 = n1875 | n1959 ;
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1208), .o (n1962) );
  assign n1963 = n1790 | n1962 ;
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  assign n1966 = ~n1793 & n1965 ;
  assign n1967 = n1760 & ~n1790 ;
  assign n1968 = n1138 & n1233 ;
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  assign n1969 = n303 & n1929 ;
  buffer buf_n1970( .i (n1969), .o (n1970) );
  buffer buf_n1971( .i (n1970), .o (n1971) );
  assign n1972 = n353 & ~n1882 ;
  assign n1973 = n1971 | n1972 ;
  buffer buf_n1974( .i (n1323), .o (n1974) );
  assign n1975 = n1320 & ~n1974 ;
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  assign n1976 = n347 & n1880 ;
  assign n1977 = n1975 | n1976 ;
  assign n1978 = n1973 | n1977 ;
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  assign n1980 = n332 & ~n1335 ;
  buffer buf_n1285( .i (n1284), .o (n1285) );
  assign n1981 = n1285 | n1472 ;
  assign n1982 = n321 & n1981 ;
  assign n1983 = ~n1980 & n1982 ;
  assign n1984 = ~n1979 & n1983 ;
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n1986( .i (n1985), .o (n1986) );
  assign n1987 = ~n435 & n1880 ;
  buffer buf_n1988( .i (n1987), .o (n1988) );
  assign n1989 = n179 & ~n1315 ;
  assign n1990 = n1988 | n1989 ;
  buffer buf_n1991( .i (n1283), .o (n1991) );
  assign n1992 = n111 | n1991 ;
  buffer buf_n1993( .i (n1992), .o (n1993) );
  buffer buf_n1994( .i (n1974), .o (n1994) );
  assign n1995 = n461 | n1994 ;
  assign n1996 = n1993 & n1995 ;
  assign n1997 = ~n1990 & n1996 ;
  buffer buf_n1998( .i (n1997), .o (n1998) );
  buffer buf_n1999( .i (n1998), .o (n1999) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n2000( .i (n1335), .o (n2000) );
  assign n2001 = n90 | n2000 ;
  buffer buf_n2002( .i (n2001), .o (n2002) );
  assign n2003 = n448 | n1991 ;
  assign n2004 = ~n320 & n2003 ;
  buffer buf_n2005( .i (n2004), .o (n2005) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  assign n2007 = ~n97 & n1929 ;
  buffer buf_n2008( .i (n2007), .o (n2008) );
  buffer buf_n2009( .i (n2008), .o (n2009) );
  buffer buf_n2010( .i (n2009), .o (n2010) );
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n168( .i (n167), .o (n168) );
  assign n2012 = n168 & ~n1994 ;
  buffer buf_n2013( .i (n2012), .o (n2013) );
  assign n2014 = n2011 | n2013 ;
  assign n2015 = n2006 & ~n2014 ;
  assign n2016 = n2002 & n2015 ;
  assign n2017 = n1999 & n2016 ;
  assign n2018 = n1986 | n2017 ;
  assign n2019 = ~n1272 & n2018 ;
  buffer buf_n2020( .i (n1242), .o (n2020) );
  assign n2021 = ~n2019 & n2020 ;
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  assign n2025 = ~n1968 & n2024 ;
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2028( .i (n2027), .o (n2028) );
  buffer buf_n2029( .i (n2028), .o (n2029) );
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n2031( .i (n2030), .o (n2031) );
  assign n2032 = n1967 | n2031 ;
  buffer buf_n2033( .i (n2032), .o (n2033) );
  buffer buf_n2034( .i (n2033), .o (n2034) );
  assign n2035 = n1966 | n2034 ;
  buffer buf_n2036( .i (n2035), .o (n2036) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  assign n2037 = ~n1179 & n1964 ;
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  assign n2040 = ~n1831 & n2039 ;
  buffer buf_n2041( .i (n2040), .o (n2041) );
  assign n2042 = n1233 & n1805 ;
  assign n2043 = n168 & ~n1315 ;
  buffer buf_n2044( .i (n447), .o (n2044) );
  assign n2045 = n1974 | n2044 ;
  assign n2046 = n98 & n434 ;
  assign n2047 = n1991 | n2046 ;
  assign n2048 = n2045 & n2047 ;
  assign n2049 = ~n2043 & n2048 ;
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  assign n2053 = n464 | n1337 ;
  buffer buf_n160( .i (n159), .o (n160) );
  assign n2054 = n160 & ~n1994 ;
  buffer buf_n2055( .i (n320), .o (n2055) );
  assign n2056 = n2054 | n2055 ;
  buffer buf_n2057( .i (n2056), .o (n2057) );
  assign n2059 = ~n85 & n1929 ;
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2063( .i (n1307), .o (n2063) );
  assign n2064 = n178 & n2063 ;
  assign n2065 = n2061 | n2064 ;
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n2067( .i (n2066), .o (n2067) );
  assign n2068 = n2057 | n2067 ;
  assign n2069 = n2053 & ~n2068 ;
  assign n2070 = n2052 & n2069 ;
  assign n2071 = n340 & n2063 ;
  assign n2072 = n325 | n348 ;
  buffer buf_n2073( .i (n2072), .o (n2073) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n2075( .i (n2074), .o (n2075) );
  buffer buf_n2076( .i (n2075), .o (n2076) );
  assign n2077 = ~n1974 & n2076 ;
  assign n2078 = n2071 | n2077 ;
  assign n2079 = n347 & ~n1882 ;
  buffer buf_n2080( .i (n1299), .o (n2080) );
  assign n2081 = ~n134 & n2080 ;
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  assign n2084 = n2079 | n2083 ;
  assign n2085 = n2078 | n2084 ;
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  assign n2089 = n309 & ~n1337 ;
  assign n2090 = n118 & ~n333 ;
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  assign n2096 = n1991 | n2094 ;
  assign n2097 = n320 & n2096 ;
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n2099( .i (n2098), .o (n2099) );
  buffer buf_n2100( .i (n2099), .o (n2100) );
  assign n2101 = ~n2089 & n2100 ;
  assign n2102 = ~n2088 & n2101 ;
  assign n2103 = n2070 | n2102 ;
  buffer buf_n2104( .i (n1271), .o (n2104) );
  assign n2105 = n2103 & ~n2104 ;
  assign n2106 = n2020 & ~n2105 ;
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  assign n2110 = ~n2042 & n2109 ;
  buffer buf_n2111( .i (n2110), .o (n2111) );
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  buffer buf_n2119( .i (n2118), .o (n2119) );
  buffer buf_n2120( .i (n2119), .o (n2120) );
  buffer buf_n2121( .i (n2120), .o (n2121) );
  assign n2122 = n1179 | n1964 ;
  assign n2123 = ~n1763 & n2122 ;
  buffer buf_n2124( .i (n2123), .o (n2124) );
  assign n2125 = n1831 & ~n2124 ;
  assign n2126 = n2121 | n2125 ;
  assign n2127 = n2041 | n2126 ;
  buffer buf_n2128( .i (n2127), .o (n2128) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  assign n2131 = n1547 & n1601 ;
  buffer buf_n2132( .i (n2131), .o (n2132) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  assign n2133 = n1546 & n1573 ;
  buffer buf_n2134( .i (n2133), .o (n2134) );
  assign n2135 = n1594 | n1636 ;
  buffer buf_n2136( .i (n2135), .o (n2136) );
  assign n2137 = ~n1638 & n2136 ;
  buffer buf_n2138( .i (n2137), .o (n2138) );
  buffer buf_n2139( .i (n2138), .o (n2139) );
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  assign n2142 = ~n2134 & n2141 ;
  assign n2143 = n2132 | n2142 ;
  buffer buf_n2144( .i (n2143), .o (n2144) );
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n1633( .i (n1632), .o (n1633) );
  assign n2151 = n1527 | n1633 ;
  buffer buf_n2152( .i (n2151), .o (n2152) );
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n1557( .i (n1556), .o (n1557) );
  buffer buf_n1558( .i (n1557), .o (n1558) );
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  assign n2155 = n1408 & n1546 ;
  assign n2156 = n1565 | n2155 ;
  assign n2157 = ~n2134 & n2156 ;
  buffer buf_n2158( .i (n2157), .o (n2158) );
  assign n2159 = n2154 | n2158 ;
  assign n2160 = n2154 & n2158 ;
  assign n2161 = n2159 & ~n2160 ;
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  assign n2163 = n1548 & ~n1614 ;
  buffer buf_n2164( .i (n2163), .o (n2164) );
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n2166( .i (n2165), .o (n2166) );
  buffer buf_n2167( .i (n2166), .o (n2167) );
  assign n2168 = n2162 | n2167 ;
  buffer buf_n2169( .i (n2168), .o (n2169) );
  assign n2170 = n1187 | n2169 ;
  assign n2171 = ~n1771 & n2170 ;
  assign n2172 = n2150 & ~n2171 ;
  buffer buf_n2173( .i (n2172), .o (n2173) );
  assign n2174 = ~n1187 & n2169 ;
  buffer buf_n2175( .i (n2174), .o (n2175) );
  assign n2176 = ~n2150 & n2175 ;
  assign n2177 = n1428 & n1591 ;
  buffer buf_n1915( .i (n1914), .o (n1915) );
  assign n2178 = n1915 | n1994 ;
  buffer buf_n2179( .i (n2178), .o (n2179) );
  buffer buf_n2180( .i (n2179), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  assign n2182 = n1339 & n2181 ;
  assign n2183 = ~n136 & n2063 ;
  buffer buf_n2184( .i (n2183), .o (n2184) );
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  assign n2186 = n1347 & ~n2062 ;
  assign n2187 = ~n2185 & n2186 ;
  assign n2188 = n306 & ~n1315 ;
  buffer buf_n2189( .i (n2188), .o (n2189) );
  assign n2190 = n1341 & n2055 ;
  assign n2191 = ~n2189 & n2190 ;
  assign n2192 = n2187 & n2191 ;
  buffer buf_n2193( .i (n2192), .o (n2193) );
  assign n2194 = n2182 & n2193 ;
  buffer buf_n140( .i (G16), .o (n140) );
  buffer buf_n2195( .i (n1323), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  assign n2197 = n140 & ~n2196 ;
  buffer buf_n141( .i (G17), .o (n141) );
  buffer buf_n2198( .i (n1313), .o (n2198) );
  assign n2199 = n141 & ~n2198 ;
  assign n2200 = n176 & n2080 ;
  buffer buf_n2201( .i (n2200), .o (n2201) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  assign n2203 = n2199 | n2202 ;
  assign n2204 = n2197 | n2203 ;
  buffer buf_n2205( .i (n2204), .o (n2205) );
  buffer buf_n2206( .i (n2205), .o (n2206) );
  buffer buf_n2207( .i (n2206), .o (n2207) );
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  assign n2208 = n170 & ~n2000 ;
  buffer buf_n151( .i (n150), .o (n151) );
  assign n2209 = n151 & n1309 ;
  assign n2210 = n1285 | n1878 ;
  assign n2211 = ~n2209 & n2210 ;
  buffer buf_n2212( .i (n2211), .o (n2212) );
  assign n2213 = ~n2208 & n2212 ;
  assign n2214 = ~n2058 & n2213 ;
  assign n2215 = ~n2207 & n2214 ;
  assign n2216 = n2194 | n2215 ;
  assign n2217 = ~n2104 & n2216 ;
  assign n2218 = n2020 & ~n2217 ;
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n2221( .i (n2220), .o (n2221) );
  assign n2222 = ~n2177 & n2221 ;
  buffer buf_n2223( .i (n2222), .o (n2223) );
  buffer buf_n2224( .i (n2223), .o (n2224) );
  buffer buf_n2225( .i (n2224), .o (n2225) );
  buffer buf_n2226( .i (n2225), .o (n2226) );
  buffer buf_n2227( .i (n2226), .o (n2227) );
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  buffer buf_n2231( .i (n2230), .o (n2231) );
  buffer buf_n2232( .i (n2231), .o (n2232) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  buffer buf_n2235( .i (n2234), .o (n2235) );
  buffer buf_n2236( .i (n2235), .o (n2236) );
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  assign n2241 = n2176 | n2240 ;
  assign n2242 = n2173 | n2241 ;
  buffer buf_n2243( .i (n2242), .o (n2243) );
  assign n2244 = n617 & n1579 ;
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  assign n2249 = n689 | n2248 ;
  assign n2250 = n689 & n2248 ;
  assign n2251 = n2249 & ~n2250 ;
  buffer buf_n2252( .i (n2251), .o (n2252) );
  assign n2260 = n1428 & n2252 ;
  assign n2261 = n143 | n171 ;
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  buffer buf_n2265( .i (n2264), .o (n2265) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  buffer buf_n2269( .i (n1283), .o (n2269) );
  assign n2270 = n2267 & ~n2269 ;
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2273( .i (n2272), .o (n2273) );
  buffer buf_n2274( .i (n2273), .o (n2274) );
  buffer buf_n2275( .i (n2274), .o (n2275) );
  buffer buf_n2276( .i (n2198), .o (n2276) );
  assign n2277 = n140 & ~n2276 ;
  buffer buf_n2278( .i (n2277), .o (n2278) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  assign n2280 = n162 & ~n2000 ;
  assign n2281 = n2279 | n2280 ;
  assign n2282 = n141 & n2063 ;
  assign n2283 = G15 | n152 ;
  assign n2284 = ~n2195 & n2283 ;
  assign n2285 = n2282 | n2284 ;
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  assign n2286 = n165 & n2080 ;
  assign n2287 = n643 & ~n2286 ;
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n2289( .i (n2288), .o (n2289) );
  assign n2290 = ~n2285 & n2289 ;
  buffer buf_n2291( .i (n2290), .o (n2291) );
  buffer buf_n2292( .i (n2291), .o (n2292) );
  assign n2293 = ~n2281 & n2292 ;
  assign n2294 = ~n2275 & n2293 ;
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  assign n2295 = n416 & n2002 ;
  assign n2296 = n137 | n2276 ;
  assign n2297 = ~n1902 & n2296 ;
  assign n2298 = ~n124 & n1309 ;
  assign n2299 = n1993 & ~n2298 ;
  assign n2300 = n2297 & n2299 ;
  buffer buf_n1463( .i (n1462), .o (n1463) );
  assign n2301 = n1463 | n2196 ;
  buffer buf_n2302( .i (n2301), .o (n2302) );
  assign n2303 = n2005 & n2302 ;
  assign n2304 = n2300 & n2303 ;
  buffer buf_n2305( .i (n2304), .o (n2305) );
  assign n2306 = n2295 & n2305 ;
  assign n2307 = n2294 | n2306 ;
  assign n2308 = ~n2104 & n2307 ;
  assign n2309 = n2020 & ~n2308 ;
  buffer buf_n2310( .i (n2309), .o (n2310) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  assign n2313 = ~n2260 & n2312 ;
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n2321( .i (n2320), .o (n2321) );
  buffer buf_n2322( .i (n2321), .o (n2322) );
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2325( .i (n2324), .o (n2325) );
  buffer buf_n2326( .i (n2325), .o (n2326) );
  buffer buf_n2327( .i (n2326), .o (n2327) );
  buffer buf_n2328( .i (n2327), .o (n2328) );
  buffer buf_n2329( .i (n2328), .o (n2329) );
  buffer buf_n2330( .i (n2329), .o (n2330) );
  buffer buf_n2331( .i (n2330), .o (n2331) );
  assign n2332 = n2162 & n2167 ;
  buffer buf_n2333( .i (n2332), .o (n2333) );
  assign n2336 = ~n2144 & n2165 ;
  assign n2337 = n1184 | n2336 ;
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  assign n2340 = n2333 | n2339 ;
  assign n2341 = ~n1771 & n2340 ;
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  assign n2342 = n1650 & ~n2259 ;
  assign n2343 = ~n1650 & n2259 ;
  assign n2344 = n2342 | n2343 ;
  buffer buf_n2345( .i (n2344), .o (n2345) );
  buffer buf_n2346( .i (n2345), .o (n2346) );
  assign n2347 = n2132 & ~n2346 ;
  assign n2348 = ~n2132 & n2346 ;
  assign n2349 = n2347 | n2348 ;
  buffer buf_n2350( .i (n2349), .o (n2350) );
  buffer buf_n2351( .i (n2350), .o (n2351) );
  buffer buf_n2352( .i (n2351), .o (n2352) );
  buffer buf_n2353( .i (n2352), .o (n2353) );
  buffer buf_n2354( .i (n2353), .o (n2354) );
  buffer buf_n2355( .i (n2354), .o (n2355) );
  assign n2356 = ~n2341 & n2355 ;
  assign n2357 = n2331 | n2356 ;
  buffer buf_n2358( .i (n2357), .o (n2358) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n2335( .i (n2334), .o (n2335) );
  assign n2360 = n2175 & ~n2335 ;
  assign n2361 = n1428 & n1556 ;
  assign n2362 = n306 & n1309 ;
  assign n2363 = n331 & ~n2276 ;
  assign n2364 = n2362 | n2363 ;
  assign n2365 = n87 & n136 ;
  assign n2366 = n1285 | n2365 ;
  assign n2367 = ~n2010 & n2366 ;
  assign n2368 = ~n2364 & n2367 ;
  buffer buf_n2369( .i (n2368), .o (n2369) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  assign n2370 = n114 | n2000 ;
  buffer buf_n2095( .i (n2094), .o (n2095) );
  assign n2371 = n2095 | n2196 ;
  assign n2372 = n2055 & n2371 ;
  buffer buf_n2373( .i (n2372), .o (n2373) );
  assign n2374 = n2370 & n2373 ;
  assign n2375 = n2369 & n2374 ;
  buffer buf_n142( .i (n141), .o (n142) );
  assign n2376 = n142 & ~n2196 ;
  buffer buf_n2377( .i (n2376), .o (n2377) );
  buffer buf_n2378( .i (n2377), .o (n2378) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n2379( .i (n1307), .o (n2379) );
  assign n2380 = n153 & n2379 ;
  buffer buf_n2381( .i (n2380), .o (n2381) );
  buffer buf_n2382( .i (n2381), .o (n2382) );
  assign n2383 = n2013 | n2382 ;
  assign n2384 = n2378 | n2383 ;
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  assign n2385 = n2268 & ~n2276 ;
  assign n2386 = n703 | n2385 ;
  assign n2387 = ~n433 & n2080 ;
  buffer buf_n2388( .i (n2387), .o (n2388) );
  buffer buf_n2389( .i (n2388), .o (n2389) );
  assign n2390 = n159 & ~n2269 ;
  assign n2391 = n2389 | n2390 ;
  buffer buf_n2392( .i (n2391), .o (n2392) );
  assign n2393 = n2386 | n2392 ;
  assign n2394 = n2006 & ~n2393 ;
  assign n2395 = ~n2384 & n2394 ;
  assign n2396 = n2375 | n2395 ;
  assign n2397 = ~n1271 & n2396 ;
  assign n2398 = n1242 & ~n2397 ;
  buffer buf_n2399( .i (n2398), .o (n2399) );
  buffer buf_n2400( .i (n2399), .o (n2400) );
  buffer buf_n2401( .i (n2400), .o (n2401) );
  buffer buf_n2402( .i (n2401), .o (n2402) );
  assign n2403 = ~n2361 & n2402 ;
  buffer buf_n2404( .i (n2403), .o (n2404) );
  buffer buf_n2405( .i (n2404), .o (n2405) );
  buffer buf_n2406( .i (n2405), .o (n2406) );
  buffer buf_n2407( .i (n2406), .o (n2407) );
  buffer buf_n2408( .i (n2407), .o (n2408) );
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  buffer buf_n2411( .i (n2410), .o (n2411) );
  buffer buf_n2412( .i (n2411), .o (n2412) );
  buffer buf_n2413( .i (n2412), .o (n2413) );
  buffer buf_n2414( .i (n2413), .o (n2414) );
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n2416( .i (n2415), .o (n2416) );
  buffer buf_n2417( .i (n2416), .o (n2417) );
  assign n2418 = n1768 & ~n2162 ;
  assign n2419 = n2417 | n2418 ;
  buffer buf_n2420( .i (n2419), .o (n2420) );
  buffer buf_n2421( .i (n2420), .o (n2421) );
  buffer buf_n2422( .i (n2421), .o (n2422) );
  assign n2423 = n2360 | n2422 ;
  buffer buf_n2424( .i (n2423), .o (n2424) );
  buffer buf_n2359( .i (n2358), .o (n2359) );
  assign n2425 = n2243 | n2359 ;
  buffer buf_n2426( .i (n2425), .o (n2426) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  assign n2427 = n1544 | n2424 ;
  buffer buf_n2428( .i (n2427), .o (n2428) );
  buffer buf_n2129( .i (n2128), .o (n2129) );
  buffer buf_n2130( .i (n2129), .o (n2130) );
  assign n2429 = n1961 | n2130 ;
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  assign n2431 = n1391 & ~n2036 ;
  buffer buf_n2432( .i (n2431), .o (n2432) );
  buffer buf_n2433( .i (n2432), .o (n2433) );
  buffer buf_n2434( .i (n2433), .o (n2434) );
  buffer buf_n2435( .i (n2434), .o (n2435) );
  buffer buf_n2436( .i (n2435), .o (n2436) );
  buffer buf_n2437( .i (n2436), .o (n2437) );
  assign n2438 = ~n2430 & n2437 ;
  buffer buf_n2439( .i (n2438), .o (n2439) );
  buffer buf_n2440( .i (n2439), .o (n2440) );
  buffer buf_n2441( .i (n2440), .o (n2441) );
  assign n2442 = ~n2428 & n2441 ;
  assign n2443 = ~n2426 & n2442 ;
  buffer buf_n2444( .i (n2443), .o (n2444) );
  inverter inv_n2497( .i (n2444), .o (n2497) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  assign n2445 = n402 & ~n2426 ;
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  assign n2448 = n239 & ~n2444 ;
  assign n2449 = n2447 | ~n2448 ;
  assign n2450 = n1544 & n2424 ;
  buffer buf_n2451( .i (n2450), .o (n2451) );
  assign n2452 = n2428 & ~n2451 ;
  buffer buf_n2453( .i (n2452), .o (n2453) );
  assign n2454 = ~n1391 & n2036 ;
  buffer buf_n2455( .i (n2454), .o (n2455) );
  assign n2456 = n2432 | n2455 ;
  buffer buf_n2457( .i (n2456), .o (n2457) );
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n2460( .i (n2459), .o (n2460) );
  buffer buf_n2461( .i (n2460), .o (n2461) );
  buffer buf_n2462( .i (n2461), .o (n2462) );
  assign n2463 = n1961 & n2130 ;
  buffer buf_n2464( .i (n2463), .o (n2464) );
  assign n2465 = n2430 & ~n2464 ;
  buffer buf_n2466( .i (n2465), .o (n2466) );
  assign n2467 = n2462 | n2466 ;
  assign n2468 = n2462 & n2466 ;
  assign n2469 = n2467 & ~n2468 ;
  buffer buf_n2470( .i (n2469), .o (n2470) );
  buffer buf_n2471( .i (n2470), .o (n2471) );
  assign n2472 = n2453 & n2471 ;
  assign n2473 = n2453 | n2471 ;
  assign n2474 = ~n2472 & n2473 ;
  buffer buf_n2475( .i (n2474), .o (n2475) );
  buffer buf_n2476( .i (n2475), .o (n2476) );
  buffer buf_n2477( .i (n2476), .o (n2477) );
  buffer buf_n417( .i (G50), .o (n417) );
  assign n2478 = n2243 & n2359 ;
  buffer buf_n2479( .i (n2478), .o (n2479) );
  assign n2480 = n2426 & ~n2479 ;
  buffer buf_n2481( .i (n2480), .o (n2481) );
  assign n2484 = n417 & n2481 ;
  buffer buf_n2485( .i (n2484), .o (n2485) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  assign n2486 = n417 | n2481 ;
  assign n2487 = ~n1112 & n2486 ;
  assign n2488 = ~n2485 & n2487 ;
  buffer buf_n2489( .i (n2488), .o (n2489) );
  assign n2490 = n2477 & n2489 ;
  assign n2491 = n2477 | n2489 ;
  assign n2492 = n2490 | ~n2491 ;
  buffer buf_n2482( .i (n2481), .o (n2482) );
  buffer buf_n2483( .i (n2482), .o (n2483) );
  assign n2493 = n2475 | n2483 ;
  assign n2494 = n2475 & n2483 ;
  assign n2495 = n2493 & ~n2494 ;
  assign G3519 = n471 ;
  assign G3520 = n474 ;
  assign G3521 = n517 ;
  assign G3522 = n544 ;
  assign G3523 = n571 ;
  assign G3524 = n1037 ;
  assign G3525 = n1068 ;
  assign G3526 = n1151 ;
  assign G3527 = n1216 ;
  assign G3528 = n2496 ;
  assign G3529 = n1537 ;
  assign G3530 = n1736 ;
  assign G3531 = n1961 ;
  assign G3532 = n2036 ;
  assign G3533 = n2128 ;
  assign G3534 = n2243 ;
  assign G3535 = n2358 ;
  assign G3536 = n2424 ;
  assign G3537 = n2497 ;
  assign G3538 = n2449 ;
  assign G3539 = n2492 ;
  assign G3540 = n2495 ;
endmodule
