module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( a_44_ , a_5_ , a_38_ , a_43_ , a_20_ , a_27_ , a_8_ , a_40_ , a_47_ , a_11_ , a_0_ , a_6_ , a_16_ , a_9_ , a_31_ , a_4_ , a_30_ , a_35_ , a_26_ , a_19_ , a_7_ , a_13_ , a_45_ , a_34_ , a_42_ , a_14_ , a_41_ , a_17_ , a_37_ , a_18_ , a_29_ , a_21_ , a_32_ , a_22_ , a_36_ , a_3_ , a_28_ , a_46_ , a_25_ , a_10_ , a_12_ , a_33_ , a_24_ , a_1_ , a_15_ , a_2_ , a_39_ , a_23_ , b_47_ , b_43_ , b_40_ , b_11_ , b_7_ , b_5_ , b_32_ , b_17_ , b_29_ , b_25_ , b_12_ , b_16_ , b_1_ , b_42_ , b_0_ , b_28_ , b_9_ , b_36_ , b_2_ , b_20_ , b_41_ , b_33_ , b_31_ , b_34_ , b_13_ , b_21_ , b_35_ , b_39_ , b_27_ , b_46_ , b_4_ , b_14_ , b_37_ , b_22_ , b_6_ , b_38_ , b_18_ , b_15_ , b_30_ , b_8_ , b_26_ , b_24_ , b_19_ , b_23_ , b_10_ , b_3_ , b_45_ , b_44_ );
  input a_44_ , a_5_ , a_38_ , a_43_ , a_20_ , a_27_ , a_8_ , a_40_ , a_47_ , a_11_ , a_0_ , a_6_ , a_16_ , a_9_ , a_31_ , a_4_ , a_30_ , a_35_ , a_26_ , a_19_ , a_7_ , a_13_ , a_45_ , a_34_ , a_42_ , a_14_ , a_41_ , a_17_ , a_37_ , a_18_ , a_29_ , a_21_ , a_32_ , a_22_ , a_36_ , a_3_ , a_28_ , a_46_ , a_25_ , a_10_ , a_12_ , a_33_ , a_24_ , a_1_ , a_15_ , a_2_ , a_39_ , a_23_ ;
  output b_47_ , b_43_ , b_40_ , b_11_ , b_7_ , b_5_ , b_32_ , b_17_ , b_29_ , b_25_ , b_12_ , b_16_ , b_1_ , b_42_ , b_0_ , b_28_ , b_9_ , b_36_ , b_2_ , b_20_ , b_41_ , b_33_ , b_31_ , b_34_ , b_13_ , b_21_ , b_35_ , b_39_ , b_27_ , b_46_ , b_4_ , b_14_ , b_37_ , b_22_ , b_6_ , b_38_ , b_18_ , b_15_ , b_30_ , b_8_ , b_26_ , b_24_ , b_19_ , b_23_ , b_10_ , b_3_ , b_45_ , b_44_ ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 ;
  assign n49 = a_35_ & a_34_ ;
  assign n50 = a_33_ & n49 ;
  buffer buf_n51( .i (n50), .o (n51) );
  assign n52 = a_31_ | a_32_ ;
  assign n53 = a_30_ | n52 ;
  buffer buf_n54( .i (n53), .o (n54) );
  assign n55 = n51 & n54 ;
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  assign n58 = a_35_ | a_34_ ;
  assign n59 = a_33_ | n58 ;
  buffer buf_n60( .i (n59), .o (n60) );
  assign n61 = a_31_ & a_32_ ;
  assign n62 = a_30_ & n61 ;
  buffer buf_n63( .i (n62), .o (n63) );
  assign n64 = n60 & n63 ;
  buffer buf_n65( .i (n64), .o (n65) );
  assign n66 = ( a_35_ & a_34_ ) | ( a_35_ & a_33_ ) | ( a_34_ & a_33_ ) ;
  buffer buf_n67( .i (n66), .o (n67) );
  assign n68 = ( a_31_ & a_30_ ) | ( a_31_ & a_32_ ) | ( a_30_ & a_32_ ) ;
  buffer buf_n69( .i (n68), .o (n69) );
  assign n70 = n67 & n69 ;
  buffer buf_n71( .i (n70), .o (n71) );
  assign n72 = n65 & n71 ;
  assign n73 = n57 & n72 ;
  buffer buf_n74( .i (n73), .o (n74) );
  assign n75 = a_29_ & a_28_ ;
  assign n76 = a_27_ & n75 ;
  buffer buf_n77( .i (n76), .o (n77) );
  assign n78 = a_26_ | a_25_ ;
  assign n79 = a_24_ | n78 ;
  buffer buf_n80( .i (n79), .o (n80) );
  assign n81 = n77 | n80 ;
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  assign n84 = ( a_27_ & a_29_ ) | ( a_27_ & a_28_ ) | ( a_29_ & a_28_ ) ;
  buffer buf_n85( .i (n84), .o (n85) );
  assign n86 = ( a_26_ & a_25_ ) | ( a_26_ & a_24_ ) | ( a_25_ & a_24_ ) ;
  buffer buf_n87( .i (n86), .o (n87) );
  assign n88 = n85 | n87 ;
  buffer buf_n89( .i (n88), .o (n89) );
  assign n90 = a_29_ | a_28_ ;
  assign n91 = a_27_ | n90 ;
  buffer buf_n92( .i (n91), .o (n92) );
  assign n93 = a_26_ & a_25_ ;
  assign n94 = a_24_ & n93 ;
  buffer buf_n95( .i (n94), .o (n95) );
  assign n96 = n92 | n95 ;
  buffer buf_n97( .i (n96), .o (n97) );
  assign n98 = n89 | n97 ;
  assign n99 = n83 | n98 ;
  buffer buf_n100( .i (n99), .o (n100) );
  assign n101 = n74 & n100 ;
  buffer buf_n102( .i (n101), .o (n102) );
  assign n103 = n51 | n54 ;
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  assign n106 = n60 | n63 ;
  buffer buf_n107( .i (n106), .o (n107) );
  assign n108 = n67 | n69 ;
  buffer buf_n109( .i (n108), .o (n109) );
  assign n110 = n107 & n109 ;
  assign n111 = n105 & n110 ;
  buffer buf_n112( .i (n111), .o (n112) );
  assign n113 = n77 & n80 ;
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  assign n116 = n85 & n87 ;
  buffer buf_n117( .i (n116), .o (n117) );
  assign n118 = n92 & n95 ;
  buffer buf_n119( .i (n118), .o (n119) );
  assign n120 = n117 | n119 ;
  assign n121 = n115 | n120 ;
  buffer buf_n122( .i (n121), .o (n122) );
  assign n123 = n112 & n122 ;
  buffer buf_n124( .i (n123), .o (n124) );
  assign n125 = n102 & n124 ;
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  assign n128 = ( n56 & n65 ) | ( n56 & n71 ) | ( n65 & n71 ) ;
  buffer buf_n129( .i (n128), .o (n129) );
  assign n130 = ( n82 & n89 ) | ( n82 & n97 ) | ( n89 & n97 ) ;
  buffer buf_n131( .i (n130), .o (n131) );
  assign n132 = n129 & n131 ;
  buffer buf_n133( .i (n132), .o (n133) );
  assign n134 = ( n104 & n107 ) | ( n104 & n109 ) | ( n107 & n109 ) ;
  buffer buf_n135( .i (n134), .o (n135) );
  assign n136 = ( n114 & n117 ) | ( n114 & n119 ) | ( n117 & n119 ) ;
  buffer buf_n137( .i (n136), .o (n137) );
  assign n138 = n135 & n137 ;
  buffer buf_n139( .i (n138), .o (n139) );
  assign n140 = n133 & n139 ;
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  assign n143 = n65 | n71 ;
  assign n144 = n57 | n143 ;
  buffer buf_n145( .i (n144), .o (n145) );
  assign n146 = n89 & n97 ;
  assign n147 = n83 & n146 ;
  buffer buf_n148( .i (n147), .o (n148) );
  assign n149 = n145 & n148 ;
  buffer buf_n150( .i (n149), .o (n150) );
  assign n151 = n107 | n109 ;
  assign n152 = n105 | n151 ;
  buffer buf_n153( .i (n152), .o (n153) );
  assign n154 = n117 & n119 ;
  assign n155 = n115 & n154 ;
  buffer buf_n156( .i (n155), .o (n156) );
  assign n157 = n153 & n156 ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n159 = n150 & n158 ;
  buffer buf_n160( .i (n159), .o (n160) );
  assign n161 = n142 & n160 ;
  assign n162 = n127 & n161 ;
  buffer buf_n163( .i (n162), .o (n163) );
  assign n164 = a_40_ & a_41_ ;
  assign n165 = a_39_ & n164 ;
  buffer buf_n166( .i (n165), .o (n166) );
  assign n167 = a_38_ | a_37_ ;
  assign n168 = a_36_ | n167 ;
  buffer buf_n169( .i (n168), .o (n169) );
  assign n170 = n166 & n169 ;
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  assign n173 = a_40_ | a_41_ ;
  assign n174 = a_39_ | n173 ;
  buffer buf_n175( .i (n174), .o (n175) );
  assign n176 = a_38_ & a_37_ ;
  assign n177 = a_36_ & n176 ;
  buffer buf_n178( .i (n177), .o (n178) );
  assign n179 = n175 & n178 ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = ( a_40_ & a_41_ ) | ( a_40_ & a_39_ ) | ( a_41_ & a_39_ ) ;
  buffer buf_n182( .i (n181), .o (n182) );
  assign n183 = ( a_38_ & a_37_ ) | ( a_38_ & a_36_ ) | ( a_37_ & a_36_ ) ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n185 = n182 & n184 ;
  buffer buf_n186( .i (n185), .o (n186) );
  assign n187 = n180 | n186 ;
  assign n188 = n172 | n187 ;
  buffer buf_n189( .i (n188), .o (n189) );
  assign n190 = ( a_44_ & a_43_ ) | ( a_44_ & a_42_ ) | ( a_43_ & a_42_ ) ;
  buffer buf_n191( .i (n190), .o (n191) );
  assign n192 = ( a_47_ & a_45_ ) | ( a_47_ & a_46_ ) | ( a_45_ & a_46_ ) ;
  buffer buf_n193( .i (n192), .o (n193) );
  assign n194 = n191 | n193 ;
  buffer buf_n195( .i (n194), .o (n195) );
  assign n196 = a_44_ & a_43_ ;
  assign n197 = a_42_ & n196 ;
  buffer buf_n198( .i (n197), .o (n198) );
  assign n199 = a_47_ | a_46_ ;
  assign n200 = a_45_ | n199 ;
  buffer buf_n201( .i (n200), .o (n201) );
  assign n202 = n198 | n201 ;
  buffer buf_n203( .i (n202), .o (n203) );
  assign n204 = n195 & n203 ;
  assign n205 = a_47_ & a_46_ ;
  assign n206 = a_45_ & n205 ;
  buffer buf_n207( .i (n206), .o (n207) );
  assign n208 = a_44_ | a_43_ ;
  assign n209 = a_42_ | n208 ;
  buffer buf_n210( .i (n209), .o (n210) );
  assign n211 = n207 | n210 ;
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  assign n214 = n204 & n213 ;
  buffer buf_n215( .i (n214), .o (n215) );
  assign n216 = n189 | n215 ;
  buffer buf_n217( .i (n216), .o (n217) );
  assign n218 = n166 | n169 ;
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  assign n221 = n175 | n178 ;
  buffer buf_n222( .i (n221), .o (n222) );
  assign n223 = n182 | n184 ;
  buffer buf_n224( .i (n223), .o (n224) );
  assign n225 = n222 | n224 ;
  assign n226 = n220 | n225 ;
  buffer buf_n227( .i (n226), .o (n227) );
  assign n228 = n191 & n193 ;
  buffer buf_n229( .i (n228), .o (n229) );
  assign n230 = n198 & n201 ;
  buffer buf_n231( .i (n230), .o (n231) );
  assign n232 = n229 & n231 ;
  assign n233 = n207 & n210 ;
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  assign n236 = n232 & n235 ;
  buffer buf_n237( .i (n236), .o (n237) );
  assign n238 = n227 | n237 ;
  buffer buf_n239( .i (n238), .o (n239) );
  assign n240 = n217 | n239 ;
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  assign n243 = n180 & n186 ;
  assign n244 = n172 & n243 ;
  buffer buf_n245( .i (n244), .o (n245) );
  assign n246 = n195 | n203 ;
  assign n247 = n213 | n246 ;
  buffer buf_n248( .i (n247), .o (n248) );
  assign n249 = n245 | n248 ;
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = n222 & n224 ;
  assign n252 = n220 & n251 ;
  buffer buf_n253( .i (n252), .o (n253) );
  assign n254 = n229 | n231 ;
  assign n255 = n235 | n254 ;
  buffer buf_n256( .i (n255), .o (n256) );
  assign n257 = n253 | n256 ;
  buffer buf_n258( .i (n257), .o (n258) );
  assign n259 = n250 | n258 ;
  buffer buf_n260( .i (n259), .o (n260) );
  assign n261 = ( n171 & n180 ) | ( n171 & n186 ) | ( n180 & n186 ) ;
  buffer buf_n262( .i (n261), .o (n262) );
  assign n263 = ( n195 & n203 ) | ( n195 & n212 ) | ( n203 & n212 ) ;
  buffer buf_n264( .i (n263), .o (n264) );
  assign n265 = n262 | n264 ;
  buffer buf_n266( .i (n265), .o (n266) );
  assign n267 = ( n219 & n222 ) | ( n219 & n224 ) | ( n222 & n224 ) ;
  buffer buf_n268( .i (n267), .o (n268) );
  assign n269 = ( n229 & n231 ) | ( n229 & n234 ) | ( n231 & n234 ) ;
  buffer buf_n270( .i (n269), .o (n270) );
  assign n271 = n268 | n270 ;
  buffer buf_n272( .i (n271), .o (n272) );
  assign n273 = n266 | n272 ;
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  assign n276 = n260 | n275 ;
  assign n277 = n242 | n276 ;
  buffer buf_n278( .i (n277), .o (n278) );
  assign n279 = n163 & n278 ;
  buffer buf_n280( .i (n279), .o (n280) );
  assign n281 = n74 | n100 ;
  buffer buf_n282( .i (n281), .o (n282) );
  assign n283 = n112 | n122 ;
  buffer buf_n284( .i (n283), .o (n284) );
  assign n285 = n282 & n284 ;
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  assign n288 = n145 | n148 ;
  buffer buf_n289( .i (n288), .o (n289) );
  assign n290 = n153 | n156 ;
  buffer buf_n291( .i (n290), .o (n291) );
  assign n292 = n289 & n291 ;
  buffer buf_n293( .i (n292), .o (n293) );
  assign n294 = n129 | n131 ;
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = n135 | n137 ;
  buffer buf_n297( .i (n296), .o (n297) );
  assign n298 = n295 & n297 ;
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  assign n301 = n293 & n300 ;
  assign n302 = n287 & n301 ;
  buffer buf_n303( .i (n302), .o (n303) );
  assign n304 = n189 & n215 ;
  buffer buf_n305( .i (n304), .o (n305) );
  assign n306 = n227 & n237 ;
  buffer buf_n307( .i (n306), .o (n307) );
  assign n308 = n305 | n307 ;
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  assign n311 = n245 & n248 ;
  buffer buf_n312( .i (n311), .o (n312) );
  assign n313 = n253 & n256 ;
  buffer buf_n314( .i (n313), .o (n314) );
  assign n315 = n312 | n314 ;
  buffer buf_n316( .i (n315), .o (n316) );
  assign n317 = n262 & n264 ;
  buffer buf_n318( .i (n317), .o (n318) );
  assign n319 = n268 & n270 ;
  buffer buf_n320( .i (n319), .o (n320) );
  assign n321 = n318 | n320 ;
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  assign n324 = n316 | n323 ;
  assign n325 = n310 | n324 ;
  buffer buf_n326( .i (n325), .o (n326) );
  assign n327 = n303 & n326 ;
  buffer buf_n328( .i (n327), .o (n328) );
  assign n329 = n280 & n328 ;
  buffer buf_n330( .i (n329), .o (n330) );
  assign n331 = n102 | n124 ;
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  assign n334 = n133 | n139 ;
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  assign n337 = n150 | n158 ;
  buffer buf_n338( .i (n337), .o (n338) );
  assign n339 = n336 & n338 ;
  assign n340 = n333 & n339 ;
  buffer buf_n341( .i (n340), .o (n341) );
  assign n342 = n217 & n239 ;
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  assign n345 = n250 & n258 ;
  buffer buf_n346( .i (n345), .o (n346) );
  assign n347 = n266 & n272 ;
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  assign n350 = n346 | n349 ;
  assign n351 = n344 | n350 ;
  buffer buf_n352( .i (n351), .o (n352) );
  assign n353 = n341 & n352 ;
  buffer buf_n354( .i (n353), .o (n354) );
  assign n355 = n282 | n284 ;
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  assign n358 = n289 | n291 ;
  buffer buf_n359( .i (n358), .o (n359) );
  assign n360 = n295 | n297 ;
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  assign n363 = n359 & n362 ;
  assign n364 = n357 & n363 ;
  buffer buf_n365( .i (n364), .o (n365) );
  assign n366 = n305 & n307 ;
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  assign n369 = n312 & n314 ;
  buffer buf_n370( .i (n369), .o (n370) );
  assign n371 = n318 & n320 ;
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  assign n374 = n370 | n373 ;
  assign n375 = n368 | n374 ;
  buffer buf_n376( .i (n375), .o (n376) );
  assign n377 = n365 & n376 ;
  buffer buf_n378( .i (n377), .o (n378) );
  assign n379 = n354 & n378 ;
  buffer buf_n380( .i (n379), .o (n380) );
  assign n381 = n330 & n380 ;
  buffer buf_n382( .i (n381), .o (n382) );
  assign n383 = ( n126 & n142 ) | ( n126 & n160 ) | ( n142 & n160 ) ;
  buffer buf_n384( .i (n383), .o (n384) );
  assign n385 = ( n241 & n260 ) | ( n241 & n275 ) | ( n260 & n275 ) ;
  buffer buf_n386( .i (n385), .o (n386) );
  assign n387 = n384 & n386 ;
  buffer buf_n388( .i (n387), .o (n388) );
  assign n389 = ( n286 & n293 ) | ( n286 & n300 ) | ( n293 & n300 ) ;
  buffer buf_n390( .i (n389), .o (n390) );
  assign n391 = ( n309 & n316 ) | ( n309 & n323 ) | ( n316 & n323 ) ;
  buffer buf_n392( .i (n391), .o (n392) );
  assign n393 = n390 & n392 ;
  buffer buf_n394( .i (n393), .o (n394) );
  assign n395 = n388 & n394 ;
  buffer buf_n396( .i (n395), .o (n396) );
  assign n397 = ( n332 & n336 ) | ( n332 & n338 ) | ( n336 & n338 ) ;
  buffer buf_n398( .i (n397), .o (n398) );
  assign n399 = ( n343 & n346 ) | ( n343 & n349 ) | ( n346 & n349 ) ;
  buffer buf_n400( .i (n399), .o (n400) );
  assign n401 = n398 & n400 ;
  buffer buf_n402( .i (n401), .o (n402) );
  assign n403 = ( n356 & n359 ) | ( n356 & n362 ) | ( n359 & n362 ) ;
  buffer buf_n404( .i (n403), .o (n404) );
  assign n405 = ( n367 & n370 ) | ( n367 & n373 ) | ( n370 & n373 ) ;
  buffer buf_n406( .i (n405), .o (n406) );
  assign n407 = n404 & n406 ;
  buffer buf_n408( .i (n407), .o (n408) );
  assign n409 = n402 & n408 ;
  buffer buf_n410( .i (n409), .o (n410) );
  assign n411 = n396 & n410 ;
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  assign n414 = n382 & n413 ;
  assign n415 = n142 | n160 ;
  assign n416 = n127 | n415 ;
  buffer buf_n417( .i (n416), .o (n417) );
  assign n418 = n260 & n275 ;
  assign n419 = n242 & n418 ;
  buffer buf_n420( .i (n419), .o (n420) );
  assign n421 = n417 & n420 ;
  buffer buf_n422( .i (n421), .o (n422) );
  assign n423 = n293 | n300 ;
  assign n424 = n287 | n423 ;
  buffer buf_n425( .i (n424), .o (n425) );
  assign n426 = n316 & n323 ;
  assign n427 = n310 & n426 ;
  buffer buf_n428( .i (n427), .o (n428) );
  assign n429 = n425 & n428 ;
  buffer buf_n430( .i (n429), .o (n430) );
  assign n431 = n422 & n430 ;
  buffer buf_n432( .i (n431), .o (n432) );
  assign n433 = n336 | n338 ;
  assign n434 = n333 | n433 ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n436 = n346 & n349 ;
  assign n437 = n344 & n436 ;
  buffer buf_n438( .i (n437), .o (n438) );
  assign n439 = n435 & n438 ;
  buffer buf_n440( .i (n439), .o (n440) );
  assign n441 = n359 | n362 ;
  assign n442 = n357 | n441 ;
  buffer buf_n443( .i (n442), .o (n443) );
  assign n444 = n370 & n373 ;
  assign n445 = n368 & n444 ;
  buffer buf_n446( .i (n445), .o (n446) );
  assign n447 = n443 & n446 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = n440 & n448 ;
  buffer buf_n450( .i (n449), .o (n450) );
  assign n451 = n432 & n450 ;
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  assign n454 = n414 & n453 ;
  buffer buf_n455( .i (n454), .o (n455) );
  assign n456 = a_11_ & a_10_ ;
  assign n457 = a_9_ & n456 ;
  buffer buf_n458( .i (n457), .o (n458) );
  assign n459 = a_8_ | a_7_ ;
  assign n460 = a_6_ | n459 ;
  buffer buf_n461( .i (n460), .o (n461) );
  assign n462 = n458 & n461 ;
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  assign n465 = a_11_ | a_10_ ;
  assign n466 = a_9_ | n465 ;
  buffer buf_n467( .i (n466), .o (n467) );
  assign n468 = a_8_ & a_7_ ;
  assign n469 = a_6_ & n468 ;
  buffer buf_n470( .i (n469), .o (n470) );
  assign n471 = n467 & n470 ;
  buffer buf_n472( .i (n471), .o (n472) );
  assign n473 = ( a_11_ & a_9_ ) | ( a_11_ & a_10_ ) | ( a_9_ & a_10_ ) ;
  buffer buf_n474( .i (n473), .o (n474) );
  assign n475 = ( a_8_ & a_6_ ) | ( a_8_ & a_7_ ) | ( a_6_ & a_7_ ) ;
  buffer buf_n476( .i (n475), .o (n476) );
  assign n477 = n474 & n476 ;
  buffer buf_n478( .i (n477), .o (n478) );
  assign n479 = n472 & n478 ;
  assign n480 = n464 & n479 ;
  buffer buf_n481( .i (n480), .o (n481) );
  assign n482 = a_5_ & a_4_ ;
  assign n483 = a_3_ & n482 ;
  buffer buf_n484( .i (n483), .o (n484) );
  assign n485 = a_1_ | a_2_ ;
  assign n486 = a_0_ | n485 ;
  buffer buf_n487( .i (n486), .o (n487) );
  assign n488 = n484 | n487 ;
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  assign n491 = a_5_ | a_4_ ;
  assign n492 = a_3_ | n491 ;
  buffer buf_n493( .i (n492), .o (n493) );
  assign n494 = a_1_ & a_2_ ;
  assign n495 = a_0_ & n494 ;
  buffer buf_n496( .i (n495), .o (n496) );
  assign n497 = n493 | n496 ;
  buffer buf_n498( .i (n497), .o (n498) );
  assign n499 = ( a_5_ & a_4_ ) | ( a_5_ & a_3_ ) | ( a_4_ & a_3_ ) ;
  buffer buf_n500( .i (n499), .o (n500) );
  assign n501 = ( a_0_ & a_1_ ) | ( a_0_ & a_2_ ) | ( a_1_ & a_2_ ) ;
  buffer buf_n502( .i (n501), .o (n502) );
  assign n503 = n500 | n502 ;
  buffer buf_n504( .i (n503), .o (n504) );
  assign n505 = n498 | n504 ;
  assign n506 = n490 | n505 ;
  buffer buf_n507( .i (n506), .o (n507) );
  assign n508 = n481 & n507 ;
  buffer buf_n509( .i (n508), .o (n509) );
  assign n510 = n458 | n461 ;
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  assign n513 = n467 | n470 ;
  buffer buf_n514( .i (n513), .o (n514) );
  assign n515 = n474 | n476 ;
  buffer buf_n516( .i (n515), .o (n516) );
  assign n517 = n514 & n516 ;
  assign n518 = n512 & n517 ;
  buffer buf_n519( .i (n518), .o (n519) );
  assign n520 = n484 & n487 ;
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  assign n523 = n493 & n496 ;
  buffer buf_n524( .i (n523), .o (n524) );
  assign n525 = n500 & n502 ;
  buffer buf_n526( .i (n525), .o (n526) );
  assign n527 = n524 | n526 ;
  assign n528 = n522 | n527 ;
  buffer buf_n529( .i (n528), .o (n529) );
  assign n530 = n519 & n529 ;
  buffer buf_n531( .i (n530), .o (n531) );
  assign n532 = n509 & n531 ;
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  assign n535 = n472 | n478 ;
  assign n536 = n464 | n535 ;
  buffer buf_n537( .i (n536), .o (n537) );
  assign n538 = n498 & n504 ;
  assign n539 = n490 & n538 ;
  buffer buf_n540( .i (n539), .o (n540) );
  assign n541 = n537 & n540 ;
  buffer buf_n542( .i (n541), .o (n542) );
  assign n543 = n514 | n516 ;
  assign n544 = n512 | n543 ;
  buffer buf_n545( .i (n544), .o (n545) );
  assign n546 = n524 & n526 ;
  assign n547 = n522 & n546 ;
  buffer buf_n548( .i (n547), .o (n548) );
  assign n549 = n545 & n548 ;
  buffer buf_n550( .i (n549), .o (n550) );
  assign n551 = n542 & n550 ;
  buffer buf_n552( .i (n551), .o (n552) );
  assign n553 = ( n463 & n472 ) | ( n463 & n478 ) | ( n472 & n478 ) ;
  buffer buf_n554( .i (n553), .o (n554) );
  assign n555 = ( n489 & n498 ) | ( n489 & n504 ) | ( n498 & n504 ) ;
  buffer buf_n556( .i (n555), .o (n556) );
  assign n557 = n554 & n556 ;
  buffer buf_n558( .i (n557), .o (n558) );
  assign n559 = ( n511 & n514 ) | ( n511 & n516 ) | ( n514 & n516 ) ;
  buffer buf_n560( .i (n559), .o (n560) );
  assign n561 = ( n521 & n524 ) | ( n521 & n526 ) | ( n524 & n526 ) ;
  buffer buf_n562( .i (n561), .o (n562) );
  assign n563 = n560 & n562 ;
  buffer buf_n564( .i (n563), .o (n564) );
  assign n565 = n558 & n564 ;
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  assign n568 = n552 & n567 ;
  assign n569 = n534 & n568 ;
  buffer buf_n570( .i (n569), .o (n570) );
  assign n571 = a_22_ & a_23_ ;
  assign n572 = a_21_ & n571 ;
  buffer buf_n573( .i (n572), .o (n573) );
  assign n574 = a_20_ | a_19_ ;
  assign n575 = a_18_ | n574 ;
  buffer buf_n576( .i (n575), .o (n576) );
  assign n577 = n573 | n576 ;
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  assign n580 = a_22_ | a_23_ ;
  assign n581 = a_21_ | n580 ;
  buffer buf_n582( .i (n581), .o (n582) );
  assign n583 = a_20_ & a_19_ ;
  assign n584 = a_18_ & n583 ;
  buffer buf_n585( .i (n584), .o (n585) );
  assign n586 = n582 | n585 ;
  buffer buf_n587( .i (n586), .o (n587) );
  assign n588 = ( a_21_ & a_22_ ) | ( a_21_ & a_23_ ) | ( a_22_ & a_23_ ) ;
  buffer buf_n589( .i (n588), .o (n589) );
  assign n590 = ( a_20_ & a_19_ ) | ( a_20_ & a_18_ ) | ( a_19_ & a_18_ ) ;
  buffer buf_n591( .i (n590), .o (n591) );
  assign n592 = n589 | n591 ;
  buffer buf_n593( .i (n592), .o (n593) );
  assign n594 = n587 & n593 ;
  assign n595 = n579 & n594 ;
  buffer buf_n596( .i (n595), .o (n596) );
  assign n597 = a_16_ & a_17_ ;
  assign n598 = a_15_ & n597 ;
  buffer buf_n599( .i (n598), .o (n599) );
  assign n600 = a_13_ | a_14_ ;
  assign n601 = a_12_ | n600 ;
  buffer buf_n602( .i (n601), .o (n602) );
  assign n603 = n599 & n602 ;
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  assign n606 = a_16_ | a_17_ ;
  assign n607 = a_15_ | n606 ;
  buffer buf_n608( .i (n607), .o (n608) );
  assign n609 = a_13_ & a_14_ ;
  assign n610 = a_12_ & n609 ;
  buffer buf_n611( .i (n610), .o (n611) );
  assign n612 = n608 & n611 ;
  buffer buf_n613( .i (n612), .o (n613) );
  assign n614 = ( a_16_ & a_17_ ) | ( a_16_ & a_15_ ) | ( a_17_ & a_15_ ) ;
  buffer buf_n615( .i (n614), .o (n615) );
  assign n616 = ( a_13_ & a_14_ ) | ( a_13_ & a_12_ ) | ( a_14_ & a_12_ ) ;
  buffer buf_n617( .i (n616), .o (n617) );
  assign n618 = n615 & n617 ;
  buffer buf_n619( .i (n618), .o (n619) );
  assign n620 = n613 | n619 ;
  assign n621 = n605 | n620 ;
  buffer buf_n622( .i (n621), .o (n622) );
  assign n623 = n596 | n622 ;
  buffer buf_n624( .i (n623), .o (n624) );
  assign n625 = n573 & n576 ;
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  assign n628 = n582 & n585 ;
  buffer buf_n629( .i (n628), .o (n629) );
  assign n630 = n589 & n591 ;
  buffer buf_n631( .i (n630), .o (n631) );
  assign n632 = n629 & n631 ;
  assign n633 = n627 & n632 ;
  buffer buf_n634( .i (n633), .o (n634) );
  assign n635 = n608 | n611 ;
  buffer buf_n636( .i (n635), .o (n636) );
  assign n637 = n615 | n617 ;
  buffer buf_n638( .i (n637), .o (n638) );
  assign n639 = n636 | n638 ;
  assign n640 = n599 | n602 ;
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  assign n643 = n639 | n642 ;
  buffer buf_n644( .i (n643), .o (n644) );
  assign n645 = n634 | n644 ;
  buffer buf_n646( .i (n645), .o (n646) );
  assign n647 = n624 | n646 ;
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  assign n650 = n587 | n593 ;
  assign n651 = n579 | n650 ;
  buffer buf_n652( .i (n651), .o (n652) );
  assign n653 = n613 & n619 ;
  assign n654 = n605 & n653 ;
  buffer buf_n655( .i (n654), .o (n655) );
  assign n656 = n652 | n655 ;
  buffer buf_n657( .i (n656), .o (n657) );
  assign n658 = n629 | n631 ;
  assign n659 = n627 | n658 ;
  buffer buf_n660( .i (n659), .o (n660) );
  assign n661 = n636 & n638 ;
  assign n662 = n642 & n661 ;
  buffer buf_n663( .i (n662), .o (n663) );
  assign n664 = n660 | n663 ;
  buffer buf_n665( .i (n664), .o (n665) );
  assign n666 = n657 | n665 ;
  buffer buf_n667( .i (n666), .o (n667) );
  assign n668 = ( n578 & n587 ) | ( n578 & n593 ) | ( n587 & n593 ) ;
  buffer buf_n669( .i (n668), .o (n669) );
  assign n670 = ( n604 & n613 ) | ( n604 & n619 ) | ( n613 & n619 ) ;
  buffer buf_n671( .i (n670), .o (n671) );
  assign n672 = n669 | n671 ;
  buffer buf_n673( .i (n672), .o (n673) );
  assign n674 = ( n626 & n629 ) | ( n626 & n631 ) | ( n629 & n631 ) ;
  buffer buf_n675( .i (n674), .o (n675) );
  assign n676 = ( n636 & n638 ) | ( n636 & n641 ) | ( n638 & n641 ) ;
  buffer buf_n677( .i (n676), .o (n677) );
  assign n678 = n675 | n677 ;
  buffer buf_n679( .i (n678), .o (n679) );
  assign n680 = n673 | n679 ;
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  assign n683 = n667 | n682 ;
  assign n684 = n649 | n683 ;
  buffer buf_n685( .i (n684), .o (n685) );
  assign n686 = n570 | n685 ;
  buffer buf_n687( .i (n686), .o (n687) );
  assign n688 = n481 | n507 ;
  buffer buf_n689( .i (n688), .o (n689) );
  assign n690 = n519 | n529 ;
  buffer buf_n691( .i (n690), .o (n691) );
  assign n692 = n689 & n691 ;
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  assign n695 = n554 | n556 ;
  buffer buf_n696( .i (n695), .o (n696) );
  assign n697 = n560 | n562 ;
  buffer buf_n698( .i (n697), .o (n698) );
  assign n699 = n696 & n698 ;
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  assign n702 = n537 | n540 ;
  buffer buf_n703( .i (n702), .o (n703) );
  assign n704 = n545 | n548 ;
  buffer buf_n705( .i (n704), .o (n705) );
  assign n706 = n703 & n705 ;
  buffer buf_n707( .i (n706), .o (n707) );
  assign n708 = n701 & n707 ;
  assign n709 = n694 & n708 ;
  buffer buf_n710( .i (n709), .o (n710) );
  assign n711 = n596 & n622 ;
  buffer buf_n712( .i (n711), .o (n712) );
  assign n713 = n634 & n644 ;
  buffer buf_n714( .i (n713), .o (n714) );
  assign n715 = n712 | n714 ;
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  assign n718 = n652 & n655 ;
  buffer buf_n719( .i (n718), .o (n719) );
  assign n720 = n660 & n663 ;
  buffer buf_n721( .i (n720), .o (n721) );
  assign n722 = n719 | n721 ;
  buffer buf_n723( .i (n722), .o (n723) );
  assign n724 = n669 & n671 ;
  buffer buf_n725( .i (n724), .o (n725) );
  assign n726 = n675 & n677 ;
  buffer buf_n727( .i (n726), .o (n727) );
  assign n728 = n725 | n727 ;
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  assign n731 = n723 | n730 ;
  assign n732 = n717 | n731 ;
  buffer buf_n733( .i (n732), .o (n733) );
  assign n734 = n710 | n733 ;
  buffer buf_n735( .i (n734), .o (n735) );
  assign n736 = n687 | n735 ;
  buffer buf_n737( .i (n736), .o (n737) );
  assign n738 = n542 | n550 ;
  buffer buf_n739( .i (n738), .o (n739) );
  assign n740 = n558 | n564 ;
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  assign n743 = n739 & n742 ;
  assign n744 = n509 | n531 ;
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  assign n747 = n743 & n746 ;
  buffer buf_n748( .i (n747), .o (n748) );
  assign n749 = n624 & n646 ;
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  assign n752 = n657 & n665 ;
  buffer buf_n753( .i (n752), .o (n753) );
  assign n754 = n673 & n679 ;
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  assign n757 = n753 | n756 ;
  assign n758 = n751 | n757 ;
  buffer buf_n759( .i (n758), .o (n759) );
  assign n760 = n748 | n759 ;
  buffer buf_n761( .i (n760), .o (n761) );
  assign n762 = n689 | n691 ;
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  assign n765 = n696 | n698 ;
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  assign n768 = n703 | n705 ;
  buffer buf_n769( .i (n768), .o (n769) );
  assign n770 = n767 & n769 ;
  assign n771 = n764 & n770 ;
  buffer buf_n772( .i (n771), .o (n772) );
  assign n773 = n712 & n714 ;
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  assign n776 = n719 & n721 ;
  buffer buf_n777( .i (n776), .o (n777) );
  assign n778 = n725 & n727 ;
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  assign n781 = n777 | n780 ;
  assign n782 = n775 | n781 ;
  buffer buf_n783( .i (n782), .o (n783) );
  assign n784 = n772 | n783 ;
  buffer buf_n785( .i (n784), .o (n785) );
  assign n786 = n761 | n785 ;
  buffer buf_n787( .i (n786), .o (n787) );
  assign n788 = n737 | n787 ;
  buffer buf_n789( .i (n788), .o (n789) );
  assign n790 = ( n533 & n552 ) | ( n533 & n567 ) | ( n552 & n567 ) ;
  buffer buf_n791( .i (n790), .o (n791) );
  assign n792 = ( n648 & n667 ) | ( n648 & n682 ) | ( n667 & n682 ) ;
  buffer buf_n793( .i (n792), .o (n793) );
  assign n794 = n791 | n793 ;
  buffer buf_n795( .i (n794), .o (n795) );
  assign n796 = ( n693 & n701 ) | ( n693 & n707 ) | ( n701 & n707 ) ;
  buffer buf_n797( .i (n796), .o (n797) );
  assign n798 = ( n716 & n723 ) | ( n716 & n730 ) | ( n723 & n730 ) ;
  buffer buf_n799( .i (n798), .o (n799) );
  assign n800 = n797 | n799 ;
  buffer buf_n801( .i (n800), .o (n801) );
  assign n802 = n795 | n801 ;
  buffer buf_n803( .i (n802), .o (n803) );
  assign n804 = ( n739 & n742 ) | ( n739 & n745 ) | ( n742 & n745 ) ;
  buffer buf_n805( .i (n804), .o (n805) );
  assign n806 = ( n750 & n753 ) | ( n750 & n756 ) | ( n753 & n756 ) ;
  buffer buf_n807( .i (n806), .o (n807) );
  assign n808 = n805 | n807 ;
  buffer buf_n809( .i (n808), .o (n809) );
  assign n810 = ( n763 & n767 ) | ( n763 & n769 ) | ( n767 & n769 ) ;
  buffer buf_n811( .i (n810), .o (n811) );
  assign n812 = ( n774 & n777 ) | ( n774 & n780 ) | ( n777 & n780 ) ;
  buffer buf_n813( .i (n812), .o (n813) );
  assign n814 = n811 | n813 ;
  buffer buf_n815( .i (n814), .o (n815) );
  assign n816 = n809 | n815 ;
  buffer buf_n817( .i (n816), .o (n817) );
  assign n818 = n803 | n817 ;
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  assign n821 = n789 | n820 ;
  assign n822 = n552 | n567 ;
  assign n823 = n534 | n822 ;
  buffer buf_n824( .i (n823), .o (n824) );
  assign n825 = n667 & n682 ;
  assign n826 = n649 & n825 ;
  buffer buf_n827( .i (n826), .o (n827) );
  assign n828 = n824 | n827 ;
  buffer buf_n829( .i (n828), .o (n829) );
  assign n830 = n701 | n707 ;
  assign n831 = n694 | n830 ;
  buffer buf_n832( .i (n831), .o (n832) );
  assign n833 = n723 & n730 ;
  assign n834 = n717 & n833 ;
  buffer buf_n835( .i (n834), .o (n835) );
  assign n836 = n832 | n835 ;
  buffer buf_n837( .i (n836), .o (n837) );
  assign n838 = n829 | n837 ;
  buffer buf_n839( .i (n838), .o (n839) );
  assign n840 = n739 | n742 ;
  assign n841 = n746 | n840 ;
  buffer buf_n842( .i (n841), .o (n842) );
  assign n843 = n753 & n756 ;
  assign n844 = n751 & n843 ;
  buffer buf_n845( .i (n844), .o (n845) );
  assign n846 = n842 | n845 ;
  buffer buf_n847( .i (n846), .o (n847) );
  assign n848 = n767 | n769 ;
  assign n849 = n764 | n848 ;
  buffer buf_n850( .i (n849), .o (n850) );
  assign n851 = n777 & n780 ;
  assign n852 = n775 & n851 ;
  buffer buf_n853( .i (n852), .o (n853) );
  assign n854 = n850 | n853 ;
  buffer buf_n855( .i (n854), .o (n855) );
  assign n856 = n847 | n855 ;
  buffer buf_n857( .i (n856), .o (n857) );
  assign n858 = n839 | n857 ;
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  assign n861 = n821 | n860 ;
  buffer buf_n862( .i (n861), .o (n862) );
  assign n863 = n455 | n862 ;
  buffer buf_n864( .i (n863), .o (n864) );
  assign n865 = n163 | n278 ;
  buffer buf_n866( .i (n865), .o (n866) );
  assign n867 = n303 | n326 ;
  buffer buf_n868( .i (n867), .o (n868) );
  assign n869 = n866 & n868 ;
  buffer buf_n870( .i (n869), .o (n870) );
  assign n871 = n341 | n352 ;
  buffer buf_n872( .i (n871), .o (n872) );
  assign n873 = n365 | n376 ;
  buffer buf_n874( .i (n873), .o (n874) );
  assign n875 = n872 & n874 ;
  buffer buf_n876( .i (n875), .o (n876) );
  assign n877 = n870 & n876 ;
  buffer buf_n878( .i (n877), .o (n878) );
  assign n879 = n384 | n386 ;
  buffer buf_n880( .i (n879), .o (n880) );
  assign n881 = n390 | n392 ;
  buffer buf_n882( .i (n881), .o (n882) );
  assign n883 = n880 & n882 ;
  buffer buf_n884( .i (n883), .o (n884) );
  assign n885 = n398 | n400 ;
  buffer buf_n886( .i (n885), .o (n886) );
  assign n887 = n404 | n406 ;
  buffer buf_n888( .i (n887), .o (n888) );
  assign n889 = n886 & n888 ;
  buffer buf_n890( .i (n889), .o (n890) );
  assign n891 = n884 & n890 ;
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  assign n894 = n878 & n893 ;
  assign n895 = n417 | n420 ;
  buffer buf_n896( .i (n895), .o (n896) );
  assign n897 = n425 | n428 ;
  buffer buf_n898( .i (n897), .o (n898) );
  assign n899 = n896 & n898 ;
  buffer buf_n900( .i (n899), .o (n900) );
  assign n901 = n435 | n438 ;
  buffer buf_n902( .i (n901), .o (n902) );
  assign n903 = n443 | n446 ;
  buffer buf_n904( .i (n903), .o (n904) );
  assign n905 = n902 & n904 ;
  buffer buf_n906( .i (n905), .o (n906) );
  assign n907 = n900 & n906 ;
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  assign n910 = n894 & n909 ;
  buffer buf_n911( .i (n910), .o (n911) );
  assign n912 = n570 & n685 ;
  buffer buf_n913( .i (n912), .o (n913) );
  assign n914 = n710 & n733 ;
  buffer buf_n915( .i (n914), .o (n915) );
  assign n916 = n913 | n915 ;
  buffer buf_n917( .i (n916), .o (n917) );
  assign n918 = n748 & n759 ;
  buffer buf_n919( .i (n918), .o (n919) );
  assign n920 = n772 & n783 ;
  buffer buf_n921( .i (n920), .o (n921) );
  assign n922 = n919 | n921 ;
  buffer buf_n923( .i (n922), .o (n923) );
  assign n924 = n917 | n923 ;
  buffer buf_n925( .i (n924), .o (n925) );
  assign n926 = n791 & n793 ;
  buffer buf_n927( .i (n926), .o (n927) );
  assign n928 = n797 & n799 ;
  buffer buf_n929( .i (n928), .o (n929) );
  assign n930 = n927 | n929 ;
  buffer buf_n931( .i (n930), .o (n931) );
  assign n932 = n805 & n807 ;
  buffer buf_n933( .i (n932), .o (n933) );
  assign n934 = n811 & n813 ;
  buffer buf_n935( .i (n934), .o (n935) );
  assign n936 = n933 | n935 ;
  buffer buf_n937( .i (n936), .o (n937) );
  assign n938 = n931 | n937 ;
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  assign n941 = n925 | n940 ;
  assign n942 = n824 & n827 ;
  buffer buf_n943( .i (n942), .o (n943) );
  assign n944 = n832 & n835 ;
  buffer buf_n945( .i (n944), .o (n945) );
  assign n946 = n943 | n945 ;
  buffer buf_n947( .i (n946), .o (n947) );
  assign n948 = n842 & n845 ;
  buffer buf_n949( .i (n948), .o (n949) );
  assign n950 = n850 & n853 ;
  buffer buf_n951( .i (n950), .o (n951) );
  assign n952 = n949 | n951 ;
  buffer buf_n953( .i (n952), .o (n953) );
  assign n954 = n947 | n953 ;
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  assign n957 = n941 | n956 ;
  buffer buf_n958( .i (n957), .o (n958) );
  assign n959 = n911 | n958 ;
  buffer buf_n960( .i (n959), .o (n960) );
  assign n961 = n864 | n960 ;
  buffer buf_n962( .i (n961), .o (n962) );
  assign n963 = n280 | n328 ;
  buffer buf_n964( .i (n963), .o (n964) );
  assign n965 = n354 | n378 ;
  buffer buf_n966( .i (n965), .o (n966) );
  assign n967 = n964 & n966 ;
  buffer buf_n968( .i (n967), .o (n968) );
  assign n969 = n388 | n394 ;
  buffer buf_n970( .i (n969), .o (n970) );
  assign n971 = n402 | n408 ;
  buffer buf_n972( .i (n971), .o (n972) );
  assign n973 = n970 & n972 ;
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  assign n976 = n968 & n975 ;
  assign n977 = n422 | n430 ;
  buffer buf_n978( .i (n977), .o (n978) );
  assign n979 = n440 | n448 ;
  buffer buf_n980( .i (n979), .o (n980) );
  assign n981 = n978 & n980 ;
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  assign n984 = n976 & n983 ;
  buffer buf_n985( .i (n984), .o (n985) );
  assign n986 = n687 & n735 ;
  buffer buf_n987( .i (n986), .o (n987) );
  assign n988 = n761 & n785 ;
  buffer buf_n989( .i (n988), .o (n989) );
  assign n990 = n987 | n989 ;
  buffer buf_n991( .i (n990), .o (n991) );
  assign n992 = n795 & n801 ;
  buffer buf_n993( .i (n992), .o (n993) );
  assign n994 = n809 & n815 ;
  buffer buf_n995( .i (n994), .o (n995) );
  assign n996 = n993 | n995 ;
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  assign n999 = n991 | n998 ;
  assign n1000 = n829 & n837 ;
  buffer buf_n1001( .i (n1000), .o (n1001) );
  assign n1002 = n847 & n855 ;
  buffer buf_n1003( .i (n1002), .o (n1003) );
  assign n1004 = n1001 | n1003 ;
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  assign n1007 = n999 | n1006 ;
  buffer buf_n1008( .i (n1007), .o (n1008) );
  assign n1009 = n985 | n1008 ;
  buffer buf_n1010( .i (n1009), .o (n1010) );
  assign n1011 = n866 | n868 ;
  buffer buf_n1012( .i (n1011), .o (n1012) );
  assign n1013 = n872 | n874 ;
  buffer buf_n1014( .i (n1013), .o (n1014) );
  assign n1015 = n1012 & n1014 ;
  buffer buf_n1016( .i (n1015), .o (n1016) );
  assign n1017 = n880 | n882 ;
  buffer buf_n1018( .i (n1017), .o (n1018) );
  assign n1019 = n886 | n888 ;
  buffer buf_n1020( .i (n1019), .o (n1020) );
  assign n1021 = n1018 & n1020 ;
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  assign n1024 = n1016 & n1023 ;
  assign n1025 = n896 | n898 ;
  buffer buf_n1026( .i (n1025), .o (n1026) );
  assign n1027 = n902 | n904 ;
  buffer buf_n1028( .i (n1027), .o (n1028) );
  assign n1029 = n1026 & n1028 ;
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  assign n1032 = n1024 & n1031 ;
  buffer buf_n1033( .i (n1032), .o (n1033) );
  assign n1034 = n913 & n915 ;
  buffer buf_n1035( .i (n1034), .o (n1035) );
  assign n1036 = n919 & n921 ;
  buffer buf_n1037( .i (n1036), .o (n1037) );
  assign n1038 = n1035 | n1037 ;
  buffer buf_n1039( .i (n1038), .o (n1039) );
  assign n1040 = n927 & n929 ;
  buffer buf_n1041( .i (n1040), .o (n1041) );
  assign n1042 = n933 & n935 ;
  buffer buf_n1043( .i (n1042), .o (n1043) );
  assign n1044 = n1041 | n1043 ;
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  assign n1047 = n1039 | n1046 ;
  assign n1048 = n943 & n945 ;
  buffer buf_n1049( .i (n1048), .o (n1049) );
  assign n1050 = n949 & n951 ;
  buffer buf_n1051( .i (n1050), .o (n1051) );
  assign n1052 = n1049 | n1051 ;
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  assign n1055 = n1047 | n1054 ;
  buffer buf_n1056( .i (n1055), .o (n1056) );
  assign n1057 = n1033 | n1056 ;
  buffer buf_n1058( .i (n1057), .o (n1058) );
  assign n1059 = n1010 | n1058 ;
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1061 = n962 | n1060 ;
  buffer buf_n1062( .i (n1061), .o (n1062) );
  assign n1063 = n330 | n380 ;
  buffer buf_n1064( .i (n1063), .o (n1064) );
  assign n1065 = n396 | n410 ;
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  assign n1068 = n1064 & n1067 ;
  assign n1069 = n432 | n450 ;
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  assign n1072 = n1068 & n1071 ;
  buffer buf_n1073( .i (n1072), .o (n1073) );
  assign n1074 = n737 & n787 ;
  buffer buf_n1075( .i (n1074), .o (n1075) );
  assign n1076 = n803 & n817 ;
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  assign n1079 = n1075 | n1078 ;
  assign n1080 = n839 & n857 ;
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  assign n1083 = n1079 | n1082 ;
  buffer buf_n1084( .i (n1083), .o (n1084) );
  assign n1085 = n1073 | n1084 ;
  buffer buf_n1086( .i (n1085), .o (n1086) );
  assign n1087 = n870 | n876 ;
  buffer buf_n1088( .i (n1087), .o (n1088) );
  assign n1089 = n884 | n890 ;
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  assign n1092 = n1088 & n1091 ;
  assign n1093 = n900 | n906 ;
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  assign n1096 = n1092 & n1095 ;
  buffer buf_n1097( .i (n1096), .o (n1097) );
  assign n1098 = n917 & n923 ;
  buffer buf_n1099( .i (n1098), .o (n1099) );
  assign n1100 = n931 & n937 ;
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  assign n1103 = n1099 | n1102 ;
  assign n1104 = n947 & n953 ;
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  assign n1107 = n1103 | n1106 ;
  buffer buf_n1108( .i (n1107), .o (n1108) );
  assign n1109 = n1097 | n1108 ;
  buffer buf_n1110( .i (n1109), .o (n1110) );
  assign n1111 = n1086 | n1110 ;
  buffer buf_n1112( .i (n1111), .o (n1112) );
  assign n1113 = n964 | n966 ;
  buffer buf_n1114( .i (n1113), .o (n1114) );
  assign n1115 = n970 | n972 ;
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  assign n1118 = n1114 & n1117 ;
  assign n1119 = n978 | n980 ;
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  assign n1122 = n1118 & n1121 ;
  buffer buf_n1123( .i (n1122), .o (n1123) );
  assign n1124 = n987 & n989 ;
  buffer buf_n1125( .i (n1124), .o (n1125) );
  assign n1126 = n993 & n995 ;
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  assign n1129 = n1125 | n1128 ;
  assign n1130 = n1001 & n1003 ;
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  assign n1133 = n1129 | n1132 ;
  buffer buf_n1134( .i (n1133), .o (n1134) );
  assign n1135 = n1123 | n1134 ;
  buffer buf_n1136( .i (n1135), .o (n1136) );
  assign n1137 = n1012 | n1014 ;
  buffer buf_n1138( .i (n1137), .o (n1138) );
  assign n1139 = n1018 | n1020 ;
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  assign n1142 = n1138 & n1141 ;
  assign n1143 = n1026 | n1028 ;
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  assign n1146 = n1142 & n1145 ;
  buffer buf_n1147( .i (n1146), .o (n1147) );
  assign n1148 = n1035 & n1037 ;
  buffer buf_n1149( .i (n1148), .o (n1149) );
  assign n1150 = n1041 & n1043 ;
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  assign n1153 = n1149 | n1152 ;
  assign n1154 = n1049 & n1051 ;
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  assign n1157 = n1153 | n1156 ;
  buffer buf_n1158( .i (n1157), .o (n1158) );
  assign n1159 = n1147 | n1158 ;
  buffer buf_n1160( .i (n1159), .o (n1160) );
  assign n1161 = n1136 | n1160 ;
  buffer buf_n1162( .i (n1161), .o (n1162) );
  assign n1163 = n1112 | n1162 ;
  buffer buf_n1164( .i (n1163), .o (n1164) );
  assign n1165 = n1062 | n1164 ;
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  assign n1168 = ( n382 & n413 ) | ( n382 & n452 ) | ( n413 & n452 ) ;
  buffer buf_n1169( .i (n1168), .o (n1169) );
  assign n1170 = ( n789 & n820 ) | ( n789 & n859 ) | ( n820 & n859 ) ;
  buffer buf_n1171( .i (n1170), .o (n1171) );
  assign n1172 = n1169 | n1171 ;
  buffer buf_n1173( .i (n1172), .o (n1173) );
  assign n1174 = ( n878 & n893 ) | ( n878 & n908 ) | ( n893 & n908 ) ;
  buffer buf_n1175( .i (n1174), .o (n1175) );
  assign n1176 = ( n925 & n940 ) | ( n925 & n955 ) | ( n940 & n955 ) ;
  buffer buf_n1177( .i (n1176), .o (n1177) );
  assign n1178 = n1175 | n1177 ;
  buffer buf_n1179( .i (n1178), .o (n1179) );
  assign n1180 = n1173 | n1179 ;
  buffer buf_n1181( .i (n1180), .o (n1181) );
  assign n1182 = ( n968 & n975 ) | ( n968 & n982 ) | ( n975 & n982 ) ;
  buffer buf_n1183( .i (n1182), .o (n1183) );
  assign n1184 = ( n991 & n998 ) | ( n991 & n1005 ) | ( n998 & n1005 ) ;
  buffer buf_n1185( .i (n1184), .o (n1185) );
  assign n1186 = n1183 | n1185 ;
  buffer buf_n1187( .i (n1186), .o (n1187) );
  assign n1188 = ( n1016 & n1023 ) | ( n1016 & n1030 ) | ( n1023 & n1030 ) ;
  buffer buf_n1189( .i (n1188), .o (n1189) );
  assign n1190 = ( n1039 & n1046 ) | ( n1039 & n1053 ) | ( n1046 & n1053 ) ;
  buffer buf_n1191( .i (n1190), .o (n1191) );
  assign n1192 = n1189 | n1191 ;
  buffer buf_n1193( .i (n1192), .o (n1193) );
  assign n1194 = n1187 | n1193 ;
  buffer buf_n1195( .i (n1194), .o (n1195) );
  assign n1196 = n1181 | n1195 ;
  buffer buf_n1197( .i (n1196), .o (n1197) );
  assign n1198 = ( n1064 & n1067 ) | ( n1064 & n1070 ) | ( n1067 & n1070 ) ;
  buffer buf_n1199( .i (n1198), .o (n1199) );
  assign n1200 = ( n1075 & n1078 ) | ( n1075 & n1081 ) | ( n1078 & n1081 ) ;
  buffer buf_n1201( .i (n1200), .o (n1201) );
  assign n1202 = n1199 | n1201 ;
  buffer buf_n1203( .i (n1202), .o (n1203) );
  assign n1204 = ( n1088 & n1091 ) | ( n1088 & n1094 ) | ( n1091 & n1094 ) ;
  buffer buf_n1205( .i (n1204), .o (n1205) );
  assign n1206 = ( n1099 & n1102 ) | ( n1099 & n1105 ) | ( n1102 & n1105 ) ;
  buffer buf_n1207( .i (n1206), .o (n1207) );
  assign n1208 = n1205 | n1207 ;
  buffer buf_n1209( .i (n1208), .o (n1209) );
  assign n1210 = n1203 | n1209 ;
  buffer buf_n1211( .i (n1210), .o (n1211) );
  assign n1212 = ( n1114 & n1117 ) | ( n1114 & n1120 ) | ( n1117 & n1120 ) ;
  buffer buf_n1213( .i (n1212), .o (n1213) );
  assign n1214 = ( n1125 & n1128 ) | ( n1125 & n1131 ) | ( n1128 & n1131 ) ;
  buffer buf_n1215( .i (n1214), .o (n1215) );
  assign n1216 = n1213 | n1215 ;
  buffer buf_n1217( .i (n1216), .o (n1217) );
  assign n1218 = ( n1138 & n1141 ) | ( n1138 & n1144 ) | ( n1141 & n1144 ) ;
  buffer buf_n1219( .i (n1218), .o (n1219) );
  assign n1220 = ( n1149 & n1152 ) | ( n1149 & n1155 ) | ( n1152 & n1155 ) ;
  buffer buf_n1221( .i (n1220), .o (n1221) );
  assign n1222 = n1219 | n1221 ;
  buffer buf_n1223( .i (n1222), .o (n1223) );
  assign n1224 = n1217 | n1223 ;
  buffer buf_n1225( .i (n1224), .o (n1225) );
  assign n1226 = n1211 | n1225 ;
  buffer buf_n1227( .i (n1226), .o (n1227) );
  assign n1228 = n1197 | n1227 ;
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  assign n1231 = n382 | n413 ;
  assign n1232 = n453 | n1231 ;
  buffer buf_n1233( .i (n1232), .o (n1233) );
  assign n1234 = n789 & n820 ;
  assign n1235 = n860 & n1234 ;
  buffer buf_n1236( .i (n1235), .o (n1236) );
  assign n1237 = n1233 | n1236 ;
  buffer buf_n1238( .i (n1237), .o (n1238) );
  assign n1239 = n878 | n893 ;
  assign n1240 = n909 | n1239 ;
  buffer buf_n1241( .i (n1240), .o (n1241) );
  assign n1242 = n925 & n940 ;
  assign n1243 = n956 & n1242 ;
  buffer buf_n1244( .i (n1243), .o (n1244) );
  assign n1245 = n1241 | n1244 ;
  buffer buf_n1246( .i (n1245), .o (n1246) );
  assign n1247 = n1238 | n1246 ;
  buffer buf_n1248( .i (n1247), .o (n1248) );
  assign n1249 = n968 | n975 ;
  assign n1250 = n983 | n1249 ;
  buffer buf_n1251( .i (n1250), .o (n1251) );
  assign n1252 = n991 & n998 ;
  assign n1253 = n1006 & n1252 ;
  buffer buf_n1254( .i (n1253), .o (n1254) );
  assign n1255 = n1251 | n1254 ;
  buffer buf_n1256( .i (n1255), .o (n1256) );
  assign n1257 = n1016 | n1023 ;
  assign n1258 = n1031 | n1257 ;
  buffer buf_n1259( .i (n1258), .o (n1259) );
  assign n1260 = n1039 & n1046 ;
  assign n1261 = n1054 & n1260 ;
  buffer buf_n1262( .i (n1261), .o (n1262) );
  assign n1263 = n1259 | n1262 ;
  buffer buf_n1264( .i (n1263), .o (n1264) );
  assign n1265 = n1256 | n1264 ;
  buffer buf_n1266( .i (n1265), .o (n1266) );
  assign n1267 = n1248 | n1266 ;
  buffer buf_n1268( .i (n1267), .o (n1268) );
  assign n1269 = n1064 | n1067 ;
  assign n1270 = n1071 | n1269 ;
  buffer buf_n1271( .i (n1270), .o (n1271) );
  assign n1272 = n1075 & n1078 ;
  assign n1273 = n1082 & n1272 ;
  buffer buf_n1274( .i (n1273), .o (n1274) );
  assign n1275 = n1271 | n1274 ;
  buffer buf_n1276( .i (n1275), .o (n1276) );
  assign n1277 = n1088 | n1091 ;
  assign n1278 = n1095 | n1277 ;
  buffer buf_n1279( .i (n1278), .o (n1279) );
  assign n1280 = n1099 & n1102 ;
  assign n1281 = n1106 & n1280 ;
  buffer buf_n1282( .i (n1281), .o (n1282) );
  assign n1283 = n1279 | n1282 ;
  buffer buf_n1284( .i (n1283), .o (n1284) );
  assign n1285 = n1276 | n1284 ;
  buffer buf_n1286( .i (n1285), .o (n1286) );
  assign n1287 = n1114 | n1117 ;
  assign n1288 = n1121 | n1287 ;
  buffer buf_n1289( .i (n1288), .o (n1289) );
  assign n1290 = n1125 & n1128 ;
  assign n1291 = n1132 & n1290 ;
  buffer buf_n1292( .i (n1291), .o (n1292) );
  assign n1293 = n1289 | n1292 ;
  buffer buf_n1294( .i (n1293), .o (n1294) );
  assign n1295 = n1138 | n1141 ;
  assign n1296 = n1145 | n1295 ;
  buffer buf_n1297( .i (n1296), .o (n1297) );
  assign n1298 = n1149 & n1152 ;
  assign n1299 = n1156 & n1298 ;
  buffer buf_n1300( .i (n1299), .o (n1300) );
  assign n1301 = n1297 | n1300 ;
  buffer buf_n1302( .i (n1301), .o (n1302) );
  assign n1303 = n1294 | n1302 ;
  buffer buf_n1304( .i (n1303), .o (n1304) );
  assign n1305 = n1286 | n1304 ;
  buffer buf_n1306( .i (n1305), .o (n1306) );
  assign n1307 = n1268 | n1306 ;
  buffer buf_n1308( .i (n1307), .o (n1308) );
  assign n1309 = n1230 | n1308 ;
  assign n1310 = n1167 | n1309 ;
  assign n1311 = n1062 & n1164 ;
  buffer buf_n1312( .i (n1311), .o (n1312) );
  assign n1314 = n1197 & n1227 ;
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  assign n1317 = n1268 & n1306 ;
  buffer buf_n1318( .i (n1317), .o (n1318) );
  assign n1319 = ( n1312 & n1316 ) | ( n1312 & n1318 ) | ( n1316 & n1318 ) ;
  buffer buf_n1320( .i (n1319), .o (n1320) );
  assign n1321 = n962 & n1060 ;
  buffer buf_n1322( .i (n1321), .o (n1322) );
  assign n1323 = n1112 & n1162 ;
  buffer buf_n1324( .i (n1323), .o (n1324) );
  assign n1325 = n1322 | n1324 ;
  buffer buf_n1326( .i (n1325), .o (n1326) );
  assign n1328 = n1181 & n1195 ;
  buffer buf_n1329( .i (n1328), .o (n1329) );
  assign n1330 = n1211 & n1225 ;
  buffer buf_n1331( .i (n1330), .o (n1331) );
  assign n1332 = n1329 | n1331 ;
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  assign n1335 = n1248 & n1266 ;
  buffer buf_n1336( .i (n1335), .o (n1336) );
  assign n1337 = n1286 & n1304 ;
  buffer buf_n1338( .i (n1337), .o (n1338) );
  assign n1339 = n1336 | n1338 ;
  buffer buf_n1340( .i (n1339), .o (n1340) );
  assign n1341 = ( n1326 & n1334 ) | ( n1326 & n1340 ) | ( n1334 & n1340 ) ;
  buffer buf_n1342( .i (n1341), .o (n1342) );
  assign n1343 = n455 & n862 ;
  buffer buf_n1344( .i (n1343), .o (n1344) );
  assign n1345 = n911 & n958 ;
  buffer buf_n1346( .i (n1345), .o (n1346) );
  assign n1347 = n1344 & n1346 ;
  buffer buf_n1348( .i (n1347), .o (n1348) );
  assign n1349 = n985 & n1008 ;
  buffer buf_n1350( .i (n1349), .o (n1350) );
  assign n1351 = n1033 & n1056 ;
  buffer buf_n1352( .i (n1351), .o (n1352) );
  assign n1353 = n1350 & n1352 ;
  buffer buf_n1354( .i (n1353), .o (n1354) );
  assign n1355 = n1348 | n1354 ;
  buffer buf_n1356( .i (n1355), .o (n1356) );
  assign n1357 = n1073 & n1084 ;
  buffer buf_n1358( .i (n1357), .o (n1358) );
  assign n1359 = n1097 & n1108 ;
  buffer buf_n1360( .i (n1359), .o (n1360) );
  assign n1361 = n1358 & n1360 ;
  buffer buf_n1362( .i (n1361), .o (n1362) );
  assign n1363 = n1123 & n1134 ;
  buffer buf_n1364( .i (n1363), .o (n1364) );
  assign n1365 = n1147 & n1158 ;
  buffer buf_n1366( .i (n1365), .o (n1366) );
  assign n1367 = n1364 & n1366 ;
  buffer buf_n1368( .i (n1367), .o (n1368) );
  assign n1369 = n1362 | n1368 ;
  buffer buf_n1370( .i (n1369), .o (n1370) );
  assign n1371 = n1356 | n1370 ;
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  assign n1374 = n1169 & n1171 ;
  buffer buf_n1375( .i (n1374), .o (n1375) );
  assign n1376 = n1175 & n1177 ;
  buffer buf_n1377( .i (n1376), .o (n1377) );
  assign n1378 = n1375 & n1377 ;
  buffer buf_n1379( .i (n1378), .o (n1379) );
  assign n1380 = n1183 & n1185 ;
  buffer buf_n1381( .i (n1380), .o (n1381) );
  assign n1382 = n1189 & n1191 ;
  buffer buf_n1383( .i (n1382), .o (n1383) );
  assign n1384 = n1381 & n1383 ;
  buffer buf_n1385( .i (n1384), .o (n1385) );
  assign n1386 = n1379 | n1385 ;
  buffer buf_n1387( .i (n1386), .o (n1387) );
  assign n1388 = n1199 & n1201 ;
  buffer buf_n1389( .i (n1388), .o (n1389) );
  assign n1390 = n1205 & n1207 ;
  buffer buf_n1391( .i (n1390), .o (n1391) );
  assign n1392 = n1389 & n1391 ;
  buffer buf_n1393( .i (n1392), .o (n1393) );
  assign n1394 = n1213 & n1215 ;
  buffer buf_n1395( .i (n1394), .o (n1395) );
  assign n1396 = n1219 & n1221 ;
  buffer buf_n1397( .i (n1396), .o (n1397) );
  assign n1398 = n1395 & n1397 ;
  buffer buf_n1399( .i (n1398), .o (n1399) );
  assign n1400 = n1393 | n1399 ;
  buffer buf_n1401( .i (n1400), .o (n1401) );
  assign n1402 = n1387 | n1401 ;
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  assign n1405 = n1233 & n1236 ;
  buffer buf_n1406( .i (n1405), .o (n1406) );
  assign n1407 = n1241 & n1244 ;
  buffer buf_n1408( .i (n1407), .o (n1408) );
  assign n1409 = n1406 & n1408 ;
  buffer buf_n1410( .i (n1409), .o (n1410) );
  assign n1411 = n1251 & n1254 ;
  buffer buf_n1412( .i (n1411), .o (n1412) );
  assign n1413 = n1259 & n1262 ;
  buffer buf_n1414( .i (n1413), .o (n1414) );
  assign n1415 = n1412 & n1414 ;
  buffer buf_n1416( .i (n1415), .o (n1416) );
  assign n1417 = n1410 | n1416 ;
  buffer buf_n1418( .i (n1417), .o (n1418) );
  assign n1419 = n1271 & n1274 ;
  buffer buf_n1420( .i (n1419), .o (n1420) );
  assign n1421 = n1279 & n1282 ;
  buffer buf_n1422( .i (n1421), .o (n1422) );
  assign n1423 = n1420 & n1422 ;
  buffer buf_n1424( .i (n1423), .o (n1424) );
  assign n1425 = n1289 & n1292 ;
  buffer buf_n1426( .i (n1425), .o (n1426) );
  assign n1427 = n1297 & n1300 ;
  buffer buf_n1428( .i (n1427), .o (n1428) );
  assign n1429 = n1426 & n1428 ;
  buffer buf_n1430( .i (n1429), .o (n1430) );
  assign n1431 = n1424 | n1430 ;
  buffer buf_n1432( .i (n1431), .o (n1432) );
  assign n1433 = n1418 | n1432 ;
  buffer buf_n1434( .i (n1433), .o (n1434) );
  assign n1435 = n1404 | n1434 ;
  assign n1436 = n1373 | n1435 ;
  assign n1437 = n1356 & n1370 ;
  buffer buf_n1438( .i (n1437), .o (n1438) );
  assign n1440 = n1387 & n1401 ;
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  assign n1443 = n1418 & n1432 ;
  buffer buf_n1444( .i (n1443), .o (n1444) );
  assign n1445 = ( n1438 & n1442 ) | ( n1438 & n1444 ) | ( n1442 & n1444 ) ;
  buffer buf_n1446( .i (n1445), .o (n1446) );
  assign n1447 = n1348 & n1354 ;
  buffer buf_n1448( .i (n1447), .o (n1448) );
  assign n1449 = n1362 & n1368 ;
  buffer buf_n1450( .i (n1449), .o (n1450) );
  assign n1451 = n1448 | n1450 ;
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  assign n1454 = n1379 & n1385 ;
  buffer buf_n1455( .i (n1454), .o (n1455) );
  assign n1456 = n1393 & n1399 ;
  buffer buf_n1457( .i (n1456), .o (n1457) );
  assign n1458 = n1455 | n1457 ;
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  assign n1461 = n1410 & n1416 ;
  buffer buf_n1462( .i (n1461), .o (n1462) );
  assign n1463 = n1424 & n1430 ;
  buffer buf_n1464( .i (n1463), .o (n1464) );
  assign n1465 = n1462 | n1464 ;
  buffer buf_n1466( .i (n1465), .o (n1466) );
  assign n1467 = n1460 | n1466 ;
  assign n1468 = n1453 | n1467 ;
  assign n1469 = n864 & n960 ;
  buffer buf_n1470( .i (n1469), .o (n1470) );
  assign n1471 = n1010 & n1058 ;
  buffer buf_n1472( .i (n1471), .o (n1472) );
  assign n1473 = n1470 | n1472 ;
  buffer buf_n1474( .i (n1473), .o (n1474) );
  assign n1475 = n1086 & n1110 ;
  buffer buf_n1476( .i (n1475), .o (n1476) );
  assign n1477 = n1136 & n1160 ;
  buffer buf_n1478( .i (n1477), .o (n1478) );
  assign n1479 = n1476 | n1478 ;
  buffer buf_n1480( .i (n1479), .o (n1480) );
  assign n1481 = n1474 & n1480 ;
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  assign n1484 = n1173 & n1179 ;
  buffer buf_n1485( .i (n1484), .o (n1485) );
  assign n1486 = n1187 & n1193 ;
  buffer buf_n1487( .i (n1486), .o (n1487) );
  assign n1488 = n1485 | n1487 ;
  buffer buf_n1489( .i (n1488), .o (n1489) );
  assign n1490 = n1203 & n1209 ;
  buffer buf_n1491( .i (n1490), .o (n1491) );
  assign n1492 = n1217 & n1223 ;
  buffer buf_n1493( .i (n1492), .o (n1493) );
  assign n1494 = n1491 | n1493 ;
  buffer buf_n1495( .i (n1494), .o (n1495) );
  assign n1496 = n1489 & n1495 ;
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  assign n1499 = n1238 & n1246 ;
  buffer buf_n1500( .i (n1499), .o (n1500) );
  assign n1501 = n1256 & n1264 ;
  buffer buf_n1502( .i (n1501), .o (n1502) );
  assign n1503 = n1500 | n1502 ;
  buffer buf_n1504( .i (n1503), .o (n1504) );
  assign n1505 = n1276 & n1284 ;
  buffer buf_n1506( .i (n1505), .o (n1506) );
  assign n1507 = n1294 & n1302 ;
  buffer buf_n1508( .i (n1507), .o (n1508) );
  assign n1509 = n1506 | n1508 ;
  buffer buf_n1510( .i (n1509), .o (n1510) );
  assign n1511 = n1504 & n1510 ;
  buffer buf_n1512( .i (n1511), .o (n1512) );
  assign n1513 = n1498 | n1512 ;
  assign n1514 = n1483 | n1513 ;
  assign n1515 = n1344 | n1346 ;
  buffer buf_n1516( .i (n1515), .o (n1516) );
  assign n1517 = n1350 | n1352 ;
  buffer buf_n1518( .i (n1517), .o (n1518) );
  assign n1519 = n1516 & n1518 ;
  buffer buf_n1520( .i (n1519), .o (n1520) );
  assign n1521 = n1358 | n1360 ;
  buffer buf_n1522( .i (n1521), .o (n1522) );
  assign n1523 = n1364 | n1366 ;
  buffer buf_n1524( .i (n1523), .o (n1524) );
  assign n1525 = n1522 & n1524 ;
  buffer buf_n1526( .i (n1525), .o (n1526) );
  assign n1527 = n1520 | n1526 ;
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  assign n1530 = n1375 | n1377 ;
  buffer buf_n1531( .i (n1530), .o (n1531) );
  assign n1532 = n1381 | n1383 ;
  buffer buf_n1533( .i (n1532), .o (n1533) );
  assign n1534 = n1531 & n1533 ;
  buffer buf_n1535( .i (n1534), .o (n1535) );
  assign n1536 = n1389 | n1391 ;
  buffer buf_n1537( .i (n1536), .o (n1537) );
  assign n1538 = n1395 | n1397 ;
  buffer buf_n1539( .i (n1538), .o (n1539) );
  assign n1540 = n1537 & n1539 ;
  buffer buf_n1541( .i (n1540), .o (n1541) );
  assign n1542 = n1535 | n1541 ;
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  assign n1545 = n1406 | n1408 ;
  buffer buf_n1546( .i (n1545), .o (n1546) );
  assign n1547 = n1412 | n1414 ;
  buffer buf_n1548( .i (n1547), .o (n1548) );
  assign n1549 = n1546 & n1548 ;
  buffer buf_n1550( .i (n1549), .o (n1550) );
  assign n1551 = n1420 | n1422 ;
  buffer buf_n1552( .i (n1551), .o (n1552) );
  assign n1553 = n1426 | n1428 ;
  buffer buf_n1554( .i (n1553), .o (n1554) );
  assign n1555 = n1552 & n1554 ;
  buffer buf_n1556( .i (n1555), .o (n1556) );
  assign n1557 = n1550 | n1556 ;
  buffer buf_n1558( .i (n1557), .o (n1558) );
  assign n1559 = n1544 | n1558 ;
  assign n1560 = n1529 | n1559 ;
  assign n1561 = n1470 & n1472 ;
  buffer buf_n1562( .i (n1561), .o (n1562) );
  assign n1563 = n1476 & n1478 ;
  buffer buf_n1564( .i (n1563), .o (n1564) );
  assign n1565 = n1562 | n1564 ;
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  assign n1568 = n1485 & n1487 ;
  buffer buf_n1569( .i (n1568), .o (n1569) );
  assign n1570 = n1491 & n1493 ;
  buffer buf_n1571( .i (n1570), .o (n1571) );
  assign n1572 = n1569 | n1571 ;
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  assign n1575 = n1500 & n1502 ;
  buffer buf_n1576( .i (n1575), .o (n1576) );
  assign n1577 = n1506 & n1508 ;
  buffer buf_n1578( .i (n1577), .o (n1578) );
  assign n1579 = n1576 | n1578 ;
  buffer buf_n1580( .i (n1579), .o (n1580) );
  assign n1581 = n1574 | n1580 ;
  assign n1582 = n1567 | n1581 ;
  assign n1583 = n1562 & n1564 ;
  buffer buf_n1584( .i (n1583), .o (n1584) );
  assign n1586 = n1569 & n1571 ;
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  assign n1589 = n1576 & n1578 ;
  buffer buf_n1590( .i (n1589), .o (n1590) );
  assign n1591 = ( n1584 & n1588 ) | ( n1584 & n1590 ) | ( n1588 & n1590 ) ;
  buffer buf_n1592( .i (n1591), .o (n1592) );
  assign n1593 = n1520 & n1526 ;
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  assign n1596 = n1535 & n1541 ;
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  assign n1599 = n1550 & n1556 ;
  buffer buf_n1600( .i (n1599), .o (n1600) );
  assign n1601 = n1598 & n1600 ;
  assign n1602 = n1595 & n1601 ;
  assign n1603 = ( n1528 & n1544 ) | ( n1528 & n1558 ) | ( n1544 & n1558 ) ;
  buffer buf_n1604( .i (n1603), .o (n1604) );
  assign n1605 = n1448 & n1450 ;
  buffer buf_n1606( .i (n1605), .o (n1606) );
  assign n1608 = n1455 & n1457 ;
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  assign n1611 = n1462 & n1464 ;
  buffer buf_n1612( .i (n1611), .o (n1612) );
  assign n1613 = ( n1606 & n1610 ) | ( n1606 & n1612 ) | ( n1610 & n1612 ) ;
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  assign n1615 = n1316 & n1318 ;
  assign n1616 = n1313 & n1615 ;
  buffer buf_n1607( .i (n1606), .o (n1607) );
  assign n1617 = n1610 & n1612 ;
  assign n1618 = n1607 & n1617 ;
  assign n1619 = ( n1566 & n1574 ) | ( n1566 & n1580 ) | ( n1574 & n1580 ) ;
  buffer buf_n1620( .i (n1619), .o (n1620) );
  assign n1621 = n1404 & n1434 ;
  assign n1622 = n1373 & n1621 ;
  assign n1623 = n1322 & n1324 ;
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  assign n1626 = n1329 & n1331 ;
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  assign n1629 = n1336 & n1338 ;
  buffer buf_n1630( .i (n1629), .o (n1630) );
  assign n1631 = n1628 & n1630 ;
  assign n1632 = n1625 & n1631 ;
  assign n1633 = n1610 | n1612 ;
  assign n1634 = n1607 | n1633 ;
  assign n1635 = n1516 | n1518 ;
  buffer buf_n1636( .i (n1635), .o (n1636) );
  assign n1637 = n1522 | n1524 ;
  buffer buf_n1638( .i (n1637), .o (n1638) );
  assign n1639 = n1636 & n1638 ;
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  assign n1642 = n1531 | n1533 ;
  buffer buf_n1643( .i (n1642), .o (n1643) );
  assign n1644 = n1537 | n1539 ;
  buffer buf_n1645( .i (n1644), .o (n1645) );
  assign n1646 = n1643 & n1645 ;
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  assign n1649 = n1546 | n1548 ;
  buffer buf_n1650( .i (n1649), .o (n1650) );
  assign n1651 = n1552 | n1554 ;
  buffer buf_n1652( .i (n1651), .o (n1652) );
  assign n1653 = n1650 & n1652 ;
  buffer buf_n1654( .i (n1653), .o (n1654) );
  assign n1655 = n1648 | n1654 ;
  assign n1656 = n1641 | n1655 ;
  buffer buf_n1327( .i (n1326), .o (n1327) );
  assign n1657 = n1334 | n1340 ;
  assign n1658 = n1327 | n1657 ;
  assign n1659 = n1474 | n1480 ;
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  assign n1662 = n1489 | n1495 ;
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  assign n1665 = n1504 | n1510 ;
  buffer buf_n1666( .i (n1665), .o (n1666) );
  assign n1667 = n1664 & n1666 ;
  assign n1668 = n1661 & n1667 ;
  assign n1669 = ( n1482 & n1498 ) | ( n1482 & n1512 ) | ( n1498 & n1512 ) ;
  buffer buf_n1670( .i (n1669), .o (n1670) );
  assign n1671 = ( n1660 & n1664 ) | ( n1660 & n1666 ) | ( n1664 & n1666 ) ;
  buffer buf_n1672( .i (n1671), .o (n1672) );
  assign n1673 = ( n1594 & n1598 ) | ( n1594 & n1600 ) | ( n1598 & n1600 ) ;
  buffer buf_n1674( .i (n1673), .o (n1674) );
  assign n1675 = n1636 | n1638 ;
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  assign n1678 = n1643 | n1645 ;
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  assign n1681 = n1650 | n1652 ;
  buffer buf_n1682( .i (n1681), .o (n1682) );
  assign n1683 = n1680 & n1682 ;
  assign n1684 = n1677 & n1683 ;
  assign n1685 = n1664 | n1666 ;
  assign n1686 = n1661 | n1685 ;
  assign n1687 = n1334 & n1340 ;
  assign n1688 = n1327 & n1687 ;
  assign n1689 = n1574 & n1580 ;
  assign n1690 = n1567 & n1689 ;
  assign n1691 = ( n1166 & n1230 ) | ( n1166 & n1308 ) | ( n1230 & n1308 ) ;
  buffer buf_n1692( .i (n1691), .o (n1692) );
  assign n1693 = ( n1452 & n1460 ) | ( n1452 & n1466 ) | ( n1460 & n1466 ) ;
  buffer buf_n1694( .i (n1693), .o (n1694) );
  assign n1695 = n1598 | n1600 ;
  assign n1696 = n1595 | n1695 ;
  assign n1697 = ( n1624 & n1628 ) | ( n1624 & n1630 ) | ( n1628 & n1630 ) ;
  buffer buf_n1698( .i (n1697), .o (n1698) );
  assign n1699 = ( n1676 & n1680 ) | ( n1676 & n1682 ) | ( n1680 & n1682 ) ;
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  assign n1701 = n1442 & n1444 ;
  assign n1702 = n1439 & n1701 ;
  assign n1703 = n1628 | n1630 ;
  assign n1704 = n1625 | n1703 ;
  assign n1705 = n1648 & n1654 ;
  assign n1706 = n1641 & n1705 ;
  assign n1707 = n1544 & n1558 ;
  assign n1708 = n1529 & n1707 ;
  assign n1709 = n1498 & n1512 ;
  assign n1710 = n1483 & n1709 ;
  assign n1711 = n1442 | n1444 ;
  assign n1712 = n1439 | n1711 ;
  buffer buf_n1585( .i (n1584), .o (n1585) );
  assign n1713 = n1588 | n1590 ;
  assign n1714 = n1585 | n1713 ;
  assign n1715 = n1588 & n1590 ;
  assign n1716 = n1585 & n1715 ;
  assign n1717 = ( n1640 & n1648 ) | ( n1640 & n1654 ) | ( n1648 & n1654 ) ;
  buffer buf_n1718( .i (n1717), .o (n1718) );
  assign n1719 = n1680 | n1682 ;
  assign n1720 = n1677 | n1719 ;
  assign n1721 = ( n1372 & n1404 ) | ( n1372 & n1434 ) | ( n1404 & n1434 ) ;
  buffer buf_n1722( .i (n1721), .o (n1722) );
  assign n1723 = n1460 & n1466 ;
  assign n1724 = n1453 & n1723 ;
  assign n1725 = n1230 & n1308 ;
  assign n1726 = n1167 & n1725 ;
  assign n1727 = n1316 | n1318 ;
  assign n1728 = n1313 | n1727 ;
  assign b_47_ = n1310 ;
  assign b_43_ = n1320 ;
  assign b_40_ = n1342 ;
  assign b_11_ = n1436 ;
  assign b_7_ = n1446 ;
  assign b_5_ = n1468 ;
  assign b_32_ = n1514 ;
  assign b_17_ = n1560 ;
  assign b_29_ = n1582 ;
  assign b_25_ = n1592 ;
  assign b_12_ = n1602 ;
  assign b_16_ = n1604 ;
  assign b_1_ = n1614 ;
  assign b_42_ = n1616 ;
  assign b_0_ = n1618 ;
  assign b_28_ = n1620 ;
  assign b_9_ = n1622 ;
  assign b_36_ = n1632 ;
  assign b_2_ = n1634 ;
  assign b_20_ = n1656 ;
  assign b_41_ = n1658 ;
  assign b_33_ = n1668 ;
  assign b_31_ = n1670 ;
  assign b_34_ = n1672 ;
  assign b_13_ = n1674 ;
  assign b_21_ = n1684 ;
  assign b_35_ = n1686 ;
  assign b_39_ = n1688 ;
  assign b_27_ = n1690 ;
  assign b_46_ = n1692 ;
  assign b_4_ = n1694 ;
  assign b_14_ = n1696 ;
  assign b_37_ = n1698 ;
  assign b_22_ = n1700 ;
  assign b_6_ = n1702 ;
  assign b_38_ = n1704 ;
  assign b_18_ = n1706 ;
  assign b_15_ = n1708 ;
  assign b_30_ = n1710 ;
  assign b_8_ = n1712 ;
  assign b_26_ = n1714 ;
  assign b_24_ = n1716 ;
  assign b_19_ = n1718 ;
  assign b_23_ = n1720 ;
  assign b_10_ = n1722 ;
  assign b_3_ = n1724 ;
  assign b_45_ = n1726 ;
  assign b_44_ = n1728 ;
endmodule
