module top( a_11_ , a_18_ , a_15_ , a_3_ , a_9_ , a_6_ , a_28_ , a_7_ , a_25_ , a_29_ , a_22_ , a_26_ , a_1_ , a_8_ , a_16_ , a_10_ , a_30_ , a_12_ , a_24_ , a_5_ , a_0_ , a_17_ , a_4_ , a_14_ , a_20_ , a_27_ , a_23_ , a_13_ , a_31_ , a_2_ , a_19_ , a_21_ , b_9_ , b_1_ , b_17_ , b_11_ , b_31_ , b_26_ , b_29_ , b_24_ , b_23_ , b_8_ , b_4_ , b_25_ , b_7_ , b_5_ , b_18_ , b_12_ , b_16_ , b_22_ , b_14_ , b_20_ , b_15_ , b_3_ , b_30_ , b_27_ , b_21_ , b_19_ , b_13_ , b_6_ , b_0_ , b_10_ , b_28_ , b_2_ );
  input a_11_ , a_18_ , a_15_ , a_3_ , a_9_ , a_6_ , a_28_ , a_7_ , a_25_ , a_29_ , a_22_ , a_26_ , a_1_ , a_8_ , a_16_ , a_10_ , a_30_ , a_12_ , a_24_ , a_5_ , a_0_ , a_17_ , a_4_ , a_14_ , a_20_ , a_27_ , a_23_ , a_13_ , a_31_ , a_2_ , a_19_ , a_21_ ;
  output b_9_ , b_1_ , b_17_ , b_11_ , b_31_ , b_26_ , b_29_ , b_24_ , b_23_ , b_8_ , b_4_ , b_25_ , b_7_ , b_5_ , b_18_ , b_12_ , b_16_ , b_22_ , b_14_ , b_20_ , b_15_ , b_3_ , b_30_ , b_27_ , b_21_ , b_19_ , b_13_ , b_6_ , b_0_ , b_10_ , b_28_ , b_2_ ;
  wire n65 , n67 , n69 , n71 , n73 , n75 , n77 , n79 , n81 , n83 , n85 , n87 , n89 , n91 , n93 , n95 , n97 , n99 , n101 , n103 , n105 , n107 , n109 , n111 , n113 , n115 , n117 , n119 , n121 , n123 , n125 , n127 , n129 , n131 , n133 , n135 , n137 , n139 , n141 , n143 , n145 , n147 , n149 , n151 , n153 , n155 , n157 , n159 , n161 , n163 , n165 , n167 , n169 , n171 , n173 , n175 , n177 , n179 , n181 , n183 , n185 , n187 , n189 , n191 , n193 , n195 , n197 , n199 , n201 , n203 , n205 , n207 , n209 , n211 , n213 , n215 , n217 , n219 , n221 , n223 , n225 , n227 , n229 , n231 , n233 , n235 , n237 , n239 , n241 , n243 , n245 , n247 , n249 , n251 , n253 , n255 , n257 , n259 , n261 , n263 , n265 , n267 , n269 , n271 , n273 , n275 , n277 , n279 , n281 , n283 , n285 , n287 , n289 , n291 , n293 , n295 , n297 , n299 , n301 , n303 , n305 , n307 , n309 , n311 , n313 , n315 , n317 , n319 , n321 , n323 , n325 , n327 , n329 , n331 , n333 , n335 , n337 , n339 , n341 , n343 , n345 , n347 , n349 , n351 , n353 , n355 , n357 , n359 , n361 , n363 , n365 , n367 , n369 , n371 , n373 , n375 , n377 , n379 , n381 , n383 , n385 , n387 , n389 , n391 , n393 , n395 , n397 , n399 , n401 , n403 , n405 , n407 , n409 , n411 , n413 , n415 , n417 , n419 , n421 , n423 , n425 , n427 , n429 , n431 , n433 , n435 , n437 , n439 , n441 , n443 , n445 , n447 , n449 , n451 , n453 , n455 , n457 , n459 , n461 , n463 , n465 , n467 , n469 , n471 , n473 , n475 , n477 , n479 , n481 , n483 , n485 , n487 , n489 , n491 , n493 , n495 , n497 , n499 , n501 , n503 , n505 , n507 , n509 , n511 , n513 , n515 , n517 , n519 , n521 , n523 , n525 , n527 , n529 , n531 , n533 , n535 , n537 , n539 , n541 , n543 , n545 , n547 , n549 , n551 , n553 , n555 , n557 , n559 , n561 , n563 , n565 , n567 , n569 , n571 , n573 , n575 , n577 , n579 , n581 , n583 , n585 , n587 , n589 , n591 , n593 , n595 , n597 , n599 , n601 , n603 , n605 , n607 , n609 , n611 , n613 , n615 , n617 , n619 , n621 , n623 , n625 , n627 , n629 , n631 , n633 , n635 , n637 , n639 , n641 , n643 , n645 , n647 , n649 , n651 , n653 , n655 , n657 , n659 , n661 , n663 , n665 , n667 , n669 , n671 , n673 , n675 , n677 , n679 , n681 , n683 , n685 , n687 , n689 , n691 , n693 , n695 , n697 , n699 , n701 , n703 , n705 , n707 , n709 , n711 , n713 , n715 , n717 , n719 , n721 , n723 , n725 , n727 , n729 , n731 , n733 , n735 , n737 , n739 , n741 , n743 , n745 , n747 , n749 , n751 , n753 , n755 , n757 , n759 , n761 , n763 , n765 , n766 , n768 , n770 , n772 , n774 , n776 , n778 , n780 , n782 , n784 , n786 , n788 , n790 , n792 , n794 , n795 , n797 , n799 , n801 , n803 , n805 , n807 , n809 , n811 , n813 , n815 , n817 , n819 , n821 , n823 , n825 , n827 , n829 , n831 , n833 , n835 , n837 , n839 , n841 , n843 , n845 , n847 , n849 , n851 , n853 , n855 , n856 , n858 , n860 , n861 , n863 , n865 , n867 , n869 , n871 , n873 , n875 , n877 , n879 , n881 , n883 , n885 , n887 , n889 , n890 , n892 , n894 , n896 , n898 , n900 , n902 , n903 , n905 , n907 , n908 , n910 , n912 , n913 , n915 , n917 , n919 , n921 , n923 , n925 , n926 , n927 , n929 , n931 , n933 , n935 , n937 , n939 , n940 , n941 , n943 , n945 , n946 , n947 , n949 , n951 , n952 , n954 , n956 , n958 , n960 , n962 , n964 , n965 , n966 , n967 , n969 , n971 , n972 , n974 , n976 , n977 , n978 , n980 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 ;
  buffer buf_n35( .i (a_15_), .o (n35) );
  buffer buf_n56( .i (a_14_), .o (n56) );
  assign n65 = n35 | n56 ;
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n50( .i (a_12_), .o (n50) );
  buffer buf_n60( .i (a_13_), .o (n60) );
  assign n67 = n50 & n60 ;
  buffer buf_n68( .i (n67), .o (n68) );
  assign n69 = n66 & n68 ;
  buffer buf_n70( .i (n69), .o (n70) );
  assign n71 = n35 & n56 ;
  buffer buf_n72( .i (n71), .o (n72) );
  assign n73 = n50 | n60 ;
  buffer buf_n74( .i (n73), .o (n74) );
  assign n75 = n72 & n74 ;
  buffer buf_n76( .i (n75), .o (n76) );
  assign n77 = n70 | n76 ;
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n33( .i (a_11_), .o (n33) );
  buffer buf_n48( .i (a_10_), .o (n48) );
  assign n79 = n33 | n48 ;
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n37( .i (a_9_), .o (n37) );
  buffer buf_n46( .i (a_8_), .o (n46) );
  assign n81 = n37 & n46 ;
  buffer buf_n82( .i (n81), .o (n82) );
  assign n83 = n80 | n82 ;
  buffer buf_n84( .i (n83), .o (n84) );
  assign n85 = n33 & n48 ;
  buffer buf_n86( .i (n85), .o (n86) );
  assign n87 = n37 | n46 ;
  buffer buf_n88( .i (n87), .o (n88) );
  assign n89 = n86 | n88 ;
  buffer buf_n90( .i (n89), .o (n90) );
  assign n91 = n84 & n90 ;
  buffer buf_n92( .i (n91), .o (n92) );
  assign n93 = n78 & n92 ;
  buffer buf_n94( .i (n93), .o (n94) );
  assign n95 = n66 | n68 ;
  buffer buf_n96( .i (n95), .o (n96) );
  assign n97 = n72 | n74 ;
  buffer buf_n98( .i (n97), .o (n98) );
  assign n99 = n96 | n98 ;
  buffer buf_n100( .i (n99), .o (n100) );
  assign n101 = n80 & n82 ;
  buffer buf_n102( .i (n101), .o (n102) );
  assign n103 = n86 & n88 ;
  buffer buf_n104( .i (n103), .o (n104) );
  assign n105 = n102 & n104 ;
  buffer buf_n106( .i (n105), .o (n106) );
  assign n107 = n100 & n106 ;
  buffer buf_n108( .i (n107), .o (n108) );
  assign n109 = n94 & n108 ;
  buffer buf_n110( .i (n109), .o (n110) );
  assign n111 = n70 & n76 ;
  buffer buf_n112( .i (n111), .o (n112) );
  assign n113 = n84 | n90 ;
  buffer buf_n114( .i (n113), .o (n114) );
  assign n115 = n112 & n114 ;
  buffer buf_n116( .i (n115), .o (n116) );
  assign n117 = n96 & n98 ;
  buffer buf_n118( .i (n117), .o (n118) );
  assign n119 = n102 | n104 ;
  buffer buf_n120( .i (n119), .o (n120) );
  assign n121 = n118 & n120 ;
  buffer buf_n122( .i (n121), .o (n122) );
  assign n123 = n116 & n122 ;
  buffer buf_n124( .i (n123), .o (n124) );
  assign n125 = n110 | n124 ;
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n36( .i (a_3_), .o (n36) );
  buffer buf_n62( .i (a_2_), .o (n62) );
  assign n127 = n36 | n62 ;
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n45( .i (a_1_), .o (n45) );
  buffer buf_n53( .i (a_0_), .o (n53) );
  assign n129 = n45 & n53 ;
  buffer buf_n130( .i (n129), .o (n130) );
  assign n131 = n128 | n130 ;
  buffer buf_n132( .i (n131), .o (n132) );
  assign n133 = n36 & n62 ;
  buffer buf_n134( .i (n133), .o (n134) );
  assign n135 = n45 | n53 ;
  buffer buf_n136( .i (n135), .o (n136) );
  assign n137 = n134 | n136 ;
  buffer buf_n138( .i (n137), .o (n138) );
  assign n139 = n132 | n138 ;
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n38( .i (a_6_), .o (n38) );
  buffer buf_n40( .i (a_7_), .o (n40) );
  assign n141 = n38 | n40 ;
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n52( .i (a_5_), .o (n52) );
  buffer buf_n55( .i (a_4_), .o (n55) );
  assign n143 = n52 & n55 ;
  buffer buf_n144( .i (n143), .o (n144) );
  assign n145 = n142 & n144 ;
  buffer buf_n146( .i (n145), .o (n146) );
  assign n147 = n38 & n40 ;
  buffer buf_n148( .i (n147), .o (n148) );
  assign n149 = n52 | n55 ;
  buffer buf_n150( .i (n149), .o (n150) );
  assign n151 = n148 & n150 ;
  buffer buf_n152( .i (n151), .o (n152) );
  assign n153 = n146 & n152 ;
  buffer buf_n154( .i (n153), .o (n154) );
  assign n155 = n140 | n154 ;
  buffer buf_n156( .i (n155), .o (n156) );
  assign n157 = n128 & n130 ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n159 = n134 & n136 ;
  buffer buf_n160( .i (n159), .o (n160) );
  assign n161 = n158 | n160 ;
  buffer buf_n162( .i (n161), .o (n162) );
  assign n163 = n142 | n144 ;
  buffer buf_n164( .i (n163), .o (n164) );
  assign n165 = n148 | n150 ;
  buffer buf_n166( .i (n165), .o (n166) );
  assign n167 = n164 & n166 ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = n162 | n168 ;
  buffer buf_n170( .i (n169), .o (n170) );
  assign n171 = n156 | n170 ;
  buffer buf_n172( .i (n171), .o (n172) );
  assign n173 = n158 & n160 ;
  buffer buf_n174( .i (n173), .o (n174) );
  assign n175 = n164 | n166 ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n177 = n174 | n176 ;
  buffer buf_n178( .i (n177), .o (n178) );
  assign n179 = n132 & n138 ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = n146 | n152 ;
  buffer buf_n182( .i (n181), .o (n182) );
  assign n183 = n180 | n182 ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n185 = n178 | n184 ;
  buffer buf_n186( .i (n185), .o (n186) );
  assign n187 = n172 & n186 ;
  buffer buf_n188( .i (n187), .o (n188) );
  assign n189 = n126 | n188 ;
  buffer buf_n190( .i (n189), .o (n190) );
  assign n191 = n78 | n92 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = n100 | n106 ;
  buffer buf_n194( .i (n193), .o (n194) );
  assign n195 = n192 & n194 ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n197 = n112 | n114 ;
  buffer buf_n198( .i (n197), .o (n198) );
  assign n199 = n118 | n120 ;
  buffer buf_n200( .i (n199), .o (n200) );
  assign n201 = n198 & n200 ;
  buffer buf_n202( .i (n201), .o (n202) );
  assign n203 = n196 | n202 ;
  buffer buf_n204( .i (n203), .o (n204) );
  assign n205 = n140 & n154 ;
  buffer buf_n206( .i (n205), .o (n206) );
  assign n207 = n162 & n168 ;
  buffer buf_n208( .i (n207), .o (n208) );
  assign n209 = n206 | n208 ;
  buffer buf_n210( .i (n209), .o (n210) );
  assign n211 = n174 & n176 ;
  buffer buf_n212( .i (n211), .o (n212) );
  assign n213 = n180 & n182 ;
  buffer buf_n214( .i (n213), .o (n214) );
  assign n215 = n212 | n214 ;
  buffer buf_n216( .i (n215), .o (n216) );
  assign n217 = n210 & n216 ;
  buffer buf_n218( .i (n217), .o (n218) );
  assign n219 = n204 | n218 ;
  buffer buf_n220( .i (n219), .o (n220) );
  assign n221 = n190 | n220 ;
  buffer buf_n222( .i (n221), .o (n222) );
  assign n223 = n94 | n108 ;
  buffer buf_n224( .i (n223), .o (n224) );
  assign n225 = n116 | n122 ;
  buffer buf_n226( .i (n225), .o (n226) );
  assign n227 = n224 | n226 ;
  buffer buf_n228( .i (n227), .o (n228) );
  assign n229 = n156 & n170 ;
  buffer buf_n230( .i (n229), .o (n230) );
  assign n231 = n178 & n184 ;
  buffer buf_n232( .i (n231), .o (n232) );
  assign n233 = n230 & n232 ;
  buffer buf_n234( .i (n233), .o (n234) );
  assign n235 = n228 | n234 ;
  buffer buf_n236( .i (n235), .o (n236) );
  assign n237 = n192 | n194 ;
  buffer buf_n238( .i (n237), .o (n238) );
  assign n239 = n198 | n200 ;
  buffer buf_n240( .i (n239), .o (n240) );
  assign n241 = n238 | n240 ;
  buffer buf_n242( .i (n241), .o (n242) );
  assign n243 = n206 & n208 ;
  buffer buf_n244( .i (n243), .o (n244) );
  assign n245 = n212 & n214 ;
  buffer buf_n246( .i (n245), .o (n246) );
  assign n247 = n244 & n246 ;
  buffer buf_n248( .i (n247), .o (n248) );
  assign n249 = n242 | n248 ;
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = n236 | n250 ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n253 = n222 & n252 ;
  buffer buf_n254( .i (n253), .o (n254) );
  assign n255 = n110 & n124 ;
  buffer buf_n256( .i (n255), .o (n256) );
  assign n257 = n172 | n186 ;
  buffer buf_n258( .i (n257), .o (n258) );
  assign n259 = n256 | n258 ;
  buffer buf_n260( .i (n259), .o (n260) );
  assign n261 = n196 & n202 ;
  buffer buf_n262( .i (n261), .o (n262) );
  assign n263 = n210 | n216 ;
  buffer buf_n264( .i (n263), .o (n264) );
  assign n265 = n262 | n264 ;
  buffer buf_n266( .i (n265), .o (n266) );
  assign n267 = n260 | n266 ;
  buffer buf_n268( .i (n267), .o (n268) );
  assign n269 = n238 & n240 ;
  buffer buf_n270( .i (n269), .o (n270) );
  assign n271 = n244 | n246 ;
  buffer buf_n272( .i (n271), .o (n272) );
  assign n273 = n270 | n272 ;
  buffer buf_n274( .i (n273), .o (n274) );
  assign n275 = n224 & n226 ;
  buffer buf_n276( .i (n275), .o (n276) );
  assign n277 = n230 | n232 ;
  buffer buf_n278( .i (n277), .o (n278) );
  assign n279 = n276 | n278 ;
  buffer buf_n280( .i (n279), .o (n280) );
  assign n281 = n274 | n280 ;
  buffer buf_n282( .i (n281), .o (n282) );
  assign n283 = n268 & n282 ;
  buffer buf_n284( .i (n283), .o (n284) );
  assign n285 = n254 & n284 ;
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n44( .i (a_26_), .o (n44) );
  buffer buf_n58( .i (a_27_), .o (n58) );
  assign n287 = n44 | n58 ;
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n41( .i (a_25_), .o (n41) );
  buffer buf_n51( .i (a_24_), .o (n51) );
  assign n289 = n41 & n51 ;
  buffer buf_n290( .i (n289), .o (n290) );
  assign n291 = n288 & n290 ;
  buffer buf_n292( .i (n291), .o (n292) );
  assign n293 = n44 & n58 ;
  buffer buf_n294( .i (n293), .o (n294) );
  assign n295 = n41 | n51 ;
  buffer buf_n296( .i (n295), .o (n296) );
  assign n297 = n294 & n296 ;
  buffer buf_n298( .i (n297), .o (n298) );
  assign n299 = n292 & n298 ;
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n49( .i (a_30_), .o (n49) );
  buffer buf_n61( .i (a_31_), .o (n61) );
  assign n301 = n49 & n61 ;
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n39( .i (a_28_), .o (n39) );
  buffer buf_n42( .i (a_29_), .o (n42) );
  assign n303 = n39 | n42 ;
  buffer buf_n304( .i (n303), .o (n304) );
  assign n305 = n302 | n304 ;
  buffer buf_n306( .i (n305), .o (n306) );
  assign n307 = n39 & n42 ;
  buffer buf_n308( .i (n307), .o (n308) );
  assign n309 = n49 | n61 ;
  buffer buf_n310( .i (n309), .o (n310) );
  assign n311 = n308 | n310 ;
  buffer buf_n312( .i (n311), .o (n312) );
  assign n313 = n306 | n312 ;
  buffer buf_n314( .i (n313), .o (n314) );
  assign n315 = n300 & n314 ;
  buffer buf_n316( .i (n315), .o (n316) );
  assign n317 = n288 | n290 ;
  buffer buf_n318( .i (n317), .o (n318) );
  assign n319 = n294 | n296 ;
  buffer buf_n320( .i (n319), .o (n320) );
  assign n321 = n318 & n320 ;
  buffer buf_n322( .i (n321), .o (n322) );
  assign n323 = n302 & n304 ;
  buffer buf_n324( .i (n323), .o (n324) );
  assign n325 = n308 & n310 ;
  buffer buf_n326( .i (n325), .o (n326) );
  assign n327 = n324 | n326 ;
  buffer buf_n328( .i (n327), .o (n328) );
  assign n329 = n322 & n328 ;
  buffer buf_n330( .i (n329), .o (n330) );
  assign n331 = n316 & n330 ;
  buffer buf_n332( .i (n331), .o (n332) );
  assign n333 = n292 | n298 ;
  buffer buf_n334( .i (n333), .o (n334) );
  assign n335 = n306 & n312 ;
  buffer buf_n336( .i (n335), .o (n336) );
  assign n337 = n334 & n336 ;
  buffer buf_n338( .i (n337), .o (n338) );
  assign n339 = n318 | n320 ;
  buffer buf_n340( .i (n339), .o (n340) );
  assign n341 = n324 & n326 ;
  buffer buf_n342( .i (n341), .o (n342) );
  assign n343 = n340 & n342 ;
  buffer buf_n344( .i (n343), .o (n344) );
  assign n345 = n338 & n344 ;
  buffer buf_n346( .i (n345), .o (n346) );
  assign n347 = n332 & n346 ;
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n43( .i (a_22_), .o (n43) );
  buffer buf_n59( .i (a_23_), .o (n59) );
  assign n349 = n43 | n59 ;
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n57( .i (a_20_), .o (n57) );
  buffer buf_n64( .i (a_21_), .o (n64) );
  assign n351 = n57 & n64 ;
  buffer buf_n352( .i (n351), .o (n352) );
  assign n353 = n350 & n352 ;
  buffer buf_n354( .i (n353), .o (n354) );
  assign n355 = n43 & n59 ;
  buffer buf_n356( .i (n355), .o (n356) );
  assign n357 = n57 | n64 ;
  buffer buf_n358( .i (n357), .o (n358) );
  assign n359 = n356 & n358 ;
  buffer buf_n360( .i (n359), .o (n360) );
  assign n361 = n354 | n360 ;
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n34( .i (a_18_), .o (n34) );
  buffer buf_n63( .i (a_19_), .o (n63) );
  assign n363 = n34 | n63 ;
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n47( .i (a_16_), .o (n47) );
  buffer buf_n54( .i (a_17_), .o (n54) );
  assign n365 = n47 & n54 ;
  buffer buf_n366( .i (n365), .o (n366) );
  assign n367 = n364 | n366 ;
  buffer buf_n368( .i (n367), .o (n368) );
  assign n369 = n34 & n63 ;
  buffer buf_n370( .i (n369), .o (n370) );
  assign n371 = n47 | n54 ;
  buffer buf_n372( .i (n371), .o (n372) );
  assign n373 = n370 | n372 ;
  buffer buf_n374( .i (n373), .o (n374) );
  assign n375 = n368 & n374 ;
  buffer buf_n376( .i (n375), .o (n376) );
  assign n377 = n362 | n376 ;
  buffer buf_n378( .i (n377), .o (n378) );
  assign n379 = n350 | n352 ;
  buffer buf_n380( .i (n379), .o (n380) );
  assign n381 = n356 | n358 ;
  buffer buf_n382( .i (n381), .o (n382) );
  assign n383 = n380 | n382 ;
  buffer buf_n384( .i (n383), .o (n384) );
  assign n385 = n364 & n366 ;
  buffer buf_n386( .i (n385), .o (n386) );
  assign n387 = n370 & n372 ;
  buffer buf_n388( .i (n387), .o (n388) );
  assign n389 = n386 & n388 ;
  buffer buf_n390( .i (n389), .o (n390) );
  assign n391 = n384 | n390 ;
  buffer buf_n392( .i (n391), .o (n392) );
  assign n393 = n378 | n392 ;
  buffer buf_n394( .i (n393), .o (n394) );
  assign n395 = n354 & n360 ;
  buffer buf_n396( .i (n395), .o (n396) );
  assign n397 = n368 | n374 ;
  buffer buf_n398( .i (n397), .o (n398) );
  assign n399 = n396 | n398 ;
  buffer buf_n400( .i (n399), .o (n400) );
  assign n401 = n380 & n382 ;
  buffer buf_n402( .i (n401), .o (n402) );
  assign n403 = n386 | n388 ;
  buffer buf_n404( .i (n403), .o (n404) );
  assign n405 = n402 | n404 ;
  buffer buf_n406( .i (n405), .o (n406) );
  assign n407 = n400 | n406 ;
  buffer buf_n408( .i (n407), .o (n408) );
  assign n409 = n394 | n408 ;
  buffer buf_n410( .i (n409), .o (n410) );
  assign n411 = n348 & n410 ;
  buffer buf_n412( .i (n411), .o (n412) );
  assign n413 = n362 & n376 ;
  buffer buf_n414( .i (n413), .o (n414) );
  assign n415 = n384 & n390 ;
  buffer buf_n416( .i (n415), .o (n416) );
  assign n417 = n414 | n416 ;
  buffer buf_n418( .i (n417), .o (n418) );
  assign n419 = n396 & n398 ;
  buffer buf_n420( .i (n419), .o (n420) );
  assign n421 = n402 & n404 ;
  buffer buf_n422( .i (n421), .o (n422) );
  assign n423 = n420 | n422 ;
  buffer buf_n424( .i (n423), .o (n424) );
  assign n425 = n418 | n424 ;
  buffer buf_n426( .i (n425), .o (n426) );
  assign n427 = n300 | n314 ;
  buffer buf_n428( .i (n427), .o (n428) );
  assign n429 = n322 | n328 ;
  buffer buf_n430( .i (n429), .o (n430) );
  assign n431 = n428 & n430 ;
  buffer buf_n432( .i (n431), .o (n432) );
  assign n433 = n334 | n336 ;
  buffer buf_n434( .i (n433), .o (n434) );
  assign n435 = n340 | n342 ;
  buffer buf_n436( .i (n435), .o (n436) );
  assign n437 = n434 & n436 ;
  buffer buf_n438( .i (n437), .o (n438) );
  assign n439 = n432 & n438 ;
  buffer buf_n440( .i (n439), .o (n440) );
  assign n441 = n426 & n440 ;
  buffer buf_n442( .i (n441), .o (n442) );
  assign n443 = n412 & n442 ;
  buffer buf_n444( .i (n443), .o (n444) );
  assign n445 = n316 | n330 ;
  buffer buf_n446( .i (n445), .o (n446) );
  assign n447 = n338 | n344 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = n446 & n448 ;
  buffer buf_n450( .i (n449), .o (n450) );
  assign n451 = n378 & n392 ;
  buffer buf_n452( .i (n451), .o (n452) );
  assign n453 = n400 & n406 ;
  buffer buf_n454( .i (n453), .o (n454) );
  assign n455 = n452 | n454 ;
  buffer buf_n456( .i (n455), .o (n456) );
  assign n457 = n450 & n456 ;
  buffer buf_n458( .i (n457), .o (n458) );
  assign n459 = n414 & n416 ;
  buffer buf_n460( .i (n459), .o (n460) );
  assign n461 = n420 & n422 ;
  buffer buf_n462( .i (n461), .o (n462) );
  assign n463 = n460 | n462 ;
  buffer buf_n464( .i (n463), .o (n464) );
  assign n465 = n428 | n430 ;
  buffer buf_n466( .i (n465), .o (n466) );
  assign n467 = n434 | n436 ;
  buffer buf_n468( .i (n467), .o (n468) );
  assign n469 = n466 & n468 ;
  buffer buf_n470( .i (n469), .o (n470) );
  assign n471 = n464 & n470 ;
  buffer buf_n472( .i (n471), .o (n472) );
  assign n473 = n458 & n472 ;
  buffer buf_n474( .i (n473), .o (n474) );
  assign n475 = n444 | n474 ;
  buffer buf_n476( .i (n475), .o (n476) );
  assign n477 = n332 | n346 ;
  buffer buf_n478( .i (n477), .o (n478) );
  assign n479 = n394 & n408 ;
  buffer buf_n480( .i (n479), .o (n480) );
  assign n481 = n478 & n480 ;
  buffer buf_n482( .i (n481), .o (n482) );
  assign n483 = n418 & n424 ;
  buffer buf_n484( .i (n483), .o (n484) );
  assign n485 = n432 | n438 ;
  buffer buf_n486( .i (n485), .o (n486) );
  assign n487 = n484 & n486 ;
  buffer buf_n488( .i (n487), .o (n488) );
  assign n489 = n482 & n488 ;
  buffer buf_n490( .i (n489), .o (n490) );
  assign n491 = n446 | n448 ;
  buffer buf_n492( .i (n491), .o (n492) );
  assign n493 = n452 & n454 ;
  buffer buf_n494( .i (n493), .o (n494) );
  assign n495 = n492 & n494 ;
  buffer buf_n496( .i (n495), .o (n496) );
  assign n497 = n460 & n462 ;
  buffer buf_n498( .i (n497), .o (n498) );
  assign n499 = n466 | n468 ;
  buffer buf_n500( .i (n499), .o (n500) );
  assign n501 = n498 & n500 ;
  buffer buf_n502( .i (n501), .o (n502) );
  assign n503 = n496 & n502 ;
  buffer buf_n504( .i (n503), .o (n504) );
  assign n505 = n490 | n504 ;
  buffer buf_n506( .i (n505), .o (n506) );
  assign n507 = n476 | n506 ;
  buffer buf_n508( .i (n507), .o (n508) );
  assign n509 = n286 & n508 ;
  buffer buf_n510( .i (n509), .o (n510) );
  assign n511 = n126 & n188 ;
  buffer buf_n512( .i (n511), .o (n512) );
  assign n513 = n204 & n218 ;
  buffer buf_n514( .i (n513), .o (n514) );
  assign n515 = n512 | n514 ;
  buffer buf_n516( .i (n515), .o (n516) );
  assign n517 = n228 & n234 ;
  buffer buf_n518( .i (n517), .o (n518) );
  assign n519 = n242 & n248 ;
  buffer buf_n520( .i (n519), .o (n520) );
  assign n521 = n518 | n520 ;
  buffer buf_n522( .i (n521), .o (n522) );
  assign n523 = n516 & n522 ;
  buffer buf_n524( .i (n523), .o (n524) );
  assign n525 = n256 & n258 ;
  buffer buf_n526( .i (n525), .o (n526) );
  assign n527 = n262 & n264 ;
  buffer buf_n528( .i (n527), .o (n528) );
  assign n529 = n526 | n528 ;
  buffer buf_n530( .i (n529), .o (n530) );
  assign n531 = n276 & n278 ;
  buffer buf_n532( .i (n531), .o (n532) );
  assign n533 = n270 & n272 ;
  buffer buf_n534( .i (n533), .o (n534) );
  assign n535 = n532 | n534 ;
  buffer buf_n536( .i (n535), .o (n536) );
  assign n537 = n530 & n536 ;
  buffer buf_n538( .i (n537), .o (n538) );
  assign n539 = n524 & n538 ;
  buffer buf_n540( .i (n539), .o (n540) );
  assign n541 = n478 | n480 ;
  buffer buf_n542( .i (n541), .o (n542) );
  assign n543 = n484 | n486 ;
  buffer buf_n544( .i (n543), .o (n544) );
  assign n545 = n542 & n544 ;
  buffer buf_n546( .i (n545), .o (n546) );
  assign n547 = n492 | n494 ;
  buffer buf_n548( .i (n547), .o (n548) );
  assign n549 = n498 | n500 ;
  buffer buf_n550( .i (n549), .o (n550) );
  assign n551 = n548 & n550 ;
  buffer buf_n552( .i (n551), .o (n552) );
  assign n553 = n546 | n552 ;
  buffer buf_n554( .i (n553), .o (n554) );
  assign n555 = n348 | n410 ;
  buffer buf_n556( .i (n555), .o (n556) );
  assign n557 = n426 | n440 ;
  buffer buf_n558( .i (n557), .o (n558) );
  assign n559 = n556 & n558 ;
  buffer buf_n560( .i (n559), .o (n560) );
  assign n561 = n450 | n456 ;
  buffer buf_n562( .i (n561), .o (n562) );
  assign n563 = n464 | n470 ;
  buffer buf_n564( .i (n563), .o (n564) );
  assign n565 = n562 & n564 ;
  buffer buf_n566( .i (n565), .o (n566) );
  assign n567 = n560 | n566 ;
  buffer buf_n568( .i (n567), .o (n568) );
  assign n569 = n554 | n568 ;
  buffer buf_n570( .i (n569), .o (n570) );
  assign n571 = n540 & n570 ;
  buffer buf_n572( .i (n571), .o (n572) );
  assign n573 = n510 | n572 ;
  buffer buf_n574( .i (n573), .o (n574) );
  assign n575 = n190 & n220 ;
  buffer buf_n576( .i (n575), .o (n576) );
  assign n577 = n236 & n250 ;
  buffer buf_n578( .i (n577), .o (n578) );
  assign n579 = n576 & n578 ;
  buffer buf_n580( .i (n579), .o (n580) );
  assign n581 = n260 & n266 ;
  buffer buf_n582( .i (n581), .o (n582) );
  assign n583 = n274 & n280 ;
  buffer buf_n584( .i (n583), .o (n584) );
  assign n585 = n582 & n584 ;
  buffer buf_n586( .i (n585), .o (n586) );
  assign n587 = n580 & n586 ;
  buffer buf_n588( .i (n587), .o (n588) );
  assign n589 = n412 | n442 ;
  buffer buf_n590( .i (n589), .o (n590) );
  assign n591 = n458 | n472 ;
  buffer buf_n592( .i (n591), .o (n592) );
  assign n593 = n590 | n592 ;
  buffer buf_n594( .i (n593), .o (n594) );
  assign n595 = n482 | n488 ;
  buffer buf_n596( .i (n595), .o (n596) );
  assign n597 = n496 | n502 ;
  buffer buf_n598( .i (n597), .o (n598) );
  assign n599 = n596 | n598 ;
  buffer buf_n600( .i (n599), .o (n600) );
  assign n601 = n594 | n600 ;
  buffer buf_n602( .i (n601), .o (n602) );
  assign n603 = n588 & n602 ;
  buffer buf_n604( .i (n603), .o (n604) );
  assign n605 = n512 & n514 ;
  buffer buf_n606( .i (n605), .o (n606) );
  assign n607 = n518 & n520 ;
  buffer buf_n608( .i (n607), .o (n608) );
  assign n609 = n606 & n608 ;
  buffer buf_n610( .i (n609), .o (n610) );
  assign n611 = n526 & n528 ;
  buffer buf_n612( .i (n611), .o (n612) );
  assign n613 = n532 & n534 ;
  buffer buf_n614( .i (n613), .o (n614) );
  assign n615 = n612 & n614 ;
  buffer buf_n616( .i (n615), .o (n616) );
  assign n617 = n610 & n616 ;
  buffer buf_n618( .i (n617), .o (n618) );
  assign n619 = n542 | n544 ;
  buffer buf_n620( .i (n619), .o (n620) );
  assign n621 = n548 | n550 ;
  buffer buf_n622( .i (n621), .o (n622) );
  assign n623 = n620 | n622 ;
  buffer buf_n624( .i (n623), .o (n624) );
  assign n625 = n556 | n558 ;
  buffer buf_n626( .i (n625), .o (n626) );
  assign n627 = n562 | n564 ;
  buffer buf_n628( .i (n627), .o (n628) );
  assign n629 = n626 | n628 ;
  buffer buf_n630( .i (n629), .o (n630) );
  assign n631 = n624 | n630 ;
  buffer buf_n632( .i (n631), .o (n632) );
  assign n633 = n618 & n632 ;
  buffer buf_n634( .i (n633), .o (n634) );
  assign n635 = n604 | n634 ;
  buffer buf_n636( .i (n635), .o (n636) );
  assign n637 = n574 & n636 ;
  buffer buf_n638( .i (n637), .o (n638) );
  assign n639 = n222 | n252 ;
  buffer buf_n640( .i (n639), .o (n640) );
  assign n641 = n268 | n282 ;
  buffer buf_n642( .i (n641), .o (n642) );
  assign n643 = n640 & n642 ;
  buffer buf_n644( .i (n643), .o (n644) );
  assign n645 = n444 & n474 ;
  buffer buf_n646( .i (n645), .o (n646) );
  assign n647 = n490 & n504 ;
  buffer buf_n648( .i (n647), .o (n648) );
  assign n649 = n646 | n648 ;
  buffer buf_n650( .i (n649), .o (n650) );
  assign n651 = n644 & n650 ;
  buffer buf_n652( .i (n651), .o (n652) );
  assign n653 = n516 | n522 ;
  buffer buf_n654( .i (n653), .o (n654) );
  assign n655 = n530 | n536 ;
  buffer buf_n656( .i (n655), .o (n656) );
  assign n657 = n654 & n656 ;
  buffer buf_n658( .i (n657), .o (n658) );
  assign n659 = n546 & n552 ;
  buffer buf_n660( .i (n659), .o (n660) );
  assign n661 = n560 & n566 ;
  buffer buf_n662( .i (n661), .o (n662) );
  assign n663 = n660 | n662 ;
  buffer buf_n664( .i (n663), .o (n664) );
  assign n665 = n658 & n664 ;
  buffer buf_n666( .i (n665), .o (n666) );
  assign n667 = n652 | n666 ;
  buffer buf_n668( .i (n667), .o (n668) );
  assign n669 = n576 | n578 ;
  buffer buf_n670( .i (n669), .o (n670) );
  assign n671 = n582 | n584 ;
  buffer buf_n672( .i (n671), .o (n672) );
  assign n673 = n670 & n672 ;
  buffer buf_n674( .i (n673), .o (n674) );
  assign n675 = n590 & n592 ;
  buffer buf_n676( .i (n675), .o (n676) );
  assign n677 = n596 & n598 ;
  buffer buf_n678( .i (n677), .o (n678) );
  assign n679 = n676 | n678 ;
  buffer buf_n680( .i (n679), .o (n680) );
  assign n681 = n674 & n680 ;
  buffer buf_n682( .i (n681), .o (n682) );
  assign n683 = n606 | n608 ;
  buffer buf_n684( .i (n683), .o (n684) );
  assign n685 = n612 | n614 ;
  buffer buf_n686( .i (n685), .o (n686) );
  assign n687 = n684 & n686 ;
  buffer buf_n688( .i (n687), .o (n688) );
  assign n689 = n620 & n622 ;
  buffer buf_n690( .i (n689), .o (n690) );
  assign n691 = n626 & n628 ;
  buffer buf_n692( .i (n691), .o (n692) );
  assign n693 = n690 | n692 ;
  buffer buf_n694( .i (n693), .o (n694) );
  assign n695 = n688 & n694 ;
  buffer buf_n696( .i (n695), .o (n696) );
  assign n697 = n682 | n696 ;
  buffer buf_n698( .i (n697), .o (n698) );
  assign n699 = n668 & n698 ;
  buffer buf_n700( .i (n699), .o (n700) );
  assign n701 = n638 & n700 ;
  buffer buf_n702( .i (n701), .o (n702) );
  assign n703 = n254 | n284 ;
  buffer buf_n704( .i (n703), .o (n704) );
  assign n705 = n476 & n506 ;
  buffer buf_n706( .i (n705), .o (n706) );
  assign n707 = n704 & n706 ;
  buffer buf_n708( .i (n707), .o (n708) );
  assign n709 = n524 | n538 ;
  buffer buf_n710( .i (n709), .o (n710) );
  assign n711 = n554 & n568 ;
  buffer buf_n712( .i (n711), .o (n712) );
  assign n713 = n710 & n712 ;
  buffer buf_n714( .i (n713), .o (n714) );
  assign n715 = n708 | n714 ;
  buffer buf_n716( .i (n715), .o (n716) );
  assign n717 = n580 | n586 ;
  buffer buf_n718( .i (n717), .o (n718) );
  assign n719 = n594 & n600 ;
  buffer buf_n720( .i (n719), .o (n720) );
  assign n721 = n718 & n720 ;
  buffer buf_n722( .i (n721), .o (n722) );
  assign n723 = n610 | n616 ;
  buffer buf_n724( .i (n723), .o (n724) );
  assign n725 = n624 & n630 ;
  buffer buf_n726( .i (n725), .o (n726) );
  assign n727 = n724 & n726 ;
  buffer buf_n728( .i (n727), .o (n728) );
  assign n729 = n722 | n728 ;
  buffer buf_n730( .i (n729), .o (n730) );
  assign n731 = n716 & n730 ;
  buffer buf_n732( .i (n731), .o (n732) );
  assign n733 = n640 | n642 ;
  buffer buf_n734( .i (n733), .o (n734) );
  assign n735 = n646 & n648 ;
  buffer buf_n736( .i (n735), .o (n736) );
  assign n737 = n734 & n736 ;
  buffer buf_n738( .i (n737), .o (n738) );
  assign n739 = n654 | n656 ;
  buffer buf_n740( .i (n739), .o (n740) );
  assign n741 = n660 & n662 ;
  buffer buf_n742( .i (n741), .o (n742) );
  assign n743 = n740 & n742 ;
  buffer buf_n744( .i (n743), .o (n744) );
  assign n745 = n738 | n744 ;
  buffer buf_n746( .i (n745), .o (n746) );
  assign n747 = n670 | n672 ;
  buffer buf_n748( .i (n747), .o (n748) );
  assign n749 = n676 & n678 ;
  buffer buf_n750( .i (n749), .o (n750) );
  assign n751 = n748 & n750 ;
  buffer buf_n752( .i (n751), .o (n752) );
  assign n753 = n684 | n686 ;
  buffer buf_n754( .i (n753), .o (n754) );
  assign n755 = n690 & n692 ;
  buffer buf_n756( .i (n755), .o (n756) );
  assign n757 = n754 & n756 ;
  buffer buf_n758( .i (n757), .o (n758) );
  assign n759 = n752 | n758 ;
  buffer buf_n760( .i (n759), .o (n760) );
  assign n761 = n746 & n760 ;
  buffer buf_n762( .i (n761), .o (n762) );
  assign n763 = n732 & n762 ;
  buffer buf_n764( .i (n763), .o (n764) );
  assign n765 = n702 | n764 ;
  assign n766 = n510 & n572 ;
  buffer buf_n767( .i (n766), .o (n767) );
  assign n768 = n604 & n634 ;
  buffer buf_n769( .i (n768), .o (n769) );
  assign n770 = n767 & n769 ;
  buffer buf_n771( .i (n770), .o (n771) );
  assign n772 = n652 & n666 ;
  buffer buf_n773( .i (n772), .o (n773) );
  assign n774 = n682 & n696 ;
  buffer buf_n775( .i (n774), .o (n775) );
  assign n776 = n773 & n775 ;
  buffer buf_n777( .i (n776), .o (n777) );
  assign n778 = n771 & n777 ;
  buffer buf_n779( .i (n778), .o (n779) );
  assign n780 = n708 & n714 ;
  buffer buf_n781( .i (n780), .o (n781) );
  assign n782 = n722 & n728 ;
  buffer buf_n783( .i (n782), .o (n783) );
  assign n784 = n781 & n783 ;
  buffer buf_n785( .i (n784), .o (n785) );
  assign n786 = n738 & n744 ;
  buffer buf_n787( .i (n786), .o (n787) );
  assign n788 = n752 & n758 ;
  buffer buf_n789( .i (n788), .o (n789) );
  assign n790 = n787 & n789 ;
  buffer buf_n791( .i (n790), .o (n791) );
  assign n792 = n785 & n791 ;
  buffer buf_n793( .i (n792), .o (n793) );
  assign n794 = n779 | n793 ;
  assign n795 = n286 | n508 ;
  buffer buf_n796( .i (n795), .o (n796) );
  assign n797 = n540 | n570 ;
  buffer buf_n798( .i (n797), .o (n798) );
  assign n799 = n796 & n798 ;
  buffer buf_n800( .i (n799), .o (n800) );
  assign n801 = n588 | n602 ;
  buffer buf_n802( .i (n801), .o (n802) );
  assign n803 = n618 | n632 ;
  buffer buf_n804( .i (n803), .o (n804) );
  assign n805 = n802 & n804 ;
  buffer buf_n806( .i (n805), .o (n806) );
  assign n807 = n800 & n806 ;
  buffer buf_n808( .i (n807), .o (n808) );
  assign n809 = n644 | n650 ;
  buffer buf_n810( .i (n809), .o (n810) );
  assign n811 = n658 | n664 ;
  buffer buf_n812( .i (n811), .o (n812) );
  assign n813 = n810 & n812 ;
  buffer buf_n814( .i (n813), .o (n814) );
  assign n815 = n674 | n680 ;
  buffer buf_n816( .i (n815), .o (n816) );
  assign n817 = n688 | n694 ;
  buffer buf_n818( .i (n817), .o (n818) );
  assign n819 = n816 & n818 ;
  buffer buf_n820( .i (n819), .o (n820) );
  assign n821 = n814 & n820 ;
  buffer buf_n822( .i (n821), .o (n822) );
  assign n823 = n808 & n822 ;
  buffer buf_n824( .i (n823), .o (n824) );
  assign n825 = n704 | n706 ;
  buffer buf_n826( .i (n825), .o (n826) );
  assign n827 = n710 | n712 ;
  buffer buf_n828( .i (n827), .o (n828) );
  assign n829 = n826 & n828 ;
  buffer buf_n830( .i (n829), .o (n830) );
  assign n831 = n718 | n720 ;
  buffer buf_n832( .i (n831), .o (n832) );
  assign n833 = n724 | n726 ;
  buffer buf_n834( .i (n833), .o (n834) );
  assign n835 = n832 & n834 ;
  buffer buf_n836( .i (n835), .o (n836) );
  assign n837 = n830 & n836 ;
  buffer buf_n838( .i (n837), .o (n838) );
  assign n839 = n734 | n736 ;
  buffer buf_n840( .i (n839), .o (n840) );
  assign n841 = n740 | n742 ;
  buffer buf_n842( .i (n841), .o (n842) );
  assign n843 = n840 & n842 ;
  buffer buf_n844( .i (n843), .o (n844) );
  assign n845 = n748 | n750 ;
  buffer buf_n846( .i (n845), .o (n846) );
  assign n847 = n754 | n756 ;
  buffer buf_n848( .i (n847), .o (n848) );
  assign n849 = n846 & n848 ;
  buffer buf_n850( .i (n849), .o (n850) );
  assign n851 = n844 & n850 ;
  buffer buf_n852( .i (n851), .o (n852) );
  assign n853 = n838 & n852 ;
  buffer buf_n854( .i (n853), .o (n854) );
  assign n855 = n824 | n854 ;
  assign n856 = n638 | n700 ;
  buffer buf_n857( .i (n856), .o (n857) );
  assign n858 = n732 | n762 ;
  buffer buf_n859( .i (n858), .o (n859) );
  assign n860 = n857 | n859 ;
  assign n861 = n796 | n798 ;
  buffer buf_n862( .i (n861), .o (n862) );
  assign n863 = n802 | n804 ;
  buffer buf_n864( .i (n863), .o (n864) );
  assign n865 = n862 | n864 ;
  buffer buf_n866( .i (n865), .o (n866) );
  assign n867 = n810 | n812 ;
  buffer buf_n868( .i (n867), .o (n868) );
  assign n869 = n816 | n818 ;
  buffer buf_n870( .i (n869), .o (n870) );
  assign n871 = n868 | n870 ;
  buffer buf_n872( .i (n871), .o (n872) );
  assign n873 = n866 | n872 ;
  buffer buf_n874( .i (n873), .o (n874) );
  assign n875 = n826 | n828 ;
  buffer buf_n876( .i (n875), .o (n876) );
  assign n877 = n832 | n834 ;
  buffer buf_n878( .i (n877), .o (n878) );
  assign n879 = n876 | n878 ;
  buffer buf_n880( .i (n879), .o (n880) );
  assign n881 = n840 | n842 ;
  buffer buf_n882( .i (n881), .o (n882) );
  assign n883 = n846 | n848 ;
  buffer buf_n884( .i (n883), .o (n884) );
  assign n885 = n882 | n884 ;
  buffer buf_n886( .i (n885), .o (n886) );
  assign n887 = n880 | n886 ;
  buffer buf_n888( .i (n887), .o (n888) );
  assign n889 = n874 | n888 ;
  assign n890 = n862 & n864 ;
  buffer buf_n891( .i (n890), .o (n891) );
  assign n892 = n868 & n870 ;
  buffer buf_n893( .i (n892), .o (n893) );
  assign n894 = n891 | n893 ;
  buffer buf_n895( .i (n894), .o (n895) );
  assign n896 = n876 & n878 ;
  buffer buf_n897( .i (n896), .o (n897) );
  assign n898 = n882 & n884 ;
  buffer buf_n899( .i (n898), .o (n899) );
  assign n900 = n897 | n899 ;
  buffer buf_n901( .i (n900), .o (n901) );
  assign n902 = n895 & n901 ;
  assign n903 = n866 & n872 ;
  buffer buf_n904( .i (n903), .o (n904) );
  assign n905 = n880 & n886 ;
  buffer buf_n906( .i (n905), .o (n906) );
  assign n907 = n904 | n906 ;
  assign n908 = n891 & n893 ;
  buffer buf_n909( .i (n908), .o (n909) );
  assign n910 = n897 & n899 ;
  buffer buf_n911( .i (n910), .o (n911) );
  assign n912 = n909 & n911 ;
  assign n913 = n800 | n806 ;
  buffer buf_n914( .i (n913), .o (n914) );
  assign n915 = n814 | n820 ;
  buffer buf_n916( .i (n915), .o (n916) );
  assign n917 = n914 | n916 ;
  buffer buf_n918( .i (n917), .o (n918) );
  assign n919 = n830 | n836 ;
  buffer buf_n920( .i (n919), .o (n920) );
  assign n921 = n844 | n850 ;
  buffer buf_n922( .i (n921), .o (n922) );
  assign n923 = n920 | n922 ;
  buffer buf_n924( .i (n923), .o (n924) );
  assign n925 = n918 | n924 ;
  assign n926 = n702 & n764 ;
  assign n927 = n767 | n769 ;
  buffer buf_n928( .i (n927), .o (n928) );
  assign n929 = n773 | n775 ;
  buffer buf_n930( .i (n929), .o (n930) );
  assign n931 = n928 & n930 ;
  buffer buf_n932( .i (n931), .o (n932) );
  assign n933 = n781 | n783 ;
  buffer buf_n934( .i (n933), .o (n934) );
  assign n935 = n787 | n789 ;
  buffer buf_n936( .i (n935), .o (n936) );
  assign n937 = n934 & n936 ;
  buffer buf_n938( .i (n937), .o (n938) );
  assign n939 = n932 & n938 ;
  assign n940 = n909 | n911 ;
  assign n941 = n928 | n930 ;
  buffer buf_n942( .i (n941), .o (n942) );
  assign n943 = n934 | n936 ;
  buffer buf_n944( .i (n943), .o (n944) );
  assign n945 = n942 | n944 ;
  assign n946 = n932 | n938 ;
  assign n947 = n808 | n822 ;
  buffer buf_n948( .i (n947), .o (n948) );
  assign n949 = n838 | n852 ;
  buffer buf_n950( .i (n949), .o (n950) );
  assign n951 = n948 & n950 ;
  assign n952 = n574 | n636 ;
  buffer buf_n953( .i (n952), .o (n953) );
  assign n954 = n668 | n698 ;
  buffer buf_n955( .i (n954), .o (n955) );
  assign n956 = n953 & n955 ;
  buffer buf_n957( .i (n956), .o (n957) );
  assign n958 = n716 | n730 ;
  buffer buf_n959( .i (n958), .o (n959) );
  assign n960 = n746 | n760 ;
  buffer buf_n961( .i (n960), .o (n961) );
  assign n962 = n959 & n961 ;
  buffer buf_n963( .i (n962), .o (n963) );
  assign n964 = n957 & n963 ;
  assign n965 = n824 & n854 ;
  assign n966 = n918 & n924 ;
  assign n967 = n953 | n955 ;
  buffer buf_n968( .i (n967), .o (n968) );
  assign n969 = n959 | n961 ;
  buffer buf_n970( .i (n969), .o (n970) );
  assign n971 = n968 & n970 ;
  assign n972 = n914 & n916 ;
  buffer buf_n973( .i (n972), .o (n973) );
  assign n974 = n920 & n922 ;
  buffer buf_n975( .i (n974), .o (n975) );
  assign n976 = n973 & n975 ;
  assign n977 = n968 | n970 ;
  assign n978 = n771 | n777 ;
  buffer buf_n979( .i (n978), .o (n979) );
  assign n980 = n785 | n791 ;
  buffer buf_n981( .i (n980), .o (n981) );
  assign n982 = n979 | n981 ;
  assign n983 = n874 & n888 ;
  assign n984 = n895 | n901 ;
  assign n985 = n973 | n975 ;
  assign n986 = n948 | n950 ;
  assign n987 = n957 | n963 ;
  assign n988 = n942 & n944 ;
  assign n989 = n779 & n793 ;
  assign n990 = n857 & n859 ;
  assign n991 = n904 & n906 ;
  assign n992 = n979 & n981 ;
  assign b_9_ = n765 ;
  assign b_1_ = n794 ;
  assign b_17_ = n855 ;
  assign b_11_ = n860 ;
  assign b_31_ = n889 ;
  assign b_26_ = n902 ;
  assign b_29_ = n907 ;
  assign b_24_ = n912 ;
  assign b_23_ = n925 ;
  assign b_8_ = n926 ;
  assign b_4_ = n939 ;
  assign b_25_ = n940 ;
  assign b_7_ = n945 ;
  assign b_5_ = n946 ;
  assign b_18_ = n951 ;
  assign b_12_ = n964 ;
  assign b_16_ = n965 ;
  assign b_22_ = n966 ;
  assign b_14_ = n971 ;
  assign b_20_ = n976 ;
  assign b_15_ = n977 ;
  assign b_3_ = n982 ;
  assign b_30_ = n983 ;
  assign b_27_ = n984 ;
  assign b_21_ = n985 ;
  assign b_19_ = n986 ;
  assign b_13_ = n987 ;
  assign b_6_ = n988 ;
  assign b_0_ = n989 ;
  assign b_10_ = n990 ;
  assign b_28_ = n991 ;
  assign b_2_ = n992 ;
endmodule
