module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G6 , G7 , G8 , G9 , G3519 , G3520 , G3521 , G3522 , G3523 , G3524 , G3525 , G3526 , G3527 , G3528 , G3529 , G3530 , G3531 , G3532 , G3533 , G3534 , G3535 , G3536 , G3537 , G3538 , G3539 , G3540 );
  input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G6 , G7 , G8 , G9 ;
  output G3519 , G3520 , G3521 , G3522 , G3523 , G3524 , G3525 , G3526 , G3527 , G3528 , G3529 , G3530 , G3531 , G3532 , G3533 , G3534 , G3535 , G3536 , G3537 , G3538 , G3539 , G3540 ;
  wire n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 ;
  buffer buf_n661( .i (G8), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n672( .i (G9), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  assign n686 = n662 | n673 ;
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n79( .i (G10), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n648( .i (G7), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  assign n688 = n80 | n649 ;
  buffer buf_n689( .i (n688), .o (n689) );
  assign n692 = ~n687 & ~n689 ;
  buffer buf_n92( .i (G11), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n104( .i (G12), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n118( .i (G13), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  assign n693 = n106 | n120 ;
  buffer buf_n694( .i (n693), .o (n694) );
  assign n695 = ~n96 | ~n694 ;
  buffer buf_n51( .i (G1), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n330( .i (G3), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  assign n696 = n56 | n335 ;
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n352( .i (G32), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  assign n698 = n355 & ~n675 ;
  buffer buf_n346( .i (G31), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  assign n699 = n349 & ~n664 ;
  assign n700 = n698 | n699 ;
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n381( .i (G36), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  assign n701 = ~n121 & n384 ;
  buffer buf_n131( .i (G14), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n389( .i (G37), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  assign n702 = ~n134 & n392 ;
  assign n703 = n701 | n702 ;
  assign n704 = n700 | n703 ;
  buffer buf_n364( .i (G34), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  assign n705 = ~n95 & n367 ;
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n373( .i (G35), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  assign n706 = ~n107 & n376 ;
  assign n707 = n705 | n706 ;
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n358( .i (G33), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  assign n708 = ~n82 & n361 ;
  buffer buf_n340( .i (G30), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  assign n709 = n343 & ~n651 ;
  assign n710 = n708 | n709 ;
  assign n711 = n707 | n710 ;
  assign n712 = n704 | n711 ;
  assign n713 = n697 & n712 ;
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n185( .i (G2), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n717 = ~n52 & n186 ;
  buffer buf_n718( .i (n717), .o (n718) );
  assign n721 = ~n333 & n718 ;
  buffer buf_n722( .i (n721), .o (n722) );
  assign n723 = ~n651 & n687 ;
  buffer buf_n724( .i (n723), .o (n724) );
  assign n731 = n722 & n724 ;
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  assign n736 = n192 | n697 ;
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  assign n738 = n380 | n388 ;
  assign n739 = n372 & n738 ;
  assign n740 = ~n737 & n739 ;
  assign n741 = n735 | n740 ;
  assign n742 = ~n716 & ~n741 ;
  assign n743 = n382 | n390 ;
  assign n744 = n382 & n390 ;
  assign n745 = n743 & ~n744 ;
  buffer buf_n746( .i (n745), .o (n746) );
  assign n747 = n365 & ~n374 ;
  assign n748 = ~n365 & n374 ;
  assign n749 = n747 | n748 ;
  buffer buf_n750( .i (n749), .o (n750) );
  assign n751 = n746 | n750 ;
  assign n752 = n746 & n750 ;
  assign n753 = n751 & ~n752 ;
  buffer buf_n754( .i (n753), .o (n754) );
  assign n755 = n341 & ~n347 ;
  assign n756 = ~n341 & n347 ;
  assign n757 = n755 | n756 ;
  buffer buf_n758( .i (n757), .o (n758) );
  assign n759 = n353 | n359 ;
  assign n760 = n353 & n359 ;
  assign n761 = n759 & ~n760 ;
  buffer buf_n762( .i (n761), .o (n762) );
  assign n763 = n758 | n762 ;
  assign n764 = n758 & n762 ;
  assign n765 = n763 & ~n764 ;
  buffer buf_n766( .i (n765), .o (n766) );
  assign n767 = n754 | n766 ;
  assign n768 = n754 & n766 ;
  assign n769 = n767 & ~n768 ;
  assign n770 = n663 & n674 ;
  assign n771 = n687 & ~n770 ;
  buffer buf_n772( .i (n771), .o (n772) );
  assign n773 = n81 & n650 ;
  assign n774 = n689 & ~n773 ;
  buffer buf_n775( .i (n774), .o (n775) );
  assign n776 = ~n772 & n775 ;
  assign n777 = n772 & ~n775 ;
  assign n778 = n776 | n777 ;
  buffer buf_n779( .i (n778), .o (n779) );
  assign n780 = ~n94 & n120 ;
  assign n781 = n94 & ~n120 ;
  assign n782 = n780 | n781 ;
  buffer buf_n783( .i (n782), .o (n783) );
  assign n784 = n106 | n133 ;
  assign n785 = n106 & n133 ;
  assign n786 = n784 & ~n785 ;
  buffer buf_n787( .i (n786), .o (n787) );
  assign n788 = n783 & ~n787 ;
  assign n789 = ~n783 & n787 ;
  assign n790 = n788 | n789 ;
  buffer buf_n791( .i (n790), .o (n791) );
  assign n792 = n779 & n791 ;
  assign n793 = n779 | n791 ;
  assign n794 = ~n792 & n793 ;
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  assign n795 = n333 & n718 ;
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  assign n801 = n657 | n800 ;
  assign n802 = ~n53 & n332 ;
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  assign n807 = n53 & n187 ;
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n418( .i (G4), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  assign n809 = n53 & n332 ;
  assign n810 = n421 & n809 ;
  assign n811 = n808 | n810 ;
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  assign n815 = n806 | n813 ;
  buffer buf_n816( .i (n815), .o (n816) );
  assign n817 = n657 & n816 ;
  assign n818 = n801 & ~n817 ;
  buffer buf_n814( .i (n813), .o (n814) );
  assign n819 = n651 | n687 ;
  assign n820 = n334 & n819 ;
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n218( .i (G21), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  assign n823 = n333 | n421 ;
  buffer buf_n824( .i (n823), .o (n824) );
  assign n825 = n223 & ~n824 ;
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  assign n826 = ~n332 & n420 ;
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  assign n829 = ~n666 & n828 ;
  assign n830 = n825 | n829 ;
  assign n831 = n822 | n830 ;
  assign n832 = n814 & n831 ;
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  assign n835 = n818 | n834 ;
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n261( .i (G25), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n264( .i (G26), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  assign n838 = n262 | n265 ;
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n572( .i (G5), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n636( .i (G6), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  assign n850 = n573 | n637 ;
  buffer buf_n851( .i (n52), .o (n851) );
  assign n852 = n850 & ~n851 ;
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n396( .i (G38), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n574( .i (n573), .o (n574) );
  assign n859 = n420 & n574 ;
  buffer buf_n860( .i (n859), .o (n860) );
  assign n865 = n808 & ~n860 ;
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  assign n869 = n403 & ~n867 ;
  buffer buf_n870( .i (n869), .o (n870) );
  assign n871 = n858 & n870 ;
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  assign n873 = n345 & ~n854 ;
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n318( .i (G28), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n569( .i (G49), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  assign n875 = n420 | n571 ;
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  assign n878 = n323 & ~n877 ;
  assign n879 = n82 & ~n421 ;
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n324( .i (G29), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n422( .i (n421), .o (n422) );
  assign n881 = n328 & n422 ;
  assign n882 = n880 | n881 ;
  assign n883 = n878 | n882 ;
  assign n884 = n874 | n883 ;
  assign n885 = ~n868 & n884 ;
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  assign n888 = n872 | n887 ;
  buffer buf_n889( .i (n888), .o (n889) );
  assign n890 = n849 & ~n889 ;
  assign n891 = n837 | n890 ;
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n241( .i (G23), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (G24), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  assign n893 = n249 | n258 ;
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  assign n898 = ~n889 & n897 ;
  assign n899 = n837 & n898 ;
  buffer buf_n900( .i (n899), .o (n900) );
  assign n902 = n892 & ~n900 ;
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  assign n904 = n670 & n816 ;
  assign n905 = n670 | n800 ;
  assign n906 = ~n904 & n905 ;
  assign n907 = n335 & n772 ;
  buffer buf_n676( .i (n675), .o (n676) );
  assign n908 = ~n676 & n827 ;
  buffer buf_n230( .i (G22), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n909( .i (n331), .o (n909) );
  assign n910 = n232 & ~n909 ;
  buffer buf_n911( .i (n910), .o (n911) );
  assign n919 = ~n422 & n911 ;
  assign n920 = n908 | n919 ;
  assign n921 = n907 | n920 ;
  assign n922 = n813 & n921 ;
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  assign n926 = n906 | n925 ;
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  assign n929 = n351 & ~n854 ;
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n329( .i (n328), .o (n329) );
  assign n931 = n329 & ~n877 ;
  buffer buf_n932( .i (n419), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  assign n934 = n95 | n933 ;
  buffer buf_n935( .i (n934), .o (n935) );
  assign n936 = ~n344 & n422 ;
  assign n937 = n935 & ~n936 ;
  assign n938 = n931 | n937 ;
  assign n939 = n930 | n938 ;
  assign n940 = ~n868 & n939 ;
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  assign n943 = n872 | n942 ;
  buffer buf_n944( .i (n943), .o (n944) );
  assign n945 = n849 & ~n944 ;
  assign n946 = n928 | n945 ;
  buffer buf_n947( .i (n946), .o (n947) );
  assign n948 = n897 & ~n944 ;
  assign n949 = n928 & n948 ;
  buffer buf_n950( .i (n949), .o (n950) );
  assign n951 = n947 & ~n950 ;
  buffer buf_n952( .i (n951), .o (n952) );
  assign n953 = n903 & n952 ;
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  assign n955 = n337 & n813 ;
  buffer buf_n956( .i (n955), .o (n956) );
  assign n957 = n816 & ~n956 ;
  assign n958 = n89 & ~n957 ;
  assign n959 = ~n86 & n798 ;
  assign n960 = n666 | n824 ;
  buffer buf_n97( .i (n96), .o (n97) );
  assign n961 = ~n97 & n828 ;
  assign n962 = n960 & ~n961 ;
  buffer buf_n963( .i (n812), .o (n963) );
  assign n964 = ~n962 & n963 ;
  assign n965 = n959 | n964 ;
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  assign n968 = n958 | n967 ;
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  assign n971 = n363 & ~n854 ;
  assign n972 = n350 & ~n876 ;
  assign n973 = n121 | n933 ;
  assign n974 = ~n355 & n933 ;
  assign n975 = n973 & ~n974 ;
  assign n976 = n972 | n975 ;
  assign n977 = n971 | n976 ;
  assign n978 = ~n867 & n977 ;
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  assign n982 = n872 | n981 ;
  buffer buf_n983( .i (n982), .o (n983) );
  assign n984 = n849 & ~n983 ;
  assign n985 = n970 | n984 ;
  buffer buf_n986( .i (n985), .o (n986) );
  assign n987 = n897 & ~n983 ;
  assign n988 = n970 & n987 ;
  buffer buf_n989( .i (n988), .o (n989) );
  assign n990 = n986 & ~n989 ;
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  assign n1002 = n800 | n956 ;
  buffer buf_n1003( .i (n1002), .o (n1003) );
  assign n1004 = ~n683 & n1003 ;
  assign n1005 = n653 & ~n824 ;
  assign n1006 = n84 & n828 ;
  assign n1007 = n1005 | n1006 ;
  assign n1008 = n963 & n1007 ;
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  assign n1011 = n681 & ~n816 ;
  assign n1012 = n1010 | n1011 ;
  buffer buf_n1013( .i (n1012), .o (n1013) );
  assign n1014 = n1004 | n1013 ;
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n1016( .i (n853), .o (n1016) );
  assign n1017 = n357 & ~n1016 ;
  buffer buf_n1018( .i (n1017), .o (n1018) );
  assign n1019 = n345 & ~n877 ;
  assign n1020 = n107 | n933 ;
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n932), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  assign n1024 = ~n350 & n1023 ;
  assign n1025 = n1021 & ~n1024 ;
  assign n1026 = n1019 | n1025 ;
  assign n1027 = n1018 | n1026 ;
  assign n1028 = ~n868 & n1027 ;
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  assign n1031 = n872 | n1030 ;
  buffer buf_n1032( .i (n1031), .o (n1032) );
  assign n1033 = n849 & ~n1032 ;
  assign n1034 = n1015 | n1033 ;
  buffer buf_n1035( .i (n1034), .o (n1035) );
  assign n1036 = n897 & ~n1032 ;
  assign n1037 = n1015 & n1036 ;
  buffer buf_n1038( .i (n1037), .o (n1038) );
  assign n1040 = n1035 & ~n1038 ;
  buffer buf_n1041( .i (n1040), .o (n1041) );
  assign n1042 = n991 & n1041 ;
  buffer buf_n1043( .i (n1042), .o (n1043) );
  assign n1044 = n954 & n1043 ;
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  assign n1052 = n96 | n694 ;
  assign n1053 = n335 & n1052 ;
  buffer buf_n1054( .i (n1053), .o (n1054) );
  assign n1055 = n677 | n824 ;
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  assign n1056 = ~n109 & n828 ;
  assign n1057 = n1055 & ~n1056 ;
  assign n1058 = ~n1054 & n1057 ;
  assign n1059 = n814 & ~n1058 ;
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n423( .i (n422), .o (n423) );
  assign n1062 = ~n56 & n423 ;
  assign n1063 = n797 | n1062 ;
  assign n1064 = n963 | n1063 ;
  buffer buf_n1065( .i (n1064), .o (n1065) );
  assign n1066 = n101 & ~n1065 ;
  assign n1067 = ~n101 & n800 ;
  assign n1068 = n1066 | n1067 ;
  assign n1069 = n1061 | n1068 ;
  buffer buf_n1070( .i (n1069), .o (n1070) );
  assign n1071 = n357 & ~n877 ;
  buffer buf_n135( .i (n134), .o (n135) );
  assign n1072 = n135 | n1023 ;
  assign n1073 = ~n362 & n1023 ;
  assign n1074 = n1072 & ~n1073 ;
  assign n1075 = n1071 | n1074 ;
  buffer buf_n638( .i (n637), .o (n638) );
  assign n1076 = n638 | n851 ;
  buffer buf_n1077( .i (n1076), .o (n1077) );
  assign n1078 = n400 | n1077 ;
  assign n1079 = ~n368 & n1077 ;
  assign n1080 = n1078 & ~n1079 ;
  buffer buf_n1081( .i (n1080), .o (n1081) );
  assign n1082 = n1075 | n1081 ;
  assign n1083 = ~n868 & n1082 ;
  buffer buf_n1084( .i (n1083), .o (n1084) );
  assign n1085 = n894 & ~n1084 ;
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  assign n1088 = n1070 & n1087 ;
  buffer buf_n1089( .i (n1088), .o (n1089) );
  assign n1092 = n846 & ~n1084 ;
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  assign n1095 = n1070 | n1094 ;
  buffer buf_n1096( .i (n1095), .o (n1096) );
  assign n1098 = ~n1089 & n1096 ;
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n1101( .i (n799), .o (n1101) );
  assign n1102 = n113 | n1101 ;
  assign n1103 = n113 & n1065 ;
  assign n1104 = n1102 & ~n1103 ;
  assign n1105 = n107 & n121 ;
  assign n1106 = n694 & ~n1105 ;
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  assign n1111 = n956 & n1110 ;
  assign n1112 = ~n334 & n808 ;
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n122( .i (n121), .o (n122) );
  assign n1114 = n122 & n1023 ;
  assign n1115 = n880 | n1114 ;
  assign n1116 = n1113 & n1115 ;
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  assign n1120 = n1111 | n1119 ;
  assign n1121 = n1104 | n1120 ;
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  assign n1124 = n576 | n1077 ;
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  assign n1129 = n870 & ~n1128 ;
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n1131 = n379 & n1125 ;
  buffer buf_n1132( .i (n876), .o (n1132) );
  assign n1133 = n363 & ~n1132 ;
  buffer buf_n404( .i (G39), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n1134( .i (n1022), .o (n1134) );
  assign n1135 = n408 | n1134 ;
  assign n1136 = ~n368 & n1134 ;
  assign n1137 = n1135 & ~n1136 ;
  assign n1138 = n1133 | n1137 ;
  assign n1139 = n1131 | n1138 ;
  buffer buf_n1140( .i (n867), .o (n1140) );
  assign n1141 = n1139 & ~n1140 ;
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  assign n1144 = n1130 | n1143 ;
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n896), .o (n1146) );
  assign n1147 = ~n1145 & n1146 ;
  assign n1148 = n1123 & n1147 ;
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n848), .o (n1150) );
  assign n1151 = ~n1145 & n1150 ;
  assign n1152 = n1123 | n1151 ;
  buffer buf_n1153( .i (n1152), .o (n1153) );
  assign n1154 = ~n1149 & n1153 ;
  buffer buf_n1155( .i (n1154), .o (n1155) );
  assign n1156 = n1100 & n1155 ;
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  assign n1158 = ~n129 & n1003 ;
  assign n1159 = n127 & ~n1065 ;
  assign n1160 = n135 & n1134 ;
  assign n1161 = n935 & ~n1160 ;
  assign n1162 = n1113 & ~n1161 ;
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  assign n1166 = n1159 | n1165 ;
  buffer buf_n1167( .i (n1166), .o (n1167) );
  assign n1168 = n1158 | n1167 ;
  buffer buf_n1169( .i (n1168), .o (n1169) );
  assign n1170 = n387 & n1125 ;
  assign n1171 = n377 & n1134 ;
  buffer buf_n438( .i (G40), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n1172( .i (n1022), .o (n1172) );
  assign n1173 = n442 & ~n1172 ;
  assign n1174 = n1171 | n1173 ;
  assign n1175 = n369 & ~n1132 ;
  assign n1176 = n1174 | n1175 ;
  assign n1177 = n1170 | n1176 ;
  assign n1178 = ~n1140 & n1177 ;
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  assign n1181 = n1130 | n1180 ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  assign n1183 = n1146 & ~n1182 ;
  assign n1184 = n1169 & n1183 ;
  buffer buf_n1185( .i (n1184), .o (n1185) );
  assign n1190 = n1150 & ~n1182 ;
  assign n1191 = n1169 | n1190 ;
  buffer buf_n1192( .i (n1191), .o (n1192) );
  assign n1193 = ~n1185 & n1192 ;
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  assign n1197 = n1157 & n1196 ;
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  assign n1199 = ~n956 & n1065 ;
  assign n1200 = n141 & ~n1199 ;
  assign n1201 = ~n137 & n797 ;
  assign n1202 = n408 & n1172 ;
  assign n1203 = n1021 & ~n1202 ;
  assign n1204 = n1113 & ~n1203 ;
  assign n1205 = n1201 | n1204 ;
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  assign n1209 = n1200 | n1208 ;
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  assign n1212 = n395 & n1125 ;
  assign n1213 = n385 & n1172 ;
  buffer buf_n449( .i (G41), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  assign n1214 = n453 & ~n1172 ;
  assign n1215 = n1213 | n1214 ;
  assign n1216 = n378 & ~n1132 ;
  assign n1217 = n1215 | n1216 ;
  assign n1218 = n1212 | n1217 ;
  assign n1219 = ~n1140 & n1218 ;
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  assign n1222 = n1130 | n1221 ;
  buffer buf_n1223( .i (n1222), .o (n1223) );
  assign n1224 = n1146 & ~n1223 ;
  assign n1225 = n1211 & n1224 ;
  buffer buf_n1226( .i (n1225), .o (n1226) );
  assign n1233 = n1150 & ~n1223 ;
  assign n1234 = n1211 | n1233 ;
  buffer buf_n1235( .i (n1234), .o (n1235) );
  assign n1236 = ~n1226 & n1235 ;
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  assign n1242 = n1198 & n1241 ;
  buffer buf_n1243( .i (n1242), .o (n1243) );
  assign n1244 = n1047 & n1243 ;
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  assign n1245 = n1198 & n1232 ;
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  assign n1246 = n1157 & n1189 ;
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  assign n1247 = n1097 & n1149 ;
  assign n1248 = n1091 | n1247 ;
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  assign n1252 = n1246 | n1251 ;
  buffer buf_n1253( .i (n1252), .o (n1253) );
  assign n1254 = n1245 | n1253 ;
  buffer buf_n1255( .i (n1254), .o (n1255) );
  assign n1256 = n1048 & n1255 ;
  buffer buf_n1039( .i (n1038), .o (n1039) );
  assign n1257 = n989 & n1035 ;
  assign n1258 = n1039 | n1257 ;
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  assign n1261 = n954 & n1260 ;
  buffer buf_n901( .i (n900), .o (n901) );
  assign n1262 = n892 & n950 ;
  assign n1263 = n901 | n1262 ;
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  assign n1267 = n1261 | n1266 ;
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  assign n1275 = n1256 | n1271 ;
  buffer buf_n269( .i (G27), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n522( .i (G48), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  assign n1276 = n276 & n529 ;
  buffer buf_n1277( .i (n1276), .o (n1277) );
  assign n1318 = ~n737 & n1277 ;
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  assign n1334 = n1169 & n1322 ;
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  assign n1338 = n1194 | n1337 ;
  assign n1339 = n1194 & n1337 ;
  assign n1340 = n1338 & ~n1339 ;
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n494( .i (G47), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  assign n1343 = n1210 & n1321 ;
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  assign n1348 = n1237 | n1347 ;
  assign n1349 = n1237 & n1347 ;
  assign n1350 = n1348 & ~n1349 ;
  buffer buf_n1351( .i (n1350), .o (n1351) );
  assign n1352 = n515 & n1351 ;
  assign n1353 = ~n1342 & n1352 ;
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  assign n1360 = n581 & ~n737 ;
  buffer buf_n1361( .i (n1360), .o (n1361) );
  assign n1389 = n730 & ~n1361 ;
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  assign n1406 = n1255 & ~n1333 ;
  buffer buf_n1407( .i (n1406), .o (n1407) );
  assign n1414 = ~n78 & n1407 ;
  assign n1415 = n1405 | n1414 ;
  buffer buf_n1416( .i (n827), .o (n1416) );
  assign n1417 = ~n190 & n1416 ;
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  assign n1433 = n1351 & n1432 ;
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  assign n1434 = ~n647 & n1361 ;
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  assign n1455 = ~n243 & n909 ;
  assign n1456 = n718 & ~n1455 ;
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n263( .i (n262), .o (n263) );
  assign n1470 = n263 & n909 ;
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  assign n1474 = n252 & n909 ;
  buffer buf_n1475( .i (n1474), .o (n1475) );
  assign n1476 = n268 & ~n1475 ;
  buffer buf_n1477( .i (n1476), .o (n1477) );
  assign n1478 = n1473 & n1477 ;
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n470( .i (G43), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  assign n1484 = n412 | n478 ;
  buffer buf_n1485( .i (n1484), .o (n1485) );
  assign n1486 = ~n1481 & n1485 ;
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  assign n1487 = ~n339 & n458 ;
  assign n1488 = n428 & ~n1487 ;
  assign n1489 = ~n1486 & n1488 ;
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  assign n1490 = n253 | n839 ;
  assign n1491 = n334 & n1490 ;
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  assign n1494 = n445 & n1493 ;
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n481( .i (G44), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  assign n1497 = n268 | n1475 ;
  buffer buf_n1498( .i (n1497), .o (n1498) );
  assign n1499 = n1473 | n1498 ;
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  assign n1502 = n490 & n1501 ;
  assign n1503 = n1496 | n1502 ;
  assign n1504 = ~n1473 & n1477 ;
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n491( .i (G45), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  assign n1508 = n450 | n492 ;
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  assign n1516 = ~n1506 & n1515 ;
  assign n1517 = n1473 & ~n1498 ;
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n460( .i (G42), .o (n460) );
  buffer buf_n493( .i (G46), .o (n493) );
  assign n1523 = n460 | n493 ;
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  assign n1532 = ~n1519 & n1531 ;
  assign n1533 = n1516 | n1532 ;
  assign n1534 = n1503 | n1533 ;
  assign n1535 = n1489 & ~n1534 ;
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  assign n1538 = n338 & n1505 ;
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  assign n1543 = n103 | n1540 ;
  buffer buf_n1544( .i (n1543), .o (n1544) );
  assign n1545 = n127 | n1480 ;
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  assign n1549 = n1544 & n1548 ;
  assign n1550 = n681 | n1480 ;
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  assign n1552 = n658 | n1507 ;
  assign n1553 = n1551 & n1552 ;
  buffer buf_n1520( .i (n1519), .o (n1520) );
  assign n1554 = n89 | n1520 ;
  assign n1555 = ~n670 & n1501 ;
  buffer buf_n1556( .i (n1555), .o (n1556) );
  assign n1557 = n1554 & ~n1556 ;
  assign n1558 = n1553 & n1557 ;
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  assign n1559 = n239 & ~n1519 ;
  assign n1560 = n428 | n1559 ;
  buffer buf_n1561( .i (n1560), .o (n1561) );
  assign n1562 = ~n111 & n1493 ;
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  assign n1567 = n1561 | n1566 ;
  assign n1568 = n1558 & ~n1567 ;
  assign n1569 = n1549 & n1568 ;
  assign n1570 = n1537 | n1569 ;
  assign n1571 = ~n1468 & n1570 ;
  assign n1572 = n1439 & ~n1571 ;
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  assign n1577 = ~n1433 & n1576 ;
  buffer buf_n1578( .i (n1577), .o (n1578) );
  assign n1579 = n515 & ~n1351 ;
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  assign n1583 = ~n515 & n1351 ;
  assign n1584 = n1444 | n1583 ;
  assign n1585 = n1580 | n1584 ;
  assign n1586 = ~n1578 & n1585 ;
  buffer buf_n1587( .i (n1586), .o (n1587) );
  inverter inv_n2635( .i (n1587), .o (n2635) );
  assign n1596 = n969 & n1321 ;
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  assign n1601 = n991 | n1600 ;
  assign n1602 = n991 & n1600 ;
  assign n1603 = n1601 & ~n1602 ;
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  assign n1613 = ~n204 & n437 ;
  buffer buf_n1614( .i (n1613), .o (n1614) );
  assign n1615 = n1604 & n1614 ;
  buffer buf_n205( .i (G20), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n1616 = n214 & n1501 ;
  assign n1617 = ~n668 & n1493 ;
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n175( .i (G19), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  assign n1619 = n183 & ~n1505 ;
  assign n1620 = n1618 | n1619 ;
  assign n1621 = n1616 | n1620 ;
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  assign n1625 = n660 | n1541 ;
  buffer buf_n165( .i (G18), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  assign n1626 = n174 & ~n1519 ;
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  assign n1627 = ~n226 & n680 ;
  assign n1628 = n1480 | n1627 ;
  assign n1629 = ~n1626 & n1628 ;
  buffer buf_n1630( .i (n1629), .o (n1630) );
  assign n1631 = ~n1561 & n1630 ;
  assign n1632 = n1625 & n1631 ;
  assign n1633 = ~n1624 & n1632 ;
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  assign n1634 = n447 & n1501 ;
  assign n1635 = n1564 | n1634 ;
  assign n1636 = n458 & ~n1506 ;
  assign n1637 = n99 & ~n411 ;
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1640( .i (n1479), .o (n1640) );
  assign n1641 = n1638 | n1640 ;
  assign n1642 = ~n1636 & n1641 ;
  assign n1643 = ~n1635 & n1642 ;
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n130( .i (n129), .o (n130) );
  assign n1646 = n130 | n1541 ;
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  assign n1647 = n138 & ~n467 ;
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1518), .o (n1649) );
  assign n1650 = n1648 | n1649 ;
  assign n1651 = n428 & n1650 ;
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  assign n1654 = n1646 & n1653 ;
  assign n1655 = n1645 & n1654 ;
  assign n1656 = n1633 | n1655 ;
  assign n1657 = ~n1468 & n1656 ;
  assign n1658 = n1439 & ~n1657 ;
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  assign n1663 = ~n1615 & n1662 ;
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  assign n1675 = n1179 | n1220 ;
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  assign n1676 = n260 | n1084 ;
  assign n1677 = n1675 | n1676 ;
  buffer buf_n1678( .i (n1677), .o (n1678) );
  assign n1679 = n1145 | n1678 ;
  buffer buf_n1680( .i (n1679), .o (n1680) );
  assign n1681 = n1182 & n1223 ;
  assign n1682 = n260 & n1084 ;
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  assign n1685 = n1145 & n1684 ;
  assign n1686 = n1681 & n1685 ;
  assign n1687 = n1680 & ~n1686 ;
  assign n1688 = n1324 | n1687 ;
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  assign n1697 = n1243 & n1332 ;
  assign n1698 = n1696 & ~n1697 ;
  buffer buf_n1699( .i (n1698), .o (n1699) );
  assign n1700 = n521 & ~n1699 ;
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  assign n1704 = ~n1407 & n1610 ;
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  assign n1706 = ~n1001 & n1408 ;
  assign n1707 = n1705 | n1706 ;
  buffer buf_n1708( .i (n1707), .o (n1708) );
  assign n1709 = n1703 | n1708 ;
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  assign n1711 = n1703 & n1708 ;
  assign n1712 = n1454 | n1711 ;
  assign n1713 = n1710 & ~n1712 ;
  assign n1714 = n1674 | n1713 ;
  buffer buf_n1715( .i (n1714), .o (n1715) );
  assign n1723 = n521 & n1699 ;
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  assign n1727 = n1015 & n1322 ;
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  assign n1731 = n1041 & ~n1730 ;
  assign n1732 = ~n1041 & n1730 ;
  assign n1733 = n1731 | n1732 ;
  buffer buf_n1734( .i (n1733), .o (n1734) );
  assign n1744 = n1604 & n1734 ;
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  assign n1752 = n278 & ~n737 ;
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  assign n1759 = n927 & n1755 ;
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  assign n1764 = n952 | n1763 ;
  assign n1765 = n952 & n1763 ;
  assign n1766 = n1764 & ~n1765 ;
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  assign n1771 = n1745 & n1769 ;
  buffer buf_n1772( .i (n1771), .o (n1772) );
  assign n1778 = n1048 & n1772 ;
  assign n1779 = n1048 | n1772 ;
  assign n1780 = ~n1778 & n1779 ;
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  assign n1784 = n1725 & ~n1783 ;
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  assign n1788 = n1051 | n1408 ;
  assign n1789 = ~n1274 & n1788 ;
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  assign n1791 = n1038 & ~n1324 ;
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  assign n1797 = n989 & ~n1324 ;
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  assign n1810 = n1734 & ~n1801 ;
  assign n1811 = n1796 | n1810 ;
  buffer buf_n1812( .i (n1811), .o (n1812) );
  assign n1813 = n1770 & n1812 ;
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  assign n1815 = n950 & ~n1758 ;
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  buffer buf_n1821( .i (n1820), .o (n1821) );
  buffer buf_n1822( .i (n1821), .o (n1822) );
  buffer buf_n1823( .i (n1822), .o (n1823) );
  buffer buf_n1824( .i (n1823), .o (n1824) );
  assign n1825 = n1814 | n1824 ;
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  assign n1830 = n1790 & n1829 ;
  assign n1831 = n1790 | n1829 ;
  assign n1832 = ~n1830 & n1831 ;
  buffer buf_n1833( .i (n1832), .o (n1833) );
  assign n1834 = n1787 & n1833 ;
  assign n1835 = n1787 | n1833 ;
  assign n1836 = ~n1834 & n1835 ;
  assign n1837 = n56 | n190 ;
  buffer buf_n1838( .i (n1837), .o (n1838) );
  assign n1839 = n697 & n1838 ;
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  buffer buf_n1846( .i (n1845), .o (n1846) );
  buffer buf_n1847( .i (n1846), .o (n1847) );
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  assign n1868 = ~n1836 & n1867 ;
  assign n1869 = n653 & ~n677 ;
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  assign n1870 = n691 | n772 ;
  assign n1871 = ~n1869 & n1870 ;
  assign n1872 = n1838 | n1871 ;
  assign n1873 = ~n136 & n722 ;
  assign n1874 = ~n1107 & n1873 ;
  buffer buf_n1875( .i (n1874), .o (n1875) );
  assign n1876 = n1872 & ~n1875 ;
  buffer buf_n1877( .i (n1876), .o (n1877) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  buffer buf_n1879( .i (n1878), .o (n1879) );
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n1888( .i (n1887), .o (n1888) );
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  assign n1905 = n1868 | ~n1904 ;
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  assign n1906 = ~n803 & n1077 ;
  assign n1907 = ~n720 & n1906 ;
  buffer buf_n1908( .i (n1907), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n1915( .i (n1914), .o (n1915) );
  buffer buf_n1916( .i (n1915), .o (n1916) );
  buffer buf_n1917( .i (n1916), .o (n1917) );
  buffer buf_n1918( .i (n1917), .o (n1918) );
  buffer buf_n1919( .i (n1918), .o (n1919) );
  buffer buf_n1920( .i (n1919), .o (n1920) );
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  buffer buf_n1930( .i (n1929), .o (n1930) );
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n1934( .i (n1933), .o (n1934) );
  buffer buf_n1935( .i (n1934), .o (n1935) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n1941( .i (n1323), .o (n1941) );
  assign n1942 = n1226 & ~n1941 ;
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  assign n1947 = n1341 | n1946 ;
  buffer buf_n1948( .i (n1947), .o (n1948) );
  assign n1949 = n1194 & n1943 ;
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  assign n1954 = n1948 & ~n1953 ;
  buffer buf_n1955( .i (n1954), .o (n1955) );
  assign n1956 = n1582 | n1955 ;
  assign n1957 = n1582 & n1955 ;
  assign n1958 = n1956 & ~n1957 ;
  buffer buf_n1959( .i (n1958), .o (n1959) );
  assign n1960 = n1408 & n1959 ;
  assign n1961 = n1379 | n1960 ;
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  assign n1966 = n1122 & n1321 ;
  buffer buf_n1967( .i (n1966), .o (n1967) );
  buffer buf_n1968( .i (n1967), .o (n1968) );
  buffer buf_n1969( .i (n1968), .o (n1969) );
  buffer buf_n1970( .i (n1969), .o (n1970) );
  assign n1971 = n1155 | n1970 ;
  assign n1972 = n1155 & n1970 ;
  assign n1973 = n1971 & ~n1972 ;
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  assign n1979 = n1185 & ~n1941 ;
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  buffer buf_n1983( .i (n1982), .o (n1983) );
  buffer buf_n1984( .i (n1983), .o (n1984) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  assign n1986 = n1948 & ~n1985 ;
  buffer buf_n1987( .i (n1986), .o (n1987) );
  assign n1988 = n1978 | n1987 ;
  buffer buf_n1989( .i (n1988), .o (n1989) );
  assign n1990 = n1978 & n1987 ;
  buffer buf_n1991( .i (n1990), .o (n1991) );
  assign n1992 = n1989 & ~n1991 ;
  buffer buf_n1993( .i (n1992), .o (n1993) );
  assign n1994 = ~n1359 & n1993 ;
  buffer buf_n1995( .i (n1994), .o (n1995) );
  assign n1996 = n1359 & ~n1993 ;
  buffer buf_n1997( .i (n1996), .o (n1997) );
  assign n1999 = n1995 | n1997 ;
  buffer buf_n2000( .i (n1999), .o (n2000) );
  assign n2001 = n1413 & ~n2000 ;
  assign n2002 = n1965 | n2001 ;
  assign n2003 = ~n1936 & n2002 ;
  buffer buf_n1998( .i (n1997), .o (n1998) );
  assign n2004 = n1149 & ~n1941 ;
  buffer buf_n2005( .i (n2004), .o (n2005) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n2007( .i (n2006), .o (n2007) );
  buffer buf_n2008( .i (n2007), .o (n2008) );
  buffer buf_n2009( .i (n2008), .o (n2009) );
  buffer buf_n2010( .i (n2009), .o (n2010) );
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n2012( .i (n2011), .o (n2012) );
  buffer buf_n2013( .i (n2012), .o (n2013) );
  buffer buf_n2014( .i (n2013), .o (n2014) );
  assign n2015 = n1989 & ~n2014 ;
  buffer buf_n2016( .i (n2015), .o (n2016) );
  buffer buf_n2017( .i (n1320), .o (n2017) );
  assign n2018 = n1070 & n2017 ;
  buffer buf_n2019( .i (n2018), .o (n2019) );
  buffer buf_n2020( .i (n2019), .o (n2020) );
  buffer buf_n2021( .i (n2020), .o (n2021) );
  assign n2022 = n1099 | n2021 ;
  assign n2023 = n1099 & n2021 ;
  assign n2024 = n2022 & ~n2023 ;
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2028( .i (n2027), .o (n2028) );
  buffer buf_n2029( .i (n2028), .o (n2029) );
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n2031( .i (n2030), .o (n2031) );
  buffer buf_n2032( .i (n2031), .o (n2032) );
  buffer buf_n2033( .i (n2032), .o (n2033) );
  buffer buf_n2034( .i (n2033), .o (n2034) );
  assign n2035 = n2016 & ~n2034 ;
  assign n2036 = ~n2016 & n2034 ;
  assign n2037 = n2035 | n2036 ;
  buffer buf_n2038( .i (n2037), .o (n2038) );
  assign n2039 = n1998 & ~n2038 ;
  assign n2040 = ~n1998 & n2038 ;
  assign n2041 = n2039 | n2040 ;
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  assign n2044 = ~n2003 & n2043 ;
  assign n2045 = n1431 & n2025 ;
  assign n2046 = ~n182 & n655 ;
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  assign n2049 = n1520 | n2048 ;
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n2050( .i (n1500), .o (n2050) );
  assign n2051 = n227 & n2050 ;
  assign n2052 = n214 & ~n1506 ;
  assign n2053 = n2051 | n2052 ;
  assign n2054 = n2049 & ~n2053 ;
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n240( .i (n239), .o (n240) );
  assign n2055 = n89 & ~n240 ;
  assign n2056 = n1482 | n2055 ;
  assign n2057 = n2054 & n2056 ;
  assign n2058 = ~n679 & n1493 ;
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n671( .i (n670), .o (n671) );
  assign n2062 = n671 | n1539 ;
  assign n2063 = ~n2061 & n2062 ;
  assign n2064 = ~n430 & n2063 ;
  assign n2065 = n2057 & n2064 ;
  assign n2066 = n1485 & ~n1520 ;
  assign n2067 = n112 & ~n446 ;
  buffer buf_n2068( .i (n2067), .o (n2068) );
  assign n2069 = n1481 | n2068 ;
  assign n2070 = ~n2066 & n2069 ;
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n2072( .i (n1505), .o (n2072) );
  assign n2073 = n469 & ~n2072 ;
  assign n2074 = n458 & n2050 ;
  assign n2075 = n2073 | n2074 ;
  buffer buf_n2076( .i (n2075), .o (n2076) );
  assign n2077 = n141 | n1539 ;
  buffer buf_n2078( .i (n1492), .o (n2078) );
  assign n2079 = ~n125 & n2078 ;
  assign n2080 = n426 & ~n2079 ;
  buffer buf_n2081( .i (n2080), .o (n2081) );
  buffer buf_n2082( .i (n2081), .o (n2082) );
  assign n2083 = n2077 & n2082 ;
  assign n2084 = ~n2076 & n2083 ;
  assign n2085 = n2071 & n2084 ;
  assign n2086 = n2065 | n2085 ;
  assign n2087 = ~n1467 & n2086 ;
  assign n2088 = n1438 & ~n2087 ;
  buffer buf_n2089( .i (n2088), .o (n2089) );
  buffer buf_n2090( .i (n2089), .o (n2090) );
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  assign n2093 = ~n2045 & n2092 ;
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n2099( .i (n2098), .o (n2099) );
  buffer buf_n2100( .i (n2099), .o (n2100) );
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n2102( .i (n2101), .o (n2102) );
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  assign n2109 = n2044 | n2108 ;
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n2111( .i (n1407), .o (n2111) );
  assign n2112 = n1959 | n2111 ;
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  assign n2115 = ~n1962 & n2114 ;
  assign n2116 = n1929 & ~n1959 ;
  assign n2117 = n1341 & n1432 ;
  buffer buf_n1469( .i (n1468), .o (n1469) );
  assign n2118 = n411 & n2078 ;
  buffer buf_n2119( .i (n2118), .o (n2119) );
  buffer buf_n2120( .i (n2119), .o (n2120) );
  assign n2121 = n490 & ~n2072 ;
  assign n2122 = n2120 | n2121 ;
  assign n2123 = n1515 & ~n1649 ;
  buffer buf_n479( .i (n478), .o (n479) );
  assign n2124 = n479 & n2050 ;
  assign n2125 = n2123 | n2124 ;
  assign n2126 = n2122 | n2125 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n2127 = n448 & ~n1539 ;
  assign n2128 = n1640 | n1648 ;
  buffer buf_n2129( .i (n427), .o (n2129) );
  assign n2130 = n2128 & n2129 ;
  assign n2131 = ~n2127 & n2130 ;
  assign n2132 = ~n2126 & n2131 ;
  buffer buf_n2133( .i (n2132), .o (n2133) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  assign n2136 = ~n657 & n2050 ;
  buffer buf_n2137( .i (n2136), .o (n2137) );
  assign n2138 = n240 & ~n1507 ;
  assign n2139 = n2137 | n2138 ;
  assign n2140 = n113 | n1640 ;
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n1649), .o (n2142) );
  assign n2143 = n682 | n2142 ;
  assign n2144 = n2141 & n2143 ;
  assign n2145 = ~n2139 & n2144 ;
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  assign n2148 = n91 | n1541 ;
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n2150( .i (n669), .o (n2150) );
  assign n2151 = n1640 | n2150 ;
  assign n2152 = ~n2129 & n2151 ;
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  assign n2155 = ~n99 & n2078 ;
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n2158( .i (n2157), .o (n2158) );
  buffer buf_n2159( .i (n2158), .o (n2159) );
  buffer buf_n228( .i (n227), .o (n228) );
  assign n2160 = n228 & ~n2142 ;
  buffer buf_n2161( .i (n2160), .o (n2161) );
  assign n2162 = n2159 | n2161 ;
  assign n2163 = n2154 & ~n2162 ;
  assign n2164 = n2149 & n2163 ;
  assign n2165 = n2147 & n2164 ;
  assign n2166 = n2135 | n2165 ;
  assign n2167 = ~n1469 & n2166 ;
  assign n2168 = n1440 & ~n2167 ;
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  buffer buf_n2171( .i (n2170), .o (n2171) );
  assign n2172 = ~n2117 & n2171 ;
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n2175( .i (n2174), .o (n2175) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n2177), .o (n2178) );
  assign n2179 = n2116 | n2178 ;
  buffer buf_n2180( .i (n2179), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  assign n2182 = n2115 | n2181 ;
  buffer buf_n2183( .i (n2182), .o (n2183) );
  buffer buf_n1380( .i (n1379), .o (n1380) );
  assign n2184 = ~n1380 & n2113 ;
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  assign n2187 = ~n2000 & n2186 ;
  buffer buf_n2188( .i (n2187), .o (n2188) );
  assign n2189 = n1432 & n1974 ;
  assign n2190 = n228 & ~n1507 ;
  assign n2191 = n1649 | n2150 ;
  assign n2192 = n100 & n656 ;
  buffer buf_n2193( .i (n1479), .o (n2193) );
  assign n2194 = n2192 | n2193 ;
  assign n2195 = n2191 & n2194 ;
  assign n2196 = ~n2190 & n2195 ;
  buffer buf_n2197( .i (n2196), .o (n2197) );
  buffer buf_n2198( .i (n2197), .o (n2198) );
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  assign n2200 = n685 | n1542 ;
  buffer buf_n215( .i (n214), .o (n215) );
  assign n2201 = n215 & ~n2142 ;
  assign n2202 = n429 | n2201 ;
  buffer buf_n2203( .i (n2202), .o (n2203) );
  assign n2204 = ~n86 & n2078 ;
  buffer buf_n2205( .i (n2204), .o (n2205) );
  buffer buf_n2206( .i (n2205), .o (n2206) );
  buffer buf_n2208( .i (n1500), .o (n2208) );
  assign n2209 = n239 & n2208 ;
  assign n2210 = n2206 | n2209 ;
  buffer buf_n2211( .i (n2210), .o (n2211) );
  buffer buf_n2212( .i (n2211), .o (n2212) );
  assign n2213 = n2203 | n2212 ;
  assign n2214 = n2200 & ~n2213 ;
  assign n2215 = n2199 & n2214 ;
  assign n2216 = n469 & n2208 ;
  buffer buf_n2217( .i (n2216), .o (n2217) );
  assign n2218 = n447 | n490 ;
  assign n2219 = ~n2142 & n2218 ;
  assign n2220 = n2217 | n2219 ;
  buffer buf_n480( .i (n479), .o (n480) );
  assign n2221 = n480 & ~n1507 ;
  buffer buf_n2222( .i (n1492), .o (n2222) );
  assign n2223 = ~n138 & n2222 ;
  buffer buf_n2224( .i (n2223), .o (n2224) );
  buffer buf_n2225( .i (n2224), .o (n2225) );
  buffer buf_n2226( .i (n2225), .o (n2226) );
  assign n2227 = n2221 | n2226 ;
  assign n2228 = n2220 | n2227 ;
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  assign n2231 = n417 & ~n1542 ;
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n459( .i (n458), .o (n459) );
  assign n2232 = n128 & ~n459 ;
  buffer buf_n2233( .i (n2232), .o (n2233) );
  assign n2234 = n1483 | n2233 ;
  assign n2235 = n431 & n2234 ;
  assign n2236 = ~n2231 & n2235 ;
  assign n2237 = ~n2230 & n2236 ;
  assign n2238 = n2215 | n2237 ;
  assign n2239 = ~n1469 & n2238 ;
  assign n2240 = n1440 & ~n2239 ;
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  assign n2244 = ~n2189 & n2243 ;
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  buffer buf_n2250( .i (n2249), .o (n2250) );
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  assign n2256 = n1380 | n2113 ;
  assign n2257 = ~n1932 & n2256 ;
  buffer buf_n2258( .i (n2257), .o (n2258) );
  assign n2259 = n2000 & ~n2258 ;
  assign n2260 = n2255 | n2259 ;
  assign n2261 = n2188 | n2260 ;
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  assign n2265 = n1725 & n1777 ;
  buffer buf_n2266( .i (n2265), .o (n2266) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  assign n2267 = n1724 & n1751 ;
  buffer buf_n2268( .i (n2267), .o (n2268) );
  assign n2269 = n1770 | n1812 ;
  buffer buf_n2270( .i (n2269), .o (n2270) );
  assign n2271 = ~n1814 & n2270 ;
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2273( .i (n2272), .o (n2273) );
  buffer buf_n2274( .i (n2273), .o (n2274) );
  buffer buf_n2275( .i (n2274), .o (n2275) );
  assign n2276 = ~n2268 & n2275 ;
  assign n2277 = n2266 | n2276 ;
  buffer buf_n2278( .i (n2277), .o (n2278) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  buffer buf_n2280( .i (n2279), .o (n2280) );
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  assign n2285 = n1705 | n1809 ;
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  assign n2289 = n1612 & n1724 ;
  assign n2290 = n1743 | n2289 ;
  assign n2291 = ~n2268 & n2290 ;
  buffer buf_n2292( .i (n2291), .o (n2292) );
  assign n2293 = n2288 | n2292 ;
  assign n2294 = n2288 & n2292 ;
  assign n2295 = n2293 & ~n2294 ;
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  assign n2297 = n1726 & ~n1790 ;
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  buffer buf_n2301( .i (n2300), .o (n2301) );
  assign n2302 = n2296 | n2301 ;
  buffer buf_n2303( .i (n2302), .o (n2303) );
  assign n2304 = n1388 | n2303 ;
  assign n2305 = ~n1940 & n2304 ;
  assign n2306 = n2284 & ~n2305 ;
  buffer buf_n2307( .i (n2306), .o (n2307) );
  assign n2308 = ~n1388 & n2303 ;
  buffer buf_n2309( .i (n2308), .o (n2309) );
  assign n2310 = ~n2284 & n2309 ;
  assign n2311 = n1614 & n1767 ;
  buffer buf_n2312( .i (n1518), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  assign n2314 = n2068 | n2313 ;
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  assign n2317 = n1544 & n2316 ;
  assign n2318 = ~n140 & n2208 ;
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n2207( .i (n2206), .o (n2207) );
  assign n2321 = n1551 & ~n2207 ;
  assign n2322 = ~n2320 & n2321 ;
  buffer buf_n2323( .i (n2072), .o (n2323) );
  assign n2324 = n414 & ~n2323 ;
  buffer buf_n2325( .i (n2324), .o (n2325) );
  assign n2326 = n429 & n1546 ;
  assign n2327 = ~n2325 & n2326 ;
  assign n2328 = n2322 & n2327 ;
  assign n2329 = n2317 & n2328 ;
  buffer buf_n143( .i (G16), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  assign n2330 = n153 & ~n2313 ;
  buffer buf_n2331( .i (n2330), .o (n2331) );
  buffer buf_n154( .i (G17), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  assign n2332 = n164 & ~n2323 ;
  assign n2333 = n237 & n2222 ;
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n2335( .i (n2334), .o (n2335) );
  buffer buf_n2336( .i (n2335), .o (n2336) );
  assign n2337 = n2332 | n2336 ;
  assign n2338 = n2331 | n2337 ;
  buffer buf_n2339( .i (n2338), .o (n2339) );
  buffer buf_n229( .i (n228), .o (n229) );
  assign n2340 = n229 & ~n1540 ;
  assign n2341 = n174 & n2208 ;
  assign n2342 = n2047 | n2193 ;
  assign n2343 = ~n2341 & n2342 ;
  buffer buf_n2344( .i (n2343), .o (n2344) );
  assign n2345 = ~n2340 & n2344 ;
  assign n2346 = ~n2203 & n2345 ;
  assign n2347 = ~n2339 & n2346 ;
  assign n2348 = n2329 | n2347 ;
  assign n2349 = ~n1468 & n2348 ;
  assign n2350 = n1439 & ~n2349 ;
  buffer buf_n2351( .i (n2350), .o (n2351) );
  buffer buf_n2352( .i (n2351), .o (n2352) );
  buffer buf_n2353( .i (n2352), .o (n2353) );
  buffer buf_n2354( .i (n2353), .o (n2354) );
  assign n2355 = ~n2311 & n2354 ;
  buffer buf_n2356( .i (n2355), .o (n2356) );
  buffer buf_n2357( .i (n2356), .o (n2357) );
  buffer buf_n2358( .i (n2357), .o (n2358) );
  buffer buf_n2359( .i (n2358), .o (n2359) );
  buffer buf_n2360( .i (n2359), .o (n2360) );
  buffer buf_n2361( .i (n2360), .o (n2361) );
  buffer buf_n2362( .i (n2361), .o (n2362) );
  buffer buf_n2363( .i (n2362), .o (n2363) );
  buffer buf_n2364( .i (n2363), .o (n2364) );
  buffer buf_n2365( .i (n2364), .o (n2365) );
  buffer buf_n2366( .i (n2365), .o (n2366) );
  buffer buf_n2367( .i (n2366), .o (n2367) );
  buffer buf_n2368( .i (n2367), .o (n2368) );
  buffer buf_n2369( .i (n2368), .o (n2369) );
  buffer buf_n2370( .i (n2369), .o (n2370) );
  buffer buf_n2371( .i (n2370), .o (n2371) );
  buffer buf_n2372( .i (n2371), .o (n2372) );
  buffer buf_n2373( .i (n2372), .o (n2373) );
  assign n2374 = n2310 | n2373 ;
  assign n2375 = n2307 | n2374 ;
  buffer buf_n2376( .i (n2375), .o (n2376) );
  assign n2377 = n836 & n1755 ;
  buffer buf_n2378( .i (n2377), .o (n2378) );
  buffer buf_n2379( .i (n2378), .o (n2379) );
  buffer buf_n2380( .i (n2379), .o (n2380) );
  buffer buf_n2381( .i (n2380), .o (n2381) );
  assign n2382 = n903 | n2381 ;
  assign n2383 = n903 & n2381 ;
  assign n2384 = n2382 & ~n2383 ;
  buffer buf_n2385( .i (n2384), .o (n2385) );
  assign n2393 = n1614 & n2385 ;
  assign n2394 = n173 | n238 ;
  buffer buf_n2395( .i (n2394), .o (n2395) );
  assign n2396 = ~n1481 & n2395 ;
  buffer buf_n2397( .i (n2396), .o (n2397) );
  buffer buf_n2398( .i (n2397), .o (n2398) );
  buffer buf_n2399( .i (n2398), .o (n2399) );
  buffer buf_n2400( .i (n2399), .o (n2400) );
  assign n2401 = n153 & ~n2323 ;
  buffer buf_n2402( .i (n2401), .o (n2402) );
  buffer buf_n2403( .i (n2402), .o (n2403) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n2404( .i (n1540), .o (n2404) );
  assign n2405 = n217 & ~n2404 ;
  assign n2406 = n2403 | n2405 ;
  buffer buf_n2407( .i (n1500), .o (n2407) );
  assign n2408 = n163 & n2407 ;
  buffer buf_n142( .i (G15), .o (n142) );
  assign n2409 = n142 | n175 ;
  buffer buf_n2410( .i (n2409), .o (n2410) );
  buffer buf_n2411( .i (n2410), .o (n2411) );
  buffer buf_n2412( .i (n2411), .o (n2412) );
  buffer buf_n2413( .i (n2412), .o (n2413) );
  buffer buf_n2414( .i (n2413), .o (n2414) );
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n2416( .i (n2415), .o (n2416) );
  buffer buf_n2417( .i (n2416), .o (n2417) );
  assign n2418 = ~n2312 & n2417 ;
  assign n2419 = n2408 | n2418 ;
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  assign n2420 = n225 & n2222 ;
  assign n2421 = n864 & ~n2420 ;
  buffer buf_n2422( .i (n2421), .o (n2422) );
  buffer buf_n2423( .i (n2422), .o (n2423) );
  assign n2424 = ~n2419 & n2423 ;
  buffer buf_n2425( .i (n2424), .o (n2425) );
  buffer buf_n2426( .i (n2425), .o (n2426) );
  assign n2427 = ~n2406 & n2426 ;
  assign n2428 = ~n2400 & n2427 ;
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  assign n2429 = n586 & n2149 ;
  assign n2430 = n141 | n2323 ;
  assign n2431 = ~n2061 & n2430 ;
  assign n2432 = ~n127 & n2407 ;
  buffer buf_n2433( .i (n2432), .o (n2433) );
  assign n2434 = n2141 & ~n2433 ;
  assign n2435 = n2431 & n2434 ;
  buffer buf_n1639( .i (n1638), .o (n1639) );
  assign n2436 = n1639 | n2313 ;
  buffer buf_n2437( .i (n2436), .o (n2437) );
  assign n2438 = n2153 & n2437 ;
  assign n2439 = n2435 & n2438 ;
  buffer buf_n2440( .i (n2439), .o (n2440) );
  assign n2441 = n2429 & n2440 ;
  assign n2442 = n2428 | n2441 ;
  assign n2443 = ~n1469 & n2442 ;
  assign n2444 = n1440 & ~n2443 ;
  buffer buf_n2445( .i (n2444), .o (n2445) );
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  assign n2448 = ~n2393 & n2447 ;
  buffer buf_n2449( .i (n2448), .o (n2449) );
  buffer buf_n2450( .i (n2449), .o (n2450) );
  buffer buf_n2451( .i (n2450), .o (n2451) );
  buffer buf_n2452( .i (n2451), .o (n2452) );
  buffer buf_n2453( .i (n2452), .o (n2453) );
  buffer buf_n2454( .i (n2453), .o (n2454) );
  buffer buf_n2455( .i (n2454), .o (n2455) );
  buffer buf_n2456( .i (n2455), .o (n2456) );
  buffer buf_n2457( .i (n2456), .o (n2457) );
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n2460( .i (n2459), .o (n2460) );
  buffer buf_n2461( .i (n2460), .o (n2461) );
  buffer buf_n2462( .i (n2461), .o (n2462) );
  buffer buf_n2463( .i (n2462), .o (n2463) );
  buffer buf_n2464( .i (n2463), .o (n2464) );
  buffer buf_n2465( .i (n2464), .o (n2465) );
  buffer buf_n2466( .i (n2465), .o (n2466) );
  assign n2467 = n2296 & n2301 ;
  buffer buf_n2468( .i (n2467), .o (n2468) );
  assign n2471 = ~n2278 & n2299 ;
  assign n2472 = n1385 | n2471 ;
  buffer buf_n2473( .i (n2472), .o (n2473) );
  buffer buf_n2474( .i (n2473), .o (n2474) );
  assign n2475 = n2468 | n2474 ;
  assign n2476 = ~n1940 & n2475 ;
  buffer buf_n2386( .i (n2385), .o (n2386) );
  buffer buf_n2387( .i (n2386), .o (n2387) );
  buffer buf_n2388( .i (n2387), .o (n2388) );
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2391( .i (n2390), .o (n2391) );
  buffer buf_n2392( .i (n2391), .o (n2392) );
  assign n2477 = n1826 & ~n2392 ;
  assign n2478 = ~n1826 & n2392 ;
  assign n2479 = n2477 | n2478 ;
  buffer buf_n2480( .i (n2479), .o (n2480) );
  buffer buf_n2481( .i (n2480), .o (n2481) );
  assign n2482 = n2266 & ~n2481 ;
  assign n2483 = ~n2266 & n2481 ;
  assign n2484 = n2482 | n2483 ;
  buffer buf_n2485( .i (n2484), .o (n2485) );
  buffer buf_n2486( .i (n2485), .o (n2486) );
  buffer buf_n2487( .i (n2486), .o (n2487) );
  buffer buf_n2488( .i (n2487), .o (n2488) );
  buffer buf_n2489( .i (n2488), .o (n2489) );
  buffer buf_n2490( .i (n2489), .o (n2490) );
  assign n2491 = ~n2476 & n2490 ;
  assign n2492 = n2466 | n2491 ;
  buffer buf_n2493( .i (n2492), .o (n2493) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  buffer buf_n2470( .i (n2469), .o (n2470) );
  assign n2495 = n2309 & ~n2470 ;
  assign n2496 = n1614 & n1734 ;
  assign n2497 = n413 & n2407 ;
  buffer buf_n2498( .i (n2497), .o (n2498) );
  buffer buf_n2499( .i (n2072), .o (n2499) );
  assign n2500 = n448 & ~n2499 ;
  assign n2501 = n2498 | n2500 ;
  assign n2502 = n87 & n139 ;
  assign n2503 = n2193 | n2502 ;
  assign n2504 = ~n2157 & n2503 ;
  buffer buf_n2505( .i (n2504), .o (n2505) );
  assign n2506 = ~n2501 & n2505 ;
  buffer buf_n2507( .i (n2506), .o (n2507) );
  buffer buf_n2508( .i (n2507), .o (n2508) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  assign n2509 = n117 | n1542 ;
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n1522( .i (n1521), .o (n1522) );
  assign n2510 = n1522 | n2233 ;
  assign n2511 = n431 & n2510 ;
  assign n2512 = n2509 & n2511 ;
  assign n2513 = n2508 & n2512 ;
  assign n2514 = n164 & ~n2313 ;
  buffer buf_n2515( .i (n2514), .o (n2515) );
  buffer buf_n2516( .i (n2515), .o (n2516) );
  buffer buf_n184( .i (n183), .o (n184) );
  assign n2517 = n184 & n2407 ;
  buffer buf_n2518( .i (n2517), .o (n2518) );
  buffer buf_n2519( .i (n2518), .o (n2519) );
  assign n2520 = n2161 | n2519 ;
  assign n2521 = n2516 | n2520 ;
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  assign n2522 = n2395 & ~n2499 ;
  assign n2523 = n918 | n2522 ;
  assign n2524 = ~n655 & n2222 ;
  buffer buf_n2525( .i (n2524), .o (n2525) );
  buffer buf_n2526( .i (n2525), .o (n2526) );
  assign n2527 = n214 & ~n2193 ;
  assign n2528 = n2526 | n2527 ;
  buffer buf_n2529( .i (n2528), .o (n2529) );
  assign n2530 = n2523 | n2529 ;
  assign n2531 = n2154 & ~n2530 ;
  assign n2532 = ~n2521 & n2531 ;
  buffer buf_n2533( .i (n2532), .o (n2533) );
  assign n2534 = n2513 | n2533 ;
  assign n2535 = ~n1469 & n2534 ;
  buffer buf_n2536( .i (n1438), .o (n2536) );
  buffer buf_n2537( .i (n2536), .o (n2537) );
  assign n2538 = ~n2535 & n2537 ;
  buffer buf_n2539( .i (n2538), .o (n2539) );
  buffer buf_n2540( .i (n2539), .o (n2540) );
  buffer buf_n2541( .i (n2540), .o (n2541) );
  assign n2542 = ~n2496 & n2541 ;
  buffer buf_n2543( .i (n2542), .o (n2543) );
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  buffer buf_n2551( .i (n2550), .o (n2551) );
  buffer buf_n2552( .i (n2551), .o (n2552) );
  buffer buf_n2553( .i (n2552), .o (n2553) );
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2555( .i (n2554), .o (n2555) );
  buffer buf_n2556( .i (n2555), .o (n2556) );
  assign n2557 = n1937 & ~n2296 ;
  assign n2558 = n2556 | n2557 ;
  buffer buf_n2559( .i (n2558), .o (n2559) );
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  assign n2562 = n2495 | n2561 ;
  buffer buf_n2563( .i (n2562), .o (n2563) );
  buffer buf_n2494( .i (n2493), .o (n2494) );
  assign n2564 = n2376 | n2494 ;
  buffer buf_n2565( .i (n2564), .o (n2565) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  assign n2566 = n1722 | n2563 ;
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  assign n2568 = n2110 | n2264 ;
  buffer buf_n2569( .i (n2568), .o (n2569) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  assign n2570 = n1595 & ~n2183 ;
  buffer buf_n2571( .i (n2570), .o (n2571) );
  buffer buf_n2572( .i (n2571), .o (n2572) );
  buffer buf_n2573( .i (n2572), .o (n2573) );
  buffer buf_n2574( .i (n2573), .o (n2574) );
  buffer buf_n2575( .i (n2574), .o (n2575) );
  buffer buf_n2576( .i (n2575), .o (n2576) );
  assign n2577 = ~n2569 & n2576 ;
  buffer buf_n2578( .i (n2577), .o (n2578) );
  buffer buf_n2579( .i (n2578), .o (n2579) );
  buffer buf_n2580( .i (n2579), .o (n2580) );
  assign n2581 = ~n2567 & n2580 ;
  assign n2582 = ~n2565 & n2581 ;
  buffer buf_n2583( .i (n2582), .o (n2583) );
  inverter inv_n2636( .i (n2583), .o (n2636) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  assign n2584 = n568 & ~n2565 ;
  buffer buf_n2585( .i (n2584), .o (n2585) );
  buffer buf_n2586( .i (n2585), .o (n2586) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  assign n2587 = n317 & ~n2583 ;
  assign n2588 = n2586 | ~n2587 ;
  assign n2589 = n1722 & n2563 ;
  buffer buf_n2590( .i (n2589), .o (n2590) );
  assign n2591 = n2567 & ~n2590 ;
  buffer buf_n2592( .i (n2591), .o (n2592) );
  assign n2593 = ~n1595 & n2183 ;
  buffer buf_n2594( .i (n2593), .o (n2594) );
  assign n2595 = n2571 | n2594 ;
  buffer buf_n2596( .i (n2595), .o (n2596) );
  buffer buf_n2597( .i (n2596), .o (n2597) );
  buffer buf_n2598( .i (n2597), .o (n2598) );
  buffer buf_n2599( .i (n2598), .o (n2599) );
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  assign n2602 = n2110 & n2264 ;
  buffer buf_n2603( .i (n2602), .o (n2603) );
  assign n2604 = n2569 & ~n2603 ;
  buffer buf_n2605( .i (n2604), .o (n2605) );
  assign n2606 = n2601 | n2605 ;
  assign n2607 = n2601 & n2605 ;
  assign n2608 = n2606 & ~n2607 ;
  buffer buf_n2609( .i (n2608), .o (n2609) );
  buffer buf_n2610( .i (n2609), .o (n2610) );
  assign n2611 = n2592 & n2610 ;
  assign n2612 = n2592 | n2610 ;
  assign n2613 = ~n2611 & n2612 ;
  buffer buf_n2614( .i (n2613), .o (n2614) );
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  buffer buf_n587( .i (G50), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  assign n2617 = n2376 & n2494 ;
  buffer buf_n2618( .i (n2617), .o (n2618) );
  assign n2619 = n2565 & ~n2618 ;
  buffer buf_n2620( .i (n2619), .o (n2620) );
  assign n2623 = n635 & n2620 ;
  buffer buf_n2624( .i (n2623), .o (n2624) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  assign n2625 = n635 | n2620 ;
  assign n2626 = ~n1317 & n2625 ;
  assign n2627 = ~n2624 & n2626 ;
  buffer buf_n2628( .i (n2627), .o (n2628) );
  assign n2629 = n2616 & n2628 ;
  assign n2630 = n2616 | n2628 ;
  assign n2631 = n2629 | ~n2630 ;
  buffer buf_n2621( .i (n2620), .o (n2621) );
  buffer buf_n2622( .i (n2621), .o (n2622) );
  assign n2632 = n2614 | n2622 ;
  assign n2633 = n2614 & n2622 ;
  assign n2634 = n2632 & ~n2633 ;
  assign G3519 = n692 ;
  assign G3520 = n695 ;
  assign G3521 = n742 ;
  assign G3522 = n769 ;
  assign G3523 = n794 ;
  assign G3524 = n1244 ;
  assign G3525 = n1275 ;
  assign G3526 = n1354 ;
  assign G3527 = n1415 ;
  assign G3528 = n2635 ;
  assign G3529 = n1715 ;
  assign G3530 = n1905 ;
  assign G3531 = n2110 ;
  assign G3532 = n2183 ;
  assign G3533 = n2262 ;
  assign G3534 = n2376 ;
  assign G3535 = n2493 ;
  assign G3536 = n2563 ;
  assign G3537 = n2636 ;
  assign G3538 = n2588 ;
  assign G3539 = n2631 ;
  assign G3540 = n2634 ;
endmodule
