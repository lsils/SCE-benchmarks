//207
module c7552(N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, N241_I, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342, N241_O);
  wire n_0000_;
  wire n_0001_;
  wire n_0002_;
  wire n_0003_;
  wire n_0004_;
  wire n_0005_;
  wire n_0006_;
  wire n_0007_;
  wire n_0008_;
  wire n_0009_;
  wire n_0010_;
  wire n_0011_;
  wire n_0012_;
  wire n_0013_;
  wire n_0014_;
  wire n_0015_;
  wire n_0016_;
  wire n_0017_;
  wire n_0018_;
  wire n_0019_;
  wire n_0020_;
  wire n_0021_;
  wire n_0022_;
  wire n_0023_;
  wire n_0024_;
  wire n_0025_;
  wire n_0026_;
  wire n_0027_;
  wire n_0028_;
  wire n_0029_;
  wire n_0030_;
  wire n_0031_;
  wire n_0032_;
  wire n_0033_;
  wire n_0034_;
  wire n_0035_;
  wire n_0036_;
  wire n_0037_;
  wire n_0038_;
  wire n_0039_;
  wire n_0040_;
  wire n_0041_;
  wire n_0042_;
  wire n_0043_;
  wire n_0044_;
  wire n_0045_;
  wire n_0046_;
  wire n_0047_;
  wire n_0048_;
  wire n_0049_;
  wire n_0050_;
  wire n_0051_;
  wire n_0052_;
  wire n_0053_;
  wire n_0054_;
  wire n_0055_;
  wire n_0056_;
  wire n_0057_;
  wire n_0058_;
  wire n_0059_;
  wire n_0060_;
  wire n_0061_;
  wire n_0062_;
  wire n_0063_;
  wire n_0064_;
  wire n_0065_;
  wire n_0066_;
  wire n_0067_;
  wire n_0068_;
  wire n_0069_;
  wire n_0070_;
  wire n_0071_;
  wire n_0072_;
  wire n_0073_;
  wire n_0074_;
  wire n_0075_;
  wire n_0076_;
  wire n_0077_;
  wire n_0078_;
  wire n_0079_;
  wire n_0080_;
  wire n_0081_;
  wire n_0082_;
  wire n_0083_;
  wire n_0084_;
  wire n_0085_;
  wire n_0086_;
  wire n_0087_;
  wire n_0088_;
  wire n_0089_;
  wire n_0090_;
  wire n_0091_;
  wire n_0092_;
  wire n_0093_;
  wire n_0094_;
  wire n_0095_;
  wire n_0096_;
  wire n_0097_;
  wire n_0098_;
  wire n_0099_;
  wire n_0100_;
  wire n_0101_;
  wire n_0102_;
  wire n_0103_;
  wire n_0104_;
  wire n_0105_;
  wire n_0106_;
  wire n_0107_;
  wire n_0108_;
  wire n_0109_;
  wire n_0110_;
  wire n_0111_;
  wire n_0112_;
  wire n_0113_;
  wire n_0114_;
  wire n_0115_;
  wire n_0116_;
  wire n_0117_;
  wire n_0118_;
  wire n_0119_;
  wire n_0120_;
  wire n_0121_;
  wire n_0122_;
  wire n_0123_;
  wire n_0124_;
  wire n_0125_;
  wire n_0126_;
  wire n_0127_;
  wire n_0128_;
  wire n_0129_;
  wire n_0130_;
  wire n_0131_;
  wire n_0132_;
  wire n_0133_;
  wire n_0134_;
  wire n_0135_;
  wire n_0136_;
  wire n_0137_;
  wire n_0138_;
  wire n_0139_;
  wire n_0140_;
  wire n_0141_;
  wire n_0142_;
  wire n_0143_;
  wire n_0144_;
  wire n_0145_;
  wire n_0146_;
  wire n_0147_;
  wire n_0148_;
  wire n_0149_;
  wire n_0150_;
  wire n_0151_;
  wire n_0152_;
  wire n_0153_;
  wire n_0154_;
  wire n_0155_;
  wire n_0156_;
  wire n_0157_;
  wire n_0158_;
  wire n_0159_;
  wire n_0160_;
  wire n_0161_;
  wire n_0162_;
  wire n_0163_;
  wire n_0164_;
  wire n_0165_;
  wire n_0166_;
  wire n_0167_;
  wire n_0168_;
  wire n_0169_;
  wire n_0170_;
  wire n_0171_;
  wire n_0172_;
  wire n_0173_;
  wire n_0174_;
  wire n_0175_;
  wire n_0176_;
  wire n_0177_;
  wire n_0178_;
  wire n_0179_;
  wire n_0180_;
  wire n_0181_;
  wire n_0182_;
  wire n_0183_;
  wire n_0184_;
  wire n_0185_;
  wire n_0186_;
  wire n_0187_;
  wire n_0188_;
  wire n_0189_;
  wire n_0190_;
  wire n_0191_;
  wire n_0192_;
  wire n_0193_;
  wire n_0194_;
  wire n_0195_;
  wire n_0196_;
  wire n_0197_;
  wire n_0198_;
  wire n_0199_;
  wire n_0200_;
  wire n_0201_;
  wire n_0202_;
  wire n_0203_;
  wire n_0204_;
  wire n_0205_;
  wire n_0206_;
  wire n_0207_;
  wire n_0208_;
  wire n_0209_;
  wire n_0210_;
  wire n_0211_;
  wire n_0212_;
  wire n_0213_;
  wire n_0214_;
  wire n_0215_;
  wire n_0216_;
  wire n_0217_;
  wire n_0218_;
  wire n_0219_;
  wire n_0220_;
  wire n_0221_;
  wire n_0222_;
  wire n_0223_;
  wire n_0224_;
  wire n_0225_;
  wire n_0226_;
  wire n_0227_;
  wire n_0228_;
  wire n_0229_;
  wire n_0230_;
  wire n_0231_;
  wire n_0232_;
  wire n_0233_;
  wire n_0234_;
  wire n_0235_;
  wire n_0236_;
  wire n_0237_;
  wire n_0238_;
  wire n_0239_;
  wire n_0240_;
  wire n_0241_;
  wire n_0242_;
  wire n_0243_;
  wire n_0244_;
  wire n_0245_;
  wire n_0246_;
  wire n_0247_;
  wire n_0248_;
  wire n_0249_;
  wire n_0250_;
  wire n_0251_;
  wire n_0252_;
  wire n_0253_;
  wire n_0254_;
  wire n_0255_;
  wire n_0256_;
  wire n_0257_;
  wire n_0258_;
  wire n_0259_;
  wire n_0260_;
  wire n_0261_;
  wire n_0262_;
  wire n_0263_;
  wire n_0264_;
  wire n_0265_;
  wire n_0266_;
  wire n_0267_;
  wire n_0268_;
  wire n_0269_;
  wire n_0270_;
  wire n_0271_;
  wire n_0272_;
  wire n_0273_;
  wire n_0274_;
  wire n_0275_;
  wire n_0276_;
  wire n_0277_;
  wire n_0278_;
  wire n_0279_;
  wire n_0280_;
  wire n_0281_;
  wire n_0282_;
  wire n_0283_;
  wire n_0284_;
  wire n_0285_;
  wire n_0286_;
  wire n_0287_;
  wire n_0288_;
  wire n_0289_;
  wire n_0290_;
  wire n_0291_;
  wire n_0292_;
  wire n_0293_;
  wire n_0294_;
  wire n_0295_;
  wire n_0296_;
  wire n_0297_;
  wire n_0298_;
  wire n_0299_;
  wire n_0300_;
  wire n_0301_;
  wire n_0302_;
  wire n_0303_;
  wire n_0304_;
  wire n_0305_;
  wire n_0306_;
  wire n_0307_;
  wire n_0308_;
  wire n_0309_;
  wire n_0310_;
  wire n_0311_;
  wire n_0312_;
  wire n_0313_;
  wire n_0314_;
  wire n_0315_;
  wire n_0316_;
  wire n_0317_;
  wire n_0318_;
  wire n_0319_;
  wire n_0320_;
  wire n_0321_;
  wire n_0322_;
  wire n_0323_;
  wire n_0324_;
  wire n_0325_;
  wire n_0326_;
  wire n_0327_;
  wire n_0328_;
  wire n_0329_;
  wire n_0330_;
  wire n_0331_;
  wire n_0332_;
  wire n_0333_;
  wire n_0334_;
  wire n_0335_;
  wire n_0336_;
  wire n_0337_;
  wire n_0338_;
  wire n_0339_;
  wire n_0340_;
  wire n_0341_;
  wire n_0342_;
  wire n_0343_;
  wire n_0344_;
  wire n_0345_;
  wire n_0346_;
  wire n_0347_;
  wire n_0348_;
  wire n_0349_;
  wire n_0350_;
  wire n_0351_;
  wire n_0352_;
  wire n_0353_;
  wire n_0354_;
  wire n_0355_;
  wire n_0356_;
  wire n_0357_;
  wire n_0358_;
  wire n_0359_;
  wire n_0360_;
  wire n_0361_;
  wire n_0362_;
  wire n_0363_;
  wire n_0364_;
  wire n_0365_;
  wire n_0366_;
  wire n_0367_;
  wire n_0368_;
  wire n_0369_;
  wire n_0370_;
  wire n_0371_;
  wire n_0372_;
  wire n_0373_;
  wire n_0374_;
  wire n_0375_;
  wire n_0376_;
  wire n_0377_;
  wire n_0378_;
  wire n_0379_;
  wire n_0380_;
  wire n_0381_;
  wire n_0382_;
  wire n_0383_;
  wire n_0384_;
  wire n_0385_;
  wire n_0386_;
  wire n_0387_;
  wire n_0388_;
  wire n_0389_;
  wire n_0390_;
  wire n_0391_;
  wire n_0392_;
  wire n_0393_;
  wire n_0394_;
  wire n_0395_;
  wire n_0396_;
  wire n_0397_;
  wire n_0398_;
  wire n_0399_;
  wire n_0400_;
  wire n_0401_;
  wire n_0402_;
  wire n_0403_;
  wire n_0404_;
  wire n_0405_;
  wire n_0406_;
  wire n_0407_;
  wire n_0408_;
  wire n_0409_;
  wire n_0410_;
  wire n_0411_;
  wire n_0412_;
  wire n_0413_;
  wire n_0414_;
  wire n_0415_;
  wire n_0416_;
  wire n_0417_;
  wire n_0418_;
  wire n_0419_;
  wire n_0420_;
  wire n_0421_;
  wire n_0422_;
  wire n_0423_;
  wire n_0424_;
  wire n_0425_;
  wire n_0426_;
  wire n_0427_;
  wire n_0428_;
  wire n_0429_;
  wire n_0430_;
  wire n_0431_;
  wire n_0432_;
  wire n_0433_;
  wire n_0434_;
  wire n_0435_;
  wire n_0436_;
  wire n_0437_;
  wire n_0438_;
  wire n_0439_;
  wire n_0440_;
  wire n_0441_;
  wire n_0442_;
  wire n_0443_;
  wire n_0444_;
  wire n_0445_;
  wire n_0446_;
  wire n_0447_;
  wire n_0448_;
  wire n_0449_;
  wire n_0450_;
  wire n_0451_;
  wire n_0452_;
  wire n_0453_;
  wire n_0454_;
  wire n_0455_;
  wire n_0456_;
  wire n_0457_;
  wire n_0458_;
  wire n_0459_;
  wire n_0460_;
  wire n_0461_;
  wire n_0462_;
  wire n_0463_;
  wire n_0464_;
  wire n_0465_;
  wire n_0466_;
  wire n_0467_;
  wire n_0468_;
  wire n_0469_;
  wire n_0470_;
  wire n_0471_;
  wire n_0472_;
  wire n_0473_;
  wire n_0474_;
  wire n_0475_;
  wire n_0476_;
  wire n_0477_;
  wire n_0478_;
  wire n_0479_;
  wire n_0480_;
  wire n_0481_;
  wire n_0482_;
  wire n_0483_;
  wire n_0484_;
  wire n_0485_;
  wire n_0486_;
  wire n_0487_;
  wire n_0488_;
  wire n_0489_;
  wire n_0490_;
  wire n_0491_;
  wire n_0492_;
  wire n_0493_;
  wire n_0494_;
  wire n_0495_;
  wire n_0496_;
  wire n_0497_;
  wire n_0498_;
  wire n_0499_;
  wire n_0500_;
  wire n_0501_;
  wire n_0502_;
  wire n_0503_;
  wire n_0504_;
  wire n_0505_;
  wire n_0506_;
  wire n_0507_;
  wire n_0508_;
  wire n_0509_;
  wire n_0510_;
  wire n_0511_;
  wire n_0512_;
  wire n_0513_;
  wire n_0514_;
  wire n_0515_;
  wire n_0516_;
  wire n_0517_;
  wire n_0518_;
  wire n_0519_;
  wire n_0520_;
  wire n_0521_;
  wire n_0522_;
  wire n_0523_;
  wire n_0524_;
  wire n_0525_;
  wire n_0526_;
  wire n_0527_;
  wire n_0528_;
  wire n_0529_;
  wire n_0530_;
  wire n_0531_;
  wire n_0532_;
  wire n_0533_;
  wire n_0534_;
  wire n_0535_;
  wire n_0536_;
  wire n_0537_;
  wire n_0538_;
  wire n_0539_;
  wire n_0540_;
  wire n_0541_;
  wire n_0542_;
  wire n_0543_;
  wire n_0544_;
  wire n_0545_;
  wire n_0546_;
  wire n_0547_;
  wire n_0548_;
  wire n_0549_;
  wire n_0550_;
  wire n_0551_;
  wire n_0552_;
  wire n_0553_;
  wire n_0554_;
  wire n_0555_;
  wire n_0556_;
  wire n_0557_;
  wire n_0558_;
  wire n_0559_;
  wire n_0560_;
  wire n_0561_;
  wire n_0562_;
  wire n_0563_;
  wire n_0564_;
  wire n_0565_;
  wire n_0566_;
  wire n_0567_;
  wire n_0568_;
  wire n_0569_;
  wire n_0570_;
  wire n_0571_;
  wire n_0572_;
  wire n_0573_;
  wire n_0574_;
  wire n_0575_;
  wire n_0576_;
  wire n_0577_;
  wire n_0578_;
  wire n_0579_;
  wire n_0580_;
  wire n_0581_;
  wire n_0582_;
  wire n_0583_;
  wire n_0584_;
  wire n_0585_;
  wire n_0586_;
  wire n_0587_;
  wire n_0588_;
  wire n_0589_;
  wire n_0590_;
  wire n_0591_;
  wire n_0592_;
  wire n_0593_;
  wire n_0594_;
  wire n_0595_;
  wire n_0596_;
  wire n_0597_;
  wire n_0598_;
  wire n_0599_;
  wire n_0600_;
  wire n_0601_;
  wire n_0602_;
  wire n_0603_;
  wire n_0604_;
  wire n_0605_;
  wire n_0606_;
  wire n_0607_;
  wire n_0608_;
  wire n_0609_;
  wire n_0610_;
  wire n_0611_;
  wire n_0612_;
  wire n_0613_;
  wire n_0614_;
  wire n_0615_;
  wire n_0616_;
  wire n_0617_;
  wire n_0618_;
  wire n_0619_;
  wire n_0620_;
  wire n_0621_;
  wire n_0622_;
  wire n_0623_;
  wire n_0624_;
  wire n_0625_;
  wire n_0626_;
  wire n_0627_;
  wire n_0628_;
  wire n_0629_;
  wire n_0630_;
  wire n_0631_;
  wire n_0632_;
  wire n_0633_;
  wire n_0634_;
  wire n_0635_;
  wire n_0636_;
  wire n_0637_;
  wire n_0638_;
  wire n_0639_;
  wire n_0640_;
  wire n_0641_;
  wire n_0642_;
  wire n_0643_;
  wire n_0644_;
  wire n_0645_;
  wire n_0646_;
  wire n_0647_;
  wire n_0648_;
  wire n_0649_;
  wire n_0650_;
  wire n_0651_;
  wire n_0652_;
  wire n_0653_;
  wire n_0654_;
  wire n_0655_;
  wire n_0656_;
  wire n_0657_;
  wire n_0658_;
  wire n_0659_;
  wire n_0660_;
  wire n_0661_;
  wire n_0662_;
  wire n_0663_;
  wire n_0664_;
  wire n_0665_;
  wire n_0666_;
  wire n_0667_;
  wire n_0668_;
  wire n_0669_;
  wire n_0670_;
  wire n_0671_;
  wire n_0672_;
  wire n_0673_;
  wire n_0674_;
  wire n_0675_;
  wire n_0676_;
  wire n_0677_;
  wire n_0678_;
  wire n_0679_;
  wire n_0680_;
  wire n_0681_;
  wire n_0682_;
  wire n_0683_;
  wire n_0684_;
  wire n_0685_;
  wire n_0686_;
  wire n_0687_;
  wire n_0688_;
  wire n_0689_;
  wire n_0690_;
  wire n_0691_;
  wire n_0692_;
  wire n_0693_;
  wire n_0694_;
  wire n_0695_;
  wire n_0696_;
  wire n_0697_;
  wire n_0698_;
  wire n_0699_;
  wire n_0700_;
  wire n_0701_;
  wire n_0702_;
  wire n_0703_;
  wire n_0704_;
  wire n_0705_;
  wire n_0706_;
  wire n_0707_;
  wire n_0708_;
  wire n_0709_;
  wire n_0710_;
  wire n_0711_;
  wire n_0712_;
  wire n_0713_;
  wire n_0714_;
  wire n_0715_;
  wire n_0716_;
  wire n_0717_;
  wire n_0718_;
  wire n_0719_;
  wire n_0720_;
  wire n_0721_;
  wire n_0722_;
  wire n_0723_;
  wire n_0724_;
  wire n_0725_;
  wire n_0726_;
  wire n_0727_;
  wire n_0728_;
  wire n_0729_;
  wire n_0730_;
  wire n_0731_;
  wire n_0732_;
  wire n_0733_;
  wire n_0734_;
  wire n_0735_;
  wire n_0736_;
  wire n_0737_;
  wire n_0738_;
  wire n_0739_;
  wire n_0740_;
  wire n_0741_;
  wire n_0742_;
  wire n_0743_;
  wire n_0744_;
  wire n_0745_;
  wire n_0746_;
  wire n_0747_;
  wire n_0748_;
  wire n_0749_;
  wire n_0750_;
  wire n_0751_;
  wire n_0752_;
  wire n_0753_;
  wire n_0754_;
  wire n_0755_;
  wire n_0756_;
  wire n_0757_;
  wire n_0758_;
  wire n_0759_;
  wire n_0760_;
  wire n_0761_;
  wire n_0762_;
  wire n_0763_;
  wire n_0764_;
  wire n_0765_;
  wire n_0766_;
  wire n_0767_;
  wire n_0768_;
  wire n_0769_;
  wire n_0770_;
  wire n_0771_;
  wire n_0772_;
  wire n_0773_;
  wire n_0774_;
  wire n_0775_;
  wire n_0776_;
  wire n_0777_;
  wire n_0778_;
  wire n_0779_;
  wire n_0780_;
  wire n_0781_;
  wire n_0782_;
  wire n_0783_;
  wire n_0784_;
  wire n_0785_;
  wire n_0786_;
  wire n_0787_;
  wire n_0788_;
  wire n_0789_;
  wire n_0790_;
  wire n_0791_;
  wire n_0792_;
  wire n_0793_;
  wire n_0794_;
  wire n_0795_;
  wire n_0796_;
  wire n_0797_;
  wire n_0798_;
  wire n_0799_;
  wire n_0800_;
  wire n_0801_;
  wire n_0802_;
  wire n_0803_;
  wire n_0804_;
  wire n_0805_;
  wire n_0806_;
  wire n_0807_;
  wire n_0808_;
  wire n_0809_;
  wire n_0810_;
  wire n_0811_;
  wire n_0812_;
  wire n_0813_;
  wire n_0814_;
  wire n_0815_;
  wire n_0816_;
  wire n_0817_;
  wire n_0818_;
  wire n_0819_;
  wire n_0820_;
  wire n_0821_;
  wire n_0822_;
  wire n_0823_;
  wire n_0824_;
  wire n_0825_;
  wire n_0826_;
  wire n_0827_;
  wire n_0828_;
  wire n_0829_;
  wire n_0830_;
  wire n_0831_;
  wire n_0832_;
  wire n_0833_;
  wire n_0834_;
  wire n_0835_;
  wire n_0836_;
  wire n_0837_;
  wire n_0838_;
  wire n_0839_;
  wire n_0840_;
  wire n_0841_;
  wire n_0842_;
  wire n_0843_;
  wire n_0844_;
  wire n_0845_;
  wire n_0846_;
  wire n_0847_;
  wire n_0848_;
  wire n_0849_;
  wire n_0850_;
  wire n_0851_;
  wire n_0852_;
  wire n_0853_;
  wire n_0854_;
  wire n_0855_;
  wire n_0856_;
  wire n_0857_;
  wire n_0858_;
  wire n_0859_;
  wire n_0860_;
  wire n_0861_;
  wire n_0862_;
  wire n_0863_;
  wire n_0864_;
  wire n_0865_;
  wire n_0866_;
  wire n_0867_;
  wire n_0868_;
  wire n_0869_;
  wire n_0870_;
  wire n_0871_;
  wire n_0872_;
  wire n_0873_;
  wire n_0874_;
  wire n_0875_;
  wire n_0876_;
  wire n_0877_;
  wire n_0878_;
  wire n_0879_;
  wire n_0880_;
  wire n_0881_;
  wire n_0882_;
  wire n_0883_;
  wire n_0884_;
  wire n_0885_;
  wire n_0886_;
  wire n_0887_;
  wire n_0888_;
  wire n_0889_;
  wire n_0890_;
  wire n_0891_;
  wire n_0892_;
  wire n_0893_;
  wire n_0894_;
  wire n_0895_;
  wire n_0896_;
  wire n_0897_;
  wire n_0898_;
  wire n_0899_;
  wire n_0900_;
  wire n_0901_;
  wire n_0902_;
  wire n_0903_;
  wire n_0904_;
  wire n_0905_;
  wire n_0906_;
  wire n_0907_;
  wire n_0908_;
  wire n_0909_;
  wire n_0910_;
  wire n_0911_;
  wire n_0912_;
  wire n_0913_;
  wire n_0914_;
  wire n_0915_;
  wire n_0916_;
  wire n_0917_;
  wire n_0918_;
  wire n_0919_;
  wire n_0920_;
  wire n_0921_;
  wire n_0922_;
  wire n_0923_;
  wire n_0924_;
  wire n_0925_;
  wire n_0926_;
  wire n_0927_;
  wire n_0928_;
  wire n_0929_;
  wire n_0930_;
  wire n_0931_;
  wire n_0932_;
  wire n_0933_;
  wire n_0934_;
  wire n_0935_;
  wire n_0936_;
  wire n_0937_;
  wire n_0938_;
  wire n_0939_;
  wire n_0940_;
  wire n_0941_;
  wire n_0942_;
  wire n_0943_;
  wire n_0944_;
  wire n_0945_;
  wire n_0946_;
  wire n_0947_;
  wire n_0948_;
  wire n_0949_;
  wire n_0950_;
  wire n_0951_;
  wire n_0952_;
  wire n_0953_;
  wire n_0954_;
  wire n_0955_;
  wire n_0956_;
  wire n_0957_;
  wire n_0958_;
  wire n_0959_;
  wire n_0960_;
  wire n_0961_;
  wire n_0962_;
  wire n_0963_;
  wire n_0964_;
  wire n_0965_;
  wire n_0966_;
  wire n_0967_;
  wire n_0968_;
  wire n_0969_;
  wire n_0970_;
  wire n_0971_;
  wire n_0972_;
  wire n_0973_;
  wire n_0974_;
  wire n_0975_;
  wire n_0976_;
  wire n_0977_;
  wire n_0978_;
  wire n_0979_;
  wire n_0980_;
  wire n_0981_;
  wire n_0982_;
  wire n_0983_;
  wire n_0984_;
  wire n_0985_;
  wire n_0986_;
  wire n_0987_;
  wire n_0988_;
  wire n_0989_;
  wire n_0990_;
  wire n_0991_;
  wire n_0992_;
  wire n_0993_;
  wire n_0994_;
  wire n_0995_;
  wire n_0996_;
  wire n_0997_;
  wire n_0998_;
  wire n_0999_;
  wire n_1000_;
  wire n_1001_;
  wire n_1002_;
  wire n_1003_;
  wire n_1004_;
  wire n_1005_;
  wire n_1006_;
  wire n_1007_;
  wire n_1008_;
  wire n_1009_;
  wire n_1010_;
  wire n_1011_;
  wire n_1012_;
  wire n_1013_;
  wire n_1014_;
  wire n_1015_;
  wire n_1016_;
  wire n_1017_;
  wire n_1018_;
  wire n_1019_;
  wire n_1020_;
  wire n_1021_;
  wire n_1022_;
  wire n_1023_;
  wire n_1024_;
  wire n_1025_;
  wire n_1026_;
  wire n_1027_;
  wire n_1028_;
  wire n_1029_;
  wire n_1030_;
  wire n_1031_;
  wire n_1032_;
  wire n_1033_;
  wire n_1034_;
  wire n_1035_;
  wire n_1036_;
  wire n_1037_;
  wire n_1038_;
  wire n_1039_;
  wire n_1040_;
  wire n_1041_;
  wire n_1042_;
  wire n_1043_;
  wire n_1044_;
  wire n_1045_;
  wire n_1046_;
  wire n_1047_;
  wire n_1048_;
  wire n_1049_;
  wire n_1050_;
  wire n_1051_;
  wire n_1052_;
  wire n_1053_;
  wire n_1054_;
  wire n_1055_;
  wire n_1056_;
  wire n_1057_;
  wire n_1058_;
  wire n_1059_;
  wire n_1060_;
  wire n_1061_;
  wire n_1062_;
  wire n_1063_;
  wire n_1064_;
  wire n_1065_;
  wire n_1066_;
  wire n_1067_;
  wire n_1068_;
  wire n_1069_;
  wire n_1070_;
  wire n_1071_;
  wire n_1072_;
  wire n_1073_;
  wire n_1074_;
  wire n_1075_;
  wire n_1076_;
  wire n_1077_;
  wire n_1078_;
  wire n_1079_;
  wire n_1080_;
  wire n_1081_;
  wire n_1082_;
  wire n_1083_;
  wire n_1084_;
  wire n_1085_;
  wire n_1086_;
  wire n_1087_;
  wire n_1088_;
  wire n_1089_;
  wire n_1090_;
  wire n_1091_;
  wire n_1092_;
  wire n_1093_;
  wire n_1094_;
  wire n_1095_;
  wire n_1096_;
  wire n_1097_;
  wire n_1098_;
  wire n_1099_;
  wire n_1100_;
  wire n_1101_;
  wire n_1102_;
  wire n_1103_;
  wire n_1104_;
  wire n_1105_;
  wire n_1106_;
  wire n_1107_;
  wire n_1108_;
  wire n_1109_;
  wire n_1110_;
  wire n_1111_;
  wire n_1112_;
  wire n_1113_;
  wire n_1114_;
  wire n_1115_;
  wire n_1116_;
  wire n_1117_;
  wire n_1118_;
  wire n_1119_;
  wire n_1120_;
  wire n_1121_;
  wire n_1122_;
  wire n_1123_;
  wire n_1124_;
  wire n_1125_;
  wire n_1126_;
  wire n_1127_;
  wire n_1128_;
  wire n_1129_;
  wire n_1130_;
  wire n_1131_;
  wire n_1132_;
  wire n_1133_;
  wire n_1134_;
  wire n_1135_;
  wire n_1136_;
  wire n_1137_;
  wire n_1138_;
  wire n_1139_;
  wire n_1140_;
  wire n_1141_;
  wire n_1142_;
  wire n_1143_;
  wire n_1144_;
  wire n_1145_;
  wire n_1146_;
  wire n_1147_;
  wire n_1148_;
  wire n_1149_;
  wire n_1150_;
  wire n_1151_;
  wire n_1152_;
  wire n_1153_;
  wire n_1154_;
  wire n_1155_;
  wire n_1156_;
  wire n_1157_;
  wire n_1158_;
  wire n_1159_;
  wire n_1160_;
  wire n_1161_;
  wire n_1162_;
  wire n_1163_;
  wire n_1164_;
  wire n_1165_;
  wire n_1166_;
  wire n_1167_;
  wire n_1168_;
  wire n_1169_;
  wire n_1170_;
  wire n_1171_;
  wire n_1172_;
  wire n_1173_;
  wire n_1174_;
  wire n_1175_;
  wire n_1176_;
  wire n_1177_;
  wire n_1178_;
  wire n_1179_;
  wire n_1180_;
  wire n_1181_;
  wire n_1182_;
  wire n_1183_;
  wire n_1184_;
  wire n_1185_;
  wire n_1186_;
  wire n_1187_;
  wire n_1188_;
  wire n_1189_;
  wire n_1190_;
  wire n_1191_;
  wire n_1192_;
  wire n_1193_;
  wire n_1194_;
  wire n_1195_;
  wire n_1196_;
  wire n_1197_;
  wire n_1198_;
  wire n_1199_;
  wire n_1200_;
  wire n_1201_;
  wire n_1202_;
  wire n_1203_;
  wire n_1204_;
  wire n_1205_;
  wire n_1206_;
  wire n_1207_;
  wire n_1208_;
  wire n_1209_;
  wire n_1210_;
  wire n_1211_;
  wire n_1212_;
  wire n_1213_;
  wire n_1214_;
  wire n_1215_;
  wire n_1216_;
  wire n_1217_;
  wire n_1218_;
  wire n_1219_;
  wire n_1220_;
  wire n_1221_;
  wire n_1222_;
  wire n_1223_;
  wire n_1224_;
  wire n_1225_;
  wire n_1226_;
  wire n_1227_;
  wire n_1228_;
  wire n_1229_;
  wire n_1230_;
  wire n_1231_;
  wire n_1232_;
  wire n_1233_;
  wire n_1234_;
  wire n_1235_;
  wire n_1236_;
  wire n_1237_;
  wire n_1238_;
  wire n_1239_;
  wire n_1240_;
  wire n_1241_;
  wire n_1242_;
  wire n_1243_;
  wire n_1244_;
  wire n_1245_;
  wire n_1246_;
  wire n_1247_;
  wire n_1248_;
  wire n_1249_;
  wire n_1250_;
  wire n_1251_;
  wire n_1252_;
  wire n_1253_;
  wire n_1254_;
  wire n_1255_;
  wire n_1256_;
  wire n_1257_;
  wire n_1258_;
  wire n_1259_;
  wire n_1260_;
  wire n_1261_;
  wire n_1262_;
  wire n_1263_;
  wire n_1264_;
  wire n_1265_;
  wire n_1266_;
  wire n_1267_;
  wire n_1268_;
  wire n_1269_;
  wire n_1270_;
  wire n_1271_;
  wire n_1272_;
  wire n_1273_;
  wire n_1274_;
  wire n_1275_;
  wire n_1276_;
  wire n_1277_;
  wire n_1278_;
  wire n_1279_;
  wire n_1280_;
  wire n_1281_;
  wire n_1282_;
  wire n_1283_;
  wire n_1284_;
  wire n_1285_;
  wire n_1286_;
  wire n_1287_;
  wire n_1288_;
  wire n_1289_;
  wire n_1290_;
  wire n_1291_;
  wire n_1292_;
  wire n_1293_;
  wire n_1294_;
  wire n_1295_;
  wire n_1296_;
  wire n_1297_;
  wire n_1298_;
  wire n_1299_;
  wire n_1300_;
  wire n_1301_;
  wire n_1302_;
  wire n_1303_;
  wire n_1304_;
  wire n_1305_;
  wire n_1306_;
  wire n_1307_;
  wire n_1308_;
  wire n_1309_;
  wire n_1310_;
  wire n_1311_;
  wire n_1312_;
  wire n_1313_;
  wire n_1314_;
  wire n_1315_;
  wire n_1316_;
  wire n_1317_;
  wire n_1318_;
  wire n_1319_;
  wire n_1320_;
  wire n_1321_;
  wire n_1322_;
  wire n_1323_;
  wire n_1324_;
  wire n_1325_;
  wire n_1326_;
  wire n_1327_;
  wire n_1328_;
  wire n_1329_;
  wire n_1330_;
  wire n_1331_;
  wire n_1332_;
  wire n_1333_;
  wire n_1334_;
  wire n_1335_;
  wire n_1336_;
  wire n_1337_;
  wire n_1338_;
  wire n_1339_;
  wire n_1340_;
  wire n_1341_;
  wire n_1342_;
  wire n_1343_;
  wire n_1344_;
  wire n_1345_;
  wire n_1346_;
  wire n_1347_;
  wire n_1348_;
  wire n_1349_;
  wire n_1350_;
  wire n_1351_;
  wire n_1352_;
  wire n_1353_;
  wire n_1354_;
  wire n_1355_;
  wire n_1356_;
  wire n_1357_;
  wire n_1358_;
  wire n_1359_;
  wire n_1360_;
  wire n_1361_;
  wire n_1362_;
  wire n_1363_;
  wire n_1364_;
  wire n_1365_;
  wire n_1366_;
  wire n_1367_;
  wire n_1368_;
  wire n_1369_;
  wire n_1370_;
  wire n_1371_;
  input N1;
  input N100;
  output N10025;
  output N10101;
  output N10102;
  output N10103;
  output N10104;
  output N10109;
  output N10110;
  output N10111;
  output N10112;
  input N103;
  output N10350;
  output N10351;
  output N10352;
  output N10353;
  output N10574;
  output N10575;
  output N10576;
  input N106;
  output N10628;
  output N10632;
  output N10641;
  output N10704;
  output N10706;
  output N10711;
  output N10712;
  output N10713;
  output N10714;
  output N10715;
  output N10716;
  output N10717;
  output N10718;
  output N10729;
  output N10759;
  output N10760;
  output N10761;
  output N10762;
  output N10763;
  output N10827;
  output N10837;
  output N10838;
  output N10839;
  output N10840;
  output N10868;
  output N10869;
  output N10870;
  output N10871;
  input N109;
  output N10905;
  output N10906;
  output N10907;
  output N10908;
  input N110;
  input N111;
  output N1110;
  output N1111;
  output N1112;
  output N1113;
  output N1114;
  input N112;
  input N113;
  output N11333;
  output N11334;
  output N11340;
  output N11342;
  input N114;
  input N115;
  input N118;
  input N12;
  input N121;
  input N124;
  input N127;
  input N130;
  input N133;
  input N134;
  input N135;
  input N138;
  input N141;
  input N144;
  input N147;
  output N1489;
  output N1490;
  input N15;
  input N150;
  input N151;
  input N152;
  input N153;
  input N154;
  input N155;
  input N156;
  input N157;
  input N158;
  input N159;
  input N160;
  input N161;
  input N162;
  input N163;
  input N164;
  input N165;
  input N166;
  input N167;
  input N168;
  input N169;
  input N170;
  input N171;
  input N172;
  input N173;
  input N174;
  input N175;
  input N176;
  input N177;
  input N178;
  output N1781;
  input N179;
  input N18;
  input N180;
  input N181;
  input N182;
  input N183;
  input N184;
  input N185;
  input N186;
  input N187;
  input N188;
  input N189;
  input N190;
  input N191;
  input N192;
  input N193;
  input N194;
  input N195;
  input N196;
  input N197;
  input N198;
  input N199;
  input N200;
  input N201;
  input N202;
  input N203;
  input N204;
  input N205;
  input N206;
  input N207;
  input N208;
  input N209;
  input N210;
  input N211;
  input N212;
  input N213;
  input N214;
  input N215;
  input N216;
  input N217;
  input N218;
  input N219;
  input N220;
  input N221;
  input N222;
  input N223;
  input N224;
  input N225;
  input N226;
  input N227;
  input N228;
  input N229;
  input N23;
  input N230;
  input N231;
  input N232;
  input N233;
  input N234;
  input N235;
  input N236;
  input N237;
  input N238;
  input N239;
  input N240;
  input N241_I;
  output N241_O;
  input N242;
  input N245;
  input N248;
  input N251;
  input N254;
  input N257;
  input N26;
  input N260;
  input N263;
  input N267;
  input N271;
  input N274;
  input N277;
  input N280;
  input N283;
  input N286;
  input N289;
  input N29;
  input N293;
  input N296;
  input N299;
  input N303;
  input N307;
  input N310;
  input N313;
  input N316;
  input N319;
  input N32;
  input N322;
  input N325;
  input N328;
  input N331;
  input N334;
  input N337;
  input N340;
  input N343;
  input N346;
  input N349;
  input N35;
  input N352;
  input N355;
  input N358;
  input N361;
  input N364;
  input N367;
  input N38;
  input N382;
  output N387;
  output N388;
  input N41;
  input N44;
  input N47;
  output N478;
  output N482;
  output N484;
  output N486;
  output N489;
  output N492;
  input N5;
  input N50;
  output N501;
  output N505;
  output N507;
  output N509;
  output N511;
  output N513;
  output N515;
  output N517;
  output N519;
  input N53;
  output N535;
  output N537;
  output N539;
  input N54;
  output N541;
  output N543;
  output N545;
  output N547;
  output N549;
  input N55;
  output N551;
  output N553;
  output N556;
  output N559;
  input N56;
  output N561;
  output N563;
  output N565;
  output N567;
  output N569;
  input N57;
  output N571;
  output N573;
  input N58;
  output N582;
  input N59;
  input N60;
  input N61;
  input N62;
  input N63;
  input N64;
  output N643;
  input N65;
  input N66;
  input N69;
  input N70;
  output N707;
  input N73;
  input N74;
  input N75;
  input N76;
  input N77;
  input N78;
  input N79;
  input N80;
  input N81;
  output N813;
  input N82;
  input N83;
  input N84;
  input N85;
  input N86;
  input N87;
  input N88;
  output N881;
  output N882;
  output N883;
  output N884;
  output N885;
  output N889;
  input N89;
  input N9;
  input N94;
  output N945;
  input N97;
  or_bb n_1372_ (
    .a(N5),
    .b(N57),
    .c(N881)
  );
  or_ii n_1373_ (
    .a(N184),
    .b(N150),
    .c(n_0653_)
  );
  or_ii n_1374_ (
    .a(N240),
    .b(N228),
    .c(n_0654_)
  );
  or_bb n_1375_ (
    .a(n_0654_),
    .b(n_0653_),
    .c(N882)
  );
  or_ii n_1376_ (
    .a(N152),
    .b(N210),
    .c(n_0655_)
  );
  or_ii n_1377_ (
    .a(N230),
    .b(N218),
    .c(n_0656_)
  );
  or_bb n_1378_ (
    .a(n_0656_),
    .b(n_0655_),
    .c(N883)
  );
  or_ii n_1379_ (
    .a(N182),
    .b(N183),
    .c(n_0657_)
  );
  or_ii n_1380_ (
    .a(N186),
    .b(N185),
    .c(n_0658_)
  );
  or_bb n_1381_ (
    .a(n_0658_),
    .b(n_0657_),
    .c(N884)
  );
  or_ii n_1382_ (
    .a(N172),
    .b(N162),
    .c(n_0659_)
  );
  or_ii n_1383_ (
    .a(N199),
    .b(N188),
    .c(n_0660_)
  );
  or_bb n_1384_ (
    .a(n_0660_),
    .b(n_0659_),
    .c(N885)
  );
  or_bi n_1385_ (
    .a(N5),
    .b(N242),
    .c(N1110)
  );
  inv n_1386_ (
    .din(N15),
    .dout(N1111)
  );
  and_bi n_1387_ (
    .a(N134),
    .b(N5),
    .c(n_0661_)
  );
  or_ii n_1388_ (
    .a(n_0661_),
    .b(N133),
    .c(N1113)
  );
  or_bi n_1389_ (
    .a(N18),
    .b(N41),
    .c(n_0662_)
  );
  or_bb n_1390_ (
    .a(n_0662_),
    .b(N310),
    .c(n_0663_)
  );
  or_bb n_1391_ (
    .a(N41),
    .b(N18),
    .c(n_0664_)
  );
  and_bi n_1392_ (
    .a(N310),
    .b(n_0664_),
    .c(n_0665_)
  );
  or_bi n_1393_ (
    .a(n_0665_),
    .b(n_0663_),
    .c(n_0666_)
  );
  and_bi n_1394_ (
    .a(N367),
    .b(n_0666_),
    .c(n_0667_)
  );
  inv n_1395_ (
    .din(N367),
    .dout(n_0668_)
  );
  or_ii n_1396_ (
    .a(n_0666_),
    .b(n_0668_),
    .c(n_0669_)
  );
  and_bi n_1397_ (
    .a(n_0669_),
    .b(n_0667_),
    .c(N10025)
  );
  inv n_1398_ (
    .din(N322),
    .dout(n_0670_)
  );
  and_bb n_1399_ (
    .a(N235),
    .b(N18),
    .c(n_0671_)
  );
  and_bi n_1400_ (
    .a(N103),
    .b(N18),
    .c(n_0672_)
  );
  and_ii n_1401_ (
    .a(n_0672_),
    .b(n_0671_),
    .c(n_0673_)
  );
  and_bi n_1402_ (
    .a(n_0670_),
    .b(n_0673_),
    .c(n_0674_)
  );
  and_bi n_1403_ (
    .a(n_0673_),
    .b(n_0670_),
    .c(n_0675_)
  );
  and_ii n_1404_ (
    .a(n_0675_),
    .b(n_0674_),
    .c(n_0676_)
  );
  or_ii n_1405_ (
    .a(N236),
    .b(N18),
    .c(n_0677_)
  );
  and_bi n_1406_ (
    .a(N23),
    .b(N18),
    .c(n_0678_)
  );
  and_bi n_1407_ (
    .a(n_0677_),
    .b(n_0678_),
    .c(n_0679_)
  );
  or_ii n_1408_ (
    .a(n_0679_),
    .b(N319),
    .c(n_0680_)
  );
  or_ii n_1409_ (
    .a(N237),
    .b(N18),
    .c(n_0681_)
  );
  and_bi n_1410_ (
    .a(N26),
    .b(N18),
    .c(n_0682_)
  );
  and_bi n_1411_ (
    .a(n_0681_),
    .b(n_0682_),
    .c(n_0683_)
  );
  or_ii n_1412_ (
    .a(n_0683_),
    .b(N316),
    .c(n_0684_)
  );
  and_ii n_1413_ (
    .a(n_0683_),
    .b(N316),
    .c(n_0685_)
  );
  and_bi n_1414_ (
    .a(n_0684_),
    .b(n_0685_),
    .c(n_0686_)
  );
  or_ii n_1415_ (
    .a(N238),
    .b(N18),
    .c(n_0687_)
  );
  and_bi n_1416_ (
    .a(N29),
    .b(N18),
    .c(n_0688_)
  );
  or_bi n_1417_ (
    .a(n_0688_),
    .b(n_0687_),
    .c(n_0689_)
  );
  and_bi n_1418_ (
    .a(N313),
    .b(n_0689_),
    .c(n_0690_)
  );
  and_bi n_1419_ (
    .a(n_0689_),
    .b(N313),
    .c(n_0691_)
  );
  or_bb n_1420_ (
    .a(n_0691_),
    .b(n_0690_),
    .c(n_0692_)
  );
  or_bb n_1421_ (
    .a(n_0692_),
    .b(n_0666_),
    .c(n_0693_)
  );
  and_bi n_1422_ (
    .a(n_0686_),
    .b(n_0693_),
    .c(n_0694_)
  );
  or_ii n_1423_ (
    .a(n_0694_),
    .b(N367),
    .c(n_0695_)
  );
  and_ii n_1424_ (
    .a(n_0679_),
    .b(N319),
    .c(n_0696_)
  );
  or_bb n_1425_ (
    .a(n_0690_),
    .b(n_0663_),
    .c(n_0697_)
  );
  or_bb n_1426_ (
    .a(n_0691_),
    .b(n_0685_),
    .c(n_0698_)
  );
  and_bi n_1427_ (
    .a(n_0697_),
    .b(n_0698_),
    .c(n_0699_)
  );
  and_bi n_1428_ (
    .a(n_0684_),
    .b(n_0699_),
    .c(n_0700_)
  );
  and_ii n_1429_ (
    .a(n_0700_),
    .b(n_0696_),
    .c(n_0701_)
  );
  and_bb n_1430_ (
    .a(n_0701_),
    .b(n_0695_),
    .c(n_0702_)
  );
  and_bi n_1431_ (
    .a(n_0680_),
    .b(n_0702_),
    .c(n_0703_)
  );
  or_ii n_1432_ (
    .a(n_0703_),
    .b(n_0676_),
    .c(n_0704_)
  );
  and_ii n_1433_ (
    .a(n_0703_),
    .b(n_0676_),
    .c(n_0705_)
  );
  and_bi n_1434_ (
    .a(n_0704_),
    .b(n_0705_),
    .c(N10109)
  );
  or_bi n_1435_ (
    .a(n_0700_),
    .b(n_0695_),
    .c(n_0706_)
  );
  or_bi n_1436_ (
    .a(n_0696_),
    .b(n_0680_),
    .c(n_0707_)
  );
  or_ii n_1437_ (
    .a(n_0707_),
    .b(n_0706_),
    .c(n_0708_)
  );
  or_bb n_1438_ (
    .a(n_0707_),
    .b(n_0706_),
    .c(n_0709_)
  );
  or_ii n_1439_ (
    .a(n_0709_),
    .b(n_0708_),
    .c(N10110)
  );
  and_bi n_1440_ (
    .a(n_0663_),
    .b(n_0691_),
    .c(n_0710_)
  );
  and_bi n_1441_ (
    .a(n_0710_),
    .b(n_0667_),
    .c(n_0711_)
  );
  and_ii n_1442_ (
    .a(n_0711_),
    .b(n_0690_),
    .c(n_0712_)
  );
  and_bi n_1443_ (
    .a(n_0712_),
    .b(n_0686_),
    .c(n_0713_)
  );
  and_bi n_1444_ (
    .a(n_0686_),
    .b(n_0712_),
    .c(n_0714_)
  );
  or_bb n_1445_ (
    .a(n_0714_),
    .b(n_0713_),
    .c(N10111)
  );
  and_bi n_1446_ (
    .a(n_0663_),
    .b(n_0667_),
    .c(n_0715_)
  );
  and_bi n_1447_ (
    .a(n_0715_),
    .b(n_0692_),
    .c(n_0716_)
  );
  and_bi n_1448_ (
    .a(n_0692_),
    .b(n_0715_),
    .c(n_0717_)
  );
  or_bb n_1449_ (
    .a(n_0717_),
    .b(n_0716_),
    .c(N10112)
  );
  and_bb n_1450_ (
    .a(N9),
    .b(N12),
    .c(n_0718_)
  );
  and_bi n_1451_ (
    .a(N18),
    .b(N154),
    .c(n_0719_)
  );
  and_ii n_1452_ (
    .a(n_0719_),
    .b(n_0718_),
    .c(n_0720_)
  );
  and_bi n_1453_ (
    .a(N18),
    .b(N153),
    .c(n_0721_)
  );
  or_ii n_1454_ (
    .a(n_0721_),
    .b(n_0720_),
    .c(n_0722_)
  );
  and_ii n_1455_ (
    .a(n_0721_),
    .b(n_0718_),
    .c(n_0723_)
  );
  and_bb n_1456_ (
    .a(n_0723_),
    .b(n_0719_),
    .c(n_0724_)
  );
  and_bi n_1457_ (
    .a(n_0722_),
    .b(n_0724_),
    .c(n_0725_)
  );
  and_bi n_1458_ (
    .a(N18),
    .b(N156),
    .c(n_0726_)
  );
  and_ii n_1459_ (
    .a(n_0726_),
    .b(n_0718_),
    .c(n_0727_)
  );
  and_bi n_1460_ (
    .a(N18),
    .b(N155),
    .c(n_0728_)
  );
  and_bb n_1461_ (
    .a(n_0728_),
    .b(n_0727_),
    .c(n_0729_)
  );
  and_ii n_1462_ (
    .a(n_0728_),
    .b(n_0718_),
    .c(n_0730_)
  );
  and_bb n_1463_ (
    .a(n_0730_),
    .b(n_0726_),
    .c(n_0731_)
  );
  or_bb n_1464_ (
    .a(n_0731_),
    .b(n_0729_),
    .c(n_0732_)
  );
  and_bi n_1465_ (
    .a(N141),
    .b(N18),
    .c(n_0733_)
  );
  and_bb n_1466_ (
    .a(N161),
    .b(N18),
    .c(n_0734_)
  );
  and_ii n_1467_ (
    .a(n_0734_),
    .b(n_0733_),
    .c(n_0735_)
  );
  and_bi n_1468_ (
    .a(N147),
    .b(N18),
    .c(n_0736_)
  );
  and_bb n_1469_ (
    .a(N151),
    .b(N18),
    .c(n_0737_)
  );
  and_ii n_1470_ (
    .a(n_0737_),
    .b(n_0736_),
    .c(n_0738_)
  );
  and_bb n_1471_ (
    .a(n_0738_),
    .b(n_0735_),
    .c(n_0739_)
  );
  and_ii n_1472_ (
    .a(n_0738_),
    .b(n_0735_),
    .c(n_0740_)
  );
  and_ii n_1473_ (
    .a(n_0740_),
    .b(n_0739_),
    .c(n_0741_)
  );
  or_bb n_1474_ (
    .a(n_0741_),
    .b(n_0732_),
    .c(n_0742_)
  );
  and_bb n_1475_ (
    .a(n_0741_),
    .b(n_0732_),
    .c(n_0743_)
  );
  and_bi n_1476_ (
    .a(n_0742_),
    .b(n_0743_),
    .c(n_0744_)
  );
  and_ii n_1477_ (
    .a(n_0744_),
    .b(n_0725_),
    .c(n_0745_)
  );
  and_bb n_1478_ (
    .a(n_0744_),
    .b(n_0725_),
    .c(n_0746_)
  );
  and_ii n_1479_ (
    .a(n_0746_),
    .b(n_0745_),
    .c(n_0747_)
  );
  and_bi n_1480_ (
    .a(N135),
    .b(N18),
    .c(n_0748_)
  );
  and_bb n_1481_ (
    .a(N158),
    .b(N18),
    .c(n_0749_)
  );
  or_bb n_1482_ (
    .a(n_0749_),
    .b(n_0748_),
    .c(n_0750_)
  );
  and_bi n_1483_ (
    .a(N18),
    .b(N157),
    .c(n_0751_)
  );
  and_ii n_1484_ (
    .a(n_0751_),
    .b(n_0718_),
    .c(n_0752_)
  );
  or_bb n_1485_ (
    .a(n_0752_),
    .b(n_0750_),
    .c(n_0753_)
  );
  and_bb n_1486_ (
    .a(n_0752_),
    .b(n_0750_),
    .c(n_0754_)
  );
  and_bi n_1487_ (
    .a(n_0753_),
    .b(n_0754_),
    .c(n_0755_)
  );
  and_bi n_1488_ (
    .a(N138),
    .b(N18),
    .c(n_0756_)
  );
  and_bb n_1489_ (
    .a(N160),
    .b(N18),
    .c(n_0757_)
  );
  and_ii n_1490_ (
    .a(n_0757_),
    .b(n_0756_),
    .c(n_0758_)
  );
  and_bi n_1491_ (
    .a(N144),
    .b(N18),
    .c(n_0759_)
  );
  and_bb n_1492_ (
    .a(N159),
    .b(N18),
    .c(n_0760_)
  );
  and_ii n_1493_ (
    .a(n_0760_),
    .b(n_0759_),
    .c(n_0761_)
  );
  and_ii n_1494_ (
    .a(n_0761_),
    .b(n_0758_),
    .c(n_0762_)
  );
  and_bb n_1495_ (
    .a(n_0761_),
    .b(n_0758_),
    .c(n_0763_)
  );
  or_bb n_1496_ (
    .a(n_0763_),
    .b(n_0762_),
    .c(n_0764_)
  );
  and_ii n_1497_ (
    .a(n_0764_),
    .b(n_0755_),
    .c(n_0765_)
  );
  and_bb n_1498_ (
    .a(n_0764_),
    .b(n_0755_),
    .c(n_0766_)
  );
  and_ii n_1499_ (
    .a(n_0766_),
    .b(n_0765_),
    .c(n_0767_)
  );
  and_bb n_1500_ (
    .a(n_0767_),
    .b(n_0747_),
    .c(n_0768_)
  );
  and_bi n_1501_ (
    .a(N18),
    .b(N209),
    .c(n_0769_)
  );
  and_bi n_1502_ (
    .a(n_0769_),
    .b(n_0718_),
    .c(n_0770_)
  );
  and_bi n_1503_ (
    .a(N18),
    .b(N214),
    .c(n_0771_)
  );
  and_ii n_1504_ (
    .a(n_0771_),
    .b(n_0718_),
    .c(n_0772_)
  );
  and_bi n_1505_ (
    .a(N18),
    .b(N213),
    .c(n_0773_)
  );
  and_bb n_1506_ (
    .a(n_0773_),
    .b(n_0772_),
    .c(n_0774_)
  );
  and_ii n_1507_ (
    .a(n_0773_),
    .b(n_0718_),
    .c(n_0775_)
  );
  and_bb n_1508_ (
    .a(n_0775_),
    .b(n_0771_),
    .c(n_0776_)
  );
  and_ii n_1509_ (
    .a(n_0776_),
    .b(n_0774_),
    .c(n_0777_)
  );
  or_bi n_1510_ (
    .a(n_0770_),
    .b(n_0777_),
    .c(n_0778_)
  );
  and_bi n_1511_ (
    .a(n_0770_),
    .b(n_0777_),
    .c(n_0779_)
  );
  and_bi n_1512_ (
    .a(n_0778_),
    .b(n_0779_),
    .c(n_0780_)
  );
  and_bi n_1513_ (
    .a(N18),
    .b(N216),
    .c(n_0781_)
  );
  and_ii n_1514_ (
    .a(n_0781_),
    .b(n_0718_),
    .c(n_0782_)
  );
  and_bi n_1515_ (
    .a(N18),
    .b(N215),
    .c(n_0783_)
  );
  and_bb n_1516_ (
    .a(n_0783_),
    .b(n_0782_),
    .c(n_0784_)
  );
  and_ii n_1517_ (
    .a(n_0783_),
    .b(n_0718_),
    .c(n_0785_)
  );
  and_bb n_1518_ (
    .a(n_0785_),
    .b(n_0781_),
    .c(n_0786_)
  );
  and_ii n_1519_ (
    .a(n_0786_),
    .b(n_0784_),
    .c(n_0787_)
  );
  or_bi n_1520_ (
    .a(n_0718_),
    .b(N18),
    .c(n_0788_)
  );
  and_ii n_1521_ (
    .a(N211),
    .b(N212),
    .c(n_0789_)
  );
  and_bb n_1522_ (
    .a(N211),
    .b(N212),
    .c(n_0790_)
  );
  or_bb n_1523_ (
    .a(n_0790_),
    .b(n_0789_),
    .c(n_0791_)
  );
  and_ii n_1524_ (
    .a(n_0791_),
    .b(n_0788_),
    .c(n_0792_)
  );
  and_bb n_1525_ (
    .a(n_0792_),
    .b(n_0787_),
    .c(n_0793_)
  );
  and_ii n_1526_ (
    .a(n_0792_),
    .b(n_0787_),
    .c(n_0794_)
  );
  and_ii n_1527_ (
    .a(n_0794_),
    .b(n_0793_),
    .c(n_0795_)
  );
  or_bi n_1528_ (
    .a(n_0780_),
    .b(n_0795_),
    .c(n_0796_)
  );
  and_bi n_1529_ (
    .a(n_0780_),
    .b(n_0795_),
    .c(n_0797_)
  );
  and_bi n_1530_ (
    .a(n_0796_),
    .b(n_0797_),
    .c(n_0798_)
  );
  and_ii n_1531_ (
    .a(n_0767_),
    .b(n_0747_),
    .c(n_0799_)
  );
  or_bb n_1532_ (
    .a(n_0799_),
    .b(n_0798_),
    .c(n_0800_)
  );
  or_bb n_1533_ (
    .a(n_0800_),
    .b(n_0768_),
    .c(n_0801_)
  );
  and_bb n_1534_ (
    .a(N232),
    .b(N18),
    .c(n_0802_)
  );
  and_bi n_1535_ (
    .a(N124),
    .b(N18),
    .c(n_0803_)
  );
  and_ii n_1536_ (
    .a(n_0803_),
    .b(n_0802_),
    .c(n_0804_)
  );
  and_bb n_1537_ (
    .a(N229),
    .b(N18),
    .c(n_0805_)
  );
  and_bi n_1538_ (
    .a(n_0662_),
    .b(n_0805_),
    .c(n_0806_)
  );
  and_bi n_1539_ (
    .a(n_0804_),
    .b(n_0806_),
    .c(n_0807_)
  );
  and_bi n_1540_ (
    .a(n_0806_),
    .b(n_0804_),
    .c(n_0808_)
  );
  and_ii n_1541_ (
    .a(n_0808_),
    .b(n_0807_),
    .c(n_0809_)
  );
  and_bb n_1542_ (
    .a(N231),
    .b(N18),
    .c(n_0810_)
  );
  and_bi n_1543_ (
    .a(N100),
    .b(N18),
    .c(n_0811_)
  );
  and_ii n_1544_ (
    .a(n_0811_),
    .b(n_0810_),
    .c(n_0812_)
  );
  and_bi n_1545_ (
    .a(n_0679_),
    .b(n_0812_),
    .c(n_0813_)
  );
  and_bi n_1546_ (
    .a(n_0812_),
    .b(n_0679_),
    .c(n_0814_)
  );
  and_ii n_1547_ (
    .a(n_0814_),
    .b(n_0813_),
    .c(n_0815_)
  );
  and_bi n_1548_ (
    .a(n_0809_),
    .b(n_0815_),
    .c(n_0816_)
  );
  and_bi n_1549_ (
    .a(n_0815_),
    .b(n_0809_),
    .c(n_0817_)
  );
  or_bb n_1550_ (
    .a(n_0817_),
    .b(n_0816_),
    .c(n_0818_)
  );
  and_bi n_1551_ (
    .a(n_0673_),
    .b(n_0683_),
    .c(n_0819_)
  );
  and_bi n_1552_ (
    .a(n_0683_),
    .b(n_0673_),
    .c(n_0820_)
  );
  or_bb n_1553_ (
    .a(n_0820_),
    .b(n_0819_),
    .c(n_0821_)
  );
  or_ii n_1554_ (
    .a(N234),
    .b(N18),
    .c(n_0822_)
  );
  and_bi n_1555_ (
    .a(N130),
    .b(N18),
    .c(n_0823_)
  );
  and_bi n_1556_ (
    .a(n_0822_),
    .b(n_0823_),
    .c(n_0824_)
  );
  or_ii n_1557_ (
    .a(N233),
    .b(N18),
    .c(n_0825_)
  );
  and_bi n_1558_ (
    .a(N127),
    .b(N18),
    .c(n_0826_)
  );
  and_bi n_1559_ (
    .a(n_0825_),
    .b(n_0826_),
    .c(n_0827_)
  );
  and_bi n_1560_ (
    .a(n_0824_),
    .b(n_0827_),
    .c(n_0828_)
  );
  and_bi n_1561_ (
    .a(n_0827_),
    .b(n_0824_),
    .c(n_0829_)
  );
  and_ii n_1562_ (
    .a(n_0829_),
    .b(n_0828_),
    .c(n_0830_)
  );
  and_bb n_1563_ (
    .a(N239),
    .b(N18),
    .c(n_0831_)
  );
  and_bi n_1564_ (
    .a(N44),
    .b(N18),
    .c(n_0832_)
  );
  and_ii n_1565_ (
    .a(n_0832_),
    .b(n_0831_),
    .c(n_0833_)
  );
  and_bi n_1566_ (
    .a(n_0833_),
    .b(n_0689_),
    .c(n_0834_)
  );
  and_bi n_1567_ (
    .a(n_0689_),
    .b(n_0833_),
    .c(n_0835_)
  );
  and_ii n_1568_ (
    .a(n_0835_),
    .b(n_0834_),
    .c(n_0836_)
  );
  and_ii n_1569_ (
    .a(n_0836_),
    .b(n_0830_),
    .c(n_0837_)
  );
  and_bb n_1570_ (
    .a(n_0836_),
    .b(n_0830_),
    .c(n_0838_)
  );
  or_bb n_1571_ (
    .a(n_0838_),
    .b(n_0837_),
    .c(n_0839_)
  );
  and_ii n_1572_ (
    .a(n_0839_),
    .b(n_0821_),
    .c(n_0840_)
  );
  and_bb n_1573_ (
    .a(n_0839_),
    .b(n_0821_),
    .c(n_0841_)
  );
  and_ii n_1574_ (
    .a(n_0841_),
    .b(n_0840_),
    .c(n_0842_)
  );
  or_bi n_1575_ (
    .a(n_0818_),
    .b(n_0842_),
    .c(n_0843_)
  );
  and_bi n_1576_ (
    .a(n_0818_),
    .b(n_0842_),
    .c(n_0844_)
  );
  and_bi n_1577_ (
    .a(n_0843_),
    .b(n_0844_),
    .c(n_0845_)
  );
  and_bb n_1578_ (
    .a(N224),
    .b(N18),
    .c(n_0846_)
  );
  and_bi n_1579_ (
    .a(N121),
    .b(N18),
    .c(n_0847_)
  );
  or_bb n_1580_ (
    .a(n_0847_),
    .b(n_0846_),
    .c(n_0848_)
  );
  and_bb n_1581_ (
    .a(N223),
    .b(N18),
    .c(n_0849_)
  );
  and_bi n_1582_ (
    .a(N47),
    .b(N18),
    .c(n_0850_)
  );
  and_ii n_1583_ (
    .a(n_0850_),
    .b(n_0849_),
    .c(n_0851_)
  );
  or_bb n_1584_ (
    .a(n_0851_),
    .b(n_0848_),
    .c(n_0852_)
  );
  and_bb n_1585_ (
    .a(n_0851_),
    .b(n_0848_),
    .c(n_0853_)
  );
  and_bi n_1586_ (
    .a(n_0852_),
    .b(n_0853_),
    .c(n_0854_)
  );
  or_ii n_1587_ (
    .a(N226),
    .b(N18),
    .c(n_0855_)
  );
  and_bi n_1588_ (
    .a(N97),
    .b(N18),
    .c(n_0856_)
  );
  and_bi n_1589_ (
    .a(n_0855_),
    .b(n_0856_),
    .c(n_0857_)
  );
  and_bb n_1590_ (
    .a(N225),
    .b(N18),
    .c(n_0858_)
  );
  and_bi n_1591_ (
    .a(N94),
    .b(N18),
    .c(n_0859_)
  );
  and_ii n_1592_ (
    .a(n_0859_),
    .b(n_0858_),
    .c(n_0860_)
  );
  and_ii n_1593_ (
    .a(n_0860_),
    .b(n_0857_),
    .c(n_0861_)
  );
  and_bb n_1594_ (
    .a(n_0860_),
    .b(n_0857_),
    .c(n_0862_)
  );
  and_ii n_1595_ (
    .a(n_0862_),
    .b(n_0861_),
    .c(n_0863_)
  );
  or_bb n_1596_ (
    .a(n_0863_),
    .b(n_0854_),
    .c(n_0864_)
  );
  and_bb n_1597_ (
    .a(n_0863_),
    .b(n_0854_),
    .c(n_0865_)
  );
  and_bi n_1598_ (
    .a(n_0864_),
    .b(n_0865_),
    .c(n_0866_)
  );
  and_bb n_1599_ (
    .a(N227),
    .b(N18),
    .c(n_0867_)
  );
  and_bi n_1600_ (
    .a(N115),
    .b(N18),
    .c(n_0868_)
  );
  and_ii n_1601_ (
    .a(n_0868_),
    .b(n_0867_),
    .c(n_0869_)
  );
  or_ii n_1602_ (
    .a(N217),
    .b(N18),
    .c(n_0870_)
  );
  and_bi n_1603_ (
    .a(N118),
    .b(N18),
    .c(n_0871_)
  );
  and_bi n_1604_ (
    .a(n_0870_),
    .b(n_0871_),
    .c(n_0872_)
  );
  and_bb n_1605_ (
    .a(n_0872_),
    .b(n_0869_),
    .c(n_0873_)
  );
  and_ii n_1606_ (
    .a(n_0872_),
    .b(n_0869_),
    .c(n_0874_)
  );
  and_ii n_1607_ (
    .a(n_0874_),
    .b(n_0873_),
    .c(n_0875_)
  );
  and_bb n_1608_ (
    .a(N220),
    .b(N18),
    .c(n_0876_)
  );
  and_bi n_1609_ (
    .a(N50),
    .b(N18),
    .c(n_0877_)
  );
  and_ii n_1610_ (
    .a(n_0877_),
    .b(n_0876_),
    .c(n_0878_)
  );
  and_bb n_1611_ (
    .a(N219),
    .b(N18),
    .c(n_0879_)
  );
  and_bi n_1612_ (
    .a(N66),
    .b(N18),
    .c(n_0880_)
  );
  and_ii n_1613_ (
    .a(n_0880_),
    .b(n_0879_),
    .c(n_0881_)
  );
  and_bi n_1614_ (
    .a(n_0878_),
    .b(n_0881_),
    .c(n_0882_)
  );
  and_bi n_1615_ (
    .a(n_0881_),
    .b(n_0878_),
    .c(n_0883_)
  );
  and_ii n_1616_ (
    .a(n_0883_),
    .b(n_0882_),
    .c(n_0884_)
  );
  or_ii n_1617_ (
    .a(N222),
    .b(N18),
    .c(n_0885_)
  );
  and_bi n_1618_ (
    .a(N35),
    .b(N18),
    .c(n_0886_)
  );
  and_bi n_1619_ (
    .a(n_0885_),
    .b(n_0886_),
    .c(n_0887_)
  );
  or_ii n_1620_ (
    .a(N221),
    .b(N18),
    .c(n_0888_)
  );
  and_bi n_1621_ (
    .a(N32),
    .b(N18),
    .c(n_0889_)
  );
  and_bi n_1622_ (
    .a(n_0888_),
    .b(n_0889_),
    .c(n_0890_)
  );
  and_ii n_1623_ (
    .a(n_0890_),
    .b(n_0887_),
    .c(n_0891_)
  );
  and_bb n_1624_ (
    .a(n_0890_),
    .b(n_0887_),
    .c(n_0892_)
  );
  and_ii n_1625_ (
    .a(n_0892_),
    .b(n_0891_),
    .c(n_0893_)
  );
  and_bi n_1626_ (
    .a(n_0884_),
    .b(n_0893_),
    .c(n_0894_)
  );
  and_bi n_1627_ (
    .a(n_0893_),
    .b(n_0884_),
    .c(n_0895_)
  );
  and_ii n_1628_ (
    .a(n_0895_),
    .b(n_0894_),
    .c(n_0896_)
  );
  and_bi n_1629_ (
    .a(n_0896_),
    .b(n_0875_),
    .c(n_0897_)
  );
  and_bi n_1630_ (
    .a(n_0875_),
    .b(n_0896_),
    .c(n_0898_)
  );
  and_ii n_1631_ (
    .a(n_0898_),
    .b(n_0897_),
    .c(n_0899_)
  );
  or_bi n_1632_ (
    .a(n_0866_),
    .b(n_0899_),
    .c(n_0900_)
  );
  and_bi n_1633_ (
    .a(n_0866_),
    .b(n_0899_),
    .c(n_0901_)
  );
  and_bi n_1634_ (
    .a(n_0900_),
    .b(n_0901_),
    .c(n_0902_)
  );
  or_bb n_1635_ (
    .a(n_0902_),
    .b(n_0845_),
    .c(n_0903_)
  );
  or_bb n_1636_ (
    .a(n_0903_),
    .b(n_0801_),
    .c(N10574)
  );
  or_bi n_1637_ (
    .a(N18),
    .b(N114),
    .c(n_0904_)
  );
  and_bi n_1638_ (
    .a(N18),
    .b(N248),
    .c(n_0905_)
  );
  and_bi n_1639_ (
    .a(n_0904_),
    .b(n_0905_),
    .c(n_0906_)
  );
  and_bi n_1640_ (
    .a(N113),
    .b(N18),
    .c(n_0907_)
  );
  and_bi n_1641_ (
    .a(N18),
    .b(N251),
    .c(n_0908_)
  );
  and_ii n_1642_ (
    .a(n_0908_),
    .b(n_0907_),
    .c(n_0909_)
  );
  and_ii n_1643_ (
    .a(n_0909_),
    .b(n_0906_),
    .c(n_0910_)
  );
  and_bb n_1644_ (
    .a(n_0909_),
    .b(n_0906_),
    .c(n_0911_)
  );
  and_ii n_1645_ (
    .a(n_0911_),
    .b(n_0910_),
    .c(n_0912_)
  );
  and_bi n_1646_ (
    .a(N112),
    .b(N18),
    .c(n_0913_)
  );
  and_bi n_1647_ (
    .a(N18),
    .b(N257),
    .c(n_0914_)
  );
  and_ii n_1648_ (
    .a(n_0914_),
    .b(n_0913_),
    .c(n_0915_)
  );
  or_bi n_1649_ (
    .a(N18),
    .b(N88),
    .c(n_0916_)
  );
  and_bi n_1650_ (
    .a(N18),
    .b(N260),
    .c(n_0917_)
  );
  and_bi n_1651_ (
    .a(n_0916_),
    .b(n_0917_),
    .c(n_0918_)
  );
  and_bi n_1652_ (
    .a(n_0915_),
    .b(n_0918_),
    .c(n_0919_)
  );
  and_bi n_1653_ (
    .a(n_0918_),
    .b(n_0915_),
    .c(n_0920_)
  );
  and_ii n_1654_ (
    .a(n_0920_),
    .b(n_0919_),
    .c(n_0921_)
  );
  and_ii n_1655_ (
    .a(n_0921_),
    .b(n_0912_),
    .c(n_0922_)
  );
  and_bb n_1656_ (
    .a(n_0921_),
    .b(n_0912_),
    .c(n_0923_)
  );
  or_bb n_1657_ (
    .a(n_0923_),
    .b(n_0922_),
    .c(n_0924_)
  );
  and_bi n_1658_ (
    .a(N111),
    .b(N18),
    .c(n_0925_)
  );
  and_bi n_1659_ (
    .a(N18),
    .b(N254),
    .c(n_0926_)
  );
  and_ii n_1660_ (
    .a(n_0926_),
    .b(n_0925_),
    .c(n_0927_)
  );
  and_bi n_1661_ (
    .a(N87),
    .b(N18),
    .c(n_0928_)
  );
  and_bi n_1662_ (
    .a(N18),
    .b(N106),
    .c(n_0929_)
  );
  and_ii n_1663_ (
    .a(n_0929_),
    .b(n_0928_),
    .c(n_0930_)
  );
  and_ii n_1664_ (
    .a(n_0930_),
    .b(n_0927_),
    .c(n_0931_)
  );
  and_bb n_1665_ (
    .a(n_0930_),
    .b(n_0927_),
    .c(n_0932_)
  );
  and_ii n_1666_ (
    .a(n_0932_),
    .b(n_0931_),
    .c(n_0933_)
  );
  or_bi n_1667_ (
    .a(N267),
    .b(N263),
    .c(n_0934_)
  );
  and_bi n_1668_ (
    .a(N267),
    .b(N263),
    .c(n_0935_)
  );
  and_bi n_1669_ (
    .a(n_0934_),
    .b(n_0935_),
    .c(n_0936_)
  );
  and_bi n_1670_ (
    .a(N18),
    .b(n_0936_),
    .c(n_0937_)
  );
  or_bb n_1671_ (
    .a(N271),
    .b(N245),
    .c(n_0938_)
  );
  and_bb n_1672_ (
    .a(N271),
    .b(N245),
    .c(n_0939_)
  );
  or_bb n_1673_ (
    .a(n_0939_),
    .b(N18),
    .c(n_0940_)
  );
  and_bi n_1674_ (
    .a(n_0938_),
    .b(n_0940_),
    .c(n_0941_)
  );
  and_ii n_1675_ (
    .a(n_0941_),
    .b(n_0937_),
    .c(n_0942_)
  );
  and_ii n_1676_ (
    .a(n_0942_),
    .b(n_0933_),
    .c(n_0943_)
  );
  and_bb n_1677_ (
    .a(n_0942_),
    .b(n_0933_),
    .c(n_0944_)
  );
  and_ii n_1678_ (
    .a(n_0944_),
    .b(n_0943_),
    .c(n_0945_)
  );
  or_bb n_1679_ (
    .a(n_0945_),
    .b(n_0924_),
    .c(n_0946_)
  );
  and_bb n_1680_ (
    .a(n_0945_),
    .b(n_0924_),
    .c(n_0947_)
  );
  and_bi n_1681_ (
    .a(n_0946_),
    .b(n_0947_),
    .c(n_0948_)
  );
  and_bb n_1682_ (
    .a(N18),
    .b(N310),
    .c(n_0949_)
  );
  and_ii n_1683_ (
    .a(N70),
    .b(N18),
    .c(n_0950_)
  );
  and_ii n_1684_ (
    .a(n_0950_),
    .b(n_0949_),
    .c(n_0951_)
  );
  and_bi n_1685_ (
    .a(N69),
    .b(N18),
    .c(n_0952_)
  );
  and_bi n_1686_ (
    .a(N18),
    .b(N307),
    .c(n_0953_)
  );
  and_ii n_1687_ (
    .a(n_0953_),
    .b(n_0952_),
    .c(n_0954_)
  );
  and_bi n_1688_ (
    .a(n_0951_),
    .b(n_0954_),
    .c(n_0955_)
  );
  and_bi n_1689_ (
    .a(n_0954_),
    .b(n_0951_),
    .c(n_0956_)
  );
  and_ii n_1690_ (
    .a(n_0956_),
    .b(n_0955_),
    .c(n_0957_)
  );
  and_bi n_1691_ (
    .a(N76),
    .b(N18),
    .c(n_0958_)
  );
  and_bi n_1692_ (
    .a(N18),
    .b(N316),
    .c(n_0959_)
  );
  and_ii n_1693_ (
    .a(n_0959_),
    .b(n_0958_),
    .c(n_0960_)
  );
  and_bi n_1694_ (
    .a(N74),
    .b(N18),
    .c(n_0961_)
  );
  and_bi n_1695_ (
    .a(N18),
    .b(N313),
    .c(n_0962_)
  );
  and_ii n_1696_ (
    .a(n_0962_),
    .b(n_0961_),
    .c(n_0963_)
  );
  and_ii n_1697_ (
    .a(n_0963_),
    .b(n_0960_),
    .c(n_0964_)
  );
  and_bb n_1698_ (
    .a(n_0963_),
    .b(n_0960_),
    .c(n_0965_)
  );
  and_ii n_1699_ (
    .a(n_0965_),
    .b(n_0964_),
    .c(n_0966_)
  );
  and_bi n_1700_ (
    .a(n_0957_),
    .b(n_0966_),
    .c(n_0967_)
  );
  and_bi n_1701_ (
    .a(n_0966_),
    .b(n_0957_),
    .c(n_0968_)
  );
  or_bb n_1702_ (
    .a(n_0968_),
    .b(n_0967_),
    .c(n_0969_)
  );
  and_bi n_1703_ (
    .a(N55),
    .b(N18),
    .c(n_0970_)
  );
  and_bi n_1704_ (
    .a(N18),
    .b(N331),
    .c(n_0971_)
  );
  and_ii n_1705_ (
    .a(n_0971_),
    .b(n_0970_),
    .c(n_0972_)
  );
  and_bi n_1706_ (
    .a(N56),
    .b(N18),
    .c(n_0973_)
  );
  and_bi n_1707_ (
    .a(N18),
    .b(N334),
    .c(n_0974_)
  );
  and_ii n_1708_ (
    .a(n_0974_),
    .b(n_0973_),
    .c(n_0975_)
  );
  and_bi n_1709_ (
    .a(n_0972_),
    .b(n_0975_),
    .c(n_0976_)
  );
  and_bi n_1710_ (
    .a(n_0975_),
    .b(n_0972_),
    .c(n_0977_)
  );
  and_ii n_1711_ (
    .a(n_0977_),
    .b(n_0976_),
    .c(n_0978_)
  );
  and_bi n_1712_ (
    .a(N54),
    .b(N18),
    .c(n_0979_)
  );
  and_bi n_1713_ (
    .a(N18),
    .b(N328),
    .c(n_0980_)
  );
  and_ii n_1714_ (
    .a(n_0980_),
    .b(n_0979_),
    .c(n_0981_)
  );
  and_bi n_1715_ (
    .a(n_0978_),
    .b(n_0981_),
    .c(n_0982_)
  );
  and_bi n_1716_ (
    .a(n_0981_),
    .b(n_0978_),
    .c(n_0983_)
  );
  or_bb n_1717_ (
    .a(n_0983_),
    .b(n_0982_),
    .c(n_0984_)
  );
  and_bi n_1718_ (
    .a(N75),
    .b(N18),
    .c(n_0985_)
  );
  and_bi n_1719_ (
    .a(N18),
    .b(N319),
    .c(n_0986_)
  );
  and_ii n_1720_ (
    .a(n_0986_),
    .b(n_0985_),
    .c(n_0987_)
  );
  and_bi n_1721_ (
    .a(N73),
    .b(N18),
    .c(n_0988_)
  );
  and_bi n_1722_ (
    .a(N18),
    .b(N322),
    .c(n_0989_)
  );
  and_ii n_1723_ (
    .a(n_0989_),
    .b(n_0988_),
    .c(n_0990_)
  );
  and_bi n_1724_ (
    .a(N53),
    .b(N18),
    .c(n_0991_)
  );
  and_bi n_1725_ (
    .a(N18),
    .b(N325),
    .c(n_0992_)
  );
  and_ii n_1726_ (
    .a(n_0992_),
    .b(n_0991_),
    .c(n_0993_)
  );
  and_ii n_1727_ (
    .a(n_0993_),
    .b(n_0990_),
    .c(n_0994_)
  );
  and_bb n_1728_ (
    .a(n_0993_),
    .b(n_0990_),
    .c(n_0995_)
  );
  or_bb n_1729_ (
    .a(n_0995_),
    .b(n_0994_),
    .c(n_0996_)
  );
  or_bb n_1730_ (
    .a(n_0996_),
    .b(n_0987_),
    .c(n_0997_)
  );
  or_ii n_1731_ (
    .a(n_0996_),
    .b(n_0987_),
    .c(n_0998_)
  );
  and_bb n_1732_ (
    .a(n_0998_),
    .b(n_0997_),
    .c(n_0999_)
  );
  and_bi n_1733_ (
    .a(n_0999_),
    .b(n_0984_),
    .c(n_1000_)
  );
  and_bi n_1734_ (
    .a(n_0984_),
    .b(n_0999_),
    .c(n_1001_)
  );
  and_ii n_1735_ (
    .a(n_1001_),
    .b(n_1000_),
    .c(n_1002_)
  );
  or_bb n_1736_ (
    .a(n_1002_),
    .b(n_0969_),
    .c(n_1003_)
  );
  and_bb n_1737_ (
    .a(n_1002_),
    .b(n_0969_),
    .c(n_1004_)
  );
  and_bi n_1738_ (
    .a(n_1003_),
    .b(n_1004_),
    .c(n_1005_)
  );
  or_bb n_1739_ (
    .a(n_1005_),
    .b(n_0948_),
    .c(n_1006_)
  );
  and_bi n_1740_ (
    .a(N81),
    .b(N18),
    .c(n_1007_)
  );
  and_bi n_1741_ (
    .a(N18),
    .b(N349),
    .c(n_1008_)
  );
  and_ii n_1742_ (
    .a(n_1008_),
    .b(n_1007_),
    .c(n_1009_)
  );
  and_bi n_1743_ (
    .a(N80),
    .b(N18),
    .c(n_1010_)
  );
  and_bi n_1744_ (
    .a(N18),
    .b(N352),
    .c(n_1011_)
  );
  and_ii n_1745_ (
    .a(n_1011_),
    .b(n_1010_),
    .c(n_1012_)
  );
  or_bb n_1746_ (
    .a(n_1012_),
    .b(n_1009_),
    .c(n_1013_)
  );
  and_bb n_1747_ (
    .a(n_1012_),
    .b(n_1009_),
    .c(n_1014_)
  );
  and_bi n_1748_ (
    .a(n_1013_),
    .b(n_1014_),
    .c(n_1015_)
  );
  and_bi n_1749_ (
    .a(N61),
    .b(N18),
    .c(n_1016_)
  );
  and_bi n_1750_ (
    .a(N18),
    .b(N361),
    .c(n_1017_)
  );
  and_ii n_1751_ (
    .a(n_1017_),
    .b(n_1016_),
    .c(n_1018_)
  );
  and_bi n_1752_ (
    .a(N62),
    .b(N18),
    .c(n_1019_)
  );
  and_bi n_1753_ (
    .a(N18),
    .b(N364),
    .c(n_1020_)
  );
  and_ii n_1754_ (
    .a(n_1020_),
    .b(n_1019_),
    .c(n_1021_)
  );
  and_bi n_1755_ (
    .a(n_1018_),
    .b(n_1021_),
    .c(n_1022_)
  );
  and_bi n_1756_ (
    .a(n_1021_),
    .b(n_1018_),
    .c(n_1023_)
  );
  and_ii n_1757_ (
    .a(n_1023_),
    .b(n_1022_),
    .c(n_1024_)
  );
  or_bi n_1758_ (
    .a(n_1015_),
    .b(n_1024_),
    .c(n_1025_)
  );
  and_bi n_1759_ (
    .a(n_1015_),
    .b(n_1024_),
    .c(n_1026_)
  );
  and_bi n_1760_ (
    .a(n_1025_),
    .b(n_1026_),
    .c(n_1027_)
  );
  and_bi n_1761_ (
    .a(N78),
    .b(N18),
    .c(n_1028_)
  );
  and_bi n_1762_ (
    .a(N18),
    .b(N343),
    .c(n_1029_)
  );
  and_ii n_1763_ (
    .a(n_1029_),
    .b(n_1028_),
    .c(n_1030_)
  );
  and_bi n_1764_ (
    .a(N59),
    .b(N18),
    .c(n_1031_)
  );
  and_bi n_1765_ (
    .a(N18),
    .b(N346),
    .c(n_1032_)
  );
  and_ii n_1766_ (
    .a(n_1032_),
    .b(n_1031_),
    .c(n_1033_)
  );
  and_ii n_1767_ (
    .a(n_1033_),
    .b(n_1030_),
    .c(n_1034_)
  );
  and_bb n_1768_ (
    .a(n_1033_),
    .b(n_1030_),
    .c(n_1035_)
  );
  and_ii n_1769_ (
    .a(n_1035_),
    .b(n_1034_),
    .c(n_1036_)
  );
  or_bi n_1770_ (
    .a(n_1027_),
    .b(n_1036_),
    .c(n_1037_)
  );
  and_bi n_1771_ (
    .a(n_1027_),
    .b(n_1036_),
    .c(n_1038_)
  );
  and_bi n_1772_ (
    .a(n_1037_),
    .b(n_1038_),
    .c(n_1039_)
  );
  and_bi n_1773_ (
    .a(N79),
    .b(N18),
    .c(n_1040_)
  );
  and_bi n_1774_ (
    .a(N18),
    .b(N355),
    .c(n_1041_)
  );
  and_ii n_1775_ (
    .a(n_1041_),
    .b(n_1040_),
    .c(n_1042_)
  );
  and_bi n_1776_ (
    .a(N60),
    .b(N18),
    .c(n_1043_)
  );
  and_bi n_1777_ (
    .a(N18),
    .b(N358),
    .c(n_1044_)
  );
  and_ii n_1778_ (
    .a(n_1044_),
    .b(n_1043_),
    .c(n_1045_)
  );
  and_ii n_1779_ (
    .a(n_1045_),
    .b(n_1042_),
    .c(n_1046_)
  );
  and_bb n_1780_ (
    .a(n_1045_),
    .b(n_1042_),
    .c(n_1047_)
  );
  and_ii n_1781_ (
    .a(n_1047_),
    .b(n_1046_),
    .c(n_1048_)
  );
  and_bi n_1782_ (
    .a(N58),
    .b(N18),
    .c(n_1049_)
  );
  and_bi n_1783_ (
    .a(N18),
    .b(N337),
    .c(n_1050_)
  );
  and_ii n_1784_ (
    .a(n_1050_),
    .b(n_1049_),
    .c(n_1051_)
  );
  and_bi n_1785_ (
    .a(N77),
    .b(N18),
    .c(n_1052_)
  );
  and_bi n_1786_ (
    .a(N18),
    .b(N340),
    .c(n_1053_)
  );
  and_ii n_1787_ (
    .a(n_1053_),
    .b(n_1052_),
    .c(n_1054_)
  );
  and_ii n_1788_ (
    .a(n_1054_),
    .b(n_1051_),
    .c(n_1055_)
  );
  and_bb n_1789_ (
    .a(n_1054_),
    .b(n_1051_),
    .c(n_1056_)
  );
  and_ii n_1790_ (
    .a(n_1056_),
    .b(n_1055_),
    .c(n_1057_)
  );
  and_ii n_1791_ (
    .a(n_1057_),
    .b(n_1048_),
    .c(n_1058_)
  );
  and_bb n_1792_ (
    .a(n_1057_),
    .b(n_1048_),
    .c(n_1059_)
  );
  and_ii n_1793_ (
    .a(n_1059_),
    .b(n_1058_),
    .c(n_1060_)
  );
  or_bb n_1794_ (
    .a(n_1060_),
    .b(n_1039_),
    .c(n_1061_)
  );
  and_bb n_1795_ (
    .a(n_1060_),
    .b(n_1039_),
    .c(n_1062_)
  );
  and_bi n_1796_ (
    .a(n_1061_),
    .b(n_1062_),
    .c(n_1063_)
  );
  and_bi n_1797_ (
    .a(N85),
    .b(N18),
    .c(n_1064_)
  );
  and_bi n_1798_ (
    .a(N18),
    .b(N286),
    .c(n_1065_)
  );
  and_ii n_1799_ (
    .a(n_1065_),
    .b(n_1064_),
    .c(n_1066_)
  );
  and_bi n_1800_ (
    .a(N64),
    .b(N18),
    .c(n_1067_)
  );
  and_bi n_1801_ (
    .a(N18),
    .b(N289),
    .c(n_1068_)
  );
  and_ii n_1802_ (
    .a(n_1068_),
    .b(n_1067_),
    .c(n_1069_)
  );
  or_bb n_1803_ (
    .a(n_1069_),
    .b(n_1066_),
    .c(n_1070_)
  );
  and_bb n_1804_ (
    .a(n_1069_),
    .b(n_1066_),
    .c(n_1071_)
  );
  and_bi n_1805_ (
    .a(n_1070_),
    .b(n_1071_),
    .c(n_1072_)
  );
  and_bi n_1806_ (
    .a(N109),
    .b(N18),
    .c(n_1073_)
  );
  and_bi n_1807_ (
    .a(N18),
    .b(N299),
    .c(n_1074_)
  );
  and_ii n_1808_ (
    .a(n_1074_),
    .b(n_1073_),
    .c(n_1075_)
  );
  and_bi n_1809_ (
    .a(N110),
    .b(N18),
    .c(n_1076_)
  );
  and_bi n_1810_ (
    .a(N18),
    .b(N303),
    .c(n_1077_)
  );
  and_ii n_1811_ (
    .a(n_1077_),
    .b(n_1076_),
    .c(n_1078_)
  );
  or_bi n_1812_ (
    .a(n_1078_),
    .b(n_1075_),
    .c(n_1079_)
  );
  and_bi n_1813_ (
    .a(n_1078_),
    .b(n_1075_),
    .c(n_1080_)
  );
  and_bi n_1814_ (
    .a(n_1079_),
    .b(n_1080_),
    .c(n_1081_)
  );
  and_ii n_1815_ (
    .a(n_1081_),
    .b(n_1072_),
    .c(n_1082_)
  );
  and_bb n_1816_ (
    .a(n_1081_),
    .b(n_1072_),
    .c(n_1083_)
  );
  and_ii n_1817_ (
    .a(n_1083_),
    .b(n_1082_),
    .c(n_1084_)
  );
  and_bi n_1818_ (
    .a(N82),
    .b(N18),
    .c(n_1085_)
  );
  and_bi n_1819_ (
    .a(N18),
    .b(N274),
    .c(n_1086_)
  );
  and_ii n_1820_ (
    .a(n_1086_),
    .b(n_1085_),
    .c(n_1087_)
  );
  and_bi n_1821_ (
    .a(N65),
    .b(N18),
    .c(n_1088_)
  );
  and_bi n_1822_ (
    .a(N18),
    .b(N277),
    .c(n_1089_)
  );
  and_ii n_1823_ (
    .a(n_1089_),
    .b(n_1088_),
    .c(n_1090_)
  );
  and_bi n_1824_ (
    .a(n_1087_),
    .b(n_1090_),
    .c(n_1091_)
  );
  and_bi n_1825_ (
    .a(n_1090_),
    .b(n_1087_),
    .c(n_1092_)
  );
  and_ii n_1826_ (
    .a(n_1092_),
    .b(n_1091_),
    .c(n_1093_)
  );
  and_bi n_1827_ (
    .a(N84),
    .b(N18),
    .c(n_1094_)
  );
  and_bi n_1828_ (
    .a(N18),
    .b(N283),
    .c(n_1095_)
  );
  and_ii n_1829_ (
    .a(n_1095_),
    .b(n_1094_),
    .c(n_1096_)
  );
  or_ii n_1830_ (
    .a(n_1096_),
    .b(n_1093_),
    .c(n_1097_)
  );
  or_bb n_1831_ (
    .a(n_1096_),
    .b(n_1093_),
    .c(n_1098_)
  );
  or_ii n_1832_ (
    .a(n_1098_),
    .b(n_1097_),
    .c(n_1099_)
  );
  and_bi n_1833_ (
    .a(N63),
    .b(N18),
    .c(n_1100_)
  );
  and_bi n_1834_ (
    .a(N18),
    .b(N293),
    .c(n_1101_)
  );
  and_ii n_1835_ (
    .a(n_1101_),
    .b(n_1100_),
    .c(n_1102_)
  );
  and_bi n_1836_ (
    .a(N86),
    .b(N18),
    .c(n_1103_)
  );
  and_bi n_1837_ (
    .a(N18),
    .b(N296),
    .c(n_1104_)
  );
  and_ii n_1838_ (
    .a(n_1104_),
    .b(n_1103_),
    .c(n_1105_)
  );
  and_bi n_1839_ (
    .a(n_1102_),
    .b(n_1105_),
    .c(n_1106_)
  );
  and_bi n_1840_ (
    .a(n_1105_),
    .b(n_1102_),
    .c(n_1107_)
  );
  and_ii n_1841_ (
    .a(n_1107_),
    .b(n_1106_),
    .c(n_1108_)
  );
  and_bi n_1842_ (
    .a(N83),
    .b(N18),
    .c(n_1109_)
  );
  and_bi n_1843_ (
    .a(N18),
    .b(N280),
    .c(n_1110_)
  );
  and_ii n_1844_ (
    .a(n_1110_),
    .b(n_1109_),
    .c(n_1111_)
  );
  or_bb n_1845_ (
    .a(n_1111_),
    .b(n_1108_),
    .c(n_1112_)
  );
  or_ii n_1846_ (
    .a(n_1111_),
    .b(n_1108_),
    .c(n_1113_)
  );
  or_ii n_1847_ (
    .a(n_1113_),
    .b(n_1112_),
    .c(n_1114_)
  );
  and_ii n_1848_ (
    .a(n_1114_),
    .b(n_1099_),
    .c(n_1115_)
  );
  and_bb n_1849_ (
    .a(n_1114_),
    .b(n_1099_),
    .c(n_1116_)
  );
  and_ii n_1850_ (
    .a(n_1116_),
    .b(n_1115_),
    .c(n_1117_)
  );
  and_bi n_1851_ (
    .a(n_1117_),
    .b(n_1084_),
    .c(n_1118_)
  );
  and_bi n_1852_ (
    .a(n_1084_),
    .b(n_1117_),
    .c(n_1119_)
  );
  or_bb n_1853_ (
    .a(n_1119_),
    .b(n_1118_),
    .c(n_1120_)
  );
  or_bb n_1854_ (
    .a(n_1120_),
    .b(n_1063_),
    .c(n_1121_)
  );
  or_bb n_1855_ (
    .a(n_1121_),
    .b(n_1006_),
    .c(N10575)
  );
  and_ii n_1856_ (
    .a(n_0788_),
    .b(N170),
    .c(n_1122_)
  );
  and_bi n_1857_ (
    .a(N18),
    .b(N167),
    .c(n_1123_)
  );
  and_ii n_1858_ (
    .a(n_1123_),
    .b(n_0718_),
    .c(n_1124_)
  );
  and_bi n_1859_ (
    .a(N18),
    .b(N166),
    .c(n_1125_)
  );
  and_bb n_1860_ (
    .a(n_1125_),
    .b(n_1124_),
    .c(n_1126_)
  );
  or_bb n_1861_ (
    .a(n_1125_),
    .b(n_0718_),
    .c(n_1127_)
  );
  and_bi n_1862_ (
    .a(n_1123_),
    .b(n_1127_),
    .c(n_1128_)
  );
  and_ii n_1863_ (
    .a(n_1128_),
    .b(n_1126_),
    .c(n_1129_)
  );
  and_ii n_1864_ (
    .a(n_1129_),
    .b(n_1122_),
    .c(n_1130_)
  );
  and_bb n_1865_ (
    .a(n_1129_),
    .b(n_1122_),
    .c(n_1131_)
  );
  or_bb n_1866_ (
    .a(n_1131_),
    .b(n_1130_),
    .c(n_1132_)
  );
  and_bi n_1867_ (
    .a(N18),
    .b(N169),
    .c(n_1133_)
  );
  and_ii n_1868_ (
    .a(n_1133_),
    .b(n_0718_),
    .c(n_1134_)
  );
  and_bi n_1869_ (
    .a(N18),
    .b(N168),
    .c(n_1135_)
  );
  and_bb n_1870_ (
    .a(n_1135_),
    .b(n_1134_),
    .c(n_1136_)
  );
  and_ii n_1871_ (
    .a(n_1135_),
    .b(n_0718_),
    .c(n_1137_)
  );
  and_bb n_1872_ (
    .a(n_1137_),
    .b(n_1133_),
    .c(n_1138_)
  );
  and_ii n_1873_ (
    .a(n_1138_),
    .b(n_1136_),
    .c(n_1139_)
  );
  or_bi n_1874_ (
    .a(N164),
    .b(N165),
    .c(n_1140_)
  );
  and_bi n_1875_ (
    .a(N164),
    .b(N165),
    .c(n_1141_)
  );
  and_bi n_1876_ (
    .a(n_1140_),
    .b(n_1141_),
    .c(n_1142_)
  );
  and_ii n_1877_ (
    .a(n_1142_),
    .b(n_0788_),
    .c(n_1143_)
  );
  and_bi n_1878_ (
    .a(n_1139_),
    .b(n_1143_),
    .c(n_1144_)
  );
  and_bi n_1879_ (
    .a(n_1143_),
    .b(n_1139_),
    .c(n_1145_)
  );
  and_ii n_1880_ (
    .a(n_1145_),
    .b(n_1144_),
    .c(n_1146_)
  );
  or_bb n_1881_ (
    .a(n_1146_),
    .b(n_1132_),
    .c(n_1147_)
  );
  and_bb n_1882_ (
    .a(n_1146_),
    .b(n_1132_),
    .c(n_1148_)
  );
  and_bi n_1883_ (
    .a(n_1147_),
    .b(n_1148_),
    .c(n_1149_)
  );
  and_bb n_1884_ (
    .a(N196),
    .b(N18),
    .c(n_1150_)
  );
  and_ii n_1885_ (
    .a(n_1150_),
    .b(n_0856_),
    .c(n_1151_)
  );
  and_bb n_1886_ (
    .a(N195),
    .b(N18),
    .c(n_1152_)
  );
  and_ii n_1887_ (
    .a(n_1152_),
    .b(n_0859_),
    .c(n_1153_)
  );
  and_ii n_1888_ (
    .a(n_1153_),
    .b(n_1151_),
    .c(n_1154_)
  );
  and_bb n_1889_ (
    .a(n_1153_),
    .b(n_1151_),
    .c(n_1155_)
  );
  and_ii n_1890_ (
    .a(n_1155_),
    .b(n_1154_),
    .c(n_1156_)
  );
  and_bb n_1891_ (
    .a(N190),
    .b(N18),
    .c(n_1157_)
  );
  and_ii n_1892_ (
    .a(n_1157_),
    .b(n_0877_),
    .c(n_1158_)
  );
  and_bb n_1893_ (
    .a(N189),
    .b(N18),
    .c(n_1159_)
  );
  and_ii n_1894_ (
    .a(n_1159_),
    .b(n_0880_),
    .c(n_1160_)
  );
  and_bi n_1895_ (
    .a(n_1158_),
    .b(n_1160_),
    .c(n_1161_)
  );
  and_bi n_1896_ (
    .a(n_1160_),
    .b(n_1158_),
    .c(n_1162_)
  );
  and_ii n_1897_ (
    .a(n_1162_),
    .b(n_1161_),
    .c(n_1163_)
  );
  and_bb n_1898_ (
    .a(N192),
    .b(N18),
    .c(n_1164_)
  );
  and_ii n_1899_ (
    .a(n_1164_),
    .b(n_0886_),
    .c(n_1165_)
  );
  and_bb n_1900_ (
    .a(N191),
    .b(N18),
    .c(n_1166_)
  );
  and_ii n_1901_ (
    .a(n_1166_),
    .b(n_0889_),
    .c(n_1167_)
  );
  and_ii n_1902_ (
    .a(n_1167_),
    .b(n_1165_),
    .c(n_1168_)
  );
  and_bb n_1903_ (
    .a(n_1167_),
    .b(n_1165_),
    .c(n_1169_)
  );
  and_ii n_1904_ (
    .a(n_1169_),
    .b(n_1168_),
    .c(n_1170_)
  );
  and_bb n_1905_ (
    .a(n_1170_),
    .b(n_1163_),
    .c(n_1171_)
  );
  and_ii n_1906_ (
    .a(n_1170_),
    .b(n_1163_),
    .c(n_1172_)
  );
  and_ii n_1907_ (
    .a(n_1172_),
    .b(n_1171_),
    .c(n_1173_)
  );
  and_bi n_1908_ (
    .a(n_1156_),
    .b(n_1173_),
    .c(n_1174_)
  );
  and_bi n_1909_ (
    .a(n_1173_),
    .b(n_1156_),
    .c(n_1175_)
  );
  and_ii n_1910_ (
    .a(n_1175_),
    .b(n_1174_),
    .c(n_1176_)
  );
  and_bb n_1911_ (
    .a(N194),
    .b(N18),
    .c(n_1177_)
  );
  and_ii n_1912_ (
    .a(n_1177_),
    .b(n_0847_),
    .c(n_1178_)
  );
  and_bb n_1913_ (
    .a(N193),
    .b(N18),
    .c(n_1179_)
  );
  and_ii n_1914_ (
    .a(n_1179_),
    .b(n_0850_),
    .c(n_1180_)
  );
  and_ii n_1915_ (
    .a(n_1180_),
    .b(n_1178_),
    .c(n_1181_)
  );
  and_bb n_1916_ (
    .a(n_1180_),
    .b(n_1178_),
    .c(n_1182_)
  );
  and_ii n_1917_ (
    .a(n_1182_),
    .b(n_1181_),
    .c(n_1183_)
  );
  and_bb n_1918_ (
    .a(N197),
    .b(N18),
    .c(n_1184_)
  );
  and_ii n_1919_ (
    .a(n_1184_),
    .b(n_0868_),
    .c(n_1185_)
  );
  and_bb n_1920_ (
    .a(N187),
    .b(N18),
    .c(n_1186_)
  );
  and_ii n_1921_ (
    .a(n_1186_),
    .b(n_0871_),
    .c(n_1187_)
  );
  and_bb n_1922_ (
    .a(n_1187_),
    .b(n_1185_),
    .c(n_1188_)
  );
  and_ii n_1923_ (
    .a(n_1187_),
    .b(n_1185_),
    .c(n_1189_)
  );
  and_ii n_1924_ (
    .a(n_1189_),
    .b(n_1188_),
    .c(n_1190_)
  );
  and_bi n_1925_ (
    .a(n_1190_),
    .b(n_1183_),
    .c(n_1191_)
  );
  and_bi n_1926_ (
    .a(n_1183_),
    .b(n_1190_),
    .c(n_1192_)
  );
  and_ii n_1927_ (
    .a(n_1192_),
    .b(n_1191_),
    .c(n_1193_)
  );
  and_bi n_1928_ (
    .a(n_1193_),
    .b(n_1176_),
    .c(n_1194_)
  );
  and_bi n_1929_ (
    .a(n_1176_),
    .b(n_1193_),
    .c(n_1195_)
  );
  or_bb n_1930_ (
    .a(n_1195_),
    .b(n_1194_),
    .c(n_1196_)
  );
  or_bb n_1931_ (
    .a(n_1196_),
    .b(n_1149_),
    .c(n_1197_)
  );
  and_bb n_1932_ (
    .a(N181),
    .b(N18),
    .c(n_1198_)
  );
  and_ii n_1933_ (
    .a(n_1198_),
    .b(n_0733_),
    .c(n_1199_)
  );
  and_bb n_1934_ (
    .a(N171),
    .b(N18),
    .c(n_1200_)
  );
  and_ii n_1935_ (
    .a(n_1200_),
    .b(n_0736_),
    .c(n_1201_)
  );
  and_bi n_1936_ (
    .a(n_1199_),
    .b(n_1201_),
    .c(n_1202_)
  );
  and_bi n_1937_ (
    .a(n_1201_),
    .b(n_1199_),
    .c(n_1203_)
  );
  or_bb n_1938_ (
    .a(n_1203_),
    .b(n_1202_),
    .c(n_1204_)
  );
  and_bi n_1939_ (
    .a(N18),
    .b(N174),
    .c(n_1205_)
  );
  and_ii n_1940_ (
    .a(n_1205_),
    .b(n_0718_),
    .c(n_1206_)
  );
  and_bi n_1941_ (
    .a(N18),
    .b(N173),
    .c(n_1207_)
  );
  and_bb n_1942_ (
    .a(n_1207_),
    .b(n_1206_),
    .c(n_1208_)
  );
  and_ii n_1943_ (
    .a(n_1207_),
    .b(n_0718_),
    .c(n_1209_)
  );
  and_bb n_1944_ (
    .a(n_1209_),
    .b(n_1205_),
    .c(n_1210_)
  );
  and_ii n_1945_ (
    .a(n_1210_),
    .b(n_1208_),
    .c(n_1211_)
  );
  and_bi n_1946_ (
    .a(N18),
    .b(N176),
    .c(n_1212_)
  );
  and_ii n_1947_ (
    .a(n_1212_),
    .b(n_0718_),
    .c(n_1213_)
  );
  and_bi n_1948_ (
    .a(N18),
    .b(N175),
    .c(n_1214_)
  );
  and_bb n_1949_ (
    .a(n_1214_),
    .b(n_1213_),
    .c(n_1215_)
  );
  and_ii n_1950_ (
    .a(n_1214_),
    .b(n_0718_),
    .c(n_1216_)
  );
  and_bb n_1951_ (
    .a(n_1216_),
    .b(n_1212_),
    .c(n_1217_)
  );
  and_ii n_1952_ (
    .a(n_1217_),
    .b(n_1215_),
    .c(n_1218_)
  );
  and_bb n_1953_ (
    .a(n_1218_),
    .b(n_1211_),
    .c(n_1219_)
  );
  and_ii n_1954_ (
    .a(n_1218_),
    .b(n_1211_),
    .c(n_1220_)
  );
  or_bb n_1955_ (
    .a(n_1220_),
    .b(n_1219_),
    .c(n_1221_)
  );
  and_ii n_1956_ (
    .a(n_1221_),
    .b(n_1204_),
    .c(n_1222_)
  );
  and_bb n_1957_ (
    .a(n_1221_),
    .b(n_1204_),
    .c(n_1223_)
  );
  and_ii n_1958_ (
    .a(n_1223_),
    .b(n_1222_),
    .c(n_1224_)
  );
  and_bb n_1959_ (
    .a(N178),
    .b(N18),
    .c(n_1225_)
  );
  and_ii n_1960_ (
    .a(n_1225_),
    .b(n_0748_),
    .c(n_1226_)
  );
  and_bi n_1961_ (
    .a(N18),
    .b(N177),
    .c(n_1227_)
  );
  and_ii n_1962_ (
    .a(n_1227_),
    .b(n_0718_),
    .c(n_1228_)
  );
  and_ii n_1963_ (
    .a(n_1228_),
    .b(n_1226_),
    .c(n_1229_)
  );
  and_bb n_1964_ (
    .a(n_1228_),
    .b(n_1226_),
    .c(n_1230_)
  );
  and_ii n_1965_ (
    .a(n_1230_),
    .b(n_1229_),
    .c(n_1231_)
  );
  and_bb n_1966_ (
    .a(N180),
    .b(N18),
    .c(n_1232_)
  );
  and_ii n_1967_ (
    .a(n_1232_),
    .b(n_0756_),
    .c(n_1233_)
  );
  and_bb n_1968_ (
    .a(N179),
    .b(N18),
    .c(n_1234_)
  );
  and_ii n_1969_ (
    .a(n_1234_),
    .b(n_0759_),
    .c(n_1235_)
  );
  and_ii n_1970_ (
    .a(n_1235_),
    .b(n_1233_),
    .c(n_1236_)
  );
  and_bb n_1971_ (
    .a(n_1235_),
    .b(n_1233_),
    .c(n_1237_)
  );
  and_ii n_1972_ (
    .a(n_1237_),
    .b(n_1236_),
    .c(n_1238_)
  );
  and_bi n_1973_ (
    .a(n_1238_),
    .b(n_1231_),
    .c(n_1239_)
  );
  and_bi n_1974_ (
    .a(n_1231_),
    .b(n_1238_),
    .c(n_1240_)
  );
  and_ii n_1975_ (
    .a(n_1240_),
    .b(n_1239_),
    .c(n_1241_)
  );
  and_bi n_1976_ (
    .a(n_1224_),
    .b(n_1241_),
    .c(n_1242_)
  );
  and_bi n_1977_ (
    .a(n_1241_),
    .b(n_1224_),
    .c(n_1243_)
  );
  or_bb n_1978_ (
    .a(n_1243_),
    .b(n_1242_),
    .c(n_1244_)
  );
  and_bb n_1979_ (
    .a(N208),
    .b(N18),
    .c(n_1245_)
  );
  and_ii n_1980_ (
    .a(n_1245_),
    .b(n_0832_),
    .c(n_1246_)
  );
  and_bb n_1981_ (
    .a(N198),
    .b(N18),
    .c(n_1247_)
  );
  and_bi n_1982_ (
    .a(n_0662_),
    .b(n_1247_),
    .c(n_1248_)
  );
  and_bb n_1983_ (
    .a(n_1248_),
    .b(n_1246_),
    .c(n_1249_)
  );
  and_ii n_1984_ (
    .a(n_1248_),
    .b(n_1246_),
    .c(n_1250_)
  );
  and_ii n_1985_ (
    .a(n_1250_),
    .b(n_1249_),
    .c(n_1251_)
  );
  and_bb n_1986_ (
    .a(N207),
    .b(N18),
    .c(n_1252_)
  );
  and_ii n_1987_ (
    .a(n_1252_),
    .b(n_0688_),
    .c(n_1253_)
  );
  and_bb n_1988_ (
    .a(N206),
    .b(N18),
    .c(n_1254_)
  );
  and_ii n_1989_ (
    .a(n_1254_),
    .b(n_0682_),
    .c(n_1255_)
  );
  and_ii n_1990_ (
    .a(n_1255_),
    .b(n_1253_),
    .c(n_1256_)
  );
  and_bb n_1991_ (
    .a(n_1255_),
    .b(n_1253_),
    .c(n_1257_)
  );
  and_ii n_1992_ (
    .a(n_1257_),
    .b(n_1256_),
    .c(n_1258_)
  );
  and_bb n_1993_ (
    .a(N205),
    .b(N18),
    .c(n_1259_)
  );
  and_ii n_1994_ (
    .a(n_1259_),
    .b(n_0678_),
    .c(n_1260_)
  );
  and_bb n_1995_ (
    .a(N204),
    .b(N18),
    .c(n_1261_)
  );
  and_ii n_1996_ (
    .a(n_1261_),
    .b(n_0672_),
    .c(n_1262_)
  );
  and_bi n_1997_ (
    .a(n_1260_),
    .b(n_1262_),
    .c(n_1263_)
  );
  and_bi n_1998_ (
    .a(n_1262_),
    .b(n_1260_),
    .c(n_1264_)
  );
  and_ii n_1999_ (
    .a(n_1264_),
    .b(n_1263_),
    .c(n_1265_)
  );
  and_bi n_2000_ (
    .a(n_1265_),
    .b(n_1258_),
    .c(n_1266_)
  );
  and_bi n_2001_ (
    .a(n_1258_),
    .b(n_1265_),
    .c(n_1267_)
  );
  and_ii n_2002_ (
    .a(n_1267_),
    .b(n_1266_),
    .c(n_1268_)
  );
  and_ii n_2003_ (
    .a(n_1268_),
    .b(n_1251_),
    .c(n_1269_)
  );
  and_bb n_2004_ (
    .a(n_1268_),
    .b(n_1251_),
    .c(n_1270_)
  );
  and_ii n_2005_ (
    .a(n_1270_),
    .b(n_1269_),
    .c(n_1271_)
  );
  and_bb n_2006_ (
    .a(N201),
    .b(N18),
    .c(n_1272_)
  );
  and_ii n_2007_ (
    .a(n_1272_),
    .b(n_0803_),
    .c(n_1273_)
  );
  and_bb n_2008_ (
    .a(N200),
    .b(N18),
    .c(n_1274_)
  );
  and_ii n_2009_ (
    .a(n_1274_),
    .b(n_0811_),
    .c(n_1275_)
  );
  and_bi n_2010_ (
    .a(n_1273_),
    .b(n_1275_),
    .c(n_1276_)
  );
  and_bi n_2011_ (
    .a(n_1275_),
    .b(n_1273_),
    .c(n_1277_)
  );
  and_ii n_2012_ (
    .a(n_1277_),
    .b(n_1276_),
    .c(n_1278_)
  );
  and_bb n_2013_ (
    .a(N203),
    .b(N18),
    .c(n_1279_)
  );
  and_ii n_2014_ (
    .a(n_1279_),
    .b(n_0823_),
    .c(n_1280_)
  );
  and_bb n_2015_ (
    .a(N202),
    .b(N18),
    .c(n_1281_)
  );
  and_ii n_2016_ (
    .a(n_1281_),
    .b(n_0826_),
    .c(n_1282_)
  );
  and_ii n_2017_ (
    .a(n_1282_),
    .b(n_1280_),
    .c(n_1283_)
  );
  and_bb n_2018_ (
    .a(n_1282_),
    .b(n_1280_),
    .c(n_1284_)
  );
  and_ii n_2019_ (
    .a(n_1284_),
    .b(n_1283_),
    .c(n_1285_)
  );
  and_bi n_2020_ (
    .a(n_1278_),
    .b(n_1285_),
    .c(n_1286_)
  );
  and_bi n_2021_ (
    .a(n_1285_),
    .b(n_1278_),
    .c(n_1287_)
  );
  and_ii n_2022_ (
    .a(n_1287_),
    .b(n_1286_),
    .c(n_1288_)
  );
  and_bb n_2023_ (
    .a(n_1288_),
    .b(n_1271_),
    .c(n_1289_)
  );
  and_ii n_2024_ (
    .a(n_1288_),
    .b(n_1271_),
    .c(n_1290_)
  );
  or_bb n_2025_ (
    .a(n_1290_),
    .b(n_1289_),
    .c(n_1291_)
  );
  or_bb n_2026_ (
    .a(n_1291_),
    .b(n_1244_),
    .c(n_1292_)
  );
  or_bb n_2027_ (
    .a(n_1292_),
    .b(n_1197_),
    .c(N10576)
  );
  inv n_2028_ (
    .din(N277),
    .dout(n_1293_)
  );
  and_bi n_2029_ (
    .a(n_1293_),
    .b(n_0738_),
    .c(n_1294_)
  );
  and_bi n_2030_ (
    .a(n_0738_),
    .b(n_1293_),
    .c(n_1295_)
  );
  and_ii n_2031_ (
    .a(n_1295_),
    .b(n_1294_),
    .c(n_1296_)
  );
  inv n_2032_ (
    .din(N364),
    .dout(n_1297_)
  );
  and_bi n_2033_ (
    .a(n_1297_),
    .b(n_0881_),
    .c(n_1298_)
  );
  and_bi n_2034_ (
    .a(n_0881_),
    .b(n_1297_),
    .c(n_1299_)
  );
  inv n_2035_ (
    .din(N361),
    .dout(n_1300_)
  );
  and_bi n_2036_ (
    .a(n_0878_),
    .b(n_1300_),
    .c(n_1301_)
  );
  and_bi n_2037_ (
    .a(n_1300_),
    .b(n_0878_),
    .c(n_1302_)
  );
  inv n_2038_ (
    .din(n_1302_),
    .dout(n_1303_)
  );
  inv n_2039_ (
    .din(N358),
    .dout(n_1304_)
  );
  and_bi n_2040_ (
    .a(n_0890_),
    .b(n_1304_),
    .c(n_1305_)
  );
  and_bi n_2041_ (
    .a(n_1304_),
    .b(n_0890_),
    .c(n_1306_)
  );
  inv n_2042_ (
    .din(N355),
    .dout(n_1307_)
  );
  and_bi n_2043_ (
    .a(n_1307_),
    .b(n_0887_),
    .c(n_1308_)
  );
  and_ii n_2044_ (
    .a(n_1308_),
    .b(n_1306_),
    .c(n_1309_)
  );
  and_ii n_2045_ (
    .a(n_1309_),
    .b(n_1305_),
    .c(n_1310_)
  );
  and_bi n_2046_ (
    .a(n_1303_),
    .b(n_1310_),
    .c(n_1311_)
  );
  or_bb n_2047_ (
    .a(n_1311_),
    .b(n_1301_),
    .c(n_1312_)
  );
  inv n_2048_ (
    .din(n_1301_),
    .dout(n_1313_)
  );
  and_ii n_2049_ (
    .a(n_1306_),
    .b(n_1305_),
    .c(n_1314_)
  );
  and_bi n_2050_ (
    .a(n_0887_),
    .b(n_1307_),
    .c(n_1315_)
  );
  or_bb n_2051_ (
    .a(n_1315_),
    .b(n_1308_),
    .c(n_1316_)
  );
  and_bi n_2052_ (
    .a(n_1314_),
    .b(n_1316_),
    .c(n_1317_)
  );
  or_ii n_2053_ (
    .a(n_1317_),
    .b(n_1313_),
    .c(n_1318_)
  );
  or_ii n_2054_ (
    .a(n_1318_),
    .b(n_1312_),
    .c(n_1319_)
  );
  or_bb n_2055_ (
    .a(n_0872_),
    .b(N340),
    .c(n_1320_)
  );
  inv n_2056_ (
    .din(N343),
    .dout(n_1321_)
  );
  and_bi n_2057_ (
    .a(n_0857_),
    .b(n_1321_),
    .c(n_1322_)
  );
  and_bi n_2058_ (
    .a(n_1320_),
    .b(n_1322_),
    .c(n_1323_)
  );
  and_bb n_2059_ (
    .a(n_0872_),
    .b(N340),
    .c(n_1324_)
  );
  and_bi n_2060_ (
    .a(n_1321_),
    .b(n_0857_),
    .c(n_1325_)
  );
  and_ii n_2061_ (
    .a(n_1325_),
    .b(n_1324_),
    .c(n_1326_)
  );
  and_bb n_2062_ (
    .a(n_1326_),
    .b(n_1323_),
    .c(n_1327_)
  );
  and_bi n_2063_ (
    .a(N349),
    .b(n_0848_),
    .c(n_1328_)
  );
  and_bi n_2064_ (
    .a(n_0848_),
    .b(N349),
    .c(n_1329_)
  );
  and_ii n_2065_ (
    .a(n_1329_),
    .b(n_1328_),
    .c(n_1330_)
  );
  inv n_2066_ (
    .din(N346),
    .dout(n_1331_)
  );
  and_bi n_2067_ (
    .a(n_0860_),
    .b(n_1331_),
    .c(n_1332_)
  );
  and_bi n_2068_ (
    .a(n_1331_),
    .b(n_0860_),
    .c(n_1333_)
  );
  and_ii n_2069_ (
    .a(n_1333_),
    .b(n_1332_),
    .c(n_1334_)
  );
  or_ii n_2070_ (
    .a(n_1334_),
    .b(n_1330_),
    .c(n_1335_)
  );
  or_bi n_2071_ (
    .a(n_1335_),
    .b(n_1327_),
    .c(n_1336_)
  );
  and_ii n_2072_ (
    .a(n_0851_),
    .b(N352),
    .c(n_1337_)
  );
  and_bb n_2073_ (
    .a(n_0851_),
    .b(N352),
    .c(n_1338_)
  );
  or_bb n_2074_ (
    .a(n_1338_),
    .b(n_1337_),
    .c(n_1339_)
  );
  and_ii n_2075_ (
    .a(n_1339_),
    .b(n_1336_),
    .c(n_1340_)
  );
  inv n_2076_ (
    .din(N334),
    .dout(n_1341_)
  );
  and_bi n_2077_ (
    .a(n_0812_),
    .b(n_1341_),
    .c(n_1342_)
  );
  and_bi n_2078_ (
    .a(n_1341_),
    .b(n_0812_),
    .c(n_1343_)
  );
  inv n_2079_ (
    .din(N331),
    .dout(n_1344_)
  );
  and_bi n_2080_ (
    .a(n_0804_),
    .b(n_1344_),
    .c(n_1345_)
  );
  inv n_2081_ (
    .din(n_1345_),
    .dout(n_1346_)
  );
  and_bi n_2082_ (
    .a(n_1344_),
    .b(n_0804_),
    .c(n_1347_)
  );
  and_bb n_2083_ (
    .a(n_0827_),
    .b(N328),
    .c(n_1348_)
  );
  or_bb n_2084_ (
    .a(n_0827_),
    .b(N328),
    .c(n_1349_)
  );
  inv n_2085_ (
    .din(N325),
    .dout(n_1350_)
  );
  and_bi n_2086_ (
    .a(n_1350_),
    .b(n_0824_),
    .c(n_1351_)
  );
  and_bi n_2087_ (
    .a(n_1349_),
    .b(n_1351_),
    .c(n_1352_)
  );
  and_ii n_2088_ (
    .a(n_1352_),
    .b(n_1348_),
    .c(n_1353_)
  );
  and_ii n_2089_ (
    .a(n_1353_),
    .b(n_1347_),
    .c(n_1354_)
  );
  and_bi n_2090_ (
    .a(n_1346_),
    .b(n_1354_),
    .c(n_1355_)
  );
  and_ii n_2091_ (
    .a(n_1355_),
    .b(n_1343_),
    .c(n_1356_)
  );
  or_bb n_2092_ (
    .a(n_1356_),
    .b(n_1342_),
    .c(n_1357_)
  );
  inv n_2093_ (
    .din(n_0675_),
    .dout(n_1358_)
  );
  or_bi n_2094_ (
    .a(n_0701_),
    .b(n_0680_),
    .c(n_1359_)
  );
  and_bi n_2095_ (
    .a(n_1358_),
    .b(n_1359_),
    .c(n_1360_)
  );
  or_bb n_2096_ (
    .a(n_1360_),
    .b(n_0674_),
    .c(n_1361_)
  );
  and_bi n_2097_ (
    .a(n_0668_),
    .b(n_1361_),
    .c(n_1362_)
  );
  and_bi n_2098_ (
    .a(n_0694_),
    .b(n_0707_),
    .c(n_1363_)
  );
  and_bi n_2099_ (
    .a(n_1359_),
    .b(n_1363_),
    .c(n_1364_)
  );
  and_bi n_2100_ (
    .a(n_1358_),
    .b(n_1364_),
    .c(n_1365_)
  );
  or_bb n_2101_ (
    .a(n_1365_),
    .b(n_0674_),
    .c(n_1366_)
  );
  and_bi n_2102_ (
    .a(n_1366_),
    .b(n_1362_),
    .c(n_1367_)
  );
  and_bi n_2103_ (
    .a(n_1349_),
    .b(n_1348_),
    .c(n_1368_)
  );
  and_bi n_2104_ (
    .a(n_0824_),
    .b(n_1350_),
    .c(n_1369_)
  );
  and_ii n_2105_ (
    .a(n_1369_),
    .b(n_1351_),
    .c(n_1370_)
  );
  or_ii n_2106_ (
    .a(n_1370_),
    .b(n_1368_),
    .c(n_1371_)
  );
  and_ii n_2107_ (
    .a(n_1347_),
    .b(n_1345_),
    .c(n_0000_)
  );
  and_ii n_2108_ (
    .a(n_1343_),
    .b(n_1342_),
    .c(n_0001_)
  );
  or_ii n_2109_ (
    .a(n_0001_),
    .b(n_0000_),
    .c(n_0002_)
  );
  or_bb n_2110_ (
    .a(n_0002_),
    .b(n_1371_),
    .c(n_0003_)
  );
  and_bi n_2111_ (
    .a(n_1367_),
    .b(n_0003_),
    .c(n_0004_)
  );
  and_bi n_2112_ (
    .a(n_1357_),
    .b(n_0004_),
    .c(n_0005_)
  );
  or_bi n_2113_ (
    .a(n_0005_),
    .b(n_1340_),
    .c(n_0006_)
  );
  and_bi n_2114_ (
    .a(n_1320_),
    .b(n_1325_),
    .c(n_0007_)
  );
  or_bb n_2115_ (
    .a(n_0007_),
    .b(n_1322_),
    .c(n_0008_)
  );
  and_ii n_2116_ (
    .a(n_0008_),
    .b(n_1332_),
    .c(n_0009_)
  );
  and_ii n_2117_ (
    .a(n_0009_),
    .b(n_1333_),
    .c(n_0010_)
  );
  and_ii n_2118_ (
    .a(n_0010_),
    .b(n_1328_),
    .c(n_0011_)
  );
  and_ii n_2119_ (
    .a(n_0011_),
    .b(n_1329_),
    .c(n_0012_)
  );
  and_ii n_2120_ (
    .a(n_0012_),
    .b(n_1338_),
    .c(n_0013_)
  );
  or_bb n_2121_ (
    .a(n_0013_),
    .b(n_1337_),
    .c(n_0014_)
  );
  or_bi n_2122_ (
    .a(n_0014_),
    .b(n_0006_),
    .c(n_0015_)
  );
  and_bi n_2123_ (
    .a(n_1312_),
    .b(n_0015_),
    .c(n_0016_)
  );
  or_bi n_2124_ (
    .a(n_0016_),
    .b(n_1319_),
    .c(n_0017_)
  );
  and_ii n_2125_ (
    .a(n_0017_),
    .b(n_1299_),
    .c(n_0018_)
  );
  and_ii n_2126_ (
    .a(n_0018_),
    .b(n_1298_),
    .c(n_0019_)
  );
  and_bi n_2127_ (
    .a(n_1296_),
    .b(n_0019_),
    .c(n_0020_)
  );
  or_bi n_2128_ (
    .a(n_1296_),
    .b(n_0019_),
    .c(n_0021_)
  );
  and_bi n_2129_ (
    .a(n_0021_),
    .b(n_0020_),
    .c(N10632)
  );
  and_ii n_2130_ (
    .a(n_0769_),
    .b(n_0718_),
    .c(n_0022_)
  );
  and_bi n_2131_ (
    .a(n_0022_),
    .b(N251),
    .c(n_0023_)
  );
  and_bi n_2132_ (
    .a(N251),
    .b(n_0022_),
    .c(n_0024_)
  );
  and_ii n_2133_ (
    .a(n_0024_),
    .b(n_0023_),
    .c(n_0025_)
  );
  and_bi n_2134_ (
    .a(N303),
    .b(n_0723_),
    .c(n_0026_)
  );
  and_bi n_2135_ (
    .a(n_0723_),
    .b(N303),
    .c(n_0027_)
  );
  and_bi n_2136_ (
    .a(N299),
    .b(n_0720_),
    .c(n_0028_)
  );
  and_bi n_2137_ (
    .a(n_0720_),
    .b(N299),
    .c(n_0029_)
  );
  and_bi n_2138_ (
    .a(N296),
    .b(n_0730_),
    .c(n_0030_)
  );
  and_bi n_2139_ (
    .a(n_0730_),
    .b(N296),
    .c(n_0031_)
  );
  and_bi n_2140_ (
    .a(n_0727_),
    .b(N293),
    .c(n_0032_)
  );
  and_ii n_2141_ (
    .a(n_0032_),
    .b(n_0031_),
    .c(n_0033_)
  );
  and_ii n_2142_ (
    .a(n_0033_),
    .b(n_0030_),
    .c(n_0034_)
  );
  and_ii n_2143_ (
    .a(n_0034_),
    .b(n_0029_),
    .c(n_0035_)
  );
  or_bb n_2144_ (
    .a(n_0035_),
    .b(n_0028_),
    .c(n_0036_)
  );
  and_bi n_2145_ (
    .a(N293),
    .b(n_0727_),
    .c(n_0037_)
  );
  and_ii n_2146_ (
    .a(n_0037_),
    .b(n_0030_),
    .c(n_0038_)
  );
  and_bb n_2147_ (
    .a(n_0033_),
    .b(n_0038_),
    .c(n_0039_)
  );
  and_ii n_2148_ (
    .a(n_0029_),
    .b(n_0028_),
    .c(n_0040_)
  );
  inv n_2149_ (
    .din(n_0040_),
    .dout(n_0041_)
  );
  and_bi n_2150_ (
    .a(n_0039_),
    .b(n_0041_),
    .c(n_0042_)
  );
  and_bi n_2151_ (
    .a(n_0036_),
    .b(n_0042_),
    .c(n_0043_)
  );
  and_bi n_2152_ (
    .a(N289),
    .b(n_0752_),
    .c(n_0044_)
  );
  and_bi n_2153_ (
    .a(n_0752_),
    .b(N289),
    .c(n_0045_)
  );
  and_bi n_2154_ (
    .a(N286),
    .b(n_0750_),
    .c(n_0046_)
  );
  and_bi n_2155_ (
    .a(n_0750_),
    .b(N286),
    .c(n_0047_)
  );
  inv n_2156_ (
    .din(N283),
    .dout(n_0048_)
  );
  and_bi n_2157_ (
    .a(n_0048_),
    .b(n_0761_),
    .c(n_0049_)
  );
  inv n_2158_ (
    .din(n_0049_),
    .dout(n_0050_)
  );
  and_bi n_2159_ (
    .a(n_0761_),
    .b(n_0048_),
    .c(n_0051_)
  );
  and_ii n_2160_ (
    .a(n_0758_),
    .b(N280),
    .c(n_0052_)
  );
  and_bb n_2161_ (
    .a(n_0758_),
    .b(N280),
    .c(n_0053_)
  );
  and_bi n_2162_ (
    .a(n_1294_),
    .b(n_0053_),
    .c(n_0054_)
  );
  and_ii n_2163_ (
    .a(n_0054_),
    .b(n_0052_),
    .c(n_0055_)
  );
  and_ii n_2164_ (
    .a(n_0055_),
    .b(n_0051_),
    .c(n_0056_)
  );
  and_bi n_2165_ (
    .a(n_0050_),
    .b(n_0056_),
    .c(n_0057_)
  );
  or_bi n_2166_ (
    .a(n_0047_),
    .b(n_0057_),
    .c(n_0058_)
  );
  and_bi n_2167_ (
    .a(n_0058_),
    .b(n_0046_),
    .c(n_0059_)
  );
  and_ii n_2168_ (
    .a(n_0059_),
    .b(n_0045_),
    .c(n_0060_)
  );
  and_ii n_2169_ (
    .a(n_0053_),
    .b(n_0052_),
    .c(n_0061_)
  );
  and_bb n_2170_ (
    .a(n_0061_),
    .b(n_1296_),
    .c(n_0062_)
  );
  and_ii n_2171_ (
    .a(n_0047_),
    .b(n_0046_),
    .c(n_0063_)
  );
  and_ii n_2172_ (
    .a(n_0051_),
    .b(n_0049_),
    .c(n_0064_)
  );
  and_bb n_2173_ (
    .a(n_0064_),
    .b(n_0063_),
    .c(n_0065_)
  );
  and_bb n_2174_ (
    .a(n_0065_),
    .b(n_0062_),
    .c(n_0066_)
  );
  or_bi n_2175_ (
    .a(n_0066_),
    .b(n_0060_),
    .c(n_0067_)
  );
  and_bi n_2176_ (
    .a(n_0067_),
    .b(n_0044_),
    .c(n_0068_)
  );
  and_bb n_2177_ (
    .a(n_0060_),
    .b(n_0019_),
    .c(n_0069_)
  );
  and_bi n_2178_ (
    .a(n_0068_),
    .b(n_0069_),
    .c(n_0070_)
  );
  and_bi n_2179_ (
    .a(n_0036_),
    .b(n_0070_),
    .c(n_0071_)
  );
  and_ii n_2180_ (
    .a(n_0071_),
    .b(n_0043_),
    .c(n_0072_)
  );
  and_ii n_2181_ (
    .a(n_0072_),
    .b(n_0027_),
    .c(n_0073_)
  );
  or_bb n_2182_ (
    .a(n_0073_),
    .b(n_0026_),
    .c(n_0074_)
  );
  and_bi n_2183_ (
    .a(n_0025_),
    .b(n_0074_),
    .c(n_0075_)
  );
  and_ii n_2184_ (
    .a(n_0073_),
    .b(n_0026_),
    .c(n_0076_)
  );
  or_bb n_2185_ (
    .a(n_0076_),
    .b(n_0025_),
    .c(n_0077_)
  );
  and_bi n_2186_ (
    .a(n_0077_),
    .b(n_0075_),
    .c(N10641)
  );
  and_ii n_2187_ (
    .a(n_0045_),
    .b(n_0044_),
    .c(n_0078_)
  );
  inv n_2188_ (
    .din(n_0078_),
    .dout(n_0079_)
  );
  inv n_2189_ (
    .din(n_0063_),
    .dout(n_0080_)
  );
  inv n_2190_ (
    .din(n_0064_),
    .dout(n_0081_)
  );
  and_bi n_2191_ (
    .a(n_0062_),
    .b(n_0081_),
    .c(n_0082_)
  );
  and_bi n_2192_ (
    .a(n_0082_),
    .b(n_0019_),
    .c(n_0083_)
  );
  and_bi n_2193_ (
    .a(n_0083_),
    .b(n_0080_),
    .c(n_0084_)
  );
  and_ii n_2194_ (
    .a(n_0084_),
    .b(n_0059_),
    .c(n_0085_)
  );
  and_bi n_2195_ (
    .a(n_0085_),
    .b(n_0079_),
    .c(n_0086_)
  );
  and_bi n_2196_ (
    .a(n_0079_),
    .b(n_0085_),
    .c(n_0087_)
  );
  or_bb n_2197_ (
    .a(n_0087_),
    .b(n_0086_),
    .c(N10711)
  );
  and_bi n_2198_ (
    .a(n_0057_),
    .b(n_0083_),
    .c(n_0088_)
  );
  and_bi n_2199_ (
    .a(n_0088_),
    .b(n_0080_),
    .c(n_0089_)
  );
  and_bi n_2200_ (
    .a(n_0080_),
    .b(n_0088_),
    .c(n_0090_)
  );
  or_bb n_2201_ (
    .a(n_0090_),
    .b(n_0089_),
    .c(N10712)
  );
  and_bi n_2202_ (
    .a(n_0062_),
    .b(n_0019_),
    .c(n_0091_)
  );
  and_bi n_2203_ (
    .a(n_0055_),
    .b(n_0091_),
    .c(n_0092_)
  );
  and_bi n_2204_ (
    .a(n_0081_),
    .b(n_0092_),
    .c(n_0093_)
  );
  and_bi n_2205_ (
    .a(n_0092_),
    .b(n_0081_),
    .c(n_0094_)
  );
  or_bb n_2206_ (
    .a(n_0094_),
    .b(n_0093_),
    .c(N10713)
  );
  and_ii n_2207_ (
    .a(n_0020_),
    .b(n_1294_),
    .c(n_0095_)
  );
  or_ii n_2208_ (
    .a(n_0095_),
    .b(n_0061_),
    .c(n_0096_)
  );
  or_bb n_2209_ (
    .a(n_0095_),
    .b(n_0061_),
    .c(n_0097_)
  );
  or_ii n_2210_ (
    .a(n_0097_),
    .b(n_0096_),
    .c(N10714)
  );
  and_bi n_2211_ (
    .a(n_0772_),
    .b(N257),
    .c(n_0098_)
  );
  and_bi n_2212_ (
    .a(N257),
    .b(n_0772_),
    .c(n_0099_)
  );
  and_bi n_2213_ (
    .a(n_0785_),
    .b(N106),
    .c(n_0100_)
  );
  inv n_2214_ (
    .din(n_0100_),
    .dout(n_0101_)
  );
  and_bi n_2215_ (
    .a(N106),
    .b(n_0785_),
    .c(n_0102_)
  );
  and_bi n_2216_ (
    .a(N254),
    .b(n_0782_),
    .c(n_0103_)
  );
  and_bi n_2217_ (
    .a(n_0782_),
    .b(N254),
    .c(n_0104_)
  );
  and_ii n_2218_ (
    .a(n_0104_),
    .b(n_0023_),
    .c(n_0105_)
  );
  or_bb n_2219_ (
    .a(n_0105_),
    .b(n_0103_),
    .c(n_0106_)
  );
  and_ii n_2220_ (
    .a(n_0106_),
    .b(n_0102_),
    .c(n_0107_)
  );
  and_bi n_2221_ (
    .a(n_0101_),
    .b(n_0107_),
    .c(n_0108_)
  );
  and_ii n_2222_ (
    .a(n_0108_),
    .b(n_0099_),
    .c(n_0109_)
  );
  and_ii n_2223_ (
    .a(n_0109_),
    .b(n_0098_),
    .c(n_0110_)
  );
  and_ii n_2224_ (
    .a(n_0102_),
    .b(n_0100_),
    .c(n_0111_)
  );
  and_ii n_2225_ (
    .a(n_0103_),
    .b(n_0104_),
    .c(n_0112_)
  );
  or_ii n_2226_ (
    .a(n_0112_),
    .b(n_0025_),
    .c(n_0113_)
  );
  and_bi n_2227_ (
    .a(n_0111_),
    .b(n_0113_),
    .c(n_0114_)
  );
  and_bi n_2228_ (
    .a(n_0114_),
    .b(n_0074_),
    .c(n_0115_)
  );
  and_ii n_2229_ (
    .a(n_0099_),
    .b(n_0098_),
    .c(n_0116_)
  );
  or_ii n_2230_ (
    .a(n_0116_),
    .b(n_0115_),
    .c(n_0117_)
  );
  or_ii n_2231_ (
    .a(n_0117_),
    .b(n_0110_),
    .c(n_0118_)
  );
  and_bi n_2232_ (
    .a(n_0775_),
    .b(N260),
    .c(n_0119_)
  );
  and_bi n_2233_ (
    .a(N260),
    .b(n_0775_),
    .c(n_0120_)
  );
  and_ii n_2234_ (
    .a(n_0120_),
    .b(n_0119_),
    .c(n_0121_)
  );
  and_bi n_2235_ (
    .a(n_0121_),
    .b(n_0118_),
    .c(n_0122_)
  );
  and_bi n_2236_ (
    .a(n_0118_),
    .b(n_0121_),
    .c(n_0123_)
  );
  or_bb n_2237_ (
    .a(n_0123_),
    .b(n_0122_),
    .c(N10715)
  );
  or_bi n_2238_ (
    .a(n_0115_),
    .b(n_0108_),
    .c(n_0124_)
  );
  and_bi n_2239_ (
    .a(n_0124_),
    .b(n_0116_),
    .c(n_0125_)
  );
  and_bi n_2240_ (
    .a(n_0116_),
    .b(n_0124_),
    .c(n_0126_)
  );
  or_bb n_2241_ (
    .a(n_0126_),
    .b(n_0125_),
    .c(N10716)
  );
  and_bi n_2242_ (
    .a(n_0076_),
    .b(n_0113_),
    .c(n_0127_)
  );
  or_bi n_2243_ (
    .a(n_0127_),
    .b(n_0106_),
    .c(n_0128_)
  );
  and_bi n_2244_ (
    .a(n_0128_),
    .b(n_0111_),
    .c(n_0129_)
  );
  and_bi n_2245_ (
    .a(n_0111_),
    .b(n_0128_),
    .c(n_0130_)
  );
  or_bb n_2246_ (
    .a(n_0130_),
    .b(n_0129_),
    .c(N10717)
  );
  and_ii n_2247_ (
    .a(n_0075_),
    .b(n_0023_),
    .c(n_0131_)
  );
  and_bi n_2248_ (
    .a(n_0131_),
    .b(n_0112_),
    .c(n_0132_)
  );
  and_bi n_2249_ (
    .a(n_0112_),
    .b(n_0131_),
    .c(n_0133_)
  );
  and_ii n_2250_ (
    .a(n_0133_),
    .b(n_0132_),
    .c(N10718)
  );
  or_bb n_2251_ (
    .a(N883),
    .b(N882),
    .c(n_0134_)
  );
  or_bb n_2252_ (
    .a(N885),
    .b(N884),
    .c(n_0135_)
  );
  or_bb n_2253_ (
    .a(n_0135_),
    .b(n_0134_),
    .c(n_0136_)
  );
  or_bb n_2254_ (
    .a(n_0136_),
    .b(N10574),
    .c(n_0137_)
  );
  or_bb n_2255_ (
    .a(N10576),
    .b(N10575),
    .c(n_0138_)
  );
  or_bb n_2256_ (
    .a(n_0138_),
    .b(n_0137_),
    .c(N10729)
  );
  and_bi n_2257_ (
    .a(n_1320_),
    .b(n_1324_),
    .c(n_0139_)
  );
  and_bi n_2258_ (
    .a(n_0139_),
    .b(n_0005_),
    .c(n_0140_)
  );
  and_bi n_2259_ (
    .a(n_0005_),
    .b(n_0139_),
    .c(n_0141_)
  );
  and_ii n_2260_ (
    .a(n_0141_),
    .b(n_0140_),
    .c(N10827)
  );
  or_bb n_2261_ (
    .a(n_0005_),
    .b(n_1336_),
    .c(n_0142_)
  );
  and_ii n_2262_ (
    .a(n_0012_),
    .b(n_1339_),
    .c(n_0143_)
  );
  and_bb n_2263_ (
    .a(n_0012_),
    .b(n_1339_),
    .c(n_0144_)
  );
  and_ii n_2264_ (
    .a(n_0144_),
    .b(n_0143_),
    .c(n_0145_)
  );
  and_bi n_2265_ (
    .a(n_0142_),
    .b(n_0145_),
    .c(n_0146_)
  );
  and_bi n_2266_ (
    .a(n_0006_),
    .b(n_0146_),
    .c(N10868)
  );
  and_bb n_2267_ (
    .a(n_1334_),
    .b(n_1327_),
    .c(n_0147_)
  );
  and_bi n_2268_ (
    .a(n_0147_),
    .b(n_0005_),
    .c(n_0148_)
  );
  and_bi n_2269_ (
    .a(n_0010_),
    .b(n_0148_),
    .c(n_0149_)
  );
  or_ii n_2270_ (
    .a(n_0149_),
    .b(n_1330_),
    .c(n_0150_)
  );
  or_bb n_2271_ (
    .a(n_0149_),
    .b(n_1330_),
    .c(n_0151_)
  );
  or_ii n_2272_ (
    .a(n_0151_),
    .b(n_0150_),
    .c(N10869)
  );
  and_ii n_2273_ (
    .a(n_1325_),
    .b(n_1322_),
    .c(n_0152_)
  );
  inv n_2274_ (
    .din(n_0152_),
    .dout(n_0153_)
  );
  and_bi n_2275_ (
    .a(n_0140_),
    .b(n_0153_),
    .c(n_0154_)
  );
  or_bi n_2276_ (
    .a(n_0154_),
    .b(n_0008_),
    .c(n_0155_)
  );
  and_bi n_2277_ (
    .a(n_0155_),
    .b(n_1334_),
    .c(n_0156_)
  );
  and_bi n_2278_ (
    .a(n_1334_),
    .b(n_0155_),
    .c(n_0157_)
  );
  or_bb n_2279_ (
    .a(n_0157_),
    .b(n_0156_),
    .c(N10870)
  );
  and_bi n_2280_ (
    .a(n_1320_),
    .b(n_0140_),
    .c(n_0158_)
  );
  and_bi n_2281_ (
    .a(n_0158_),
    .b(n_0153_),
    .c(n_0159_)
  );
  and_bi n_2282_ (
    .a(n_0153_),
    .b(n_0158_),
    .c(n_0160_)
  );
  or_bb n_2283_ (
    .a(n_0160_),
    .b(n_0159_),
    .c(N10871)
  );
  and_bb n_2284_ (
    .a(N1),
    .b(N163),
    .c(N1781)
  );
  inv n_2285_ (
    .din(N38),
    .dout(n_0161_)
  );
  and_bb n_2286_ (
    .a(N382),
    .b(N267),
    .c(n_0162_)
  );
  or_ii n_2287_ (
    .a(n_0162_),
    .b(n_0161_),
    .c(n_0163_)
  );
  and_bb n_2288_ (
    .a(n_0162_),
    .b(N263),
    .c(n_0164_)
  );
  and_bi n_2289_ (
    .a(N38),
    .b(n_0164_),
    .c(n_0165_)
  );
  and_bb n_2290_ (
    .a(N382),
    .b(N263),
    .c(n_0166_)
  );
  and_bi n_2291_ (
    .a(n_0166_),
    .b(n_0161_),
    .c(n_0167_)
  );
  and_bi n_2292_ (
    .a(n_0161_),
    .b(n_0166_),
    .c(n_0168_)
  );
  and_ii n_2293_ (
    .a(n_0168_),
    .b(n_0167_),
    .c(n_0169_)
  );
  and_bi n_2294_ (
    .a(n_0098_),
    .b(n_0120_),
    .c(n_0170_)
  );
  and_ii n_2295_ (
    .a(n_0170_),
    .b(n_0119_),
    .c(n_0171_)
  );
  or_ii n_2296_ (
    .a(n_0121_),
    .b(n_0116_),
    .c(n_0172_)
  );
  and_ii n_2297_ (
    .a(n_0172_),
    .b(n_0108_),
    .c(n_0173_)
  );
  and_bi n_2298_ (
    .a(n_0171_),
    .b(n_0173_),
    .c(n_0174_)
  );
  and_bi n_2299_ (
    .a(n_0115_),
    .b(n_0172_),
    .c(n_0175_)
  );
  and_bi n_2300_ (
    .a(n_0174_),
    .b(n_0175_),
    .c(n_0176_)
  );
  or_bb n_2301_ (
    .a(n_0176_),
    .b(n_0169_),
    .c(n_0177_)
  );
  and_bi n_2302_ (
    .a(n_0177_),
    .b(n_0165_),
    .c(n_0178_)
  );
  and_bi n_2303_ (
    .a(n_0163_),
    .b(n_0178_),
    .c(N10101)
  );
  or_bi n_2304_ (
    .a(N38),
    .b(N382),
    .c(n_0179_)
  );
  or_bb n_2305_ (
    .a(n_0179_),
    .b(n_0939_),
    .c(n_0180_)
  );
  and_bb n_2306_ (
    .a(n_1280_),
    .b(n_0993_),
    .c(n_0181_)
  );
  or_bb n_2307_ (
    .a(n_1262_),
    .b(n_0990_),
    .c(n_0182_)
  );
  and_ii n_2308_ (
    .a(n_1253_),
    .b(n_0963_),
    .c(n_0183_)
  );
  or_bb n_2309_ (
    .a(N89),
    .b(N70),
    .c(n_0184_)
  );
  and_bi n_2310_ (
    .a(n_0184_),
    .b(n_0662_),
    .c(n_0185_)
  );
  and_bi n_2311_ (
    .a(N89),
    .b(n_0950_),
    .c(n_0186_)
  );
  or_bb n_2312_ (
    .a(n_0186_),
    .b(n_0185_),
    .c(n_0187_)
  );
  or_bb n_2313_ (
    .a(n_0187_),
    .b(n_0183_),
    .c(n_0188_)
  );
  and_bb n_2314_ (
    .a(n_1255_),
    .b(n_0960_),
    .c(n_0189_)
  );
  and_bb n_2315_ (
    .a(n_1253_),
    .b(n_0963_),
    .c(n_0190_)
  );
  or_bb n_2316_ (
    .a(n_0190_),
    .b(n_0189_),
    .c(n_0191_)
  );
  and_bi n_2317_ (
    .a(n_0188_),
    .b(n_0191_),
    .c(n_0192_)
  );
  and_ii n_2318_ (
    .a(n_1255_),
    .b(n_0960_),
    .c(n_0193_)
  );
  and_ii n_2319_ (
    .a(n_1260_),
    .b(n_0987_),
    .c(n_0194_)
  );
  or_bb n_2320_ (
    .a(n_0194_),
    .b(n_0193_),
    .c(n_0195_)
  );
  or_bb n_2321_ (
    .a(n_0195_),
    .b(n_0192_),
    .c(n_0196_)
  );
  and_bb n_2322_ (
    .a(n_1262_),
    .b(n_0990_),
    .c(n_0197_)
  );
  and_bb n_2323_ (
    .a(n_1260_),
    .b(n_0987_),
    .c(n_0198_)
  );
  or_bb n_2324_ (
    .a(n_0198_),
    .b(n_0197_),
    .c(n_0199_)
  );
  and_bi n_2325_ (
    .a(n_0196_),
    .b(n_0199_),
    .c(n_0200_)
  );
  and_bi n_2326_ (
    .a(n_0182_),
    .b(n_0200_),
    .c(n_0201_)
  );
  and_ii n_2327_ (
    .a(n_0201_),
    .b(n_0181_),
    .c(n_0202_)
  );
  and_ii n_2328_ (
    .a(n_1282_),
    .b(n_0981_),
    .c(n_0203_)
  );
  and_ii n_2329_ (
    .a(n_1280_),
    .b(n_0993_),
    .c(n_0204_)
  );
  or_bb n_2330_ (
    .a(n_0204_),
    .b(n_0203_),
    .c(n_0205_)
  );
  and_ii n_2331_ (
    .a(n_0205_),
    .b(n_0202_),
    .c(n_0206_)
  );
  and_bb n_2332_ (
    .a(n_1275_),
    .b(n_0975_),
    .c(n_0207_)
  );
  and_ii n_2333_ (
    .a(n_1273_),
    .b(n_0972_),
    .c(n_0208_)
  );
  or_bb n_2334_ (
    .a(n_0208_),
    .b(n_0207_),
    .c(n_0209_)
  );
  and_bb n_2335_ (
    .a(n_1282_),
    .b(n_0981_),
    .c(n_0210_)
  );
  and_bb n_2336_ (
    .a(n_1273_),
    .b(n_0972_),
    .c(n_0211_)
  );
  or_bb n_2337_ (
    .a(n_0211_),
    .b(n_0210_),
    .c(n_0212_)
  );
  or_bb n_2338_ (
    .a(n_0212_),
    .b(n_0209_),
    .c(n_0213_)
  );
  and_ii n_2339_ (
    .a(n_0213_),
    .b(n_0206_),
    .c(n_0214_)
  );
  and_bi n_2340_ (
    .a(n_0208_),
    .b(n_0207_),
    .c(n_0215_)
  );
  and_ii n_2341_ (
    .a(n_1275_),
    .b(n_0975_),
    .c(n_0216_)
  );
  and_ii n_2342_ (
    .a(n_1187_),
    .b(n_1054_),
    .c(n_0217_)
  );
  or_bb n_2343_ (
    .a(n_0217_),
    .b(n_0216_),
    .c(n_0218_)
  );
  or_bb n_2344_ (
    .a(n_0218_),
    .b(n_0215_),
    .c(n_0219_)
  );
  and_ii n_2345_ (
    .a(n_0219_),
    .b(n_0214_),
    .c(n_0220_)
  );
  and_ii n_2346_ (
    .a(n_1178_),
    .b(n_1009_),
    .c(n_0221_)
  );
  and_ii n_2347_ (
    .a(n_1180_),
    .b(n_1012_),
    .c(n_0222_)
  );
  or_bb n_2348_ (
    .a(n_0222_),
    .b(n_0221_),
    .c(n_0223_)
  );
  and_bb n_2349_ (
    .a(n_1153_),
    .b(n_1033_),
    .c(n_0224_)
  );
  and_bb n_2350_ (
    .a(n_1178_),
    .b(n_1009_),
    .c(n_0225_)
  );
  and_bb n_2351_ (
    .a(n_1180_),
    .b(n_1012_),
    .c(n_0226_)
  );
  or_bb n_2352_ (
    .a(n_0226_),
    .b(n_0225_),
    .c(n_0227_)
  );
  or_bb n_2353_ (
    .a(n_0227_),
    .b(n_0224_),
    .c(n_0228_)
  );
  and_ii n_2354_ (
    .a(n_0228_),
    .b(n_0223_),
    .c(n_0229_)
  );
  and_ii n_2355_ (
    .a(n_1151_),
    .b(n_1030_),
    .c(n_0230_)
  );
  and_ii n_2356_ (
    .a(n_1153_),
    .b(n_1033_),
    .c(n_0231_)
  );
  and_ii n_2357_ (
    .a(n_0231_),
    .b(n_0230_),
    .c(n_0232_)
  );
  and_bb n_2358_ (
    .a(n_1187_),
    .b(n_1054_),
    .c(n_0233_)
  );
  and_bb n_2359_ (
    .a(n_1151_),
    .b(n_1030_),
    .c(n_0234_)
  );
  and_ii n_2360_ (
    .a(n_0234_),
    .b(n_0233_),
    .c(n_0235_)
  );
  and_bb n_2361_ (
    .a(n_0235_),
    .b(n_0232_),
    .c(n_0236_)
  );
  or_ii n_2362_ (
    .a(n_0236_),
    .b(n_0229_),
    .c(n_0237_)
  );
  and_ii n_2363_ (
    .a(n_0237_),
    .b(n_0220_),
    .c(n_0238_)
  );
  and_bi n_2364_ (
    .a(n_0229_),
    .b(n_0232_),
    .c(n_0239_)
  );
  and_bi n_2365_ (
    .a(n_0223_),
    .b(n_0226_),
    .c(n_0240_)
  );
  or_bb n_2366_ (
    .a(n_0240_),
    .b(n_0239_),
    .c(n_0241_)
  );
  and_ii n_2367_ (
    .a(n_0241_),
    .b(n_0238_),
    .c(n_0242_)
  );
  and_bb n_2368_ (
    .a(n_1160_),
    .b(n_1021_),
    .c(n_0243_)
  );
  and_ii n_2369_ (
    .a(n_1158_),
    .b(n_1018_),
    .c(n_0244_)
  );
  and_ii n_2370_ (
    .a(n_0244_),
    .b(n_0243_),
    .c(n_0245_)
  );
  and_ii n_2371_ (
    .a(n_1160_),
    .b(n_1021_),
    .c(n_0246_)
  );
  and_bb n_2372_ (
    .a(n_1158_),
    .b(n_1018_),
    .c(n_0247_)
  );
  or_bb n_2373_ (
    .a(n_0247_),
    .b(n_0246_),
    .c(n_0248_)
  );
  and_bi n_2374_ (
    .a(n_0245_),
    .b(n_0248_),
    .c(n_0249_)
  );
  and_ii n_2375_ (
    .a(n_1167_),
    .b(n_1045_),
    .c(n_0250_)
  );
  and_ii n_2376_ (
    .a(n_1165_),
    .b(n_1042_),
    .c(n_0251_)
  );
  and_ii n_2377_ (
    .a(n_0251_),
    .b(n_0250_),
    .c(n_0252_)
  );
  and_bb n_2378_ (
    .a(n_1167_),
    .b(n_1045_),
    .c(n_0253_)
  );
  and_bb n_2379_ (
    .a(n_1165_),
    .b(n_1042_),
    .c(n_0254_)
  );
  and_ii n_2380_ (
    .a(n_0254_),
    .b(n_0253_),
    .c(n_0255_)
  );
  and_bb n_2381_ (
    .a(n_0255_),
    .b(n_0252_),
    .c(n_0256_)
  );
  or_ii n_2382_ (
    .a(n_0256_),
    .b(n_0249_),
    .c(n_0257_)
  );
  and_ii n_2383_ (
    .a(n_0257_),
    .b(n_0242_),
    .c(n_0258_)
  );
  or_bb n_2384_ (
    .a(n_0253_),
    .b(n_0252_),
    .c(n_0259_)
  );
  and_bi n_2385_ (
    .a(n_0249_),
    .b(n_0259_),
    .c(n_0260_)
  );
  and_bi n_2386_ (
    .a(n_0244_),
    .b(n_0243_),
    .c(n_0261_)
  );
  or_bb n_2387_ (
    .a(n_0261_),
    .b(n_0246_),
    .c(n_0262_)
  );
  or_bb n_2388_ (
    .a(n_0262_),
    .b(n_0260_),
    .c(n_0263_)
  );
  and_ii n_2389_ (
    .a(n_0263_),
    .b(n_0258_),
    .c(n_0264_)
  );
  and_bi n_2390_ (
    .a(n_1228_),
    .b(n_1069_),
    .c(n_0265_)
  );
  and_ii n_2391_ (
    .a(n_1226_),
    .b(n_1066_),
    .c(n_0266_)
  );
  or_bb n_2392_ (
    .a(n_0266_),
    .b(n_0265_),
    .c(n_0267_)
  );
  and_bi n_2393_ (
    .a(n_1069_),
    .b(n_1228_),
    .c(n_0268_)
  );
  and_bb n_2394_ (
    .a(n_1226_),
    .b(n_1066_),
    .c(n_0269_)
  );
  or_bb n_2395_ (
    .a(n_0269_),
    .b(n_0268_),
    .c(n_0270_)
  );
  and_ii n_2396_ (
    .a(n_0270_),
    .b(n_0267_),
    .c(n_0271_)
  );
  and_ii n_2397_ (
    .a(n_1235_),
    .b(n_1096_),
    .c(n_0272_)
  );
  and_ii n_2398_ (
    .a(n_1233_),
    .b(n_1111_),
    .c(n_0273_)
  );
  and_ii n_2399_ (
    .a(n_0273_),
    .b(n_0272_),
    .c(n_0274_)
  );
  and_bb n_2400_ (
    .a(n_1235_),
    .b(n_1096_),
    .c(n_0275_)
  );
  and_bb n_2401_ (
    .a(n_1233_),
    .b(n_1111_),
    .c(n_0276_)
  );
  and_ii n_2402_ (
    .a(n_0276_),
    .b(n_0275_),
    .c(n_0277_)
  );
  or_ii n_2403_ (
    .a(n_0277_),
    .b(n_0274_),
    .c(n_0278_)
  );
  and_bi n_2404_ (
    .a(n_0271_),
    .b(n_0278_),
    .c(n_0279_)
  );
  and_ii n_2405_ (
    .a(n_1201_),
    .b(n_1090_),
    .c(n_0280_)
  );
  and_bb n_2406_ (
    .a(n_1201_),
    .b(n_1090_),
    .c(n_0281_)
  );
  and_ii n_2407_ (
    .a(n_0281_),
    .b(n_0280_),
    .c(n_0282_)
  );
  or_ii n_2408_ (
    .a(n_0282_),
    .b(n_0279_),
    .c(n_0283_)
  );
  or_bb n_2409_ (
    .a(n_0283_),
    .b(n_0264_),
    .c(n_0284_)
  );
  and_bb n_2410_ (
    .a(n_0280_),
    .b(n_0279_),
    .c(n_0285_)
  );
  or_bb n_2411_ (
    .a(n_0275_),
    .b(n_0274_),
    .c(n_0286_)
  );
  and_bi n_2412_ (
    .a(n_0271_),
    .b(n_0286_),
    .c(n_0287_)
  );
  and_bi n_2413_ (
    .a(n_0267_),
    .b(n_0268_),
    .c(n_0288_)
  );
  or_bb n_2414_ (
    .a(n_0288_),
    .b(n_0287_),
    .c(n_0289_)
  );
  or_bb n_2415_ (
    .a(n_0289_),
    .b(n_0285_),
    .c(n_0290_)
  );
  and_bi n_2416_ (
    .a(n_0284_),
    .b(n_0290_),
    .c(n_0291_)
  );
  and_bi n_2417_ (
    .a(n_1206_),
    .b(n_1075_),
    .c(n_0292_)
  );
  and_bi n_2418_ (
    .a(n_1209_),
    .b(n_1078_),
    .c(n_0293_)
  );
  or_bb n_2419_ (
    .a(n_0293_),
    .b(n_0292_),
    .c(n_0294_)
  );
  and_bi n_2420_ (
    .a(n_1075_),
    .b(n_1206_),
    .c(n_0295_)
  );
  and_bi n_2421_ (
    .a(n_1078_),
    .b(n_1209_),
    .c(n_0296_)
  );
  and_ii n_2422_ (
    .a(n_0296_),
    .b(n_0295_),
    .c(n_0297_)
  );
  and_bi n_2423_ (
    .a(n_0297_),
    .b(n_0294_),
    .c(n_0298_)
  );
  and_bi n_2424_ (
    .a(n_1216_),
    .b(n_1105_),
    .c(n_0299_)
  );
  and_bi n_2425_ (
    .a(n_1213_),
    .b(n_1102_),
    .c(n_0300_)
  );
  and_ii n_2426_ (
    .a(n_0300_),
    .b(n_0299_),
    .c(n_0301_)
  );
  and_bi n_2427_ (
    .a(n_1105_),
    .b(n_1216_),
    .c(n_0302_)
  );
  and_bi n_2428_ (
    .a(n_1102_),
    .b(n_1213_),
    .c(n_0303_)
  );
  and_ii n_2429_ (
    .a(n_0303_),
    .b(n_0302_),
    .c(n_0304_)
  );
  and_bb n_2430_ (
    .a(n_0304_),
    .b(n_0301_),
    .c(n_0305_)
  );
  or_ii n_2431_ (
    .a(n_0305_),
    .b(n_0298_),
    .c(n_0306_)
  );
  or_bb n_2432_ (
    .a(n_0306_),
    .b(n_0291_),
    .c(n_0307_)
  );
  or_bb n_2433_ (
    .a(n_0302_),
    .b(n_0301_),
    .c(n_0308_)
  );
  and_bi n_2434_ (
    .a(n_0298_),
    .b(n_0308_),
    .c(n_0309_)
  );
  and_bi n_2435_ (
    .a(n_0294_),
    .b(n_0296_),
    .c(n_0310_)
  );
  or_bb n_2436_ (
    .a(n_0310_),
    .b(n_0309_),
    .c(n_0311_)
  );
  and_bi n_2437_ (
    .a(n_0307_),
    .b(n_0311_),
    .c(n_0312_)
  );
  and_bi n_2438_ (
    .a(n_0930_),
    .b(n_1137_),
    .c(n_0313_)
  );
  and_bb n_2439_ (
    .a(n_1127_),
    .b(n_0918_),
    .c(n_0314_)
  );
  and_ii n_2440_ (
    .a(n_1127_),
    .b(n_0918_),
    .c(n_0315_)
  );
  or_bb n_2441_ (
    .a(n_0315_),
    .b(n_0314_),
    .c(n_0316_)
  );
  and_bi n_2442_ (
    .a(n_1124_),
    .b(n_0915_),
    .c(n_0317_)
  );
  and_bi n_2443_ (
    .a(n_0915_),
    .b(n_1124_),
    .c(n_0318_)
  );
  or_bb n_2444_ (
    .a(n_0318_),
    .b(n_0317_),
    .c(n_0319_)
  );
  or_bb n_2445_ (
    .a(n_0319_),
    .b(n_0316_),
    .c(n_0320_)
  );
  and_ii n_2446_ (
    .a(n_0320_),
    .b(n_0313_),
    .c(n_0321_)
  );
  and_ii n_2447_ (
    .a(n_0909_),
    .b(n_0718_),
    .c(n_0322_)
  );
  and_bi n_2448_ (
    .a(n_1134_),
    .b(n_0927_),
    .c(n_0323_)
  );
  or_bb n_2449_ (
    .a(n_0323_),
    .b(n_0322_),
    .c(n_0324_)
  );
  and_bb n_2450_ (
    .a(n_0909_),
    .b(n_0718_),
    .c(n_0325_)
  );
  and_bi n_2451_ (
    .a(n_1137_),
    .b(n_0930_),
    .c(n_0326_)
  );
  and_bi n_2452_ (
    .a(n_0927_),
    .b(n_1134_),
    .c(n_0327_)
  );
  or_bb n_2453_ (
    .a(n_0327_),
    .b(n_0326_),
    .c(n_0328_)
  );
  or_bb n_2454_ (
    .a(n_0328_),
    .b(n_0325_),
    .c(n_0329_)
  );
  and_ii n_2455_ (
    .a(n_0329_),
    .b(n_0324_),
    .c(n_0330_)
  );
  or_ii n_2456_ (
    .a(n_0330_),
    .b(n_0321_),
    .c(n_0331_)
  );
  or_bb n_2457_ (
    .a(n_0331_),
    .b(n_0312_),
    .c(n_0332_)
  );
  or_bi n_2458_ (
    .a(n_0327_),
    .b(n_0324_),
    .c(n_0333_)
  );
  and_bi n_2459_ (
    .a(n_0333_),
    .b(n_0326_),
    .c(n_0334_)
  );
  and_bi n_2460_ (
    .a(n_0321_),
    .b(n_0334_),
    .c(n_0335_)
  );
  and_bi n_2461_ (
    .a(N382),
    .b(n_0938_),
    .c(n_0336_)
  );
  and_bi n_2462_ (
    .a(N38),
    .b(n_0336_),
    .c(n_0337_)
  );
  or_bb n_2463_ (
    .a(n_0317_),
    .b(n_0315_),
    .c(n_0338_)
  );
  and_bi n_2464_ (
    .a(n_0338_),
    .b(n_0314_),
    .c(n_0339_)
  );
  or_bb n_2465_ (
    .a(n_0339_),
    .b(n_0337_),
    .c(n_0340_)
  );
  or_bb n_2466_ (
    .a(n_0340_),
    .b(n_0335_),
    .c(n_0341_)
  );
  and_bi n_2467_ (
    .a(n_0332_),
    .b(n_0341_),
    .c(n_0342_)
  );
  and_bi n_2468_ (
    .a(n_0180_),
    .b(n_0342_),
    .c(N10102)
  );
  inv n_2469_ (
    .din(n_0000_),
    .dout(n_0343_)
  );
  or_bb n_2470_ (
    .a(n_0343_),
    .b(n_1371_),
    .c(n_0344_)
  );
  or_bi n_2471_ (
    .a(n_0344_),
    .b(n_1367_),
    .c(n_0345_)
  );
  and_bi n_2472_ (
    .a(n_0345_),
    .b(n_1355_),
    .c(n_0346_)
  );
  or_ii n_2473_ (
    .a(n_0346_),
    .b(n_0001_),
    .c(n_0347_)
  );
  or_bb n_2474_ (
    .a(n_0346_),
    .b(n_0001_),
    .c(n_0348_)
  );
  or_ii n_2475_ (
    .a(n_0348_),
    .b(n_0347_),
    .c(N10350)
  );
  and_bi n_2476_ (
    .a(n_1367_),
    .b(n_1369_),
    .c(n_0349_)
  );
  or_ii n_2477_ (
    .a(n_0349_),
    .b(n_1368_),
    .c(n_0350_)
  );
  and_bi n_2478_ (
    .a(n_0350_),
    .b(n_1353_),
    .c(n_0351_)
  );
  and_bi n_2479_ (
    .a(n_0351_),
    .b(n_0343_),
    .c(n_0352_)
  );
  and_bi n_2480_ (
    .a(n_0343_),
    .b(n_0351_),
    .c(n_0353_)
  );
  or_bb n_2481_ (
    .a(n_0353_),
    .b(n_0352_),
    .c(N10351)
  );
  inv n_2482_ (
    .din(n_1368_),
    .dout(n_0354_)
  );
  and_ii n_2483_ (
    .a(n_0349_),
    .b(n_1351_),
    .c(n_0355_)
  );
  and_bi n_2484_ (
    .a(n_0355_),
    .b(n_0354_),
    .c(n_0356_)
  );
  and_bi n_2485_ (
    .a(n_0354_),
    .b(n_0355_),
    .c(n_0357_)
  );
  or_bb n_2486_ (
    .a(n_0357_),
    .b(n_0356_),
    .c(N10352)
  );
  and_bi n_2487_ (
    .a(n_1367_),
    .b(n_1370_),
    .c(n_0358_)
  );
  and_bi n_2488_ (
    .a(n_1370_),
    .b(n_1367_),
    .c(n_0359_)
  );
  or_bb n_2489_ (
    .a(n_0359_),
    .b(n_0358_),
    .c(N10353)
  );
  inv n_2490_ (
    .din(n_0264_),
    .dout(N10704)
  );
  and_ii n_2491_ (
    .a(n_0027_),
    .b(n_0026_),
    .c(n_0360_)
  );
  and_bi n_2492_ (
    .a(n_0072_),
    .b(n_0360_),
    .c(n_0361_)
  );
  and_bi n_2493_ (
    .a(n_0360_),
    .b(n_0072_),
    .c(n_0362_)
  );
  or_bb n_2494_ (
    .a(n_0362_),
    .b(n_0361_),
    .c(N10760)
  );
  and_bb n_2495_ (
    .a(n_0070_),
    .b(n_0039_),
    .c(n_0363_)
  );
  and_ii n_2496_ (
    .a(n_0363_),
    .b(n_0034_),
    .c(n_0364_)
  );
  and_bi n_2497_ (
    .a(n_0364_),
    .b(n_0041_),
    .c(n_0365_)
  );
  and_bi n_2498_ (
    .a(n_0041_),
    .b(n_0364_),
    .c(n_0366_)
  );
  or_bb n_2499_ (
    .a(n_0366_),
    .b(n_0365_),
    .c(N10761)
  );
  and_ii n_2500_ (
    .a(n_0031_),
    .b(n_0030_),
    .c(n_0367_)
  );
  and_bi n_2501_ (
    .a(n_0070_),
    .b(n_0037_),
    .c(n_0368_)
  );
  or_bb n_2502_ (
    .a(n_0368_),
    .b(n_0032_),
    .c(n_0369_)
  );
  or_ii n_2503_ (
    .a(n_0369_),
    .b(n_0367_),
    .c(n_0370_)
  );
  and_ii n_2504_ (
    .a(n_0369_),
    .b(n_0367_),
    .c(n_0371_)
  );
  and_bi n_2505_ (
    .a(n_0370_),
    .b(n_0371_),
    .c(N10762)
  );
  and_ii n_2506_ (
    .a(n_0032_),
    .b(n_0037_),
    .c(n_0372_)
  );
  or_ii n_2507_ (
    .a(n_0070_),
    .b(n_0372_),
    .c(n_0373_)
  );
  and_ii n_2508_ (
    .a(n_0070_),
    .b(n_0372_),
    .c(n_0374_)
  );
  and_bi n_2509_ (
    .a(n_0373_),
    .b(n_0374_),
    .c(N10763)
  );
  or_ii n_2510_ (
    .a(n_0176_),
    .b(n_0167_),
    .c(n_0375_)
  );
  and_bi n_2511_ (
    .a(n_0168_),
    .b(n_0176_),
    .c(n_0376_)
  );
  and_bi n_2512_ (
    .a(n_0375_),
    .b(n_0376_),
    .c(n_0377_)
  );
  or_ii n_2513_ (
    .a(n_0377_),
    .b(n_0162_),
    .c(n_0378_)
  );
  inv n_2514_ (
    .din(n_0162_),
    .dout(n_0379_)
  );
  and_bi n_2515_ (
    .a(n_0379_),
    .b(n_0377_),
    .c(n_0380_)
  );
  and_bi n_2516_ (
    .a(n_0378_),
    .b(n_0380_),
    .c(N10837)
  );
  and_bb n_2517_ (
    .a(n_0176_),
    .b(n_0169_),
    .c(n_0381_)
  );
  and_bi n_2518_ (
    .a(n_0177_),
    .b(n_0381_),
    .c(N10839)
  );
  and_ii n_2519_ (
    .a(n_1298_),
    .b(n_1299_),
    .c(n_0382_)
  );
  or_bi n_2520_ (
    .a(n_0382_),
    .b(n_0017_),
    .c(n_0383_)
  );
  and_bi n_2521_ (
    .a(n_0382_),
    .b(n_0017_),
    .c(n_0384_)
  );
  and_bi n_2522_ (
    .a(n_0383_),
    .b(n_0384_),
    .c(N10905)
  );
  and_ii n_2523_ (
    .a(n_1301_),
    .b(n_1302_),
    .c(n_0385_)
  );
  and_bb n_2524_ (
    .a(n_0015_),
    .b(n_1317_),
    .c(n_0386_)
  );
  and_ii n_2525_ (
    .a(n_0386_),
    .b(n_1310_),
    .c(n_0387_)
  );
  or_ii n_2526_ (
    .a(n_0387_),
    .b(n_0385_),
    .c(n_0388_)
  );
  or_bb n_2527_ (
    .a(n_0387_),
    .b(n_0385_),
    .c(n_0389_)
  );
  or_ii n_2528_ (
    .a(n_0389_),
    .b(n_0388_),
    .c(N10906)
  );
  inv n_2529_ (
    .din(n_1314_),
    .dout(n_0390_)
  );
  and_ii n_2530_ (
    .a(n_0015_),
    .b(n_1308_),
    .c(n_0391_)
  );
  or_bb n_2531_ (
    .a(n_0391_),
    .b(n_1315_),
    .c(n_0392_)
  );
  or_ii n_2532_ (
    .a(n_0392_),
    .b(n_0390_),
    .c(n_0393_)
  );
  and_bi n_2533_ (
    .a(n_1314_),
    .b(n_0392_),
    .c(n_0394_)
  );
  and_bi n_2534_ (
    .a(n_0393_),
    .b(n_0394_),
    .c(N10907)
  );
  or_bi n_2535_ (
    .a(n_1316_),
    .b(n_0015_),
    .c(n_0395_)
  );
  and_bi n_2536_ (
    .a(n_1316_),
    .b(n_0015_),
    .c(n_0396_)
  );
  and_bi n_2537_ (
    .a(n_0395_),
    .b(n_0396_),
    .c(N10908)
  );
  and_ii n_2538_ (
    .a(n_0061_),
    .b(n_1296_),
    .c(n_0397_)
  );
  or_bb n_2539_ (
    .a(n_0397_),
    .b(n_0062_),
    .c(n_0398_)
  );
  and_bi n_2540_ (
    .a(n_0059_),
    .b(n_0398_),
    .c(n_0399_)
  );
  and_bi n_2541_ (
    .a(n_0398_),
    .b(n_0059_),
    .c(n_0400_)
  );
  and_ii n_2542_ (
    .a(n_0400_),
    .b(n_0399_),
    .c(n_0401_)
  );
  and_ii n_2543_ (
    .a(n_0401_),
    .b(n_0066_),
    .c(n_0402_)
  );
  and_bi n_2544_ (
    .a(n_0057_),
    .b(n_0082_),
    .c(n_0403_)
  );
  and_bi n_2545_ (
    .a(n_1295_),
    .b(n_0052_),
    .c(n_0404_)
  );
  and_ii n_2546_ (
    .a(n_0053_),
    .b(n_1295_),
    .c(n_0405_)
  );
  and_ii n_2547_ (
    .a(n_0405_),
    .b(n_0404_),
    .c(n_0406_)
  );
  and_bi n_2548_ (
    .a(n_0078_),
    .b(n_0406_),
    .c(n_0407_)
  );
  and_bi n_2549_ (
    .a(n_0406_),
    .b(n_0078_),
    .c(n_0408_)
  );
  and_ii n_2550_ (
    .a(n_0408_),
    .b(n_0407_),
    .c(n_0409_)
  );
  and_bb n_2551_ (
    .a(n_0409_),
    .b(n_0403_),
    .c(n_0410_)
  );
  and_ii n_2552_ (
    .a(n_0409_),
    .b(n_0403_),
    .c(n_0411_)
  );
  or_bb n_2553_ (
    .a(n_0411_),
    .b(n_0410_),
    .c(n_0412_)
  );
  or_bb n_2554_ (
    .a(n_0412_),
    .b(n_0402_),
    .c(n_0413_)
  );
  and_bb n_2555_ (
    .a(n_0412_),
    .b(n_0402_),
    .c(n_0414_)
  );
  and_bi n_2556_ (
    .a(n_0413_),
    .b(n_0414_),
    .c(n_0415_)
  );
  or_bb n_2557_ (
    .a(n_0415_),
    .b(n_0019_),
    .c(n_0416_)
  );
  and_ii n_2558_ (
    .a(n_0052_),
    .b(n_1294_),
    .c(n_0417_)
  );
  and_ii n_2559_ (
    .a(n_0417_),
    .b(n_0054_),
    .c(n_0418_)
  );
  and_bi n_2560_ (
    .a(n_0418_),
    .b(n_0079_),
    .c(n_0419_)
  );
  and_bi n_2561_ (
    .a(n_0079_),
    .b(n_0418_),
    .c(n_0420_)
  );
  and_ii n_2562_ (
    .a(n_0420_),
    .b(n_0419_),
    .c(n_0421_)
  );
  and_bi n_2563_ (
    .a(n_0057_),
    .b(n_0421_),
    .c(n_0422_)
  );
  and_bi n_2564_ (
    .a(n_0421_),
    .b(n_0057_),
    .c(n_0423_)
  );
  and_ii n_2565_ (
    .a(n_0423_),
    .b(n_0422_),
    .c(n_0424_)
  );
  and_bb n_2566_ (
    .a(n_0424_),
    .b(n_0401_),
    .c(n_0425_)
  );
  and_ii n_2567_ (
    .a(n_0424_),
    .b(n_0401_),
    .c(n_0426_)
  );
  or_bb n_2568_ (
    .a(n_0426_),
    .b(n_0425_),
    .c(n_0427_)
  );
  and_bi n_2569_ (
    .a(n_0019_),
    .b(n_0427_),
    .c(n_0428_)
  );
  and_bi n_2570_ (
    .a(n_0416_),
    .b(n_0428_),
    .c(n_0429_)
  );
  and_ii n_2571_ (
    .a(n_0064_),
    .b(n_0063_),
    .c(n_0430_)
  );
  or_bb n_2572_ (
    .a(n_0430_),
    .b(n_0065_),
    .c(n_0431_)
  );
  or_bi n_2573_ (
    .a(n_0429_),
    .b(n_0431_),
    .c(n_0432_)
  );
  and_bi n_2574_ (
    .a(n_0429_),
    .b(n_0431_),
    .c(n_0433_)
  );
  and_bi n_2575_ (
    .a(n_0432_),
    .b(n_0433_),
    .c(n_0434_)
  );
  and_bi n_2576_ (
    .a(n_0034_),
    .b(n_0028_),
    .c(n_0435_)
  );
  and_ii n_2577_ (
    .a(n_0435_),
    .b(n_0035_),
    .c(n_0436_)
  );
  and_bi n_2578_ (
    .a(n_0038_),
    .b(n_0031_),
    .c(n_0437_)
  );
  and_bi n_2579_ (
    .a(n_0037_),
    .b(n_0367_),
    .c(n_0438_)
  );
  or_bb n_2580_ (
    .a(n_0438_),
    .b(n_0437_),
    .c(n_0439_)
  );
  and_bi n_2581_ (
    .a(n_0360_),
    .b(n_0040_),
    .c(n_0440_)
  );
  and_bi n_2582_ (
    .a(n_0040_),
    .b(n_0360_),
    .c(n_0441_)
  );
  or_bb n_2583_ (
    .a(n_0441_),
    .b(n_0440_),
    .c(n_0442_)
  );
  and_ii n_2584_ (
    .a(n_0442_),
    .b(n_0439_),
    .c(n_0443_)
  );
  and_bb n_2585_ (
    .a(n_0442_),
    .b(n_0439_),
    .c(n_0444_)
  );
  and_ii n_2586_ (
    .a(n_0444_),
    .b(n_0443_),
    .c(n_0445_)
  );
  and_bi n_2587_ (
    .a(n_0445_),
    .b(n_0436_),
    .c(n_0446_)
  );
  and_bi n_2588_ (
    .a(n_0436_),
    .b(n_0445_),
    .c(n_0447_)
  );
  or_bb n_2589_ (
    .a(n_0447_),
    .b(n_0446_),
    .c(n_0448_)
  );
  and_ii n_2590_ (
    .a(n_0448_),
    .b(n_0070_),
    .c(n_0449_)
  );
  and_bi n_2591_ (
    .a(n_0037_),
    .b(n_0031_),
    .c(n_0450_)
  );
  and_ii n_2592_ (
    .a(n_0450_),
    .b(n_0038_),
    .c(n_0451_)
  );
  and_bi n_2593_ (
    .a(n_0451_),
    .b(n_0040_),
    .c(n_0452_)
  );
  and_bi n_2594_ (
    .a(n_0040_),
    .b(n_0451_),
    .c(n_0453_)
  );
  and_ii n_2595_ (
    .a(n_0453_),
    .b(n_0452_),
    .c(n_0454_)
  );
  and_ii n_2596_ (
    .a(n_0372_),
    .b(n_0367_),
    .c(n_0455_)
  );
  and_ii n_2597_ (
    .a(n_0455_),
    .b(n_0039_),
    .c(n_0456_)
  );
  or_ii n_2598_ (
    .a(n_0456_),
    .b(n_0360_),
    .c(n_0457_)
  );
  and_ii n_2599_ (
    .a(n_0456_),
    .b(n_0360_),
    .c(n_0458_)
  );
  and_bi n_2600_ (
    .a(n_0457_),
    .b(n_0458_),
    .c(n_0459_)
  );
  and_ii n_2601_ (
    .a(n_0459_),
    .b(n_0043_),
    .c(n_0460_)
  );
  and_bb n_2602_ (
    .a(n_0459_),
    .b(n_0043_),
    .c(n_0461_)
  );
  and_ii n_2603_ (
    .a(n_0461_),
    .b(n_0460_),
    .c(n_0462_)
  );
  and_bi n_2604_ (
    .a(n_0462_),
    .b(n_0454_),
    .c(n_0463_)
  );
  and_bi n_2605_ (
    .a(n_0454_),
    .b(n_0462_),
    .c(n_0464_)
  );
  or_bb n_2606_ (
    .a(n_0464_),
    .b(n_0463_),
    .c(n_0465_)
  );
  and_bi n_2607_ (
    .a(n_0070_),
    .b(n_0465_),
    .c(n_0466_)
  );
  and_ii n_2608_ (
    .a(n_0466_),
    .b(n_0449_),
    .c(n_0467_)
  );
  or_bi n_2609_ (
    .a(n_0434_),
    .b(n_0467_),
    .c(n_0468_)
  );
  and_bi n_2610_ (
    .a(n_0434_),
    .b(n_0467_),
    .c(n_0469_)
  );
  and_bi n_2611_ (
    .a(n_0468_),
    .b(n_0469_),
    .c(N11333)
  );
  and_bi n_2612_ (
    .a(n_0176_),
    .b(n_0168_),
    .c(n_0470_)
  );
  or_bb n_2613_ (
    .a(n_0470_),
    .b(n_0167_),
    .c(n_0471_)
  );
  and_bi n_2614_ (
    .a(n_0111_),
    .b(n_0116_),
    .c(n_0472_)
  );
  and_bi n_2615_ (
    .a(n_0116_),
    .b(n_0111_),
    .c(n_0473_)
  );
  and_ii n_2616_ (
    .a(n_0473_),
    .b(n_0472_),
    .c(n_0474_)
  );
  and_bi n_2617_ (
    .a(n_0379_),
    .b(n_0474_),
    .c(n_0475_)
  );
  and_bi n_2618_ (
    .a(n_0474_),
    .b(n_0379_),
    .c(n_0476_)
  );
  or_bb n_2619_ (
    .a(n_0476_),
    .b(n_0475_),
    .c(n_0477_)
  );
  and_ii n_2620_ (
    .a(n_0112_),
    .b(n_0025_),
    .c(n_0478_)
  );
  and_bi n_2621_ (
    .a(n_0113_),
    .b(n_0478_),
    .c(n_0479_)
  );
  and_bi n_2622_ (
    .a(n_0110_),
    .b(n_0479_),
    .c(n_0480_)
  );
  and_bi n_2623_ (
    .a(n_0479_),
    .b(n_0110_),
    .c(n_0481_)
  );
  and_ii n_2624_ (
    .a(n_0481_),
    .b(n_0480_),
    .c(n_0482_)
  );
  and_bb n_2625_ (
    .a(n_0116_),
    .b(n_0114_),
    .c(n_0483_)
  );
  and_ii n_2626_ (
    .a(n_0483_),
    .b(n_0482_),
    .c(n_0484_)
  );
  and_bi n_2627_ (
    .a(n_0108_),
    .b(n_0114_),
    .c(n_0485_)
  );
  and_ii n_2628_ (
    .a(n_0103_),
    .b(n_0024_),
    .c(n_0486_)
  );
  and_bi n_2629_ (
    .a(n_0024_),
    .b(n_0104_),
    .c(n_0487_)
  );
  or_bb n_2630_ (
    .a(n_0487_),
    .b(n_0486_),
    .c(n_0488_)
  );
  and_bi n_2631_ (
    .a(n_0121_),
    .b(n_0488_),
    .c(n_0489_)
  );
  and_bi n_2632_ (
    .a(n_0488_),
    .b(n_0121_),
    .c(n_0490_)
  );
  or_bb n_2633_ (
    .a(n_0490_),
    .b(n_0489_),
    .c(n_0491_)
  );
  and_ii n_2634_ (
    .a(n_0491_),
    .b(n_0485_),
    .c(n_0492_)
  );
  and_bb n_2635_ (
    .a(n_0491_),
    .b(n_0485_),
    .c(n_0493_)
  );
  and_ii n_2636_ (
    .a(n_0493_),
    .b(n_0492_),
    .c(n_0494_)
  );
  and_bb n_2637_ (
    .a(n_0494_),
    .b(n_0484_),
    .c(n_0495_)
  );
  and_ii n_2638_ (
    .a(n_0494_),
    .b(n_0484_),
    .c(n_0496_)
  );
  or_bb n_2639_ (
    .a(n_0496_),
    .b(n_0495_),
    .c(n_0497_)
  );
  and_bi n_2640_ (
    .a(n_0076_),
    .b(n_0497_),
    .c(n_0498_)
  );
  and_bi n_2641_ (
    .a(n_0023_),
    .b(n_0103_),
    .c(n_0499_)
  );
  and_ii n_2642_ (
    .a(n_0105_),
    .b(n_0499_),
    .c(n_0500_)
  );
  and_bi n_2643_ (
    .a(n_0500_),
    .b(n_0121_),
    .c(n_0501_)
  );
  and_bi n_2644_ (
    .a(n_0121_),
    .b(n_0500_),
    .c(n_0502_)
  );
  and_ii n_2645_ (
    .a(n_0502_),
    .b(n_0501_),
    .c(n_0503_)
  );
  and_bi n_2646_ (
    .a(n_0503_),
    .b(n_0108_),
    .c(n_0504_)
  );
  and_bi n_2647_ (
    .a(n_0108_),
    .b(n_0503_),
    .c(n_0505_)
  );
  and_ii n_2648_ (
    .a(n_0505_),
    .b(n_0504_),
    .c(n_0506_)
  );
  and_bi n_2649_ (
    .a(n_0506_),
    .b(n_0482_),
    .c(n_0507_)
  );
  and_bi n_2650_ (
    .a(n_0482_),
    .b(n_0506_),
    .c(n_0508_)
  );
  or_bb n_2651_ (
    .a(n_0508_),
    .b(n_0507_),
    .c(n_0509_)
  );
  and_bi n_2652_ (
    .a(n_0074_),
    .b(n_0509_),
    .c(n_0510_)
  );
  or_bb n_2653_ (
    .a(n_0510_),
    .b(n_0498_),
    .c(n_0511_)
  );
  or_bb n_2654_ (
    .a(n_0511_),
    .b(n_0477_),
    .c(n_0512_)
  );
  and_bb n_2655_ (
    .a(n_0511_),
    .b(n_0477_),
    .c(n_0513_)
  );
  and_bi n_2656_ (
    .a(n_0512_),
    .b(n_0513_),
    .c(n_0514_)
  );
  or_bi n_2657_ (
    .a(n_0471_),
    .b(n_0514_),
    .c(n_0515_)
  );
  and_bi n_2658_ (
    .a(n_0471_),
    .b(n_0514_),
    .c(n_0516_)
  );
  and_bi n_2659_ (
    .a(n_0515_),
    .b(n_0516_),
    .c(N11334)
  );
  and_bb n_2660_ (
    .a(n_1308_),
    .b(n_1306_),
    .c(n_0517_)
  );
  and_ii n_2661_ (
    .a(n_0517_),
    .b(n_1309_),
    .c(n_0518_)
  );
  and_bb n_2662_ (
    .a(n_1315_),
    .b(n_1314_),
    .c(n_0519_)
  );
  or_bb n_2663_ (
    .a(n_0519_),
    .b(n_0518_),
    .c(n_0520_)
  );
  and_bi n_2664_ (
    .a(n_0382_),
    .b(n_0385_),
    .c(n_0521_)
  );
  and_bi n_2665_ (
    .a(n_0385_),
    .b(n_0382_),
    .c(n_0522_)
  );
  and_ii n_2666_ (
    .a(n_0522_),
    .b(n_0521_),
    .c(n_0523_)
  );
  and_bb n_2667_ (
    .a(n_0523_),
    .b(n_0520_),
    .c(n_0524_)
  );
  and_ii n_2668_ (
    .a(n_0523_),
    .b(n_0520_),
    .c(n_0525_)
  );
  and_ii n_2669_ (
    .a(n_0525_),
    .b(n_0524_),
    .c(n_0526_)
  );
  or_bb n_2670_ (
    .a(n_0526_),
    .b(n_1319_),
    .c(n_0527_)
  );
  and_bb n_2671_ (
    .a(n_0526_),
    .b(n_1319_),
    .c(n_0528_)
  );
  and_bi n_2672_ (
    .a(n_0527_),
    .b(n_0528_),
    .c(n_0529_)
  );
  and_bi n_2673_ (
    .a(n_0015_),
    .b(n_0529_),
    .c(n_0530_)
  );
  and_bi n_2674_ (
    .a(n_1313_),
    .b(n_1310_),
    .c(n_0531_)
  );
  and_bi n_2675_ (
    .a(n_1303_),
    .b(n_0531_),
    .c(n_0532_)
  );
  and_bi n_2676_ (
    .a(n_0390_),
    .b(n_0532_),
    .c(n_0533_)
  );
  and_bi n_2677_ (
    .a(n_0532_),
    .b(n_0390_),
    .c(n_0534_)
  );
  or_bb n_2678_ (
    .a(n_0534_),
    .b(n_0533_),
    .c(n_0535_)
  );
  and_bi n_2679_ (
    .a(n_1310_),
    .b(n_1315_),
    .c(n_0536_)
  );
  and_bi n_2680_ (
    .a(n_1315_),
    .b(n_1306_),
    .c(n_0537_)
  );
  and_ii n_2681_ (
    .a(n_0537_),
    .b(n_0536_),
    .c(n_0538_)
  );
  and_bi n_2682_ (
    .a(n_0538_),
    .b(n_0382_),
    .c(n_0539_)
  );
  and_bi n_2683_ (
    .a(n_0382_),
    .b(n_0538_),
    .c(n_0540_)
  );
  and_ii n_2684_ (
    .a(n_0540_),
    .b(n_0539_),
    .c(n_0541_)
  );
  or_bi n_2685_ (
    .a(n_0535_),
    .b(n_0541_),
    .c(n_0542_)
  );
  and_bi n_2686_ (
    .a(n_0535_),
    .b(n_0541_),
    .c(n_0543_)
  );
  or_bi n_2687_ (
    .a(n_0543_),
    .b(n_0542_),
    .c(n_0544_)
  );
  and_bi n_2688_ (
    .a(n_0544_),
    .b(n_0015_),
    .c(n_0545_)
  );
  and_ii n_2689_ (
    .a(n_0545_),
    .b(n_0530_),
    .c(n_0546_)
  );
  and_bi n_2690_ (
    .a(n_0008_),
    .b(n_1333_),
    .c(n_0547_)
  );
  and_ii n_2691_ (
    .a(n_0547_),
    .b(n_0009_),
    .c(n_0548_)
  );
  and_bi n_2692_ (
    .a(n_0152_),
    .b(n_1324_),
    .c(n_0549_)
  );
  and_bi n_2693_ (
    .a(n_1324_),
    .b(n_0152_),
    .c(n_0550_)
  );
  and_ii n_2694_ (
    .a(n_0550_),
    .b(n_0549_),
    .c(n_0551_)
  );
  and_bb n_2695_ (
    .a(n_0551_),
    .b(n_0548_),
    .c(n_0552_)
  );
  and_ii n_2696_ (
    .a(n_0551_),
    .b(n_0548_),
    .c(n_0553_)
  );
  and_ii n_2697_ (
    .a(n_0553_),
    .b(n_0552_),
    .c(n_0554_)
  );
  and_bi n_2698_ (
    .a(n_0145_),
    .b(n_0554_),
    .c(n_0555_)
  );
  and_bi n_2699_ (
    .a(n_0554_),
    .b(n_0145_),
    .c(n_0556_)
  );
  and_ii n_2700_ (
    .a(n_0556_),
    .b(n_0555_),
    .c(n_0557_)
  );
  and_bi n_2701_ (
    .a(n_0005_),
    .b(n_0557_),
    .c(n_0558_)
  );
  and_bi n_2702_ (
    .a(n_1336_),
    .b(n_0145_),
    .c(n_0559_)
  );
  or_bb n_2703_ (
    .a(n_0559_),
    .b(n_1340_),
    .c(n_0560_)
  );
  and_bi n_2704_ (
    .a(n_0010_),
    .b(n_0147_),
    .c(n_0561_)
  );
  and_ii n_2705_ (
    .a(n_1325_),
    .b(n_1320_),
    .c(n_0562_)
  );
  and_bi n_2706_ (
    .a(n_1323_),
    .b(n_1326_),
    .c(n_0563_)
  );
  or_bb n_2707_ (
    .a(n_0563_),
    .b(n_0562_),
    .c(n_0564_)
  );
  and_ii n_2708_ (
    .a(n_0564_),
    .b(n_0561_),
    .c(n_0565_)
  );
  and_bb n_2709_ (
    .a(n_0564_),
    .b(n_0561_),
    .c(n_0566_)
  );
  and_ii n_2710_ (
    .a(n_0566_),
    .b(n_0565_),
    .c(n_0567_)
  );
  or_bb n_2711_ (
    .a(n_0567_),
    .b(n_0560_),
    .c(n_0568_)
  );
  and_bb n_2712_ (
    .a(n_0567_),
    .b(n_0560_),
    .c(n_0569_)
  );
  or_bi n_2713_ (
    .a(n_0569_),
    .b(n_0568_),
    .c(n_0570_)
  );
  and_bi n_2714_ (
    .a(n_0570_),
    .b(n_0005_),
    .c(n_0571_)
  );
  and_ii n_2715_ (
    .a(n_0571_),
    .b(n_0558_),
    .c(n_0572_)
  );
  and_ii n_2716_ (
    .a(n_1334_),
    .b(n_1330_),
    .c(n_0573_)
  );
  or_bi n_2717_ (
    .a(n_0573_),
    .b(n_1335_),
    .c(n_0574_)
  );
  and_bb n_2718_ (
    .a(n_0574_),
    .b(n_0572_),
    .c(n_0575_)
  );
  and_ii n_2719_ (
    .a(n_0574_),
    .b(n_0572_),
    .c(n_0576_)
  );
  and_ii n_2720_ (
    .a(n_0576_),
    .b(n_0575_),
    .c(n_0577_)
  );
  and_ii n_2721_ (
    .a(n_0577_),
    .b(n_0546_),
    .c(n_0578_)
  );
  and_bb n_2722_ (
    .a(n_0577_),
    .b(n_0546_),
    .c(n_0579_)
  );
  or_bb n_2723_ (
    .a(n_0579_),
    .b(n_0578_),
    .c(N11340)
  );
  and_ii n_2724_ (
    .a(n_1369_),
    .b(n_1353_),
    .c(n_0580_)
  );
  and_bi n_2725_ (
    .a(n_1369_),
    .b(n_1349_),
    .c(n_0581_)
  );
  and_ii n_2726_ (
    .a(n_0581_),
    .b(n_0580_),
    .c(n_0582_)
  );
  and_ii n_2727_ (
    .a(n_0582_),
    .b(n_1355_),
    .c(n_0583_)
  );
  and_bb n_2728_ (
    .a(n_0582_),
    .b(n_1355_),
    .c(n_0584_)
  );
  or_bb n_2729_ (
    .a(n_0584_),
    .b(n_0583_),
    .c(n_0585_)
  );
  and_ii n_2730_ (
    .a(n_0001_),
    .b(n_0000_),
    .c(n_0586_)
  );
  and_bi n_2731_ (
    .a(n_0002_),
    .b(n_0586_),
    .c(n_0587_)
  );
  or_bb n_2732_ (
    .a(n_0587_),
    .b(n_1368_),
    .c(n_0588_)
  );
  and_bi n_2733_ (
    .a(n_0587_),
    .b(n_0354_),
    .c(n_0589_)
  );
  and_bi n_2734_ (
    .a(n_0588_),
    .b(n_0589_),
    .c(n_0590_)
  );
  and_ii n_2735_ (
    .a(n_0590_),
    .b(n_0585_),
    .c(n_0591_)
  );
  and_bb n_2736_ (
    .a(n_0590_),
    .b(n_0585_),
    .c(n_0592_)
  );
  and_ii n_2737_ (
    .a(n_0592_),
    .b(n_0591_),
    .c(n_0593_)
  );
  or_bb n_2738_ (
    .a(n_0593_),
    .b(n_1366_),
    .c(n_0594_)
  );
  and_bi n_2739_ (
    .a(n_1348_),
    .b(n_1351_),
    .c(n_0595_)
  );
  and_bi n_2740_ (
    .a(n_1351_),
    .b(n_1349_),
    .c(n_0596_)
  );
  or_bb n_2741_ (
    .a(n_0596_),
    .b(n_0595_),
    .c(n_0597_)
  );
  or_bi n_2742_ (
    .a(n_0597_),
    .b(n_1371_),
    .c(n_0598_)
  );
  and_bi n_2743_ (
    .a(n_1355_),
    .b(n_0598_),
    .c(n_0599_)
  );
  and_bb n_2744_ (
    .a(n_0598_),
    .b(n_0344_),
    .c(n_0600_)
  );
  and_bi n_2745_ (
    .a(n_0600_),
    .b(n_1355_),
    .c(n_0601_)
  );
  and_ii n_2746_ (
    .a(n_0601_),
    .b(n_0599_),
    .c(n_0602_)
  );
  and_ii n_2747_ (
    .a(n_0602_),
    .b(n_0587_),
    .c(n_0603_)
  );
  and_bb n_2748_ (
    .a(n_0602_),
    .b(n_0587_),
    .c(n_0604_)
  );
  or_bb n_2749_ (
    .a(n_0604_),
    .b(n_0603_),
    .c(n_0605_)
  );
  and_bi n_2750_ (
    .a(n_1366_),
    .b(n_0605_),
    .c(n_0606_)
  );
  or_bb n_2751_ (
    .a(n_0606_),
    .b(n_0668_),
    .c(n_0607_)
  );
  and_bi n_2752_ (
    .a(n_0594_),
    .b(n_0607_),
    .c(n_0608_)
  );
  and_bb n_2753_ (
    .a(n_0593_),
    .b(n_1362_),
    .c(n_0609_)
  );
  or_ii n_2754_ (
    .a(n_1361_),
    .b(n_0668_),
    .c(n_0610_)
  );
  and_bi n_2755_ (
    .a(n_0605_),
    .b(n_0610_),
    .c(n_0611_)
  );
  or_bb n_2756_ (
    .a(n_0611_),
    .b(n_0609_),
    .c(n_0612_)
  );
  or_bb n_2757_ (
    .a(n_0612_),
    .b(n_0608_),
    .c(n_0613_)
  );
  and_bb n_2758_ (
    .a(n_0700_),
    .b(n_0680_),
    .c(n_0614_)
  );
  or_bb n_2759_ (
    .a(n_0614_),
    .b(n_0701_),
    .c(n_0615_)
  );
  and_bi n_2760_ (
    .a(n_0697_),
    .b(n_0710_),
    .c(n_0616_)
  );
  and_bb n_2761_ (
    .a(n_0692_),
    .b(n_0666_),
    .c(n_0617_)
  );
  and_bi n_2762_ (
    .a(n_0693_),
    .b(n_0617_),
    .c(n_0618_)
  );
  and_bi n_2763_ (
    .a(n_0618_),
    .b(n_0676_),
    .c(n_0619_)
  );
  and_bi n_2764_ (
    .a(n_0676_),
    .b(n_0618_),
    .c(n_0620_)
  );
  and_ii n_2765_ (
    .a(n_0620_),
    .b(n_0619_),
    .c(n_0621_)
  );
  and_bi n_2766_ (
    .a(n_0621_),
    .b(n_0616_),
    .c(n_0622_)
  );
  and_bi n_2767_ (
    .a(n_0616_),
    .b(n_0621_),
    .c(n_0623_)
  );
  or_bb n_2768_ (
    .a(n_0623_),
    .b(n_0622_),
    .c(n_0624_)
  );
  and_ii n_2769_ (
    .a(n_0624_),
    .b(n_0615_),
    .c(n_0625_)
  );
  and_bb n_2770_ (
    .a(n_0624_),
    .b(n_0615_),
    .c(n_0626_)
  );
  or_bb n_2771_ (
    .a(n_0626_),
    .b(N367),
    .c(n_0627_)
  );
  or_bb n_2772_ (
    .a(n_0627_),
    .b(n_0625_),
    .c(n_0628_)
  );
  and_ii n_2773_ (
    .a(n_0700_),
    .b(n_0694_),
    .c(n_0629_)
  );
  and_ii n_2774_ (
    .a(n_0690_),
    .b(n_0665_),
    .c(n_0630_)
  );
  or_bi n_2775_ (
    .a(n_0691_),
    .b(n_0697_),
    .c(n_0631_)
  );
  and_bi n_2776_ (
    .a(n_0665_),
    .b(n_0631_),
    .c(n_0632_)
  );
  and_ii n_2777_ (
    .a(n_0632_),
    .b(n_0630_),
    .c(n_0633_)
  );
  or_bi n_2778_ (
    .a(n_0629_),
    .b(n_0633_),
    .c(n_0634_)
  );
  and_bi n_2779_ (
    .a(n_0629_),
    .b(n_0633_),
    .c(n_0635_)
  );
  and_bi n_2780_ (
    .a(n_0634_),
    .b(n_0635_),
    .c(n_0636_)
  );
  and_bi n_2781_ (
    .a(n_1364_),
    .b(n_0621_),
    .c(n_0637_)
  );
  and_bi n_2782_ (
    .a(n_0621_),
    .b(n_1364_),
    .c(n_0638_)
  );
  or_bb n_2783_ (
    .a(n_0638_),
    .b(n_0637_),
    .c(n_0639_)
  );
  or_bi n_2784_ (
    .a(n_0636_),
    .b(n_0639_),
    .c(n_0640_)
  );
  and_bi n_2785_ (
    .a(n_0636_),
    .b(n_0639_),
    .c(n_0641_)
  );
  or_bb n_2786_ (
    .a(n_0641_),
    .b(n_0668_),
    .c(n_0642_)
  );
  and_bi n_2787_ (
    .a(n_0640_),
    .b(n_0642_),
    .c(n_0643_)
  );
  and_bi n_2788_ (
    .a(n_0628_),
    .b(n_0643_),
    .c(n_0644_)
  );
  or_bi n_2789_ (
    .a(n_0686_),
    .b(n_0707_),
    .c(n_0645_)
  );
  and_bi n_2790_ (
    .a(n_0686_),
    .b(n_0707_),
    .c(n_0646_)
  );
  and_bi n_2791_ (
    .a(n_0645_),
    .b(n_0646_),
    .c(n_0647_)
  );
  and_ii n_2792_ (
    .a(n_0647_),
    .b(n_0644_),
    .c(n_0648_)
  );
  and_bb n_2793_ (
    .a(n_0647_),
    .b(n_0644_),
    .c(n_0649_)
  );
  and_ii n_2794_ (
    .a(n_0649_),
    .b(n_0648_),
    .c(n_0650_)
  );
  or_bb n_2795_ (
    .a(n_0650_),
    .b(n_0613_),
    .c(n_0651_)
  );
  and_bb n_2796_ (
    .a(n_0650_),
    .b(n_0613_),
    .c(n_0652_)
  );
  and_bi n_2797_ (
    .a(n_0651_),
    .b(n_0652_),
    .c(N11342)
  );
  and_bi n_2798_ (
    .a(n_0163_),
    .b(n_0178_),
    .c(N10104)
  );
  and_bi n_2799_ (
    .a(n_0180_),
    .b(n_0342_),
    .c(N10628)
  );
  and_bi n_2800_ (
    .a(n_0163_),
    .b(n_0178_),
    .c(N10706)
  );
  and_bi n_2801_ (
    .a(n_0163_),
    .b(n_0178_),
    .c(N10759)
  );
  assign N10103 = N10102;
  assign N10838 = N10837;
  assign N10840 = N10839;
  assign N1112 = N1110;
  assign N1114 = N1111;
  assign N1489 = N1113;
  assign N1490 = N1;
  assign N241_O = N241_I;
  assign N387 = N1;
  assign N388 = N1;
  assign N478 = N248;
  assign N482 = N254;
  assign N484 = N257;
  assign N486 = N260;
  assign N489 = N263;
  assign N492 = N267;
  assign N501 = N274;
  assign N505 = N280;
  assign N507 = N283;
  assign N509 = N286;
  assign N511 = N289;
  assign N513 = N293;
  assign N515 = N296;
  assign N517 = N299;
  assign N519 = N303;
  assign N535 = N307;
  assign N537 = N310;
  assign N539 = N313;
  assign N541 = N316;
  assign N543 = N319;
  assign N545 = N322;
  assign N547 = N325;
  assign N549 = N328;
  assign N551 = N331;
  assign N553 = N334;
  assign N556 = N337;
  assign N559 = N343;
  assign N561 = N346;
  assign N563 = N349;
  assign N565 = N352;
  assign N567 = N355;
  assign N569 = N358;
  assign N571 = N361;
  assign N573 = N364;
  assign N582 = N1111;
  assign N643 = N251;
  assign N707 = N277;
  assign N813 = N340;
  assign N889 = N1;
  assign N945 = N106;
endmodule
