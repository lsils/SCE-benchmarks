module apc64bits(in_15_,in_0_,in_4_,in_29_,in_38_,in_53_,in_42_,in_11_,in_59_,in_48_,in_54_,in_16_,in_43_,in_37_,in_61_,in_14_,in_62_,in_60_,in_40_,in_5_,in_28_,in_7_,in_6_,in_34_,in_57_,in_3_,in_56_,in_45_,in_10_,in_27_,in_21_,in_25_,in_22_,in_12_,in_58_,in_36_,in_51_,in_18_,in_9_,in_39_,in_24_,in_26_,in_8_,in_41_,in_55_,in_2_,in_49_,in_19_,in_35_,in_50_,in_32_,in_30_,in_33_,in_17_,in_31_,in_44_,in_1_,in_23_,in_52_,in_20_,in_46_,in_13_,in_63_,in_47_,out_1_,out_3_,out_6_,out_2_,out_0_,out_4_,out_5_);
    wire jinkela_wire_0;
    wire jinkela_wire_1;
    wire jinkela_wire_2;
    wire jinkela_wire_3;
    wire jinkela_wire_4;
    wire jinkela_wire_5;
    wire jinkela_wire_6;
    wire jinkela_wire_7;
    wire jinkela_wire_8;
    wire jinkela_wire_9;
    wire jinkela_wire_10;
    wire jinkela_wire_11;
    wire jinkela_wire_12;
    wire jinkela_wire_13;
    wire jinkela_wire_14;
    wire jinkela_wire_15;
    wire jinkela_wire_16;
    wire jinkela_wire_17;
    wire jinkela_wire_18;
    wire jinkela_wire_19;
    wire jinkela_wire_20;
    wire jinkela_wire_21;
    wire jinkela_wire_22;
    wire jinkela_wire_23;
    wire jinkela_wire_24;
    wire jinkela_wire_25;
    wire jinkela_wire_26;
    wire jinkela_wire_27;
    wire jinkela_wire_28;
    wire jinkela_wire_29;
    wire jinkela_wire_30;
    wire jinkela_wire_31;
    wire jinkela_wire_32;
    wire jinkela_wire_33;
    wire jinkela_wire_34;
    wire jinkela_wire_35;
    wire jinkela_wire_36;
    wire jinkela_wire_37;
    wire jinkela_wire_38;
    wire jinkela_wire_39;
    wire jinkela_wire_40;
    wire jinkela_wire_41;
    wire jinkela_wire_42;
    wire jinkela_wire_43;
    wire jinkela_wire_44;
    wire jinkela_wire_45;
    wire jinkela_wire_46;
    wire jinkela_wire_47;
    wire jinkela_wire_48;
    wire jinkela_wire_49;
    wire jinkela_wire_50;
    wire jinkela_wire_51;
    wire jinkela_wire_52;
    wire jinkela_wire_53;
    wire jinkela_wire_54;
    wire jinkela_wire_55;
    wire jinkela_wire_56;
    wire jinkela_wire_57;
    wire jinkela_wire_58;
    wire jinkela_wire_59;
    wire jinkela_wire_60;
    wire jinkela_wire_61;
    wire jinkela_wire_62;
    wire jinkela_wire_63;
    wire jinkela_wire_64;
    wire jinkela_wire_65;
    wire jinkela_wire_66;
    wire jinkela_wire_67;
    wire jinkela_wire_68;
    wire jinkela_wire_69;
    wire jinkela_wire_70;
    wire jinkela_wire_71;
    wire jinkela_wire_72;
    wire jinkela_wire_73;
    wire jinkela_wire_74;
    wire jinkela_wire_75;
    wire jinkela_wire_76;
    wire jinkela_wire_77;
    wire jinkela_wire_78;
    wire jinkela_wire_79;
    wire jinkela_wire_80;
    wire jinkela_wire_81;
    wire jinkela_wire_82;
    wire jinkela_wire_83;
    wire jinkela_wire_84;
    wire jinkela_wire_85;
    wire jinkela_wire_86;
    wire jinkela_wire_87;
    wire jinkela_wire_88;
    wire jinkela_wire_89;
    wire jinkela_wire_90;
    wire jinkela_wire_91;
    wire jinkela_wire_92;
    wire jinkela_wire_93;
    wire jinkela_wire_94;
    wire jinkela_wire_95;
    wire jinkela_wire_96;
    wire jinkela_wire_97;
    wire jinkela_wire_98;
    wire jinkela_wire_99;
    wire jinkela_wire_100;
    wire jinkela_wire_101;
    wire jinkela_wire_102;
    wire jinkela_wire_103;
    wire jinkela_wire_104;
    wire jinkela_wire_105;
    wire jinkela_wire_106;
    wire jinkela_wire_107;
    wire jinkela_wire_108;
    wire jinkela_wire_109;
    wire jinkela_wire_110;
    wire jinkela_wire_111;
    wire jinkela_wire_112;
    wire jinkela_wire_113;
    wire jinkela_wire_114;
    wire jinkela_wire_115;
    wire jinkela_wire_116;
    wire jinkela_wire_117;
    wire jinkela_wire_118;
    wire jinkela_wire_119;
    wire jinkela_wire_120;
    wire jinkela_wire_121;
    wire jinkela_wire_122;
    wire jinkela_wire_123;
    wire jinkela_wire_124;
    wire jinkela_wire_125;
    wire jinkela_wire_126;
    wire jinkela_wire_127;
    wire jinkela_wire_128;
    wire jinkela_wire_129;
    wire jinkela_wire_130;
    wire jinkela_wire_131;
    wire jinkela_wire_132;
    wire jinkela_wire_133;
    wire jinkela_wire_134;
    wire jinkela_wire_135;
    wire jinkela_wire_136;
    wire jinkela_wire_137;
    wire jinkela_wire_138;
    wire jinkela_wire_139;
    wire jinkela_wire_140;
    wire jinkela_wire_141;
    wire jinkela_wire_142;
    wire jinkela_wire_143;
    wire jinkela_wire_144;
    wire jinkela_wire_145;
    wire jinkela_wire_146;
    wire jinkela_wire_147;
    wire jinkela_wire_148;
    wire jinkela_wire_149;
    wire jinkela_wire_150;
    wire jinkela_wire_151;
    wire jinkela_wire_152;
    wire jinkela_wire_153;
    wire jinkela_wire_154;
    wire jinkela_wire_155;
    wire jinkela_wire_156;
    wire jinkela_wire_157;
    wire jinkela_wire_158;
    wire jinkela_wire_159;
    wire jinkela_wire_160;
    wire jinkela_wire_161;
    wire jinkela_wire_162;
    wire jinkela_wire_163;
    wire jinkela_wire_164;
    wire jinkela_wire_165;
    wire jinkela_wire_166;
    wire jinkela_wire_167;
    wire jinkela_wire_168;
    wire jinkela_wire_169;
    wire jinkela_wire_170;
    wire jinkela_wire_171;
    wire jinkela_wire_172;
    wire jinkela_wire_173;
    wire jinkela_wire_174;
    wire jinkela_wire_175;
    wire jinkela_wire_176;
    wire jinkela_wire_177;
    wire jinkela_wire_178;
    wire jinkela_wire_179;
    wire jinkela_wire_180;
    wire jinkela_wire_181;
    wire jinkela_wire_182;
    wire jinkela_wire_183;
    wire jinkela_wire_184;
    wire jinkela_wire_185;
    wire jinkela_wire_186;
    wire jinkela_wire_187;
    wire jinkela_wire_188;
    wire jinkela_wire_189;
    wire jinkela_wire_190;
    wire jinkela_wire_191;
    wire jinkela_wire_192;
    wire jinkela_wire_193;
    wire jinkela_wire_194;
    wire jinkela_wire_195;
    wire jinkela_wire_196;
    wire jinkela_wire_197;
    wire jinkela_wire_198;
    wire jinkela_wire_199;
    wire jinkela_wire_200;
    wire jinkela_wire_201;
    wire jinkela_wire_202;
    wire jinkela_wire_203;
    wire jinkela_wire_204;
    wire jinkela_wire_205;
    wire jinkela_wire_206;
    wire jinkela_wire_207;
    wire jinkela_wire_208;
    input in_15_;
    input in_0_;
    input in_4_;
    input in_29_;
    input in_38_;
    input in_53_;
    input in_42_;
    input in_11_;
    input in_59_;
    input in_48_;
    input in_54_;
    input in_16_;
    input in_43_;
    input in_37_;
    input in_61_;
    input in_14_;
    input in_62_;
    input in_60_;
    input in_40_;
    input in_5_;
    input in_28_;
    input in_7_;
    input in_6_;
    input in_34_;
    input in_57_;
    input in_3_;
    input in_56_;
    input in_45_;
    input in_10_;
    input in_27_;
    input in_21_;
    input in_25_;
    input in_22_;
    input in_12_;
    input in_58_;
    input in_36_;
    input in_51_;
    input in_18_;
    input in_9_;
    input in_39_;
    input in_24_;
    input in_26_;
    input in_8_;
    input in_41_;
    input in_55_;
    input in_2_;
    input in_49_;
    input in_19_;
    input in_35_;
    input in_50_;
    input in_32_;
    input in_30_;
    input in_33_;
    input in_17_;
    input in_31_;
    input in_44_;
    input in_1_;
    input in_23_;
    input in_52_;
    input in_20_;
    input in_46_;
    input in_13_;
    input in_63_;
    input in_47_;
    output out_1_;
    output out_3_;
    output out_6_;
    output out_2_;
    output out_0_;
    output out_4_;
    output out_5_;

    and_bi _099_ (
        .b(jinkela_wire_73),
        .a(jinkela_wire_65),
        .c(out_1_)
    );

    or_bb _183_ (
        .b(jinkela_wire_166),
        .a(jinkela_wire_145),
        .c(jinkela_wire_160)
    );

    and_bi _225_ (
        .b(jinkela_wire_55),
        .a(jinkela_wire_43),
        .c(jinkela_wire_125)
    );

    maj_bbi _270_ (
        .b(jinkela_wire_151),
        .a(jinkela_wire_188),
        .c(jinkela_wire_46),
        .d(jinkela_wire_13)
    );

    maj_bii _100_ (
        .b(jinkela_wire_20),
        .a(jinkela_wire_94),
        .c(jinkela_wire_70),
        .d(jinkela_wire_163)
    );

    and_bi _184_ (
        .b(jinkela_wire_63),
        .a(jinkela_wire_160),
        .c(jinkela_wire_186)
    );

    and_bi _226_ (
        .b(jinkela_wire_125),
        .a(jinkela_wire_191),
        .c(jinkela_wire_20)
    );

    and_bb _271_ (
        .b(jinkela_wire_146),
        .a(jinkela_wire_13),
        .c(jinkela_wire_9)
    );

    or_ii _101_ (
        .b(jinkela_wire_114),
        .a(jinkela_wire_92),
        .c(jinkela_wire_30)
    );

    and_bb _185_ (
        .b(jinkela_wire_66),
        .a(jinkela_wire_63),
        .c(jinkela_wire_201)
    );

    maj_bii _227_ (
        .b(jinkela_wire_95),
        .a(jinkela_wire_43),
        .c(jinkela_wire_11),
        .d(jinkela_wire_135)
    );

    or_bb _272_ (
        .b(jinkela_wire_146),
        .a(jinkela_wire_13),
        .c(jinkela_wire_80)
    );

    and_ii _102_ (
        .b(jinkela_wire_114),
        .a(jinkela_wire_92),
        .c(jinkela_wire_78)
    );

    or_bb _186_ (
        .b(jinkela_wire_66),
        .a(jinkela_wire_63),
        .c(jinkela_wire_27)
    );

    or_ii _228_ (
        .b(jinkela_wire_48),
        .a(jinkela_wire_77),
        .c(jinkela_wire_158)
    );

    and_bi _273_ (
        .b(jinkela_wire_9),
        .a(jinkela_wire_80),
        .c(jinkela_wire_11)
    );

    and_bi _103_ (
        .b(jinkela_wire_78),
        .a(jinkela_wire_30),
        .c(jinkela_wire_10)
    );

    and_bi _187_ (
        .b(jinkela_wire_201),
        .a(jinkela_wire_27),
        .c(jinkela_wire_204)
    );

    and_ii _229_ (
        .b(jinkela_wire_48),
        .a(jinkela_wire_77),
        .c(jinkela_wire_162)
    );

    and_bb _274_ (
        .b(jinkela_wire_177),
        .a(jinkela_wire_9),
        .c(jinkela_wire_111)
    );

    or_bi _104_ (
        .b(jinkela_wire_10),
        .a(jinkela_wire_163),
        .c(jinkela_wire_33)
    );

    and_bb _188_ (
        .b(jinkela_wire_84),
        .a(jinkela_wire_201),
        .c(jinkela_wire_90)
    );

    and_bi _230_ (
        .b(jinkela_wire_162),
        .a(jinkela_wire_158),
        .c(jinkela_wire_183)
    );

    or_bb _275_ (
        .b(jinkela_wire_177),
        .a(jinkela_wire_9),
        .c(jinkela_wire_124)
    );

    and_bi _105_ (
        .b(jinkela_wire_10),
        .a(jinkela_wire_163),
        .c(jinkela_wire_82)
    );

    or_bb _189_ (
        .b(jinkela_wire_84),
        .a(jinkela_wire_201),
        .c(jinkela_wire_89)
    );

    or_bi _231_ (
        .b(jinkela_wire_183),
        .a(jinkela_wire_135),
        .c(jinkela_wire_148)
    );

    and_bi _276_ (
        .b(jinkela_wire_111),
        .a(jinkela_wire_124),
        .c(jinkela_wire_48)
    );

    and_bi _106_ (
        .b(jinkela_wire_82),
        .a(jinkela_wire_33),
        .c(out_2_)
    );

    and_bi _190_ (
        .b(jinkela_wire_90),
        .a(jinkela_wire_89),
        .c(jinkela_wire_187)
    );

    and_bi _232_ (
        .b(jinkela_wire_183),
        .a(jinkela_wire_135),
        .c(jinkela_wire_181)
    );

    and_bb _277_ (
        .b(jinkela_wire_60),
        .a(jinkela_wire_111),
        .c(jinkela_wire_32)
    );

    maj_bii _107_ (
        .b(jinkela_wire_92),
        .a(jinkela_wire_163),
        .c(jinkela_wire_114),
        .d(jinkela_wire_156)
    );

    or_bb _191_ (
        .b(in_32_),
        .a(in_33_),
        .c(jinkela_wire_68)
    );

    and_bi _233_ (
        .b(jinkela_wire_181),
        .a(jinkela_wire_148),
        .c(jinkela_wire_92)
    );

    or_bb _278_ (
        .b(jinkela_wire_60),
        .a(jinkela_wire_111),
        .c(jinkela_wire_21)
    );

    or_ii _108_ (
        .b(jinkela_wire_81),
        .a(jinkela_wire_42),
        .c(jinkela_wire_40)
    );

    and_bb _192_ (
        .b(in_34_),
        .a(in_35_),
        .c(jinkela_wire_140)
    );

    maj_bii _234_ (
        .b(jinkela_wire_77),
        .a(jinkela_wire_135),
        .c(jinkela_wire_48),
        .d(jinkela_wire_87)
    );

    and_bi _279_ (
        .b(jinkela_wire_32),
        .a(jinkela_wire_21),
        .c(jinkela_wire_98)
    );

    and_ii _109_ (
        .b(jinkela_wire_81),
        .a(jinkela_wire_42),
        .c(jinkela_wire_7)
    );

    or_bb _193_ (
        .b(in_36_),
        .a(in_37_),
        .c(jinkela_wire_28)
    );

    or_ii _235_ (
        .b(jinkela_wire_98),
        .a(jinkela_wire_123),
        .c(jinkela_wire_149)
    );

    or_bb _280_ (
        .b(in_0_),
        .a(in_1_),
        .c(jinkela_wire_192)
    );

    and_bi _110_ (
        .b(jinkela_wire_7),
        .a(jinkela_wire_40),
        .c(jinkela_wire_35)
    );

    and_bb _194_ (
        .b(in_38_),
        .a(in_39_),
        .c(jinkela_wire_45)
    );

    and_ii _236_ (
        .b(jinkela_wire_98),
        .a(jinkela_wire_123),
        .c(jinkela_wire_22)
    );

    and_bb _281_ (
        .b(in_2_),
        .a(in_3_),
        .c(jinkela_wire_88)
    );

    or_bi _111_ (
        .b(jinkela_wire_35),
        .a(jinkela_wire_156),
        .c(jinkela_wire_171)
    );

    or_bb _195_ (
        .b(in_40_),
        .a(in_41_),
        .c(jinkela_wire_6)
    );

    and_bi _237_ (
        .b(jinkela_wire_22),
        .a(jinkela_wire_149),
        .c(jinkela_wire_189)
    );

    or_bb _282_ (
        .b(in_4_),
        .a(in_5_),
        .c(jinkela_wire_34)
    );

    maj_bbi _181_ (
        .b(jinkela_wire_144),
        .a(jinkela_wire_19),
        .c(jinkela_wire_133),
        .d(jinkela_wire_145)
    );

    and_bi _112_ (
        .b(jinkela_wire_35),
        .a(jinkela_wire_156),
        .c(jinkela_wire_23)
    );

    and_bb _196_ (
        .b(in_42_),
        .a(in_43_),
        .c(jinkela_wire_105)
    );

    or_bi _238_ (
        .b(jinkela_wire_189),
        .a(jinkela_wire_87),
        .c(jinkela_wire_52)
    );

    and_bb _283_ (
        .b(in_6_),
        .a(in_7_),
        .c(jinkela_wire_157)
    );

    and_bi _113_ (
        .b(jinkela_wire_23),
        .a(jinkela_wire_171),
        .c(out_3_)
    );

    or_bb _197_ (
        .b(in_44_),
        .a(in_45_),
        .c(jinkela_wire_179)
    );

    and_bi _239_ (
        .b(jinkela_wire_189),
        .a(jinkela_wire_87),
        .c(jinkela_wire_12)
    );

    or_bb _284_ (
        .b(in_8_),
        .a(in_9_),
        .c(jinkela_wire_16)
    );

    maj_bii _114_ (
        .b(jinkela_wire_42),
        .a(jinkela_wire_156),
        .c(jinkela_wire_81),
        .d(jinkela_wire_128)
    );

    and_bb _198_ (
        .b(in_46_),
        .a(in_47_),
        .c(jinkela_wire_37)
    );

    and_bi _240_ (
        .b(jinkela_wire_12),
        .a(jinkela_wire_52),
        .c(jinkela_wire_42)
    );

    and_bb _285_ (
        .b(in_10_),
        .a(in_11_),
        .c(jinkela_wire_74)
    );

    or_ii _115_ (
        .b(jinkela_wire_180),
        .a(jinkela_wire_99),
        .c(jinkela_wire_153)
    );

    maj_bbb _199_ (
        .b(jinkela_wire_140),
        .a(jinkela_wire_28),
        .c(jinkela_wire_68),
        .d(jinkela_wire_101)
    );

    maj_bii _241_ (
        .b(jinkela_wire_123),
        .a(jinkela_wire_87),
        .c(jinkela_wire_98),
        .d(jinkela_wire_141)
    );

    or_bb _286_ (
        .b(in_12_),
        .a(in_13_),
        .c(jinkela_wire_93)
    );

    and_ii _116_ (
        .b(jinkela_wire_180),
        .a(jinkela_wire_99),
        .c(jinkela_wire_36)
    );

    maj_bbi _200_ (
        .b(jinkela_wire_68),
        .a(jinkela_wire_140),
        .c(jinkela_wire_28),
        .d(jinkela_wire_196)
    );

    or_ii _242_ (
        .b(jinkela_wire_32),
        .a(jinkela_wire_197),
        .c(jinkela_wire_117)
    );

    and_bb _287_ (
        .b(in_14_),
        .a(in_15_),
        .c(jinkela_wire_49)
    );

    and_bb _182_ (
        .b(jinkela_wire_166),
        .a(jinkela_wire_145),
        .c(jinkela_wire_63)
    );

    and_bi _117_ (
        .b(jinkela_wire_36),
        .a(jinkela_wire_153),
        .c(jinkela_wire_104)
    );

    maj_bbi _201_ (
        .b(jinkela_wire_28),
        .a(jinkela_wire_196),
        .c(jinkela_wire_101),
        .d(jinkela_wire_122)
    );

    and_ii _243_ (
        .b(jinkela_wire_32),
        .a(jinkela_wire_197),
        .c(jinkela_wire_0)
    );

    maj_bbb _288_ (
        .b(jinkela_wire_88),
        .a(jinkela_wire_34),
        .c(jinkela_wire_192),
        .d(jinkela_wire_53)
    );

    or_bi _118_ (
        .b(jinkela_wire_104),
        .a(jinkela_wire_128),
        .c(jinkela_wire_86)
    );

    maj_bbb _202_ (
        .b(jinkela_wire_159),
        .a(jinkela_wire_164),
        .c(jinkela_wire_101),
        .d(jinkela_wire_109)
    );

    and_bi _247_ (
        .b(jinkela_wire_150),
        .a(jinkela_wire_167),
        .c(jinkela_wire_99)
    );

    maj_bbi _289_ (
        .b(jinkela_wire_192),
        .a(jinkela_wire_88),
        .c(jinkela_wire_34),
        .d(jinkela_wire_155)
    );

    and_bi _119_ (
        .b(jinkela_wire_104),
        .a(jinkela_wire_128),
        .c(jinkela_wire_56)
    );

    maj_bbi _203_ (
        .b(jinkela_wire_101),
        .a(jinkela_wire_159),
        .c(jinkela_wire_164),
        .d(jinkela_wire_44)
    );

    and_ii _248_ (
        .b(1'b0),
        .a(1'b0),
        .c(jinkela_wire_5)
    );

    maj_bbi _290_ (
        .b(jinkela_wire_34),
        .a(jinkela_wire_155),
        .c(jinkela_wire_53),
        .d(jinkela_wire_29)
    );

    and_bi _120_ (
        .b(jinkela_wire_56),
        .a(jinkela_wire_86),
        .c(out_4_)
    );

    maj_bbi _204_ (
        .b(jinkela_wire_164),
        .a(jinkela_wire_44),
        .c(jinkela_wire_109),
        .d(jinkela_wire_112)
    );

    and_bi _249_ (
        .b(jinkela_wire_5),
        .a(jinkela_wire_43),
        .c(jinkela_wire_17)
    );

    maj_bbb _291_ (
        .b(jinkela_wire_147),
        .a(jinkela_wire_62),
        .c(jinkela_wire_53),
        .d(jinkela_wire_72)
    );

    maj_bii _121_ (
        .b(jinkela_wire_99),
        .a(jinkela_wire_128),
        .c(jinkela_wire_180),
        .d(jinkela_wire_75)
    );

    maj_bbb _205_ (
        .b(jinkela_wire_6),
        .a(jinkela_wire_105),
        .c(jinkela_wire_45),
        .d(jinkela_wire_159)
    );

    maj_bbi _250_ (
        .b(jinkela_wire_32),
        .a(jinkela_wire_197),
        .c(jinkela_wire_141),
        .d(jinkela_wire_107)
    );

    maj_bbi _292_ (
        .b(jinkela_wire_53),
        .a(jinkela_wire_147),
        .c(jinkela_wire_62),
        .d(jinkela_wire_184)
    );

    or_ii _122_ (
        .b(jinkela_wire_190),
        .a(jinkela_wire_107),
        .c(jinkela_wire_18)
    );

    maj_bbi _206_ (
        .b(jinkela_wire_45),
        .a(jinkela_wire_6),
        .c(jinkela_wire_105),
        .d(jinkela_wire_202)
    );

    or_bb _251_ (
        .b(in_16_),
        .a(in_17_),
        .c(jinkela_wire_121)
    );

    maj_bbi _293_ (
        .b(jinkela_wire_62),
        .a(jinkela_wire_184),
        .c(jinkela_wire_72),
        .d(jinkela_wire_8)
    );

    and_ii _123_ (
        .b(jinkela_wire_190),
        .a(jinkela_wire_107),
        .c(jinkela_wire_54)
    );

    maj_bbi _207_ (
        .b(jinkela_wire_105),
        .a(jinkela_wire_202),
        .c(jinkela_wire_159),
        .d(jinkela_wire_203)
    );

    and_bb _252_ (
        .b(in_18_),
        .a(in_19_),
        .c(jinkela_wire_207)
    );

    maj_bbb _294_ (
        .b(jinkela_wire_16),
        .a(jinkela_wire_74),
        .c(jinkela_wire_157),
        .d(jinkela_wire_147)
    );

    and_bi _124_ (
        .b(jinkela_wire_54),
        .a(jinkela_wire_18),
        .c(jinkela_wire_174)
    );

    maj_bbb _208_ (
        .b(jinkela_wire_203),
        .a(jinkela_wire_179),
        .c(jinkela_wire_122),
        .d(jinkela_wire_164)
    );

    or_bb _253_ (
        .b(in_20_),
        .a(in_21_),
        .c(jinkela_wire_50)
    );

    maj_bbi _295_ (
        .b(jinkela_wire_157),
        .a(jinkela_wire_16),
        .c(jinkela_wire_74),
        .d(jinkela_wire_208)
    );

    or_bi _125_ (
        .b(jinkela_wire_174),
        .a(jinkela_wire_75),
        .c(jinkela_wire_57)
    );

    maj_bbi _209_ (
        .b(jinkela_wire_122),
        .a(jinkela_wire_203),
        .c(jinkela_wire_179),
        .d(jinkela_wire_195)
    );

    and_bb _254_ (
        .b(in_22_),
        .a(in_23_),
        .c(jinkela_wire_106)
    );

    maj_bbi _296_ (
        .b(jinkela_wire_74),
        .a(jinkela_wire_208),
        .c(jinkela_wire_147),
        .d(jinkela_wire_64)
    );

    and_bi _126_ (
        .b(jinkela_wire_174),
        .a(jinkela_wire_75),
        .c(jinkela_wire_170)
    );

    maj_bbi _210_ (
        .b(jinkela_wire_179),
        .a(jinkela_wire_195),
        .c(jinkela_wire_164),
        .d(jinkela_wire_59)
    );

    or_bb _255_ (
        .b(in_24_),
        .a(in_25_),
        .c(jinkela_wire_58)
    );

    maj_bbb _297_ (
        .b(jinkela_wire_64),
        .a(jinkela_wire_93),
        .c(jinkela_wire_29),
        .d(jinkela_wire_62)
    );

    and_bi _127_ (
        .b(jinkela_wire_170),
        .a(jinkela_wire_57),
        .c(out_5_)
    );

    and_bb _211_ (
        .b(jinkela_wire_37),
        .a(jinkela_wire_59),
        .c(jinkela_wire_119)
    );

    and_bb _256_ (
        .b(in_26_),
        .a(in_27_),
        .c(jinkela_wire_205)
    );

    maj_bbi _298_ (
        .b(jinkela_wire_29),
        .a(jinkela_wire_64),
        .c(jinkela_wire_93),
        .d(jinkela_wire_173)
    );

    maj_bbi _128_ (
        .b(jinkela_wire_190),
        .a(jinkela_wire_107),
        .c(jinkela_wire_75),
        .d(out_6_)
    );

    or_bb _212_ (
        .b(jinkela_wire_37),
        .a(jinkela_wire_59),
        .c(jinkela_wire_199)
    );

    or_bb _257_ (
        .b(in_28_),
        .a(in_29_),
        .c(jinkela_wire_151)
    );

    maj_bbi _299_ (
        .b(jinkela_wire_93),
        .a(jinkela_wire_173),
        .c(jinkela_wire_62),
        .d(jinkela_wire_130)
    );

    and_ii _129_ (
        .b(jinkela_wire_193),
        .a(jinkela_wire_17),
        .c(jinkela_wire_161)
    );

    and_bi _213_ (
        .b(jinkela_wire_119),
        .a(jinkela_wire_199),
        .c(jinkela_wire_113)
    );

    and_bb _258_ (
        .b(in_30_),
        .a(in_31_),
        .c(jinkela_wire_146)
    );

    and_bb _300_ (
        .b(jinkela_wire_49),
        .a(jinkela_wire_130),
        .c(jinkela_wire_138)
    );

    and_bi _130_ (
        .b(jinkela_wire_161),
        .a(jinkela_wire_94),
        .c(out_0_)
    );

    and_bb _214_ (
        .b(jinkela_wire_112),
        .a(jinkela_wire_119),
        .c(jinkela_wire_137)
    );

    maj_bbb _259_ (
        .b(jinkela_wire_207),
        .a(jinkela_wire_50),
        .c(jinkela_wire_121),
        .d(jinkela_wire_136)
    );

    or_bb _301_ (
        .b(jinkela_wire_49),
        .a(jinkela_wire_130),
        .c(jinkela_wire_2)
    );

    or_ii _131_ (
        .b(1'b0),
        .a(1'b0),
        .c(jinkela_wire_142)
    );

    or_bb _215_ (
        .b(jinkela_wire_112),
        .a(jinkela_wire_119),
        .c(jinkela_wire_175)
    );

    maj_bbi _260_ (
        .b(jinkela_wire_121),
        .a(jinkela_wire_207),
        .c(jinkela_wire_50),
        .d(jinkela_wire_97)
    );

    and_bi _302_ (
        .b(jinkela_wire_138),
        .a(jinkela_wire_2),
        .c(jinkela_wire_95)
    );

    or_ii _132_ (
        .b(jinkela_wire_186),
        .a(jinkela_wire_113),
        .c(jinkela_wire_178)
    );

    and_bi _216_ (
        .b(jinkela_wire_137),
        .a(jinkela_wire_175),
        .c(jinkela_wire_143)
    );

    maj_bbi _261_ (
        .b(jinkela_wire_50),
        .a(jinkela_wire_97),
        .c(jinkela_wire_136),
        .d(jinkela_wire_61)
    );

    and_bb _303_ (
        .b(jinkela_wire_8),
        .a(jinkela_wire_138),
        .c(jinkela_wire_3)
    );

    and_ii _133_ (
        .b(jinkela_wire_186),
        .a(jinkela_wire_113),
        .c(jinkela_wire_79)
    );

    and_bb _217_ (
        .b(jinkela_wire_109),
        .a(jinkela_wire_137),
        .c(jinkela_wire_69)
    );

    maj_bbb _262_ (
        .b(jinkela_wire_110),
        .a(jinkela_wire_46),
        .c(jinkela_wire_136),
        .d(jinkela_wire_60)
    );

    or_bb _304_ (
        .b(jinkela_wire_8),
        .a(jinkela_wire_138),
        .c(jinkela_wire_1)
    );

    and_bi _134_ (
        .b(jinkela_wire_79),
        .a(jinkela_wire_178),
        .c(jinkela_wire_103)
    );

    or_bb _218_ (
        .b(jinkela_wire_109),
        .a(jinkela_wire_137),
        .c(jinkela_wire_127)
    );

    maj_bbi _263_ (
        .b(jinkela_wire_136),
        .a(jinkela_wire_110),
        .c(jinkela_wire_46),
        .d(jinkela_wire_132)
    );

    and_bi _305_ (
        .b(jinkela_wire_3),
        .a(jinkela_wire_1),
        .c(jinkela_wire_77)
    );

    or_bi _135_ (
        .b(jinkela_wire_103),
        .a(jinkela_wire_142),
        .c(jinkela_wire_118)
    );

    and_bi _219_ (
        .b(jinkela_wire_69),
        .a(jinkela_wire_127),
        .c(jinkela_wire_139)
    );

    maj_bbi _264_ (
        .b(jinkela_wire_46),
        .a(jinkela_wire_132),
        .c(jinkela_wire_60),
        .d(jinkela_wire_177)
    );

    and_bb _306_ (
        .b(jinkela_wire_72),
        .a(jinkela_wire_3),
        .c(jinkela_wire_197)
    );

    and_bi _136_ (
        .b(jinkela_wire_103),
        .a(jinkela_wire_142),
        .c(jinkela_wire_131)
    );

    or_ii _220_ (
        .b(1'b0),
        .a(1'b0),
        .c(jinkela_wire_43)
    );

    maj_bbb _265_ (
        .b(jinkela_wire_58),
        .a(jinkela_wire_205),
        .c(jinkela_wire_106),
        .d(jinkela_wire_110)
    );

    or_bb _307_ (
        .b(jinkela_wire_72),
        .a(jinkela_wire_3),
        .c(jinkela_wire_108)
    );

    and_bi _137_ (
        .b(jinkela_wire_131),
        .a(jinkela_wire_118),
        .c(jinkela_wire_70)
    );

    or_ii _221_ (
        .b(jinkela_wire_11),
        .a(jinkela_wire_95),
        .c(jinkela_wire_206)
    );

    maj_bbi _266_ (
        .b(jinkela_wire_106),
        .a(jinkela_wire_58),
        .c(jinkela_wire_205),
        .d(jinkela_wire_200)
    );

    and_bi _308_ (
        .b(jinkela_wire_197),
        .a(jinkela_wire_108),
        .c(jinkela_wire_123)
    );

    maj_bii _138_ (
        .b(jinkela_wire_113),
        .a(jinkela_wire_142),
        .c(jinkela_wire_186),
        .d(jinkela_wire_85)
    );

    and_ii _222_ (
        .b(jinkela_wire_11),
        .a(jinkela_wire_95),
        .c(jinkela_wire_172)
    );

    maj_bbi _267_ (
        .b(jinkela_wire_205),
        .a(jinkela_wire_200),
        .c(jinkela_wire_110),
        .d(jinkela_wire_116)
    );

    or_ii _139_ (
        .b(jinkela_wire_204),
        .a(jinkela_wire_143),
        .c(jinkela_wire_26)
    );

    and_bi _223_ (
        .b(jinkela_wire_172),
        .a(jinkela_wire_206),
        .c(jinkela_wire_55)
    );

    maj_bbb _268_ (
        .b(jinkela_wire_116),
        .a(jinkela_wire_151),
        .c(jinkela_wire_61),
        .d(jinkela_wire_46)
    );

    and_ii _140_ (
        .b(jinkela_wire_204),
        .a(jinkela_wire_143),
        .c(jinkela_wire_176)
    );

    or_bi _224_ (
        .b(jinkela_wire_55),
        .a(jinkela_wire_43),
        .c(jinkela_wire_191)
    );

    maj_bbi _269_ (
        .b(jinkela_wire_61),
        .a(jinkela_wire_116),
        .c(jinkela_wire_151),
        .d(jinkela_wire_188)
    );

    and_bi _141_ (
        .b(jinkela_wire_176),
        .a(jinkela_wire_26),
        .c(jinkela_wire_41)
    );

    or_bi _142_ (
        .b(jinkela_wire_41),
        .a(jinkela_wire_85),
        .c(jinkela_wire_134)
    );

    and_bi _143_ (
        .b(jinkela_wire_41),
        .a(jinkela_wire_85),
        .c(jinkela_wire_51)
    );

    and_bi _144_ (
        .b(jinkela_wire_51),
        .a(jinkela_wire_134),
        .c(jinkela_wire_114)
    );

    maj_bii _145_ (
        .b(jinkela_wire_143),
        .a(jinkela_wire_85),
        .c(jinkela_wire_204),
        .d(jinkela_wire_91)
    );

    or_ii _146_ (
        .b(jinkela_wire_187),
        .a(jinkela_wire_139),
        .c(jinkela_wire_115)
    );

    and_ii _147_ (
        .b(jinkela_wire_187),
        .a(jinkela_wire_139),
        .c(jinkela_wire_83)
    );

    and_bi _148_ (
        .b(jinkela_wire_83),
        .a(jinkela_wire_115),
        .c(jinkela_wire_152)
    );

    or_bi _149_ (
        .b(jinkela_wire_152),
        .a(jinkela_wire_91),
        .c(jinkela_wire_76)
    );

    or_bi _245_ (
        .b(jinkela_wire_126),
        .a(jinkela_wire_141),
        .c(jinkela_wire_167)
    );

    and_bi _150_ (
        .b(jinkela_wire_152),
        .a(jinkela_wire_91),
        .c(jinkela_wire_67)
    );

    and_bi _151_ (
        .b(jinkela_wire_67),
        .a(jinkela_wire_76),
        .c(jinkela_wire_81)
    );

    and_bi _246_ (
        .b(jinkela_wire_126),
        .a(jinkela_wire_141),
        .c(jinkela_wire_150)
    );

    maj_bii _152_ (
        .b(jinkela_wire_139),
        .a(jinkela_wire_91),
        .c(jinkela_wire_187),
        .d(jinkela_wire_165)
    );

    and_bi _244_ (
        .b(jinkela_wire_0),
        .a(jinkela_wire_117),
        .c(jinkela_wire_126)
    );

    or_ii _153_ (
        .b(jinkela_wire_90),
        .a(jinkela_wire_69),
        .c(jinkela_wire_38)
    );

    and_ii _154_ (
        .b(jinkela_wire_90),
        .a(jinkela_wire_69),
        .c(jinkela_wire_100)
    );

    and_bi _155_ (
        .b(jinkela_wire_100),
        .a(jinkela_wire_38),
        .c(jinkela_wire_194)
    );

    or_bi _156_ (
        .b(jinkela_wire_194),
        .a(jinkela_wire_165),
        .c(jinkela_wire_129)
    );

    and_bi _157_ (
        .b(jinkela_wire_194),
        .a(jinkela_wire_165),
        .c(jinkela_wire_47)
    );

    and_bi _158_ (
        .b(jinkela_wire_47),
        .a(jinkela_wire_129),
        .c(jinkela_wire_180)
    );

    and_ii _159_ (
        .b(1'b0),
        .a(1'b0),
        .c(jinkela_wire_25)
    );

    and_bi _160_ (
        .b(jinkela_wire_25),
        .a(jinkela_wire_142),
        .c(jinkela_wire_193)
    );

    maj_bbi _161_ (
        .b(jinkela_wire_90),
        .a(jinkela_wire_69),
        .c(jinkela_wire_165),
        .d(jinkela_wire_190)
    );

    or_bb _162_ (
        .b(in_48_),
        .a(in_49_),
        .c(jinkela_wire_168)
    );

    and_bb _163_ (
        .b(in_50_),
        .a(in_51_),
        .c(jinkela_wire_198)
    );

    or_bb _164_ (
        .b(in_52_),
        .a(in_53_),
        .c(jinkela_wire_102)
    );

    and_bb _165_ (
        .b(in_54_),
        .a(in_55_),
        .c(jinkela_wire_15)
    );

    or_bb _166_ (
        .b(in_56_),
        .a(in_57_),
        .c(jinkela_wire_4)
    );

    and_bb _167_ (
        .b(in_58_),
        .a(in_59_),
        .c(jinkela_wire_169)
    );

    or_bb _168_ (
        .b(in_60_),
        .a(in_61_),
        .c(jinkela_wire_144)
    );

    and_bb _169_ (
        .b(in_62_),
        .a(in_63_),
        .c(jinkela_wire_166)
    );

    maj_bbb _170_ (
        .b(jinkela_wire_198),
        .a(jinkela_wire_102),
        .c(jinkela_wire_168),
        .d(jinkela_wire_39)
    );

    maj_bbi _171_ (
        .b(jinkela_wire_168),
        .a(jinkela_wire_198),
        .c(jinkela_wire_102),
        .d(jinkela_wire_96)
    );

    maj_bbi _172_ (
        .b(jinkela_wire_102),
        .a(jinkela_wire_96),
        .c(jinkela_wire_39),
        .d(jinkela_wire_14)
    );

    maj_bbb _173_ (
        .b(jinkela_wire_154),
        .a(jinkela_wire_133),
        .c(jinkela_wire_39),
        .d(jinkela_wire_84)
    );

    maj_bbi _174_ (
        .b(jinkela_wire_39),
        .a(jinkela_wire_154),
        .c(jinkela_wire_133),
        .d(jinkela_wire_185)
    );

    maj_bbi _175_ (
        .b(jinkela_wire_133),
        .a(jinkela_wire_185),
        .c(jinkela_wire_84),
        .d(jinkela_wire_66)
    );

    maj_bbb _176_ (
        .b(jinkela_wire_4),
        .a(jinkela_wire_169),
        .c(jinkela_wire_15),
        .d(jinkela_wire_154)
    );

    maj_bbi _177_ (
        .b(jinkela_wire_15),
        .a(jinkela_wire_4),
        .c(jinkela_wire_169),
        .d(jinkela_wire_31)
    );

    maj_bbi _178_ (
        .b(jinkela_wire_169),
        .a(jinkela_wire_31),
        .c(jinkela_wire_154),
        .d(jinkela_wire_182)
    );

    and_bi _096_ (
        .b(jinkela_wire_24),
        .a(jinkela_wire_71),
        .c(jinkela_wire_120)
    );

    or_ii _094_ (
        .b(jinkela_wire_70),
        .a(jinkela_wire_20),
        .c(jinkela_wire_71)
    );

    maj_bbb _179_ (
        .b(jinkela_wire_182),
        .a(jinkela_wire_144),
        .c(jinkela_wire_14),
        .d(jinkela_wire_133)
    );

    and_ii _095_ (
        .b(jinkela_wire_70),
        .a(jinkela_wire_20),
        .c(jinkela_wire_24)
    );

    maj_bbi _180_ (
        .b(jinkela_wire_14),
        .a(jinkela_wire_182),
        .c(jinkela_wire_144),
        .d(jinkela_wire_19)
    );

    or_ii _093_ (
        .b(jinkela_wire_193),
        .a(jinkela_wire_17),
        .c(jinkela_wire_94)
    );

    or_bi _097_ (
        .b(jinkela_wire_120),
        .a(jinkela_wire_94),
        .c(jinkela_wire_65)
    );

    and_bi _098_ (
        .b(jinkela_wire_120),
        .a(jinkela_wire_94),
        .c(jinkela_wire_73)
    );

endmodule
