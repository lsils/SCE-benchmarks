module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 ;
  buffer buf_n354( .i (x13), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n105( .i (x3), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n132( .i (x4), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n25( .i (x0), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n288( .i (x10), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n53( .i (x1), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n309( .i (x11), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  assign n616 = n58 & n314 ;
  assign n617 = ( n31 & n294 ) | ( n31 & n616 ) | ( n294 & n616 ) ;
  assign n618 = ~n32 & n617 ;
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n260( .i (x9), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  assign n622 = ( n62 & n269 ) | ( n62 & ~n619 ) | ( n269 & ~n619 ) ;
  assign n623 = n115 & n622 ;
  assign n624 = ( n116 & n621 ) | ( n116 & ~n623 ) | ( n621 & ~n623 ) ;
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n382( .i (x14), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n426( .i (x16), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n447( .i (x17), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n473( .i (x18), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  assign n633 = ~n457 & n483 ;
  buffer buf_n634( .i (n633), .o (n634) );
  assign n645 = n438 & ~n634 ;
  buffer buf_n646( .i (n645), .o (n646) );
  assign n647 = ( n396 & ~n626 ) | ( n396 & n646 ) | ( ~n626 & n646 ) ;
  assign n648 = n627 & n647 ;
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n160( .i (x5), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n79( .i (x2), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  assign n651 = ~n34 & n88 ;
  assign n652 = n63 & n651 ;
  buffer buf_n653( .i (n652), .o (n653) );
  assign n666 = n117 & n653 ;
  assign n667 = ( n173 & n486 ) | ( n173 & n666 ) | ( n486 & n666 ) ;
  assign n668 = ~n487 & n667 ;
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  assign n672 = ( n95 & n176 ) | ( n95 & ~n669 ) | ( n176 & ~n669 ) ;
  assign n673 = n649 & n672 ;
  assign n674 = ( n650 & n671 ) | ( n650 & ~n673 ) | ( n671 & ~n673 ) ;
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n399( .i (x15), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  assign n677 = ~n419 & n675 ;
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  assign n678 = n67 & n119 ;
  assign n679 = ( n40 & n94 ) | ( n40 & n678 ) | ( n94 & n678 ) ;
  assign n680 = ~n41 & n679 ;
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  assign n681 = n459 | n485 ;
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  assign n690 = n680 & ~n685 ;
  assign n691 = ( n178 & n417 ) | ( n178 & n690 ) | ( n417 & n690 ) ;
  assign n692 = ~n418 & n691 ;
  assign n693 = n390 & n434 ;
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n270( .i (n269), .o (n270) );
  assign n704 = n169 | n482 ;
  assign n705 = n270 | n704 ;
  assign n706 = ~n89 & n115 ;
  assign n707 = ( n64 & ~n705 ) | ( n64 & n706 ) | ( ~n705 & n706 ) ;
  assign n708 = ~n65 & n707 ;
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  assign n712 = n297 & ~n482 ;
  assign n713 = n319 & n712 ;
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  assign n716 = n112 & n454 ;
  assign n717 = ( ~n87 & n168 ) | ( ~n87 & n716 ) | ( n168 & n716 ) ;
  assign n718 = n88 & n717 ;
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  assign n722 = ( n90 & n171 ) | ( n90 & ~n719 ) | ( n171 & ~n719 ) ;
  assign n723 = n714 & n722 ;
  assign n724 = ( n715 & n721 ) | ( n715 & ~n723 ) | ( n721 & ~n723 ) ;
  assign n725 = ( ~n39 & n709 ) | ( ~n39 & n724 ) | ( n709 & n724 ) ;
  assign n726 = n68 & ~n725 ;
  assign n727 = ( n69 & n711 ) | ( n69 & ~n726 ) | ( n711 & ~n726 ) ;
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  assign n730 = ~n417 & n728 ;
  assign n731 = ( ~n703 & n729 ) | ( ~n703 & n730 ) | ( n729 & n730 ) ;
  assign n732 = n692 | n731 ;
  assign n733 = ( n676 & ~n677 ) | ( n676 & n732 ) | ( ~n677 & n732 ) ;
  assign n734 = n154 & n733 ;
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n210( .i (x7), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  assign n737 = n68 & n175 ;
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  assign n742 = ( n99 & n642 ) | ( n99 & n741 ) | ( n642 & n741 ) ;
  assign n743 = ~n643 & n742 ;
  assign n744 = ( n47 & n232 ) | ( n47 & n743 ) | ( n232 & n743 ) ;
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  assign n745 = n70 | n277 ;
  assign n746 = n97 | n745 ;
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  assign n750 = n232 & ~n749 ;
  assign n751 = ( ~n48 & n744 ) | ( ~n48 & n750 ) | ( n744 & n750 ) ;
  assign n752 = n735 | n751 ;
  assign n753 = ( n130 & n736 ) | ( n130 & n752 ) | ( n736 & n752 ) ;
  assign n754 = n380 & ~n753 ;
  buffer buf_n500( .i (x19), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n551( .i (x21), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n526( .i (x20), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n576( .i (x22), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  assign n755 = ~n549 & n599 ;
  assign n756 = n575 & n755 ;
  assign n757 = ~n525 & n756 ;
  assign n758 = n380 | n757 ;
  assign n759 = ~n754 & n758 ;
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  assign n760 = ~n107 & n384 ;
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  assign n765 = n387 & ~n478 ;
  assign n766 = n111 & n765 ;
  assign n767 = ( n112 & n764 ) | ( n112 & ~n766 ) | ( n764 & ~n766 ) ;
  buffer buf_n768( .i (n767), .o (n768) );
  assign n773 = n435 & ~n768 ;
  assign n774 = n409 & n773 ;
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  assign n782 = n406 & n433 ;
  assign n783 = ( n390 & n434 ) | ( n390 & n782 ) | ( n434 & n782 ) ;
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  assign n796 = n387 & n404 ;
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  assign n803 = ~n115 & n784 ;
  assign n804 = ( n785 & n801 ) | ( n785 & n803 ) | ( n801 & n803 ) ;
  assign n805 = ( n459 & ~n775 ) | ( n459 & n804 ) | ( ~n775 & n804 ) ;
  assign n806 = ~n486 & n805 ;
  assign n807 = ( n487 & ~n777 ) | ( n487 & n806 ) | ( ~n777 & n806 ) ;
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  assign n810 = ( n148 & n176 ) | ( n148 & n808 ) | ( n176 & n808 ) ;
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  assign n811 = n116 & ~n221 ;
  buffer buf_n188( .i (x6), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  assign n812 = ~n116 & n199 ;
  assign n813 = ( n117 & ~n811 ) | ( n117 & n812 ) | ( ~n811 & n812 ) ;
  buffer buf_n814( .i (n813), .o (n814) );
  assign n822 = ( n461 & ~n487 ) | ( n461 & n814 ) | ( ~n487 & n814 ) ;
  assign n823 = ( n413 & ~n461 ) | ( n413 & n814 ) | ( ~n461 & n814 ) ;
  assign n824 = n822 & n823 ;
  assign n825 = n176 & n824 ;
  assign n826 = ( ~n809 & n810 ) | ( ~n809 & n825 ) | ( n810 & n825 ) ;
  assign n827 = n97 & ~n826 ;
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  assign n828 = ( n437 & n458 ) | ( n437 & ~n484 ) | ( n458 & ~n484 ) ;
  assign n829 = n394 & ~n828 ;
  assign n830 = ( ~n395 & n486 ) | ( ~n395 & n829 ) | ( n486 & n829 ) ;
  assign n831 = ( ~n323 & n413 ) | ( ~n323 & n830 ) | ( n413 & n830 ) ;
  buffer buf_n832( .i (n485), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  assign n834 = ( n323 & n413 ) | ( n323 & ~n833 ) | ( n413 & ~n833 ) ;
  assign n835 = ~n831 & n834 ;
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  assign n836 = n147 & n303 ;
  buffer buf_n837( .i (n175), .o (n837) );
  assign n838 = ( n835 & n836 ) | ( n835 & n837 ) | ( n836 & n837 ) ;
  assign n839 = ~n177 & n838 ;
  assign n840 = ~n97 & n839 ;
  assign n841 = ( n98 & ~n827 ) | ( n98 & n840 ) | ( ~n827 & n840 ) ;
  assign n842 = n73 & ~n841 ;
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n843( .i (n412), .o (n843) );
  assign n844 = ( n440 & ~n636 ) | ( n440 & n843 ) | ( ~n636 & n843 ) ;
  assign n845 = ( n637 & n699 ) | ( n637 & n844 ) | ( n699 & n844 ) ;
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  assign n848 = ~n173 & n301 ;
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  assign n852 = ( n149 & n846 ) | ( n149 & n851 ) | ( n846 & n851 ) ;
  assign n853 = ~n847 & n852 ;
  assign n854 = n98 & n853 ;
  assign n855 = n73 | n854 ;
  assign n856 = ~n842 & n855 ;
  assign n857 = ~n47 & n856 ;
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n860( .i (n114), .o (n860) );
  assign n861 = ~n270 & n860 ;
  buffer buf_n862( .i (n861), .o (n862) );
  assign n869 = ( ~n485 & n696 ) | ( ~n485 & n862 ) | ( n696 & n862 ) ;
  assign n870 = ~n697 & n869 ;
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  assign n874 = n386 & ~n761 ;
  buffer buf_n875( .i (n874), .o (n875) );
  assign n876 = ~n266 & n875 ;
  assign n877 = ( n31 & ~n763 ) | ( n31 & n875 ) | ( ~n763 & n875 ) ;
  assign n878 = ( ~n112 & n876 ) | ( ~n112 & n877 ) | ( n876 & n877 ) ;
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  assign n886 = ( ~n637 & n871 ) | ( ~n637 & n885 ) | ( n871 & n885 ) ;
  assign n887 = n442 & ~n886 ;
  assign n888 = ( n443 & n873 ) | ( n443 & ~n887 ) | ( n873 & ~n887 ) ;
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n179( .i (n178), .o (n179) );
  assign n891 = ( n179 & ~n418 ) | ( n179 & n889 ) | ( ~n418 & n889 ) ;
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  assign n892 = n39 & ~n788 ;
  assign n893 = ~n120 & n892 ;
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  assign n897 = n120 & ~n414 ;
  assign n898 = ( n276 & ~n489 ) | ( n276 & n897 ) | ( ~n489 & n897 ) ;
  assign n899 = ~n277 & n898 ;
  assign n900 = n895 | n899 ;
  assign n901 = ~n179 & n900 ;
  assign n902 = ( n890 & ~n891 ) | ( n890 & n901 ) | ( ~n891 & n901 ) ;
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  assign n905 = ( n101 & ~n154 ) | ( n101 & n903 ) | ( ~n154 & n903 ) ;
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n278( .i (n277), .o (n278) );
  assign n906 = ~n206 & n278 ;
  assign n907 = n38 & ~n118 ;
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  assign n913 = ( n207 & n906 ) | ( n207 & n912 ) | ( n906 & n912 ) ;
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  assign n914 = n228 & n868 ;
  buffer buf_n915( .i (n914), .o (n915) );
  assign n917 = n913 | n915 ;
  buffer buf_n918( .i (n917), .o (n918) );
  assign n920 = ~n101 & n918 ;
  assign n921 = ( n904 & ~n905 ) | ( n904 & n920 ) | ( ~n905 & n920 ) ;
  assign n922 = n858 | n921 ;
  assign n923 = ( ~n78 & n859 ) | ( ~n78 & n922 ) | ( n859 & n922 ) ;
  assign n924 = n380 & n923 ;
  assign n925 = ( ~n523 & n549 ) | ( ~n523 & n599 ) | ( n549 & n599 ) ;
  buffer buf_n926( .i (n925), .o (n926) );
  assign n927 = ( ~n520 & n546 ) | ( ~n520 & n571 ) | ( n546 & n571 ) ;
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  assign n932 = n926 & ~n931 ;
  buffer buf_n933( .i (n379), .o (n933) );
  assign n934 = n932 | n933 ;
  assign n935 = ( ~n381 & n924 ) | ( ~n381 & n934 ) | ( n924 & n934 ) ;
  assign n936 = ~n548 & n928 ;
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n600( .i (n599), .o (n600) );
  assign n939 = ( n575 & n600 ) | ( n575 & ~n937 ) | ( n600 & ~n937 ) ;
  assign n940 = ( n931 & n938 ) | ( n931 & ~n939 ) | ( n938 & ~n939 ) ;
  assign n941 = ~n933 & n940 ;
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n942( .i (n484), .o (n942) );
  assign n943 = n411 | n942 ;
  assign n944 = ( n697 & n832 ) | ( n697 & n943 ) | ( n832 & n943 ) ;
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  assign n950 = ( n122 & ~n277 ) | ( n122 & n894 ) | ( ~n277 & n894 ) ;
  assign n951 = n948 | n950 ;
  assign n952 = ( n896 & ~n949 ) | ( n896 & n951 ) | ( ~n949 & n951 ) ;
  assign n953 = n152 & n952 ;
  assign n954 = ~n181 & n953 ;
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n919( .i (n918), .o (n919) );
  assign n957 = n919 & ~n955 ;
  buffer buf_n102( .i (n101), .o (n102) );
  assign n958 = n76 | n102 ;
  assign n959 = ( n956 & n957 ) | ( n956 & ~n958 ) | ( n957 & ~n958 ) ;
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  assign n960 = ( ~n114 & n391 ) | ( ~n114 & n408 ) | ( n391 & n408 ) ;
  assign n961 = n436 & n960 ;
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  assign n964 = ( n172 & n459 ) | ( n172 & n962 ) | ( n459 & n962 ) ;
  assign n965 = n114 & ~n456 ;
  assign n966 = ( ~n483 & n800 ) | ( ~n483 & n965 ) | ( n800 & n965 ) ;
  assign n967 = ~n801 & n966 ;
  assign n968 = n172 & n967 ;
  assign n969 = ( ~n963 & n964 ) | ( ~n963 & n968 ) | ( n964 & n968 ) ;
  assign n970 = n67 & n969 ;
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  assign n973 = ~n63 & n170 ;
  buffer buf_n974( .i (n973), .o (n974) );
  assign n977 = n172 & ~n974 ;
  buffer buf_n978( .i (n977), .o (n978) );
  assign n979 = ~n682 & n978 ;
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  assign n980 = ( n302 & ~n976 ) | ( n302 & n978 ) | ( ~n976 & n978 ) ;
  assign n981 = ( ~n68 & n979 ) | ( ~n68 & n980 ) | ( n979 & n980 ) ;
  assign n982 = n971 | n981 ;
  assign n983 = ( ~n791 & n972 ) | ( ~n791 & n982 ) | ( n972 & n982 ) ;
  assign n984 = n150 & n983 ;
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n462( .i (n461), .o (n462) );
  assign n987 = ~n412 & n460 ;
  buffer buf_n988( .i (n987), .o (n988) );
  assign n995 = ( n462 & n637 ) | ( n462 & ~n988 ) | ( n637 & ~n988 ) ;
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  assign n999 = n178 & n818 ;
  assign n1000 = ~n998 & n999 ;
  assign n1001 = n985 | n1000 ;
  assign n1002 = ( n74 & n986 ) | ( n74 & n1001 ) | ( n986 & n1001 ) ;
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  assign n1005 = ( n48 & ~n102 ) | ( n48 & n1003 ) | ( ~n102 & n1003 ) ;
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n324( .i (n323), .o (n324) );
  assign n1006 = n324 & ~n945 ;
  assign n1007 = ( n304 & n837 ) | ( n304 & n1006 ) | ( n837 & n1006 ) ;
  assign n1008 = ~n177 & n1007 ;
  assign n1009 = n70 & n149 ;
  buffer buf_n1010( .i (n96), .o (n1010) );
  assign n1011 = ( n1008 & n1009 ) | ( n1008 & n1010 ) | ( n1009 & n1010 ) ;
  assign n1012 = ~n98 & n1011 ;
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  assign n1016 = ~n48 & n1015 ;
  assign n1017 = ( n1004 & ~n1005 ) | ( n1004 & n1016 ) | ( ~n1005 & n1016 ) ;
  assign n1018 = n959 | n1017 ;
  assign n1019 = n933 & n1018 ;
  assign n1020 = n941 | n1019 ;
  buffer buf_n550( .i (n549), .o (n550) );
  assign n1021 = ( n550 & n575 ) | ( n550 & n600 ) | ( n575 & n600 ) ;
  assign n1022 = ~n926 & n1021 ;
  assign n1023 = n933 | n1022 ;
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n233( .i (x8), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  assign n1024 = n126 & n330 ;
  assign n1025 = n255 & n1024 ;
  assign n1026 = n44 & n72 ;
  buffer buf_n1027( .i (n1026), .o (n1027) );
  assign n1030 = n46 & ~n1027 ;
  buffer buf_n1031( .i (n1030), .o (n1031) );
  assign n1032 = n1025 & n1031 ;
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  assign n1033 = ( n181 & n643 ) | ( n181 & n821 ) | ( n643 & n821 ) ;
  assign n1034 = n117 | n394 ;
  assign n1035 = n411 | n634 ;
  assign n1036 = ( ~n118 & n1034 ) | ( ~n118 & n1035 ) | ( n1034 & n1035 ) ;
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n397( .i (n396), .o (n397) );
  assign n1040 = ( ~n120 & n397 ) | ( ~n120 & n1037 ) | ( n397 & n1037 ) ;
  assign n1041 = ~n684 & n1040 ;
  assign n1042 = ( n685 & n1039 ) | ( n685 & n1041 ) | ( n1039 & n1041 ) ;
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  assign n1045 = n443 | n996 ;
  assign n1046 = ( n150 & n781 ) | ( n150 & ~n1045 ) | ( n781 & ~n1045 ) ;
  assign n1047 = n1043 & n1046 ;
  assign n1048 = ( n152 & ~n1044 ) | ( n152 & n1047 ) | ( ~n1044 & n1047 ) ;
  assign n1049 = n181 & n1048 ;
  assign n1050 = ( ~n644 & n1033 ) | ( ~n644 & n1049 ) | ( n1033 & n1049 ) ;
  assign n1051 = ( ~n1029 & n1031 ) | ( ~n1029 & n1050 ) | ( n1031 & n1050 ) ;
  assign n1052 = ( n77 & n1032 ) | ( n77 & n1051 ) | ( n1032 & n1051 ) ;
  assign n1053 = n104 & n1052 ;
  buffer buf_n1054( .i (n379), .o (n1054) );
  assign n1055 = ~n1053 & n1054 ;
  assign n1056 = n1023 & ~n1055 ;
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  assign n1057 = ( n415 & n442 ) | ( n415 & n463 ) | ( n442 & n463 ) ;
  assign n1058 = ( ~n464 & n701 ) | ( ~n464 & n1057 ) | ( n701 & n1057 ) ;
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  assign n1063 = ~n73 & n308 ;
  assign n1064 = ( n100 & n1061 ) | ( n100 & n1063 ) | ( n1061 & n1063 ) ;
  assign n1065 = ~n1062 & n1064 ;
  buffer buf_n1066( .i (n47), .o (n1066) );
  assign n1067 = ( n377 & n1065 ) | ( n377 & n1066 ) | ( n1065 & n1066 ) ;
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  assign n1068 = ( n419 & ~n493 ) | ( n419 & n632 ) | ( ~n493 & n632 ) ;
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n444( .i (n443), .o (n444) );
  assign n1069 = ~n397 & n441 ;
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  assign n1072 = ( n444 & n491 ) | ( n444 & ~n1071 ) | ( n491 & ~n1071 ) ;
  assign n1073 = ( ~n444 & n465 ) | ( ~n444 & n1071 ) | ( n465 & n1071 ) ;
  assign n1074 = ( ~n466 & n1072 ) | ( ~n466 & n1073 ) | ( n1072 & n1073 ) ;
  assign n1075 = ( n419 & ~n632 ) | ( n419 & n1074 ) | ( ~n632 & n1074 ) ;
  assign n1076 = n1068 & ~n1075 ;
  assign n1077 = n43 & ~n71 ;
  assign n1078 = ( ~n124 & n1059 ) | ( ~n124 & n1077 ) | ( n1059 & n1077 ) ;
  assign n1079 = ~n1060 & n1078 ;
  assign n1080 = ~n100 & n1079 ;
  assign n1081 = ( ~n101 & n1076 ) | ( ~n101 & n1080 ) | ( n1076 & n1080 ) ;
  assign n1082 = n377 & n1081 ;
  assign n1083 = ( ~n49 & n1067 ) | ( ~n49 & n1082 ) | ( n1067 & n1082 ) ;
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n331( .i (x12), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  assign n1086 = n353 & n495 ;
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  assign n1091 = ( n157 & ~n185 ) | ( n157 & n1088 ) | ( ~n185 & n1088 ) ;
  assign n1092 = n1084 & ~n1091 ;
  assign n1093 = ( n1085 & n1090 ) | ( n1085 & ~n1092 ) | ( n1090 & ~n1092 ) ;
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  assign n1094 = n440 | n833 ;
  assign n1095 = ( n441 & ~n462 ) | ( n441 & n1094 ) | ( ~n462 & n1094 ) ;
  buffer buf_n1096( .i (n1095), .o (n1096) );
  assign n1097 = ( n122 & ~n1070 ) | ( n122 & n1096 ) | ( ~n1070 & n1096 ) ;
  buffer buf_n398( .i (n397), .o (n398) );
  assign n1098 = ( n398 & n489 ) | ( n398 & n638 ) | ( n489 & n638 ) ;
  assign n1099 = ( ~n122 & n1096 ) | ( ~n122 & n1098 ) | ( n1096 & n1098 ) ;
  assign n1100 = n1097 & n1099 ;
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  assign n1103 = ( n99 & n741 ) | ( n99 & n1101 ) | ( n741 & n1101 ) ;
  assign n1104 = ~n1102 & n1103 ;
  buffer buf_n1105( .i (n46), .o (n1105) );
  assign n1106 = ( n421 & n1104 ) | ( n421 & n1105 ) | ( n1104 & n1105 ) ;
  assign n1107 = ~n88 & n879 ;
  assign n1108 = ~n63 & n1107 ;
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n87), .o (n1112) );
  assign n1113 = ~n62 & n1112 ;
  assign n1114 = n62 & n391 ;
  assign n1115 = ~n86 & n316 ;
  buffer buf_n1116( .i (n1115), .o (n1116) );
  assign n1120 = n391 & ~n1116 ;
  assign n1121 = ( n1113 & n1114 ) | ( n1113 & ~n1120 ) | ( n1114 & ~n1120 ) ;
  buffer buf_n1122( .i (n1121), .o (n1122) );
  assign n1125 = ( ~n37 & n1109 ) | ( ~n37 & n1122 ) | ( n1109 & n1122 ) ;
  assign n1126 = n301 & ~n1125 ;
  assign n1127 = ( n302 & n1111 ) | ( n302 & ~n1126 ) | ( n1111 & ~n1126 ) ;
  buffer buf_n1128( .i (n636), .o (n1128) );
  assign n1129 = n1127 & ~n1128 ;
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  assign n1135 = ( n180 & ~n446 ) | ( n180 & n1133 ) | ( ~n446 & n1133 ) ;
  buffer buf_n1136( .i (n67), .o (n1136) );
  assign n1137 = ( ~n441 & n908 ) | ( ~n441 & n1136 ) | ( n908 & n1136 ) ;
  assign n1138 = ~n69 & n1137 ;
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  assign n1141 = ~n489 & n628 ;
  assign n1142 = ~n701 & n1141 ;
  assign n1143 = n92 & ~n439 ;
  assign n1144 = n302 & n1143 ;
  assign n1145 = ~n40 & n1144 ;
  assign n1146 = ~n69 & n1145 ;
  buffer buf_n1147( .i (n1146), .o (n1147) );
  assign n1148 = ( ~n1139 & n1142 ) | ( ~n1139 & n1147 ) | ( n1142 & n1147 ) ;
  assign n1149 = n1010 & ~n1147 ;
  assign n1150 = ( n1140 & n1148 ) | ( n1140 & ~n1149 ) | ( n1148 & ~n1149 ) ;
  assign n1151 = ~n180 & n1150 ;
  assign n1152 = ( n1134 & ~n1135 ) | ( n1134 & n1151 ) | ( ~n1135 & n1151 ) ;
  assign n1153 = n421 & n1152 ;
  assign n1154 = ( ~n1066 & n1106 ) | ( ~n1066 & n1153 ) | ( n1106 & n1153 ) ;
  assign n1155 = ( n156 & n1087 ) | ( n156 & n1154 ) | ( n1087 & n1154 ) ;
  assign n1156 = n379 & ~n1155 ;
  assign n1157 = ( n1054 & n1089 ) | ( n1054 & ~n1156 ) | ( n1089 & ~n1156 ) ;
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  assign n1159 = ( ~n123 & n206 ) | ( ~n123 & n251 ) | ( n206 & n251 ) ;
  assign n1160 = ~n279 & n1159 ;
  assign n1161 = ( ~n125 & n280 ) | ( ~n125 & n1160 ) | ( n280 & n1160 ) ;
  assign n1162 = n45 | n915 ;
  assign n1163 = ( n916 & n1161 ) | ( n916 & n1162 ) | ( n1161 & n1162 ) ;
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  assign n1166 = ~n75 & n376 ;
  assign n1167 = ( n102 & n1164 ) | ( n102 & ~n1166 ) | ( n1164 & ~n1166 ) ;
  assign n1168 = n1165 & ~n1167 ;
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  assign n1172 = ( n445 & n687 ) | ( n445 & n703 ) | ( n687 & n703 ) ;
  assign n1173 = ( n437 & n458 ) | ( n437 & n484 ) | ( n458 & n484 ) ;
  assign n1174 = n394 & ~n1173 ;
  assign n1175 = ( n395 & n832 ) | ( n395 & ~n1174 ) | ( n832 & ~n1174 ) ;
  buffer buf_n1176( .i (n1175), .o (n1176) );
  assign n1179 = n275 | n1176 ;
  assign n1180 = ( n95 & n121 ) | ( n95 & ~n1179 ) | ( n121 & ~n1179 ) ;
  assign n1181 = ~n96 & n1180 ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  assign n1184 = n38 & n92 ;
  buffer buf_n1185( .i (n1184), .o (n1185) );
  assign n1188 = n94 & ~n1185 ;
  buffer buf_n1189( .i (n1188), .o (n1189) );
  assign n1190 = n305 & n1189 ;
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1191( .i (n121), .o (n1191) );
  assign n1192 = ( n1187 & ~n1189 ) | ( n1187 & n1191 ) | ( ~n1189 & n1191 ) ;
  assign n1193 = ( n43 & n1190 ) | ( n43 & ~n1192 ) | ( n1190 & ~n1192 ) ;
  assign n1194 = n1182 | n1193 ;
  assign n1195 = ( ~n1172 & n1183 ) | ( ~n1172 & n1194 ) | ( n1183 & n1194 ) ;
  assign n1196 = n74 | n1195 ;
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  assign n1197 = n326 & ~n1178 ;
  assign n1198 = ( n306 & n1010 ) | ( n306 & n1197 ) | ( n1010 & n1197 ) ;
  buffer buf_n1199( .i (n1010), .o (n1199) );
  assign n1200 = n1198 & ~n1199 ;
  assign n1201 = ~n45 & n1200 ;
  assign n1202 = n74 & ~n1201 ;
  assign n1203 = n1196 & ~n1202 ;
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n422( .i (n421), .o (n422) );
  assign n1206 = ~n183 & n422 ;
  assign n1207 = ( n378 & ~n1204 ) | ( n378 & n1206 ) | ( ~n1204 & n1206 ) ;
  assign n1208 = n1205 & n1207 ;
  assign n1209 = n1089 | n1208 ;
  assign n1210 = ( n159 & n1090 ) | ( n159 & n1209 ) | ( n1090 & n1209 ) ;
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  assign n1211 = ( ~n204 & n790 ) | ( ~n204 & n837 ) | ( n790 & n837 ) ;
  assign n1212 = n149 & n1211 ;
  assign n1213 = ( n150 & n206 ) | ( n150 & ~n1212 ) | ( n206 & ~n1212 ) ;
  assign n1214 = ( n72 & ~n1199 ) | ( n72 & n1213 ) | ( ~n1199 & n1213 ) ;
  assign n1215 = n252 & ~n1199 ;
  buffer buf_n1216( .i (n72), .o (n1216) );
  assign n1217 = ( n1214 & n1215 ) | ( n1214 & ~n1216 ) | ( n1215 & ~n1216 ) ;
  assign n1218 = n46 & n1217 ;
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  assign n1221 = n209 & ~n689 ;
  assign n1222 = n182 & n1221 ;
  assign n1223 = n1219 | n1222 ;
  assign n1224 = ( n665 & n1220 ) | ( n665 & n1223 ) | ( n1220 & n1223 ) ;
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n131( .i (n130), .o (n131) );
  assign n1227 = ( n131 & ~n1054 ) | ( n131 & n1225 ) | ( ~n1054 & n1225 ) ;
  buffer buf_n50( .i (n49), .o (n50) );
  assign n1228 = n177 & ~n685 ;
  assign n1229 = n659 & n1228 ;
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  assign n1232 = ~n410 & n695 ;
  assign n1233 = n171 | n271 ;
  assign n1234 = ( n696 & ~n1232 ) | ( n696 & n1233 ) | ( ~n1232 & n1233 ) ;
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  assign n1237 = n167 & ~n797 ;
  assign n1238 = ~n455 & n1237 ;
  assign n1239 = n1112 & n1238 ;
  buffer buf_n1240( .i (n61), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  assign n1242 = ( n35 & n1239 ) | ( n35 & n1241 ) | ( n1239 & n1241 ) ;
  assign n1243 = ~n36 & n1242 ;
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  assign n1247 = ( n66 & n92 ) | ( n66 & ~n1244 ) | ( n92 & ~n1244 ) ;
  assign n1248 = ~n1235 & n1247 ;
  assign n1249 = ( n1236 & ~n1246 ) | ( n1236 & n1248 ) | ( ~n1246 & n1248 ) ;
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  buffer buf_n1252( .i (n148), .o (n1252) );
  assign n1253 = ( ~n490 & n1250 ) | ( ~n490 & n1252 ) | ( n1250 & n1252 ) ;
  buffer buf_n601( .i (x23), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n802( .i (n801), .o (n802) );
  assign n1254 = n613 & ~n802 ;
  assign n1255 = n173 & n1254 ;
  assign n1256 = n93 & n1255 ;
  assign n1257 = ( n40 & n1136 ) | ( n40 & n1256 ) | ( n1136 & n1256 ) ;
  assign n1258 = ~n41 & n1257 ;
  assign n1259 = ~n490 & n1258 ;
  assign n1260 = ( ~n1251 & n1253 ) | ( ~n1251 & n1259 ) | ( n1253 & n1259 ) ;
  buffer buf_n1261( .i (n1260), .o (n1261) );
  assign n1262 = ( n747 & n1230 ) | ( n747 & ~n1261 ) | ( n1230 & ~n1261 ) ;
  assign n1263 = n230 | n1261 ;
  assign n1264 = ( n1231 & ~n1262 ) | ( n1231 & n1263 ) | ( ~n1262 & n1263 ) ;
  assign n1265 = n127 & n1264 ;
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  assign n1268 = ( n147 & n849 ) | ( n147 & n1136 ) | ( n849 & n1136 ) ;
  buffer buf_n1269( .i (n1136), .o (n1269) );
  assign n1270 = n1268 & ~n1269 ;
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n488), .o (n1274) );
  assign n1275 = ( n148 & n463 ) | ( n148 & ~n1274 ) | ( n463 & ~n1274 ) ;
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  assign n1276 = n615 & ~n833 ;
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  assign n1279 = ( ~n464 & n1275 ) | ( ~n464 & n1278 ) | ( n1275 & n1278 ) ;
  assign n1280 = ( n71 & n1271 ) | ( n71 & n1279 ) | ( n1271 & n1279 ) ;
  assign n1281 = n179 & ~n1280 ;
  assign n1282 = ( n180 & n1273 ) | ( n180 & ~n1281 ) | ( n1273 & ~n1281 ) ;
  assign n1283 = ( ~n795 & n1013 ) | ( ~n795 & n1282 ) | ( n1013 & n1282 ) ;
  buffer buf_n1284( .i (n100), .o (n1284) );
  assign n1285 = ~n1283 & n1284 ;
  buffer buf_n1286( .i (n1284), .o (n1286) );
  assign n1287 = ( n1015 & ~n1285 ) | ( n1015 & n1286 ) | ( ~n1285 & n1286 ) ;
  assign n1288 = n1266 | n1287 ;
  assign n1289 = ( ~n50 & n1267 ) | ( ~n50 & n1288 ) | ( n1267 & n1288 ) ;
  assign n1290 = n1054 & n1289 ;
  assign n1291 = ( n1226 & ~n1227 ) | ( n1226 & n1290 ) | ( ~n1227 & n1290 ) ;
  assign n1292 = ( n119 & n396 ) | ( n119 & n461 ) | ( n396 & n461 ) ;
  buffer buf_n1293( .i (n460), .o (n1293) );
  assign n1294 = ~n440 & n1293 ;
  assign n1295 = ( ~n397 & n1292 ) | ( ~n397 & n1294 ) | ( n1292 & n1294 ) ;
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  assign n1298 = ( n96 & n738 ) | ( n96 & ~n1296 ) | ( n738 & ~n1296 ) ;
  assign n1299 = n1297 & n1298 ;
  assign n1300 = ( n44 & n151 ) | ( n44 & n1299 ) | ( n151 & n1299 ) ;
  buffer buf_n1301( .i (n837), .o (n1301) );
  assign n1302 = ( n443 & n1130 ) | ( n443 & n1301 ) | ( n1130 & n1301 ) ;
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n1303( .i (n171), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  assign n1305 = ~n772 & n1304 ;
  assign n1306 = n93 & n1305 ;
  buffer buf_n1307( .i (n39), .o (n1307) );
  buffer buf_n1308( .i (n66), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  assign n1310 = ( n1306 & n1307 ) | ( n1306 & n1309 ) | ( n1307 & n1309 ) ;
  assign n1311 = ~n41 & n1310 ;
  buffer buf_n1312( .i (n442), .o (n1312) );
  assign n1313 = n1311 & n1312 ;
  assign n1314 = ( ~n178 & n1302 ) | ( ~n178 & n1313 ) | ( n1302 & n1313 ) ;
  assign n1315 = n151 & n1314 ;
  assign n1316 = ( ~n45 & n1300 ) | ( ~n45 & n1315 ) | ( n1300 & n1315 ) ;
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  assign n1320 = ( ~n227 & n464 ) | ( ~n227 & n1191 ) | ( n464 & n1191 ) ;
  assign n1321 = n700 & n1277 ;
  assign n1322 = n1191 & n1321 ;
  assign n1323 = ( n228 & n1320 ) | ( n228 & n1322 ) | ( n1320 & n1322 ) ;
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n205), .o (n1326) );
  assign n1327 = ( n123 & ~n465 ) | ( n123 & n1326 ) | ( ~n465 & n1326 ) ;
  assign n1328 = n1070 & n1278 ;
  assign n1329 = ~n123 & n1328 ;
  assign n1330 = ( n207 & ~n1327 ) | ( n207 & n1329 ) | ( ~n1327 & n1329 ) ;
  assign n1331 = ~n1324 & n1330 ;
  buffer buf_n1332( .i (n1301), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  assign n1335 = n99 & n1334 ;
  assign n1336 = ( n1325 & n1331 ) | ( n1325 & n1335 ) | ( n1331 & n1335 ) ;
  assign n1337 = ( ~n1105 & n1317 ) | ( ~n1105 & n1336 ) | ( n1317 & n1336 ) ;
  assign n1338 = n76 & ~n1337 ;
  assign n1339 = ( n77 & n1319 ) | ( n77 & ~n1338 ) | ( n1319 & ~n1338 ) ;
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n1342( .i (n378), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  assign n1344 = ( n425 & ~n1340 ) | ( n425 & n1343 ) | ( ~n1340 & n1343 ) ;
  assign n1345 = n145 & ~n697 ;
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  assign n1348 = n203 | n1346 ;
  assign n1349 = ( ~n121 & n1347 ) | ( ~n121 & n1348 ) | ( n1347 & n1348 ) ;
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1252), .o (n1351) );
  assign n1352 = ( n228 & n1350 ) | ( n228 & ~n1351 ) | ( n1350 & ~n1351 ) ;
  buffer buf_n1353( .i (n1191), .o (n1353) );
  assign n1354 = n1350 | n1353 ;
  assign n1355 = ( n151 & n1352 ) | ( n151 & n1354 ) | ( n1352 & n1354 ) ;
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n1358( .i (n1334), .o (n1358) );
  assign n1359 = ( n994 & ~n1356 ) | ( n994 & n1358 ) | ( ~n1356 & n1358 ) ;
  assign n1360 = n1357 & n1359 ;
  assign n1361 = n1286 & n1360 ;
  assign n1362 = ( n49 & n77 ) | ( n49 & n1361 ) | ( n77 & n1361 ) ;
  assign n1363 = ~n50 & n1362 ;
  assign n1364 = n1343 & n1363 ;
  assign n1365 = ( n1341 & n1344 ) | ( n1341 & n1364 ) | ( n1344 & n1364 ) ;
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  assign n1366 = ( n696 & ~n942 ) | ( n696 & n1119 ) | ( ~n942 & n1119 ) ;
  buffer buf_n1367( .i (n695), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  assign n1369 = n1366 & ~n1368 ;
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  assign n1372 = ( n414 & n1309 ) | ( n414 & ~n1370 ) | ( n1309 & ~n1370 ) ;
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  assign n1373 = n646 & n1124 ;
  assign n1374 = n414 & n1373 ;
  assign n1375 = ( n1371 & n1372 ) | ( n1371 & n1374 ) | ( n1372 & n1374 ) ;
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  assign n1378 = n323 & ~n843 ;
  assign n1379 = ~n488 & n1378 ;
  assign n1380 = n65 & n91 ;
  buffer buf_n1381( .i (n1380), .o (n1381) );
  assign n1384 = n1308 & ~n1381 ;
  buffer buf_n1385( .i (n1384), .o (n1385) );
  assign n1386 = n1379 & n1385 ;
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  assign n1387 = ( n790 & n1383 ) | ( n790 & ~n1385 ) | ( n1383 & ~n1385 ) ;
  buffer buf_n1388( .i (n95), .o (n1388) );
  assign n1389 = ( n1386 & ~n1387 ) | ( n1386 & n1388 ) | ( ~n1387 & n1388 ) ;
  assign n1390 = ~n1376 & n1389 ;
  assign n1391 = n306 & n372 ;
  assign n1392 = ( n1377 & n1390 ) | ( n1377 & n1391 ) | ( n1390 & n1391 ) ;
  assign n1393 = ~n1334 & n1392 ;
  buffer buf_n1394( .i (n44), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  assign n1396 = ( n153 & n1393 ) | ( n153 & n1395 ) | ( n1393 & n1395 ) ;
  assign n1397 = ~n1105 & n1396 ;
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  assign n1403 = n1066 & ~n1286 ;
  buffer buf_n1404( .i (n76), .o (n1404) );
  assign n1405 = ( ~n129 & n1403 ) | ( ~n129 & n1404 ) | ( n1403 & n1404 ) ;
  assign n1406 = ~n78 & n1405 ;
  assign n1407 = n1343 & n1406 ;
  assign n1408 = n287 & n1407 ;
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  assign n1409 = ( n103 & ~n378 ) | ( n103 & n1404 ) | ( ~n378 & n1404 ) ;
  buffer buf_n1410( .i (n377), .o (n1410) );
  assign n1411 = ( n103 & ~n129 ) | ( n103 & n1410 ) | ( ~n129 & n1410 ) ;
  assign n1412 = ~n1409 & n1411 ;
  assign n1413 = n259 & n1412 ;
  assign n1414 = n52 & n1413 ;
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  assign n1415 = n424 & ~n472 ;
  assign n1416 = ( n186 & ~n499 ) | ( n186 & n1415 ) | ( ~n499 & n1415 ) ;
  assign n1417 = ~n187 & n1416 ;
  assign y0 = n759 ;
  assign y1 = n935 ;
  assign y2 = n1020 ;
  assign y3 = n1056 ;
  assign y4 = n1093 ;
  assign y5 = n1158 ;
  assign y6 = n1171 ;
  assign y7 = n1210 ;
  assign y8 = n1291 ;
  assign y9 = n1365 ;
  assign y10 = n1402 ;
  assign y11 = n1408 ;
  assign y12 = n1414 ;
  assign y13 = n1417 ;
endmodule
