module sorter32(a_11_,a_18_,a_15_,a_3_,a_9_,a_6_,a_28_,a_7_,a_25_,a_29_,a_22_,a_26_,a_1_,a_8_,a_16_,a_10_,a_30_,a_12_,a_24_,a_5_,a_0_,a_17_,a_4_,a_14_,a_20_,a_27_,a_23_,a_13_,a_31_,a_2_,a_19_,a_21_,b_9_,b_1_,b_17_,b_11_,b_31_,b_26_,b_29_,b_24_,b_23_,b_8_,b_4_,b_25_,b_7_,b_5_,b_18_,b_12_,b_16_,b_22_,b_14_,b_20_,b_15_,b_3_,b_30_,b_27_,b_21_,b_19_,b_13_,b_6_,b_0_,b_10_,b_28_,b_2_);
    wire jinkela_wire_0;
    wire jinkela_wire_1;
    wire jinkela_wire_2;
    wire jinkela_wire_3;
    wire jinkela_wire_4;
    wire jinkela_wire_5;
    wire jinkela_wire_6;
    wire jinkela_wire_7;
    wire jinkela_wire_8;
    wire jinkela_wire_9;
    wire jinkela_wire_10;
    wire jinkela_wire_11;
    wire jinkela_wire_12;
    wire jinkela_wire_13;
    wire jinkela_wire_14;
    wire jinkela_wire_15;
    wire jinkela_wire_16;
    wire jinkela_wire_17;
    wire jinkela_wire_18;
    wire jinkela_wire_19;
    wire jinkela_wire_20;
    wire jinkela_wire_21;
    wire jinkela_wire_22;
    wire jinkela_wire_23;
    wire jinkela_wire_24;
    wire jinkela_wire_25;
    wire jinkela_wire_26;
    wire jinkela_wire_27;
    wire jinkela_wire_28;
    wire jinkela_wire_29;
    wire jinkela_wire_30;
    wire jinkela_wire_31;
    wire jinkela_wire_32;
    wire jinkela_wire_33;
    wire jinkela_wire_34;
    wire jinkela_wire_35;
    wire jinkela_wire_36;
    wire jinkela_wire_37;
    wire jinkela_wire_38;
    wire jinkela_wire_39;
    wire jinkela_wire_40;
    wire jinkela_wire_41;
    wire jinkela_wire_42;
    wire jinkela_wire_43;
    wire jinkela_wire_44;
    wire jinkela_wire_45;
    wire jinkela_wire_46;
    wire jinkela_wire_47;
    wire jinkela_wire_48;
    wire jinkela_wire_49;
    wire jinkela_wire_50;
    wire jinkela_wire_51;
    wire jinkela_wire_52;
    wire jinkela_wire_53;
    wire jinkela_wire_54;
    wire jinkela_wire_55;
    wire jinkela_wire_56;
    wire jinkela_wire_57;
    wire jinkela_wire_58;
    wire jinkela_wire_59;
    wire jinkela_wire_60;
    wire jinkela_wire_61;
    wire jinkela_wire_62;
    wire jinkela_wire_63;
    wire jinkela_wire_64;
    wire jinkela_wire_65;
    wire jinkela_wire_66;
    wire jinkela_wire_67;
    wire jinkela_wire_68;
    wire jinkela_wire_69;
    wire jinkela_wire_70;
    wire jinkela_wire_71;
    wire jinkela_wire_72;
    wire jinkela_wire_73;
    wire jinkela_wire_74;
    wire jinkela_wire_75;
    wire jinkela_wire_76;
    wire jinkela_wire_77;
    wire jinkela_wire_78;
    wire jinkela_wire_79;
    wire jinkela_wire_80;
    wire jinkela_wire_81;
    wire jinkela_wire_82;
    wire jinkela_wire_83;
    wire jinkela_wire_84;
    wire jinkela_wire_85;
    wire jinkela_wire_86;
    wire jinkela_wire_87;
    wire jinkela_wire_88;
    wire jinkela_wire_89;
    wire jinkela_wire_90;
    wire jinkela_wire_91;
    wire jinkela_wire_92;
    wire jinkela_wire_93;
    wire jinkela_wire_94;
    wire jinkela_wire_95;
    wire jinkela_wire_96;
    wire jinkela_wire_97;
    wire jinkela_wire_98;
    wire jinkela_wire_99;
    wire jinkela_wire_100;
    wire jinkela_wire_101;
    wire jinkela_wire_102;
    wire jinkela_wire_103;
    wire jinkela_wire_104;
    wire jinkela_wire_105;
    wire jinkela_wire_106;
    wire jinkela_wire_107;
    wire jinkela_wire_108;
    wire jinkela_wire_109;
    wire jinkela_wire_110;
    wire jinkela_wire_111;
    wire jinkela_wire_112;
    wire jinkela_wire_113;
    wire jinkela_wire_114;
    wire jinkela_wire_115;
    wire jinkela_wire_116;
    wire jinkela_wire_117;
    wire jinkela_wire_118;
    wire jinkela_wire_119;
    wire jinkela_wire_120;
    wire jinkela_wire_121;
    wire jinkela_wire_122;
    wire jinkela_wire_123;
    wire jinkela_wire_124;
    wire jinkela_wire_125;
    wire jinkela_wire_126;
    wire jinkela_wire_127;
    wire jinkela_wire_128;
    wire jinkela_wire_129;
    wire jinkela_wire_130;
    wire jinkela_wire_131;
    wire jinkela_wire_132;
    wire jinkela_wire_133;
    wire jinkela_wire_134;
    wire jinkela_wire_135;
    wire jinkela_wire_136;
    wire jinkela_wire_137;
    wire jinkela_wire_138;
    wire jinkela_wire_139;
    wire jinkela_wire_140;
    wire jinkela_wire_141;
    wire jinkela_wire_142;
    wire jinkela_wire_143;
    wire jinkela_wire_144;
    wire jinkela_wire_145;
    wire jinkela_wire_146;
    wire jinkela_wire_147;
    wire jinkela_wire_148;
    wire jinkela_wire_149;
    wire jinkela_wire_150;
    wire jinkela_wire_151;
    wire jinkela_wire_152;
    wire jinkela_wire_153;
    wire jinkela_wire_154;
    wire jinkela_wire_155;
    wire jinkela_wire_156;
    wire jinkela_wire_157;
    wire jinkela_wire_158;
    wire jinkela_wire_159;
    wire jinkela_wire_160;
    wire jinkela_wire_161;
    wire jinkela_wire_162;
    wire jinkela_wire_163;
    wire jinkela_wire_164;
    wire jinkela_wire_165;
    wire jinkela_wire_166;
    wire jinkela_wire_167;
    wire jinkela_wire_168;
    wire jinkela_wire_169;
    wire jinkela_wire_170;
    wire jinkela_wire_171;
    wire jinkela_wire_172;
    wire jinkela_wire_173;
    wire jinkela_wire_174;
    wire jinkela_wire_175;
    wire jinkela_wire_176;
    wire jinkela_wire_177;
    wire jinkela_wire_178;
    wire jinkela_wire_179;
    wire jinkela_wire_180;
    wire jinkela_wire_181;
    wire jinkela_wire_182;
    wire jinkela_wire_183;
    wire jinkela_wire_184;
    wire jinkela_wire_185;
    wire jinkela_wire_186;
    wire jinkela_wire_187;
    wire jinkela_wire_188;
    wire jinkela_wire_189;
    wire jinkela_wire_190;
    wire jinkela_wire_191;
    wire jinkela_wire_192;
    wire jinkela_wire_193;
    wire jinkela_wire_194;
    wire jinkela_wire_195;
    wire jinkela_wire_196;
    wire jinkela_wire_197;
    wire jinkela_wire_198;
    wire jinkela_wire_199;
    wire jinkela_wire_200;
    wire jinkela_wire_201;
    wire jinkela_wire_202;
    wire jinkela_wire_203;
    wire jinkela_wire_204;
    wire jinkela_wire_205;
    wire jinkela_wire_206;
    wire jinkela_wire_207;
    wire jinkela_wire_208;
    wire jinkela_wire_209;
    wire jinkela_wire_210;
    wire jinkela_wire_211;
    wire jinkela_wire_212;
    wire jinkela_wire_213;
    wire jinkela_wire_214;
    wire jinkela_wire_215;
    wire jinkela_wire_216;
    wire jinkela_wire_217;
    wire jinkela_wire_218;
    wire jinkela_wire_219;
    wire jinkela_wire_220;
    wire jinkela_wire_221;
    wire jinkela_wire_222;
    wire jinkela_wire_223;
    wire jinkela_wire_224;
    wire jinkela_wire_225;
    wire jinkela_wire_226;
    wire jinkela_wire_227;
    wire jinkela_wire_228;
    wire jinkela_wire_229;
    wire jinkela_wire_230;
    wire jinkela_wire_231;
    wire jinkela_wire_232;
    wire jinkela_wire_233;
    wire jinkela_wire_234;
    wire jinkela_wire_235;
    wire jinkela_wire_236;
    wire jinkela_wire_237;
    wire jinkela_wire_238;
    wire jinkela_wire_239;
    wire jinkela_wire_240;
    wire jinkela_wire_241;
    wire jinkela_wire_242;
    wire jinkela_wire_243;
    wire jinkela_wire_244;
    wire jinkela_wire_245;
    wire jinkela_wire_246;
    wire jinkela_wire_247;
    wire jinkela_wire_248;
    wire jinkela_wire_249;
    wire jinkela_wire_250;
    wire jinkela_wire_251;
    wire jinkela_wire_252;
    wire jinkela_wire_253;
    wire jinkela_wire_254;
    wire jinkela_wire_255;
    wire jinkela_wire_256;
    wire jinkela_wire_257;
    wire jinkela_wire_258;
    wire jinkela_wire_259;
    wire jinkela_wire_260;
    wire jinkela_wire_261;
    wire jinkela_wire_262;
    wire jinkela_wire_263;
    wire jinkela_wire_264;
    wire jinkela_wire_265;
    wire jinkela_wire_266;
    wire jinkela_wire_267;
    wire jinkela_wire_268;
    wire jinkela_wire_269;
    wire jinkela_wire_270;
    wire jinkela_wire_271;
    wire jinkela_wire_272;
    wire jinkela_wire_273;
    wire jinkela_wire_274;
    wire jinkela_wire_275;
    wire jinkela_wire_276;
    wire jinkela_wire_277;
    wire jinkela_wire_278;
    wire jinkela_wire_279;
    wire jinkela_wire_280;
    wire jinkela_wire_281;
    wire jinkela_wire_282;
    wire jinkela_wire_283;
    wire jinkela_wire_284;
    wire jinkela_wire_285;
    wire jinkela_wire_286;
    wire jinkela_wire_287;
    wire jinkela_wire_288;
    wire jinkela_wire_289;
    wire jinkela_wire_290;
    wire jinkela_wire_291;
    wire jinkela_wire_292;
    wire jinkela_wire_293;
    wire jinkela_wire_294;
    wire jinkela_wire_295;
    wire jinkela_wire_296;
    wire jinkela_wire_297;
    wire jinkela_wire_298;
    wire jinkela_wire_299;
    wire jinkela_wire_300;
    wire jinkela_wire_301;
    wire jinkela_wire_302;
    wire jinkela_wire_303;
    wire jinkela_wire_304;
    wire jinkela_wire_305;
    wire jinkela_wire_306;
    wire jinkela_wire_307;
    wire jinkela_wire_308;
    wire jinkela_wire_309;
    wire jinkela_wire_310;
    wire jinkela_wire_311;
    wire jinkela_wire_312;
    wire jinkela_wire_313;
    wire jinkela_wire_314;
    wire jinkela_wire_315;
    wire jinkela_wire_316;
    wire jinkela_wire_317;
    wire jinkela_wire_318;
    wire jinkela_wire_319;
    wire jinkela_wire_320;
    wire jinkela_wire_321;
    wire jinkela_wire_322;
    wire jinkela_wire_323;
    wire jinkela_wire_324;
    wire jinkela_wire_325;
    wire jinkela_wire_326;
    wire jinkela_wire_327;
    wire jinkela_wire_328;
    wire jinkela_wire_329;
    wire jinkela_wire_330;
    wire jinkela_wire_331;
    wire jinkela_wire_332;
    wire jinkela_wire_333;
    wire jinkela_wire_334;
    wire jinkela_wire_335;
    wire jinkela_wire_336;
    wire jinkela_wire_337;
    wire jinkela_wire_338;
    wire jinkela_wire_339;
    wire jinkela_wire_340;
    wire jinkela_wire_341;
    wire jinkela_wire_342;
    wire jinkela_wire_343;
    wire jinkela_wire_344;
    wire jinkela_wire_345;
    wire jinkela_wire_346;
    wire jinkela_wire_347;
    wire jinkela_wire_348;
    wire jinkela_wire_349;
    wire jinkela_wire_350;
    wire jinkela_wire_351;
    wire jinkela_wire_352;
    wire jinkela_wire_353;
    wire jinkela_wire_354;
    wire jinkela_wire_355;
    wire jinkela_wire_356;
    wire jinkela_wire_357;
    wire jinkela_wire_358;
    wire jinkela_wire_359;
    wire jinkela_wire_360;
    wire jinkela_wire_361;
    wire jinkela_wire_362;
    wire jinkela_wire_363;
    wire jinkela_wire_364;
    wire jinkela_wire_365;
    wire jinkela_wire_366;
    wire jinkela_wire_367;
    wire jinkela_wire_368;
    wire jinkela_wire_369;
    wire jinkela_wire_370;
    wire jinkela_wire_371;
    wire jinkela_wire_372;
    wire jinkela_wire_373;
    wire jinkela_wire_374;
    wire jinkela_wire_375;
    wire jinkela_wire_376;
    wire jinkela_wire_377;
    wire jinkela_wire_378;
    wire jinkela_wire_379;
    wire jinkela_wire_380;
    wire jinkela_wire_381;
    wire jinkela_wire_382;
    wire jinkela_wire_383;
    wire jinkela_wire_384;
    wire jinkela_wire_385;
    wire jinkela_wire_386;
    wire jinkela_wire_387;
    wire jinkela_wire_388;
    wire jinkela_wire_389;
    wire jinkela_wire_390;
    wire jinkela_wire_391;
    wire jinkela_wire_392;
    wire jinkela_wire_393;
    wire jinkela_wire_394;
    wire jinkela_wire_395;
    wire jinkela_wire_396;
    wire jinkela_wire_397;
    wire jinkela_wire_398;
    wire jinkela_wire_399;
    wire jinkela_wire_400;
    wire jinkela_wire_401;
    wire jinkela_wire_402;
    wire jinkela_wire_403;
    wire jinkela_wire_404;
    wire jinkela_wire_405;
    wire jinkela_wire_406;
    wire jinkela_wire_407;
    wire jinkela_wire_408;
    wire jinkela_wire_409;
    wire jinkela_wire_410;
    wire jinkela_wire_411;
    wire jinkela_wire_412;
    wire jinkela_wire_413;
    wire jinkela_wire_414;
    wire jinkela_wire_415;
    wire jinkela_wire_416;
    wire jinkela_wire_417;
    wire jinkela_wire_418;
    wire jinkela_wire_419;
    wire jinkela_wire_420;
    wire jinkela_wire_421;
    wire jinkela_wire_422;
    wire jinkela_wire_423;
    wire jinkela_wire_424;
    wire jinkela_wire_425;
    wire jinkela_wire_426;
    wire jinkela_wire_427;
    wire jinkela_wire_428;
    wire jinkela_wire_429;
    wire jinkela_wire_430;
    wire jinkela_wire_431;
    wire jinkela_wire_432;
    wire jinkela_wire_433;
    wire jinkela_wire_434;
    wire jinkela_wire_435;
    wire jinkela_wire_436;
    wire jinkela_wire_437;
    wire jinkela_wire_438;
    wire jinkela_wire_439;
    wire jinkela_wire_440;
    wire jinkela_wire_441;
    wire jinkela_wire_442;
    wire jinkela_wire_443;
    wire jinkela_wire_444;
    wire jinkela_wire_445;
    wire jinkela_wire_446;
    wire jinkela_wire_447;
    input a_11_;
    input a_18_;
    input a_15_;
    input a_3_;
    input a_9_;
    input a_6_;
    input a_28_;
    input a_7_;
    input a_25_;
    input a_29_;
    input a_22_;
    input a_26_;
    input a_1_;
    input a_8_;
    input a_16_;
    input a_10_;
    input a_30_;
    input a_12_;
    input a_24_;
    input a_5_;
    input a_0_;
    input a_17_;
    input a_4_;
    input a_14_;
    input a_20_;
    input a_27_;
    input a_23_;
    input a_13_;
    input a_31_;
    input a_2_;
    input a_19_;
    input a_21_;
    output b_9_;
    output b_1_;
    output b_17_;
    output b_11_;
    output b_31_;
    output b_26_;
    output b_29_;
    output b_24_;
    output b_23_;
    output b_8_;
    output b_4_;
    output b_25_;
    output b_7_;
    output b_5_;
    output b_18_;
    output b_12_;
    output b_16_;
    output b_22_;
    output b_14_;
    output b_20_;
    output b_15_;
    output b_3_;
    output b_30_;
    output b_27_;
    output b_21_;
    output b_19_;
    output b_13_;
    output b_6_;
    output b_0_;
    output b_10_;
    output b_28_;
    output b_2_;

    or_bb _006_ (
        .b(jinkela_wire_153),
        .a(jinkela_wire_0),
        .c(jinkela_wire_271)
    );

    or_bb _048_ (
        .b(a_23_),
        .a(a_22_),
        .c(jinkela_wire_76)
    );

    and_bb _007_ (
        .b(jinkela_wire_153),
        .a(jinkela_wire_0),
        .c(jinkela_wire_229)
    );

    and_bb _049_ (
        .b(a_23_),
        .a(a_22_),
        .c(jinkela_wire_280)
    );

    or_bb _008_ (
        .b(jinkela_wire_106),
        .a(jinkela_wire_271),
        .c(jinkela_wire_249)
    );

    or_bb _050_ (
        .b(a_21_),
        .a(a_20_),
        .c(jinkela_wire_165)
    );

    and_bb _009_ (
        .b(jinkela_wire_106),
        .a(jinkela_wire_271),
        .c(jinkela_wire_391)
    );

    and_bb _051_ (
        .b(a_21_),
        .a(a_20_),
        .c(jinkela_wire_227)
    );

    or_bb _010_ (
        .b(jinkela_wire_309),
        .a(jinkela_wire_229),
        .c(jinkela_wire_158)
    );

    or_bb _052_ (
        .b(jinkela_wire_76),
        .a(jinkela_wire_227),
        .c(jinkela_wire_105)
    );

    and_bb _011_ (
        .b(jinkela_wire_309),
        .a(jinkela_wire_229),
        .c(jinkela_wire_327)
    );

    and_bb _053_ (
        .b(jinkela_wire_76),
        .a(jinkela_wire_227),
        .c(jinkela_wire_94)
    );

    or_bb _012_ (
        .b(a_27_),
        .a(a_26_),
        .c(jinkela_wire_374)
    );

    or_bb _054_ (
        .b(jinkela_wire_280),
        .a(jinkela_wire_165),
        .c(jinkela_wire_211)
    );

    and_bb _013_ (
        .b(a_27_),
        .a(a_26_),
        .c(jinkela_wire_263)
    );

    and_bb _055_ (
        .b(jinkela_wire_280),
        .a(jinkela_wire_165),
        .c(jinkela_wire_295)
    );

    or_bb _014_ (
        .b(a_25_),
        .a(a_24_),
        .c(jinkela_wire_378)
    );

    or_bb _056_ (
        .b(jinkela_wire_105),
        .a(jinkela_wire_211),
        .c(jinkela_wire_144)
    );

    and_bb _015_ (
        .b(a_25_),
        .a(a_24_),
        .c(jinkela_wire_232)
    );

    and_bb _057_ (
        .b(jinkela_wire_105),
        .a(jinkela_wire_211),
        .c(jinkela_wire_253)
    );

    or_bb _016_ (
        .b(jinkela_wire_374),
        .a(jinkela_wire_232),
        .c(jinkela_wire_99)
    );

    or_bb _058_ (
        .b(jinkela_wire_94),
        .a(jinkela_wire_295),
        .c(jinkela_wire_416)
    );

    and_bb _017_ (
        .b(jinkela_wire_374),
        .a(jinkela_wire_232),
        .c(jinkela_wire_191)
    );

    and_bb _059_ (
        .b(jinkela_wire_94),
        .a(jinkela_wire_295),
        .c(jinkela_wire_369)
    );

    or_bb _018_ (
        .b(jinkela_wire_263),
        .a(jinkela_wire_378),
        .c(jinkela_wire_421)
    );

    or_bb _060_ (
        .b(a_19_),
        .a(a_18_),
        .c(jinkela_wire_282)
    );

    and_bb _019_ (
        .b(jinkela_wire_263),
        .a(jinkela_wire_378),
        .c(jinkela_wire_167)
    );

    and_bb _061_ (
        .b(a_19_),
        .a(a_18_),
        .c(jinkela_wire_304)
    );

    or_bb _020_ (
        .b(jinkela_wire_99),
        .a(jinkela_wire_421),
        .c(jinkela_wire_200)
    );

    or_bb _062_ (
        .b(a_17_),
        .a(a_16_),
        .c(jinkela_wire_390)
    );

    and_bb _021_ (
        .b(jinkela_wire_99),
        .a(jinkela_wire_421),
        .c(jinkela_wire_149)
    );

    and_bb _063_ (
        .b(a_17_),
        .a(a_16_),
        .c(jinkela_wire_231)
    );

    or_bb _022_ (
        .b(jinkela_wire_191),
        .a(jinkela_wire_167),
        .c(jinkela_wire_342)
    );

    or_bb _064_ (
        .b(jinkela_wire_282),
        .a(jinkela_wire_231),
        .c(jinkela_wire_267)
    );

    and_bb _023_ (
        .b(jinkela_wire_191),
        .a(jinkela_wire_167),
        .c(jinkela_wire_201)
    );

    and_bb _065_ (
        .b(jinkela_wire_282),
        .a(jinkela_wire_231),
        .c(jinkela_wire_399)
    );

    or_bb _024_ (
        .b(jinkela_wire_327),
        .a(jinkela_wire_200),
        .c(jinkela_wire_181)
    );

    or_bb _066_ (
        .b(jinkela_wire_304),
        .a(jinkela_wire_390),
        .c(jinkela_wire_392)
    );

    and_bb _067_ (
        .b(jinkela_wire_304),
        .a(jinkela_wire_390),
        .c(jinkela_wire_434)
    );

    and_bb _025_ (
        .b(jinkela_wire_327),
        .a(jinkela_wire_200),
        .c(jinkela_wire_289)
    );

    or_bb _068_ (
        .b(jinkela_wire_267),
        .a(jinkela_wire_392),
        .c(jinkela_wire_433)
    );

    or_bb _026_ (
        .b(jinkela_wire_158),
        .a(jinkela_wire_149),
        .c(jinkela_wire_250)
    );

    and_bb _027_ (
        .b(jinkela_wire_158),
        .a(jinkela_wire_149),
        .c(jinkela_wire_364)
    );

    and_bb _069_ (
        .b(jinkela_wire_267),
        .a(jinkela_wire_392),
        .c(jinkela_wire_160)
    );

    or_bb _028_ (
        .b(jinkela_wire_391),
        .a(jinkela_wire_342),
        .c(jinkela_wire_426)
    );

    or_bb _070_ (
        .b(jinkela_wire_399),
        .a(jinkela_wire_434),
        .c(jinkela_wire_339)
    );

    and_bb _029_ (
        .b(jinkela_wire_391),
        .a(jinkela_wire_342),
        .c(jinkela_wire_68)
    );

    and_bb _071_ (
        .b(jinkela_wire_399),
        .a(jinkela_wire_434),
        .c(jinkela_wire_236)
    );

    or_bb _030_ (
        .b(jinkela_wire_249),
        .a(jinkela_wire_201),
        .c(jinkela_wire_377)
    );

    or_bb _072_ (
        .b(jinkela_wire_369),
        .a(jinkela_wire_433),
        .c(jinkela_wire_446)
    );

    and_bb _031_ (
        .b(jinkela_wire_249),
        .a(jinkela_wire_201),
        .c(jinkela_wire_317)
    );

    and_bb _073_ (
        .b(jinkela_wire_369),
        .a(jinkela_wire_433),
        .c(jinkela_wire_38)
    );

    or_bb _032_ (
        .b(jinkela_wire_317),
        .a(jinkela_wire_364),
        .c(jinkela_wire_408)
    );

    or_bb _074_ (
        .b(jinkela_wire_416),
        .a(jinkela_wire_160),
        .c(jinkela_wire_21)
    );

    and_bb _033_ (
        .b(jinkela_wire_317),
        .a(jinkela_wire_364),
        .c(jinkela_wire_198)
    );

    and_bb _075_ (
        .b(jinkela_wire_416),
        .a(jinkela_wire_160),
        .c(jinkela_wire_27)
    );

    or_bb _034_ (
        .b(jinkela_wire_68),
        .a(jinkela_wire_289),
        .c(jinkela_wire_387)
    );

    or_bb _076_ (
        .b(jinkela_wire_253),
        .a(jinkela_wire_339),
        .c(jinkela_wire_80)
    );

    and_bb _035_ (
        .b(jinkela_wire_68),
        .a(jinkela_wire_289),
        .c(jinkela_wire_344)
    );

    and_bb _077_ (
        .b(jinkela_wire_253),
        .a(jinkela_wire_339),
        .c(jinkela_wire_351)
    );

    or_bb _036_ (
        .b(jinkela_wire_408),
        .a(jinkela_wire_387),
        .c(jinkela_wire_302)
    );

    or_bb _078_ (
        .b(jinkela_wire_144),
        .a(jinkela_wire_236),
        .c(jinkela_wire_116)
    );

    and_bb _037_ (
        .b(jinkela_wire_408),
        .a(jinkela_wire_387),
        .c(jinkela_wire_361)
    );

    and_bb _079_ (
        .b(jinkela_wire_144),
        .a(jinkela_wire_236),
        .c(jinkela_wire_242)
    );

    or_bb _038_ (
        .b(jinkela_wire_198),
        .a(jinkela_wire_344),
        .c(jinkela_wire_273)
    );

    or_bb _080_ (
        .b(jinkela_wire_242),
        .a(jinkela_wire_27),
        .c(jinkela_wire_15)
    );

    and_bb _039_ (
        .b(jinkela_wire_198),
        .a(jinkela_wire_344),
        .c(jinkela_wire_297)
    );

    and_bb _081_ (
        .b(jinkela_wire_242),
        .a(jinkela_wire_27),
        .c(jinkela_wire_60)
    );

    or_bb _040_ (
        .b(jinkela_wire_377),
        .a(jinkela_wire_250),
        .c(jinkela_wire_203)
    );

    or_bb _082_ (
        .b(jinkela_wire_351),
        .a(jinkela_wire_38),
        .c(jinkela_wire_34)
    );

    and_bb _041_ (
        .b(jinkela_wire_377),
        .a(jinkela_wire_250),
        .c(jinkela_wire_48)
    );

    and_bb _083_ (
        .b(jinkela_wire_351),
        .a(jinkela_wire_38),
        .c(jinkela_wire_11)
    );

    or_bb _042_ (
        .b(jinkela_wire_426),
        .a(jinkela_wire_181),
        .c(jinkela_wire_65)
    );

    or_bb _084_ (
        .b(jinkela_wire_15),
        .a(jinkela_wire_34),
        .c(jinkela_wire_243)
    );

    and_bb _043_ (
        .b(jinkela_wire_426),
        .a(jinkela_wire_181),
        .c(jinkela_wire_111)
    );

    and_bb _085_ (
        .b(jinkela_wire_15),
        .a(jinkela_wire_34),
        .c(jinkela_wire_212)
    );

    or_bb _044_ (
        .b(jinkela_wire_203),
        .a(jinkela_wire_65),
        .c(jinkela_wire_381)
    );

    or_bb _086_ (
        .b(jinkela_wire_60),
        .a(jinkela_wire_11),
        .c(jinkela_wire_395)
    );

    and_bb _045_ (
        .b(jinkela_wire_203),
        .a(jinkela_wire_65),
        .c(jinkela_wire_190)
    );

    and_bb _087_ (
        .b(jinkela_wire_60),
        .a(jinkela_wire_11),
        .c(jinkela_wire_16)
    );

    or_bb _046_ (
        .b(jinkela_wire_48),
        .a(jinkela_wire_111),
        .c(jinkela_wire_445)
    );

    or_bb _088_ (
        .b(jinkela_wire_116),
        .a(jinkela_wire_21),
        .c(jinkela_wire_53)
    );

    and_bb _047_ (
        .b(jinkela_wire_48),
        .a(jinkela_wire_111),
        .c(jinkela_wire_206)
    );

    and_bb _089_ (
        .b(jinkela_wire_116),
        .a(jinkela_wire_21),
        .c(jinkela_wire_171)
    );

    or_bb _132_ (
        .b(jinkela_wire_81),
        .a(jinkela_wire_46),
        .c(jinkela_wire_194)
    );

    and_bb _429_ (
        .b(jinkela_wire_222),
        .a(jinkela_wire_110),
        .c(jinkela_wire_41)
    );

    and_bb _133_ (
        .b(jinkela_wire_81),
        .a(jinkela_wire_46),
        .c(jinkela_wire_183)
    );

    or_bb _430_ (
        .b(jinkela_wire_40),
        .a(jinkela_wire_248),
        .c(jinkela_wire_96)
    );

    or_bb _134_ (
        .b(jinkela_wire_58),
        .a(jinkela_wire_354),
        .c(jinkela_wire_85)
    );

    and_bb _431_ (
        .b(jinkela_wire_40),
        .a(jinkela_wire_248),
        .c(jinkela_wire_285)
    );

    and_bb _135_ (
        .b(jinkela_wire_58),
        .a(jinkela_wire_354),
        .c(jinkela_wire_274)
    );

    or_bb _432_ (
        .b(jinkela_wire_428),
        .a(jinkela_wire_447),
        .c(jinkela_wire_100)
    );

    or_bb _136_ (
        .b(jinkela_wire_308),
        .a(jinkela_wire_319),
        .c(jinkela_wire_143)
    );

    and_bb _433_ (
        .b(jinkela_wire_428),
        .a(jinkela_wire_447),
        .c(jinkela_wire_427)
    );

    and_bb _137_ (
        .b(jinkela_wire_308),
        .a(jinkela_wire_319),
        .c(jinkela_wire_237)
    );

    or_bb _434_ (
        .b(jinkela_wire_95),
        .a(jinkela_wire_70),
        .c(jinkela_wire_388)
    );

    or_bb _138_ (
        .b(jinkela_wire_260),
        .a(jinkela_wire_33),
        .c(jinkela_wire_420)
    );

    and_bb _435_ (
        .b(jinkela_wire_95),
        .a(jinkela_wire_70),
        .c(jinkela_wire_365)
    );

    and_bb _139_ (
        .b(jinkela_wire_260),
        .a(jinkela_wire_33),
        .c(jinkela_wire_367)
    );

    or_bb _436_ (
        .b(jinkela_wire_150),
        .a(jinkela_wire_87),
        .c(jinkela_wire_166)
    );

    or_bb _140_ (
        .b(jinkela_wire_169),
        .a(jinkela_wire_135),
        .c(jinkela_wire_66)
    );

    and_bb _437_ (
        .b(jinkela_wire_150),
        .a(jinkela_wire_87),
        .c(jinkela_wire_257)
    );

    or_bb _152_ (
        .b(jinkela_wire_440),
        .a(jinkela_wire_420),
        .c(jinkela_wire_301)
    );

    and_bb _141_ (
        .b(jinkela_wire_169),
        .a(jinkela_wire_135),
        .c(jinkela_wire_315)
    );

    or_bb _438_ (
        .b(jinkela_wire_96),
        .a(jinkela_wire_247),
        .c(jinkela_wire_189)
    );

    or_bb _142_ (
        .b(jinkela_wire_346),
        .a(jinkela_wire_196),
        .c(jinkela_wire_440)
    );

    and_bb _439_ (
        .b(jinkela_wire_96),
        .a(jinkela_wire_247),
        .c(jinkela_wire_352)
    );

    and_bb _153_ (
        .b(jinkela_wire_440),
        .a(jinkela_wire_420),
        .c(jinkela_wire_375)
    );

    and_bb _143_ (
        .b(jinkela_wire_346),
        .a(jinkela_wire_196),
        .c(jinkela_wire_286)
    );

    or_bb _440_ (
        .b(jinkela_wire_352),
        .a(jinkela_wire_365),
        .c(jinkela_wire_400)
    );

    and_bb _151_ (
        .b(jinkela_wire_438),
        .a(jinkela_wire_357),
        .c(jinkela_wire_370)
    );

    or_bb _144_ (
        .b(jinkela_wire_286),
        .a(jinkela_wire_367),
        .c(jinkela_wire_230)
    );

    and_bb _441_ (
        .b(jinkela_wire_352),
        .a(jinkela_wire_365),
        .c(jinkela_wire_305)
    );

    and_bb _145_ (
        .b(jinkela_wire_286),
        .a(jinkela_wire_367),
        .c(jinkela_wire_438)
    );

    or_bb _442_ (
        .b(jinkela_wire_257),
        .a(jinkela_wire_427),
        .c(jinkela_wire_63)
    );

    or_bb _146_ (
        .b(jinkela_wire_315),
        .a(jinkela_wire_237),
        .c(jinkela_wire_164)
    );

    and_bb _443_ (
        .b(jinkela_wire_257),
        .a(jinkela_wire_427),
        .c(jinkela_wire_251)
    );

    and_bb _147_ (
        .b(jinkela_wire_315),
        .a(jinkela_wire_237),
        .c(jinkela_wire_357)
    );

    or_bb _444_ (
        .b(jinkela_wire_400),
        .a(jinkela_wire_63),
        .c(b_27_)
    );

    or_bb _148_ (
        .b(jinkela_wire_230),
        .a(jinkela_wire_164),
        .c(jinkela_wire_413)
    );

    and_bb _445_ (
        .b(jinkela_wire_400),
        .a(jinkela_wire_63),
        .c(b_26_)
    );

    and_bb _149_ (
        .b(jinkela_wire_230),
        .a(jinkela_wire_164),
        .c(jinkela_wire_118)
    );

    or_bb _446_ (
        .b(jinkela_wire_305),
        .a(jinkela_wire_251),
        .c(b_25_)
    );

    or_bb _150_ (
        .b(jinkela_wire_438),
        .a(jinkela_wire_357),
        .c(jinkela_wire_73)
    );

    and_bb _447_ (
        .b(jinkela_wire_305),
        .a(jinkela_wire_251),
        .c(b_24_)
    );

    or_bb _154_ (
        .b(jinkela_wire_66),
        .a(jinkela_wire_143),
        .c(jinkela_wire_3)
    );

    or_bb _448_ (
        .b(jinkela_wire_189),
        .a(jinkela_wire_388),
        .c(jinkela_wire_17)
    );

    and_bb _155_ (
        .b(jinkela_wire_66),
        .a(jinkela_wire_143),
        .c(jinkela_wire_170)
    );

    and_bb _449_ (
        .b(jinkela_wire_189),
        .a(jinkela_wire_388),
        .c(jinkela_wire_207)
    );

    or_bb _156_ (
        .b(jinkela_wire_301),
        .a(jinkela_wire_3),
        .c(jinkela_wire_441)
    );

    or_bb _450_ (
        .b(jinkela_wire_166),
        .a(jinkela_wire_100),
        .c(jinkela_wire_410)
    );

    and_bb _157_ (
        .b(jinkela_wire_301),
        .a(jinkela_wire_3),
        .c(jinkela_wire_213)
    );

    and_bb _451_ (
        .b(jinkela_wire_166),
        .a(jinkela_wire_100),
        .c(jinkela_wire_35)
    );

    or_bb _158_ (
        .b(jinkela_wire_375),
        .a(jinkela_wire_170),
        .c(jinkela_wire_147)
    );

    or_bb _452_ (
        .b(jinkela_wire_17),
        .a(jinkela_wire_410),
        .c(b_31_)
    );

    and_bb _159_ (
        .b(jinkela_wire_375),
        .a(jinkela_wire_170),
        .c(jinkela_wire_424)
    );

    and_bb _453_ (
        .b(jinkela_wire_17),
        .a(jinkela_wire_410),
        .c(b_30_)
    );

    or_bb _160_ (
        .b(a_15_),
        .a(a_14_),
        .c(jinkela_wire_320)
    );

    or_bb _454_ (
        .b(jinkela_wire_207),
        .a(jinkela_wire_35),
        .c(b_29_)
    );

    and_bb _161_ (
        .b(a_15_),
        .a(a_14_),
        .c(jinkela_wire_29)
    );

    and_bb _455_ (
        .b(jinkela_wire_207),
        .a(jinkela_wire_35),
        .c(b_28_)
    );

    or_bb _162_ (
        .b(a_13_),
        .a(a_12_),
        .c(jinkela_wire_356)
    );

    or_bb _456_ (
        .b(jinkela_wire_72),
        .a(jinkela_wire_125),
        .c(jinkela_wire_350)
    );

    and_bb _163_ (
        .b(a_13_),
        .a(a_12_),
        .c(jinkela_wire_360)
    );

    and_bb _457_ (
        .b(jinkela_wire_72),
        .a(jinkela_wire_125),
        .c(jinkela_wire_405)
    );

    or_bb _164_ (
        .b(jinkela_wire_320),
        .a(jinkela_wire_360),
        .c(jinkela_wire_36)
    );

    or_bb _458_ (
        .b(jinkela_wire_137),
        .a(jinkela_wire_89),
        .c(jinkela_wire_414)
    );

    and_bb _165_ (
        .b(jinkela_wire_320),
        .a(jinkela_wire_360),
        .c(jinkela_wire_218)
    );

    and_bb _459_ (
        .b(jinkela_wire_137),
        .a(jinkela_wire_89),
        .c(jinkela_wire_403)
    );

    or_bb _166_ (
        .b(jinkela_wire_29),
        .a(jinkela_wire_356),
        .c(jinkela_wire_425)
    );

    or_bb _460_ (
        .b(jinkela_wire_41),
        .a(jinkela_wire_379),
        .c(jinkela_wire_359)
    );

    and_bb _167_ (
        .b(jinkela_wire_29),
        .a(jinkela_wire_356),
        .c(jinkela_wire_419)
    );

    and_bb _461_ (
        .b(jinkela_wire_41),
        .a(jinkela_wire_379),
        .c(jinkela_wire_288)
    );

    or_bb _168_ (
        .b(jinkela_wire_36),
        .a(jinkela_wire_425),
        .c(jinkela_wire_376)
    );

    or_bb _462_ (
        .b(jinkela_wire_285),
        .a(jinkela_wire_57),
        .c(jinkela_wire_383)
    );

    and_bb _169_ (
        .b(jinkela_wire_36),
        .a(jinkela_wire_425),
        .c(jinkela_wire_173)
    );

    and_bb _463_ (
        .b(jinkela_wire_285),
        .a(jinkela_wire_57),
        .c(jinkela_wire_124)
    );

    or_bb _170_ (
        .b(jinkela_wire_218),
        .a(jinkela_wire_419),
        .c(jinkela_wire_97)
    );

    or_bb _464_ (
        .b(jinkela_wire_124),
        .a(jinkela_wire_403),
        .c(jinkela_wire_324)
    );

    and_bb _171_ (
        .b(jinkela_wire_218),
        .a(jinkela_wire_419),
        .c(jinkela_wire_238)
    );

    and_bb _465_ (
        .b(jinkela_wire_124),
        .a(jinkela_wire_403),
        .c(jinkela_wire_208)
    );

    or_bb _172_ (
        .b(a_11_),
        .a(a_10_),
        .c(jinkela_wire_154)
    );

    or_bb _466_ (
        .b(jinkela_wire_288),
        .a(jinkela_wire_405),
        .c(jinkela_wire_432)
    );

    and_bb _173_ (
        .b(a_11_),
        .a(a_10_),
        .c(jinkela_wire_122)
    );

    and_bb _467_ (
        .b(jinkela_wire_288),
        .a(jinkela_wire_405),
        .c(jinkela_wire_62)
    );

    or_bb _174_ (
        .b(a_9_),
        .a(a_8_),
        .c(jinkela_wire_382)
    );

    or_bb _468_ (
        .b(jinkela_wire_324),
        .a(jinkela_wire_432),
        .c(b_19_)
    );

    and_bb _175_ (
        .b(a_9_),
        .a(a_8_),
        .c(jinkela_wire_162)
    );

    and_bb _469_ (
        .b(jinkela_wire_324),
        .a(jinkela_wire_432),
        .c(b_18_)
    );

    or_bb _176_ (
        .b(jinkela_wire_154),
        .a(jinkela_wire_162),
        .c(jinkela_wire_366)
    );

    or_bb _470_ (
        .b(jinkela_wire_208),
        .a(jinkela_wire_62),
        .c(b_17_)
    );

    and_bb _261_ (
        .b(jinkela_wire_180),
        .a(jinkela_wire_98),
        .c(jinkela_wire_313)
    );

    or_bb _262_ (
        .b(jinkela_wire_223),
        .a(jinkela_wire_56),
        .c(jinkela_wire_355)
    );

    and_bb _263_ (
        .b(jinkela_wire_223),
        .a(jinkela_wire_56),
        .c(jinkela_wire_261)
    );

    or_bb _264_ (
        .b(jinkela_wire_343),
        .a(jinkela_wire_24),
        .c(jinkela_wire_77)
    );

    and_bb _265_ (
        .b(jinkela_wire_343),
        .a(jinkela_wire_24),
        .c(jinkela_wire_259)
    );

    or_bb _266_ (
        .b(jinkela_wire_415),
        .a(jinkela_wire_22),
        .c(jinkela_wire_184)
    );

    and_bb _267_ (
        .b(jinkela_wire_415),
        .a(jinkela_wire_22),
        .c(jinkela_wire_234)
    );

    or_bb _268_ (
        .b(jinkela_wire_215),
        .a(jinkela_wire_43),
        .c(jinkela_wire_6)
    );

    and_bb _269_ (
        .b(jinkela_wire_215),
        .a(jinkela_wire_43),
        .c(jinkela_wire_74)
    );

    or_bb _270_ (
        .b(jinkela_wire_217),
        .a(jinkela_wire_83),
        .c(jinkela_wire_321)
    );

    and_bb _271_ (
        .b(jinkela_wire_217),
        .a(jinkela_wire_83),
        .c(jinkela_wire_362)
    );

    or_bb _272_ (
        .b(jinkela_wire_77),
        .a(jinkela_wire_192),
        .c(jinkela_wire_130)
    );

    and_bb _273_ (
        .b(jinkela_wire_77),
        .a(jinkela_wire_192),
        .c(jinkela_wire_119)
    );

    or_bb _274_ (
        .b(jinkela_wire_184),
        .a(jinkela_wire_368),
        .c(jinkela_wire_155)
    );

    and_bb _275_ (
        .b(jinkela_wire_184),
        .a(jinkela_wire_368),
        .c(jinkela_wire_133)
    );

    or_bb _276_ (
        .b(jinkela_wire_6),
        .a(jinkela_wire_283),
        .c(jinkela_wire_193)
    );

    and_bb _277_ (
        .b(jinkela_wire_6),
        .a(jinkela_wire_283),
        .c(jinkela_wire_67)
    );

    or_bb _278_ (
        .b(jinkela_wire_321),
        .a(jinkela_wire_355),
        .c(jinkela_wire_172)
    );

    and_bb _279_ (
        .b(jinkela_wire_321),
        .a(jinkela_wire_355),
        .c(jinkela_wire_209)
    );

    or_bb _280_ (
        .b(jinkela_wire_209),
        .a(jinkela_wire_133),
        .c(jinkela_wire_422)
    );

    and_bb _281_ (
        .b(jinkela_wire_209),
        .a(jinkela_wire_133),
        .c(jinkela_wire_69)
    );

    or_bb _282_ (
        .b(jinkela_wire_67),
        .a(jinkela_wire_119),
        .c(jinkela_wire_330)
    );

    and_bb _283_ (
        .b(jinkela_wire_67),
        .a(jinkela_wire_119),
        .c(jinkela_wire_396)
    );

    or_bb _284_ (
        .b(jinkela_wire_422),
        .a(jinkela_wire_330),
        .c(jinkela_wire_269)
    );

    and_bb _285_ (
        .b(jinkela_wire_422),
        .a(jinkela_wire_330),
        .c(jinkela_wire_54)
    );

    or_bb _286_ (
        .b(jinkela_wire_69),
        .a(jinkela_wire_396),
        .c(jinkela_wire_127)
    );

    and_bb _287_ (
        .b(jinkela_wire_69),
        .a(jinkela_wire_396),
        .c(jinkela_wire_140)
    );

    or_bb _288_ (
        .b(jinkela_wire_172),
        .a(jinkela_wire_155),
        .c(jinkela_wire_91)
    );

    and_bb _289_ (
        .b(jinkela_wire_172),
        .a(jinkela_wire_155),
        .c(jinkela_wire_39)
    );

    or_bb _290_ (
        .b(jinkela_wire_193),
        .a(jinkela_wire_130),
        .c(jinkela_wire_318)
    );

    and_bb _291_ (
        .b(jinkela_wire_193),
        .a(jinkela_wire_130),
        .c(jinkela_wire_353)
    );

    or_bb _292_ (
        .b(jinkela_wire_91),
        .a(jinkela_wire_318),
        .c(jinkela_wire_252)
    );

    and_bb _293_ (
        .b(jinkela_wire_91),
        .a(jinkela_wire_318),
        .c(jinkela_wire_437)
    );

    or_bb _294_ (
        .b(jinkela_wire_39),
        .a(jinkela_wire_353),
        .c(jinkela_wire_78)
    );

    and_bb _295_ (
        .b(jinkela_wire_39),
        .a(jinkela_wire_353),
        .c(jinkela_wire_389)
    );

    or_bb _296_ (
        .b(jinkela_wire_259),
        .a(jinkela_wire_132),
        .c(jinkela_wire_1)
    );

    and_bb _297_ (
        .b(jinkela_wire_259),
        .a(jinkela_wire_132),
        .c(jinkela_wire_423)
    );

    or_bb _298_ (
        .b(jinkela_wire_234),
        .a(jinkela_wire_228),
        .c(jinkela_wire_10)
    );

    and_bb _299_ (
        .b(jinkela_wire_234),
        .a(jinkela_wire_228),
        .c(jinkela_wire_107)
    );

    or_bb _300_ (
        .b(jinkela_wire_74),
        .a(jinkela_wire_313),
        .c(jinkela_wire_50)
    );

    and_bb _301_ (
        .b(jinkela_wire_74),
        .a(jinkela_wire_313),
        .c(jinkela_wire_287)
    );

    or_bb _302_ (
        .b(jinkela_wire_362),
        .a(jinkela_wire_261),
        .c(jinkela_wire_59)
    );

    and_bb _177_ (
        .b(jinkela_wire_154),
        .a(jinkela_wire_162),
        .c(jinkela_wire_23)
    );

    and_bb _219_ (
        .b(jinkela_wire_93),
        .a(jinkela_wire_266),
        .c(jinkela_wire_156)
    );

    or_bb _178_ (
        .b(jinkela_wire_122),
        .a(jinkela_wire_382),
        .c(jinkela_wire_244)
    );

    or_bb _220_ (
        .b(a_3_),
        .a(a_2_),
        .c(jinkela_wire_328)
    );

    and_bb _179_ (
        .b(jinkela_wire_122),
        .a(jinkela_wire_382),
        .c(jinkela_wire_270)
    );

    and_bb _221_ (
        .b(a_3_),
        .a(a_2_),
        .c(jinkela_wire_265)
    );

    or_bb _180_ (
        .b(jinkela_wire_366),
        .a(jinkela_wire_244),
        .c(jinkela_wire_163)
    );

    or_bb _222_ (
        .b(a_1_),
        .a(a_0_),
        .c(jinkela_wire_442)
    );

    and_bb _181_ (
        .b(jinkela_wire_366),
        .a(jinkela_wire_244),
        .c(jinkela_wire_272)
    );

    and_bb _223_ (
        .b(a_1_),
        .a(a_0_),
        .c(jinkela_wire_373)
    );

    or_bb _182_ (
        .b(jinkela_wire_23),
        .a(jinkela_wire_270),
        .c(jinkela_wire_136)
    );

    or_bb _224_ (
        .b(jinkela_wire_328),
        .a(jinkela_wire_373),
        .c(jinkela_wire_115)
    );

    and_bb _183_ (
        .b(jinkela_wire_23),
        .a(jinkela_wire_270),
        .c(jinkela_wire_18)
    );

    and_bb _225_ (
        .b(jinkela_wire_328),
        .a(jinkela_wire_373),
        .c(jinkela_wire_19)
    );

    or_bb _184_ (
        .b(jinkela_wire_238),
        .a(jinkela_wire_163),
        .c(jinkela_wire_430)
    );

    or_bb _226_ (
        .b(jinkela_wire_265),
        .a(jinkela_wire_442),
        .c(jinkela_wire_210)
    );

    and_bb _185_ (
        .b(jinkela_wire_238),
        .a(jinkela_wire_163),
        .c(jinkela_wire_28)
    );

    and_bb _227_ (
        .b(jinkela_wire_265),
        .a(jinkela_wire_442),
        .c(jinkela_wire_90)
    );

    or_bb _186_ (
        .b(jinkela_wire_97),
        .a(jinkela_wire_272),
        .c(jinkela_wire_42)
    );

    or_bb _228_ (
        .b(jinkela_wire_115),
        .a(jinkela_wire_210),
        .c(jinkela_wire_314)
    );

    and_bb _187_ (
        .b(jinkela_wire_97),
        .a(jinkela_wire_272),
        .c(jinkela_wire_182)
    );

    and_bb _229_ (
        .b(jinkela_wire_115),
        .a(jinkela_wire_210),
        .c(jinkela_wire_131)
    );

    or_bb _188_ (
        .b(jinkela_wire_173),
        .a(jinkela_wire_136),
        .c(jinkela_wire_254)
    );

    or_bb _230_ (
        .b(jinkela_wire_19),
        .a(jinkela_wire_90),
        .c(jinkela_wire_79)
    );

    and_bb _189_ (
        .b(jinkela_wire_173),
        .a(jinkela_wire_136),
        .c(jinkela_wire_246)
    );

    and_bb _231_ (
        .b(jinkela_wire_19),
        .a(jinkela_wire_90),
        .c(jinkela_wire_187)
    );

    or_bb _190_ (
        .b(jinkela_wire_376),
        .a(jinkela_wire_18),
        .c(jinkela_wire_202)
    );

    or_bb _232_ (
        .b(jinkela_wire_156),
        .a(jinkela_wire_314),
        .c(jinkela_wire_340)
    );

    and_bb _191_ (
        .b(jinkela_wire_376),
        .a(jinkela_wire_18),
        .c(jinkela_wire_64)
    );

    and_bb _233_ (
        .b(jinkela_wire_156),
        .a(jinkela_wire_314),
        .c(jinkela_wire_331)
    );

    or_bb _192_ (
        .b(jinkela_wire_64),
        .a(jinkela_wire_182),
        .c(jinkela_wire_332)
    );

    or_bb _234_ (
        .b(jinkela_wire_75),
        .a(jinkela_wire_131),
        .c(jinkela_wire_264)
    );

    and_bb _193_ (
        .b(jinkela_wire_64),
        .a(jinkela_wire_182),
        .c(jinkela_wire_168)
    );

    and_bb _235_ (
        .b(jinkela_wire_75),
        .a(jinkela_wire_131),
        .c(jinkela_wire_436)
    );

    or_bb _194_ (
        .b(jinkela_wire_246),
        .a(jinkela_wire_28),
        .c(jinkela_wire_152)
    );

    or_bb _236_ (
        .b(jinkela_wire_30),
        .a(jinkela_wire_79),
        .c(jinkela_wire_307)
    );

    and_bb _195_ (
        .b(jinkela_wire_246),
        .a(jinkela_wire_28),
        .c(jinkela_wire_114)
    );

    and_bb _237_ (
        .b(jinkela_wire_30),
        .a(jinkela_wire_79),
        .c(jinkela_wire_296)
    );

    or_bb _196_ (
        .b(jinkela_wire_332),
        .a(jinkela_wire_152),
        .c(jinkela_wire_223)
    );

    or_bb _238_ (
        .b(jinkela_wire_26),
        .a(jinkela_wire_187),
        .c(jinkela_wire_84)
    );

    and_bb _197_ (
        .b(jinkela_wire_332),
        .a(jinkela_wire_152),
        .c(jinkela_wire_180)
    );

    and_bb _239_ (
        .b(jinkela_wire_26),
        .a(jinkela_wire_187),
        .c(jinkela_wire_412)
    );

    or_bb _198_ (
        .b(jinkela_wire_168),
        .a(jinkela_wire_114),
        .c(jinkela_wire_117)
    );

    or_bb _240_ (
        .b(jinkela_wire_412),
        .a(jinkela_wire_436),
        .c(jinkela_wire_404)
    );

    and_bb _199_ (
        .b(jinkela_wire_168),
        .a(jinkela_wire_114),
        .c(jinkela_wire_341)
    );

    and_bb _241_ (
        .b(jinkela_wire_412),
        .a(jinkela_wire_436),
        .c(jinkela_wire_284)
    );

    or_bb _200_ (
        .b(jinkela_wire_202),
        .a(jinkela_wire_42),
        .c(jinkela_wire_402)
    );

    or_bb _242_ (
        .b(jinkela_wire_296),
        .a(jinkela_wire_331),
        .c(jinkela_wire_245)
    );

    and_bb _201_ (
        .b(jinkela_wire_202),
        .a(jinkela_wire_42),
        .c(jinkela_wire_101)
    );

    and_bb _243_ (
        .b(jinkela_wire_296),
        .a(jinkela_wire_331),
        .c(jinkela_wire_92)
    );

    or_bb _202_ (
        .b(jinkela_wire_254),
        .a(jinkela_wire_430),
        .c(jinkela_wire_294)
    );

    or_bb _244_ (
        .b(jinkela_wire_404),
        .a(jinkela_wire_245),
        .c(jinkela_wire_24)
    );

    and_bb _203_ (
        .b(jinkela_wire_254),
        .a(jinkela_wire_430),
        .c(jinkela_wire_8)
    );

    and_bb _245_ (
        .b(jinkela_wire_404),
        .a(jinkela_wire_245),
        .c(jinkela_wire_22)
    );

    or_bb _204_ (
        .b(jinkela_wire_402),
        .a(jinkela_wire_294),
        .c(jinkela_wire_217)
    );

    or_bb _246_ (
        .b(jinkela_wire_284),
        .a(jinkela_wire_92),
        .c(jinkela_wire_43)
    );

    and_bb _205_ (
        .b(jinkela_wire_402),
        .a(jinkela_wire_294),
        .c(jinkela_wire_215)
    );

    and_bb _247_ (
        .b(jinkela_wire_284),
        .a(jinkela_wire_92),
        .c(jinkela_wire_83)
    );

    or_bb _206_ (
        .b(jinkela_wire_101),
        .a(jinkela_wire_8),
        .c(jinkela_wire_415)
    );

    or_bb _248_ (
        .b(jinkela_wire_84),
        .a(jinkela_wire_264),
        .c(jinkela_wire_179)
    );

    and_bb _207_ (
        .b(jinkela_wire_101),
        .a(jinkela_wire_8),
        .c(jinkela_wire_343)
    );

    and_bb _249_ (
        .b(jinkela_wire_84),
        .a(jinkela_wire_264),
        .c(jinkela_wire_88)
    );

    or_bb _208_ (
        .b(a_7_),
        .a(a_6_),
        .c(jinkela_wire_325)
    );

    or_bb _250_ (
        .b(jinkela_wire_307),
        .a(jinkela_wire_340),
        .c(jinkela_wire_45)
    );

    and_bb _209_ (
        .b(a_7_),
        .a(a_6_),
        .c(jinkela_wire_112)
    );

    and_bb _251_ (
        .b(jinkela_wire_307),
        .a(jinkela_wire_340),
        .c(jinkela_wire_335)
    );

    or_bb _210_ (
        .b(a_5_),
        .a(a_4_),
        .c(jinkela_wire_151)
    );

    or_bb _252_ (
        .b(jinkela_wire_179),
        .a(jinkela_wire_45),
        .c(jinkela_wire_219)
    );

    and_bb _211_ (
        .b(a_5_),
        .a(a_4_),
        .c(jinkela_wire_49)
    );

    and_bb _253_ (
        .b(jinkela_wire_179),
        .a(jinkela_wire_45),
        .c(jinkela_wire_185)
    );

    or_bb _212_ (
        .b(jinkela_wire_325),
        .a(jinkela_wire_49),
        .c(jinkela_wire_276)
    );

    or_bb _254_ (
        .b(jinkela_wire_88),
        .a(jinkela_wire_335),
        .c(jinkela_wire_98)
    );

    and_bb _213_ (
        .b(jinkela_wire_325),
        .a(jinkela_wire_49),
        .c(jinkela_wire_93)
    );

    and_bb _255_ (
        .b(jinkela_wire_88),
        .a(jinkela_wire_335),
        .c(jinkela_wire_56)
    );

    or_bb _214_ (
        .b(jinkela_wire_112),
        .a(jinkela_wire_151),
        .c(jinkela_wire_439)
    );

    or_bb _256_ (
        .b(jinkela_wire_341),
        .a(jinkela_wire_219),
        .c(jinkela_wire_192)
    );

    and_bb _215_ (
        .b(jinkela_wire_112),
        .a(jinkela_wire_151),
        .c(jinkela_wire_266)
    );

    and_bb _257_ (
        .b(jinkela_wire_341),
        .a(jinkela_wire_219),
        .c(jinkela_wire_132)
    );

    or_bb _216_ (
        .b(jinkela_wire_276),
        .a(jinkela_wire_439),
        .c(jinkela_wire_26)
    );

    or_bb _258_ (
        .b(jinkela_wire_117),
        .a(jinkela_wire_185),
        .c(jinkela_wire_368)
    );

    and_bb _217_ (
        .b(jinkela_wire_276),
        .a(jinkela_wire_439),
        .c(jinkela_wire_30)
    );

    and_bb _259_ (
        .b(jinkela_wire_117),
        .a(jinkela_wire_185),
        .c(jinkela_wire_228)
    );

    or_bb _218_ (
        .b(jinkela_wire_93),
        .a(jinkela_wire_266),
        .c(jinkela_wire_75)
    );

    or_bb _260_ (
        .b(jinkela_wire_180),
        .a(jinkela_wire_98),
        .c(jinkela_wire_283)
    );

    and_bb _303_ (
        .b(jinkela_wire_362),
        .a(jinkela_wire_261),
        .c(jinkela_wire_277)
    );

    and_bb _345_ (
        .b(jinkela_wire_274),
        .a(jinkela_wire_224),
        .c(jinkela_wire_300)
    );

    and_bb _471_ (
        .b(jinkela_wire_208),
        .a(jinkela_wire_62),
        .c(b_16_)
    );

    or_bb _304_ (
        .b(jinkela_wire_277),
        .a(jinkela_wire_107),
        .c(jinkela_wire_334)
    );

    or_bb _346_ (
        .b(jinkela_wire_85),
        .a(jinkela_wire_298),
        .c(jinkela_wire_371)
    );

    or_bb _472_ (
        .b(jinkela_wire_383),
        .a(jinkela_wire_414),
        .c(jinkela_wire_199)
    );

    and_bb _305_ (
        .b(jinkela_wire_277),
        .a(jinkela_wire_107),
        .c(jinkela_wire_121)
    );

    and_bb _347_ (
        .b(jinkela_wire_85),
        .a(jinkela_wire_298),
        .c(jinkela_wire_326)
    );

    and_bb _473_ (
        .b(jinkela_wire_383),
        .a(jinkela_wire_414),
        .c(jinkela_wire_429)
    );

    or_bb _306_ (
        .b(jinkela_wire_287),
        .a(jinkela_wire_423),
        .c(jinkela_wire_444)
    );

    or_bb _348_ (
        .b(jinkela_wire_183),
        .a(jinkela_wire_4),
        .c(jinkela_wire_222)
    );

    or_bb _474_ (
        .b(jinkela_wire_359),
        .a(jinkela_wire_350),
        .c(jinkela_wire_401)
    );

    and_bb _307_ (
        .b(jinkela_wire_287),
        .a(jinkela_wire_423),
        .c(jinkela_wire_177)
    );

    and_bb _349_ (
        .b(jinkela_wire_183),
        .a(jinkela_wire_4),
        .c(jinkela_wire_37)
    );

    and_bb _475_ (
        .b(jinkela_wire_359),
        .a(jinkela_wire_350),
        .c(jinkela_wire_262)
    );

    or_bb _308_ (
        .b(jinkela_wire_334),
        .a(jinkela_wire_444),
        .c(jinkela_wire_224)
    );

    or_bb _350_ (
        .b(jinkela_wire_194),
        .a(jinkela_wire_293),
        .c(jinkela_wire_40)
    );

    or_bb _476_ (
        .b(jinkela_wire_199),
        .a(jinkela_wire_401),
        .c(b_23_)
    );

    and_bb _309_ (
        .b(jinkela_wire_334),
        .a(jinkela_wire_444),
        .c(jinkela_wire_298)
    );

    and_bb _351_ (
        .b(jinkela_wire_194),
        .a(jinkela_wire_293),
        .c(jinkela_wire_407)
    );

    and_bb _477_ (
        .b(jinkela_wire_199),
        .a(jinkela_wire_401),
        .c(b_22_)
    );

    or_bb _310_ (
        .b(jinkela_wire_121),
        .a(jinkela_wire_177),
        .c(jinkela_wire_4)
    );

    or_bb _352_ (
        .b(jinkela_wire_235),
        .a(jinkela_wire_138),
        .c(jinkela_wire_275)
    );

    or_bb _478_ (
        .b(jinkela_wire_429),
        .a(jinkela_wire_262),
        .c(b_21_)
    );

    and_bb _311_ (
        .b(jinkela_wire_121),
        .a(jinkela_wire_177),
        .c(jinkela_wire_293)
    );

    and_bb _353_ (
        .b(jinkela_wire_235),
        .a(jinkela_wire_138),
        .c(jinkela_wire_103)
    );

    and_bb _479_ (
        .b(jinkela_wire_429),
        .a(jinkela_wire_262),
        .c(b_20_)
    );

    or_bb _312_ (
        .b(jinkela_wire_59),
        .a(jinkela_wire_10),
        .c(jinkela_wire_363)
    );

    or_bb _354_ (
        .b(jinkela_wire_61),
        .a(jinkela_wire_55),
        .c(jinkela_wire_82)
    );

    and_bb _313_ (
        .b(jinkela_wire_59),
        .a(jinkela_wire_10),
        .c(jinkela_wire_32)
    );

    and_bb _355_ (
        .b(jinkela_wire_61),
        .a(jinkela_wire_55),
        .c(jinkela_wire_268)
    );

    or_bb _314_ (
        .b(jinkela_wire_50),
        .a(jinkela_wire_1),
        .c(jinkela_wire_349)
    );

    or_bb _356_ (
        .b(jinkela_wire_109),
        .a(jinkela_wire_12),
        .c(jinkela_wire_178)
    );

    and_bb _315_ (
        .b(jinkela_wire_50),
        .a(jinkela_wire_1),
        .c(jinkela_wire_312)
    );

    and_bb _357_ (
        .b(jinkela_wire_109),
        .a(jinkela_wire_12),
        .c(jinkela_wire_175)
    );

    or_bb _316_ (
        .b(jinkela_wire_363),
        .a(jinkela_wire_349),
        .c(jinkela_wire_258)
    );

    or_bb _358_ (
        .b(jinkela_wire_323),
        .a(jinkela_wire_233),
        .c(jinkela_wire_176)
    );

    and_bb _317_ (
        .b(jinkela_wire_363),
        .a(jinkela_wire_349),
        .c(jinkela_wire_142)
    );

    and_bb _359_ (
        .b(jinkela_wire_323),
        .a(jinkela_wire_233),
        .c(jinkela_wire_134)
    );

    or_bb _318_ (
        .b(jinkela_wire_32),
        .a(jinkela_wire_312),
        .c(jinkela_wire_139)
    );

    or_bb _360_ (
        .b(jinkela_wire_300),
        .a(jinkela_wire_7),
        .c(jinkela_wire_347)
    );

    and_bb _319_ (
        .b(jinkela_wire_32),
        .a(jinkela_wire_312),
        .c(jinkela_wire_291)
    );

    and_bb _361_ (
        .b(jinkela_wire_300),
        .a(jinkela_wire_7),
        .c(jinkela_wire_104)
    );

    or_bb _320_ (
        .b(jinkela_wire_370),
        .a(jinkela_wire_252),
        .c(jinkela_wire_397)
    );

    or_bb _362_ (
        .b(jinkela_wire_326),
        .a(jinkela_wire_216),
        .c(jinkela_wire_290)
    );

    and_bb _321_ (
        .b(jinkela_wire_370),
        .a(jinkela_wire_252),
        .c(jinkela_wire_138)
    );

    and_bb _363_ (
        .b(jinkela_wire_326),
        .a(jinkela_wire_216),
        .c(jinkela_wire_123)
    );

    or_bb _322_ (
        .b(jinkela_wire_73),
        .a(jinkela_wire_437),
        .c(jinkela_wire_393)
    );

    or_bb _364_ (
        .b(jinkela_wire_37),
        .a(jinkela_wire_148),
        .c(jinkela_wire_14)
    );

    and_bb _323_ (
        .b(jinkela_wire_73),
        .a(jinkela_wire_437),
        .c(jinkela_wire_55)
    );

    and_bb _365_ (
        .b(jinkela_wire_37),
        .a(jinkela_wire_148),
        .c(jinkela_wire_329)
    );

    or_bb _324_ (
        .b(jinkela_wire_118),
        .a(jinkela_wire_78),
        .c(jinkela_wire_226)
    );

    or_bb _366_ (
        .b(jinkela_wire_407),
        .a(jinkela_wire_322),
        .c(jinkela_wire_13)
    );

    and_bb _325_ (
        .b(jinkela_wire_118),
        .a(jinkela_wire_78),
        .c(jinkela_wire_12)
    );

    and_bb _367_ (
        .b(jinkela_wire_407),
        .a(jinkela_wire_322),
        .c(jinkela_wire_240)
    );

    or_bb _326_ (
        .b(jinkela_wire_413),
        .a(jinkela_wire_389),
        .c(jinkela_wire_195)
    );

    or_bb _368_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_275),
        .c(jinkela_wire_51)
    );

    and_bb _327_ (
        .b(jinkela_wire_413),
        .a(jinkela_wire_389),
        .c(jinkela_wire_233)
    );

    and_bb _369_ (
        .b(jinkela_wire_347),
        .a(jinkela_wire_275),
        .c(jinkela_wire_31)
    );

    or_bb _328_ (
        .b(jinkela_wire_424),
        .a(jinkela_wire_269),
        .c(jinkela_wire_126)
    );

    or_bb _370_ (
        .b(jinkela_wire_290),
        .a(jinkela_wire_82),
        .c(jinkela_wire_52)
    );

    and_bb _329_ (
        .b(jinkela_wire_424),
        .a(jinkela_wire_269),
        .c(jinkela_wire_7)
    );

    and_bb _371_ (
        .b(jinkela_wire_290),
        .a(jinkela_wire_82),
        .c(jinkela_wire_108)
    );

    or_bb _330_ (
        .b(jinkela_wire_147),
        .a(jinkela_wire_54),
        .c(jinkela_wire_197)
    );

    or_bb _372_ (
        .b(jinkela_wire_14),
        .a(jinkela_wire_178),
        .c(jinkela_wire_225)
    );

    and_bb _331_ (
        .b(jinkela_wire_147),
        .a(jinkela_wire_54),
        .c(jinkela_wire_216)
    );

    and_bb _373_ (
        .b(jinkela_wire_14),
        .a(jinkela_wire_178),
        .c(jinkela_wire_443)
    );

    or_bb _332_ (
        .b(jinkela_wire_213),
        .a(jinkela_wire_127),
        .c(jinkela_wire_110)
    );

    or_bb _374_ (
        .b(jinkela_wire_13),
        .a(jinkela_wire_176),
        .c(jinkela_wire_146)
    );

    and_bb _333_ (
        .b(jinkela_wire_213),
        .a(jinkela_wire_127),
        .c(jinkela_wire_148)
    );

    and_bb _375_ (
        .b(jinkela_wire_13),
        .a(jinkela_wire_176),
        .c(jinkela_wire_221)
    );

    or_bb _334_ (
        .b(jinkela_wire_441),
        .a(jinkela_wire_140),
        .c(jinkela_wire_248)
    );

    or_bb _376_ (
        .b(jinkela_wire_221),
        .a(jinkela_wire_108),
        .c(jinkela_wire_71)
    );

    and_bb _335_ (
        .b(jinkela_wire_441),
        .a(jinkela_wire_140),
        .c(jinkela_wire_322)
    );

    and_bb _377_ (
        .b(jinkela_wire_221),
        .a(jinkela_wire_108),
        .c(jinkela_wire_299)
    );

    or_bb _336_ (
        .b(jinkela_wire_47),
        .a(jinkela_wire_258),
        .c(jinkela_wire_310)
    );

    or_bb _378_ (
        .b(jinkela_wire_443),
        .a(jinkela_wire_31),
        .c(jinkela_wire_188)
    );

    and_bb _337_ (
        .b(jinkela_wire_47),
        .a(jinkela_wire_258),
        .c(jinkela_wire_235)
    );

    and_bb _379_ (
        .b(jinkela_wire_443),
        .a(jinkela_wire_31),
        .c(jinkela_wire_204)
    );

    or_bb _338_ (
        .b(jinkela_wire_386),
        .a(jinkela_wire_142),
        .c(jinkela_wire_345)
    );

    or_bb _380_ (
        .b(jinkela_wire_71),
        .a(jinkela_wire_188),
        .c(b_11_)
    );

    and_bb _339_ (
        .b(jinkela_wire_386),
        .a(jinkela_wire_142),
        .c(jinkela_wire_61)
    );

    and_bb _381_ (
        .b(jinkela_wire_71),
        .a(jinkela_wire_188),
        .c(b_10_)
    );

    or_bb _340_ (
        .b(jinkela_wire_311),
        .a(jinkela_wire_139),
        .c(jinkela_wire_358)
    );

    or_bb _382_ (
        .b(jinkela_wire_299),
        .a(jinkela_wire_204),
        .c(b_9_)
    );

    and_bb _341_ (
        .b(jinkela_wire_311),
        .a(jinkela_wire_139),
        .c(jinkela_wire_109)
    );

    and_bb _383_ (
        .b(jinkela_wire_299),
        .a(jinkela_wire_204),
        .c(b_8_)
    );

    or_bb _342_ (
        .b(jinkela_wire_338),
        .a(jinkela_wire_291),
        .c(jinkela_wire_2)
    );

    or_bb _384_ (
        .b(jinkela_wire_146),
        .a(jinkela_wire_52),
        .c(jinkela_wire_159)
    );

    and_bb _343_ (
        .b(jinkela_wire_338),
        .a(jinkela_wire_291),
        .c(jinkela_wire_323)
    );

    and_bb _385_ (
        .b(jinkela_wire_146),
        .a(jinkela_wire_52),
        .c(jinkela_wire_113)
    );

    or_bb _344_ (
        .b(jinkela_wire_274),
        .a(jinkela_wire_224),
        .c(jinkela_wire_9)
    );

    or_bb _386_ (
        .b(jinkela_wire_225),
        .a(jinkela_wire_51),
        .c(jinkela_wire_161)
    );

    and_bb _003_ (
        .b(a_29_),
        .a(a_28_),
        .c(jinkela_wire_25)
    );

    and_bb _001_ (
        .b(a_31_),
        .a(a_30_),
        .c(jinkela_wire_153)
    );

    or_bb _002_ (
        .b(a_29_),
        .a(a_28_),
        .c(jinkela_wire_0)
    );

    or_bb _000_ (
        .b(a_31_),
        .a(a_30_),
        .c(jinkela_wire_256)
    );

    or_bb _004_ (
        .b(jinkela_wire_256),
        .a(jinkela_wire_25),
        .c(jinkela_wire_106)
    );

    and_bb _005_ (
        .b(jinkela_wire_256),
        .a(jinkela_wire_25),
        .c(jinkela_wire_309)
    );

    and_bb _387_ (
        .b(jinkela_wire_225),
        .a(jinkela_wire_51),
        .c(jinkela_wire_279)
    );

    or_bb _388_ (
        .b(jinkela_wire_159),
        .a(jinkela_wire_161),
        .c(b_15_)
    );

    and_bb _389_ (
        .b(jinkela_wire_159),
        .a(jinkela_wire_161),
        .c(b_14_)
    );

    or_bb _390_ (
        .b(jinkela_wire_113),
        .a(jinkela_wire_279),
        .c(b_13_)
    );

    and_bb _391_ (
        .b(jinkela_wire_113),
        .a(jinkela_wire_279),
        .c(b_12_)
    );

    or_bb _392_ (
        .b(jinkela_wire_104),
        .a(jinkela_wire_103),
        .c(jinkela_wire_44)
    );

    and_bb _393_ (
        .b(jinkela_wire_104),
        .a(jinkela_wire_103),
        .c(jinkela_wire_348)
    );

    or_bb _394_ (
        .b(jinkela_wire_123),
        .a(jinkela_wire_268),
        .c(jinkela_wire_281)
    );

    and_bb _395_ (
        .b(jinkela_wire_123),
        .a(jinkela_wire_268),
        .c(jinkela_wire_255)
    );

    or_bb _396_ (
        .b(jinkela_wire_329),
        .a(jinkela_wire_175),
        .c(jinkela_wire_174)
    );

    and_bb _397_ (
        .b(jinkela_wire_329),
        .a(jinkela_wire_175),
        .c(jinkela_wire_337)
    );

    or_bb _398_ (
        .b(jinkela_wire_240),
        .a(jinkela_wire_134),
        .c(jinkela_wire_157)
    );

    and_bb _399_ (
        .b(jinkela_wire_240),
        .a(jinkela_wire_134),
        .c(jinkela_wire_205)
    );

    or_bb _400_ (
        .b(jinkela_wire_205),
        .a(jinkela_wire_255),
        .c(jinkela_wire_278)
    );

    and_bb _401_ (
        .b(jinkela_wire_205),
        .a(jinkela_wire_255),
        .c(jinkela_wire_435)
    );

    or_bb _402_ (
        .b(jinkela_wire_337),
        .a(jinkela_wire_348),
        .c(jinkela_wire_241)
    );

    and_bb _403_ (
        .b(jinkela_wire_337),
        .a(jinkela_wire_348),
        .c(jinkela_wire_20)
    );

    or_bb _404_ (
        .b(jinkela_wire_278),
        .a(jinkela_wire_241),
        .c(b_3_)
    );

    and_bb _405_ (
        .b(jinkela_wire_278),
        .a(jinkela_wire_241),
        .c(b_2_)
    );

    or_bb _406_ (
        .b(jinkela_wire_435),
        .a(jinkela_wire_20),
        .c(b_1_)
    );

    and_bb _407_ (
        .b(jinkela_wire_435),
        .a(jinkela_wire_20),
        .c(b_0_)
    );

    or_bb _408_ (
        .b(jinkela_wire_157),
        .a(jinkela_wire_281),
        .c(jinkela_wire_186)
    );

    and_bb _409_ (
        .b(jinkela_wire_157),
        .a(jinkela_wire_281),
        .c(jinkela_wire_333)
    );

    or_bb _410_ (
        .b(jinkela_wire_174),
        .a(jinkela_wire_44),
        .c(jinkela_wire_380)
    );

    and_bb _411_ (
        .b(jinkela_wire_174),
        .a(jinkela_wire_44),
        .c(jinkela_wire_145)
    );

    or_bb _412_ (
        .b(jinkela_wire_186),
        .a(jinkela_wire_380),
        .c(b_7_)
    );

    and_bb _413_ (
        .b(jinkela_wire_186),
        .a(jinkela_wire_380),
        .c(b_6_)
    );

    or_bb _414_ (
        .b(jinkela_wire_333),
        .a(jinkela_wire_145),
        .c(b_5_)
    );

    and_bb _415_ (
        .b(jinkela_wire_333),
        .a(jinkela_wire_145),
        .c(b_4_)
    );

    or_bb _416_ (
        .b(jinkela_wire_310),
        .a(jinkela_wire_397),
        .c(jinkela_wire_447)
    );

    and_bb _417_ (
        .b(jinkela_wire_310),
        .a(jinkela_wire_397),
        .c(jinkela_wire_125)
    );

    or_bb _418_ (
        .b(jinkela_wire_345),
        .a(jinkela_wire_393),
        .c(jinkela_wire_70)
    );

    and_bb _419_ (
        .b(jinkela_wire_345),
        .a(jinkela_wire_393),
        .c(jinkela_wire_89)
    );

    or_bb _420_ (
        .b(jinkela_wire_358),
        .a(jinkela_wire_226),
        .c(jinkela_wire_87)
    );

    and_bb _421_ (
        .b(jinkela_wire_358),
        .a(jinkela_wire_226),
        .c(jinkela_wire_379)
    );

    or_bb _422_ (
        .b(jinkela_wire_2),
        .a(jinkela_wire_195),
        .c(jinkela_wire_247)
    );

    and_bb _423_ (
        .b(jinkela_wire_2),
        .a(jinkela_wire_195),
        .c(jinkela_wire_57)
    );

    or_bb _424_ (
        .b(jinkela_wire_9),
        .a(jinkela_wire_126),
        .c(jinkela_wire_428)
    );

    and_bb _425_ (
        .b(jinkela_wire_9),
        .a(jinkela_wire_126),
        .c(jinkela_wire_72)
    );

    or_bb _426_ (
        .b(jinkela_wire_371),
        .a(jinkela_wire_197),
        .c(jinkela_wire_95)
    );

    and_bb _427_ (
        .b(jinkela_wire_371),
        .a(jinkela_wire_197),
        .c(jinkela_wire_137)
    );

    or_bb _428_ (
        .b(jinkela_wire_222),
        .a(jinkela_wire_110),
        .c(jinkela_wire_150)
    );

    or_bb _090_ (
        .b(jinkela_wire_80),
        .a(jinkela_wire_446),
        .c(jinkela_wire_214)
    );

    and_bb _091_ (
        .b(jinkela_wire_80),
        .a(jinkela_wire_446),
        .c(jinkela_wire_292)
    );

    or_bb _092_ (
        .b(jinkela_wire_53),
        .a(jinkela_wire_214),
        .c(jinkela_wire_220)
    );

    and_bb _093_ (
        .b(jinkela_wire_53),
        .a(jinkela_wire_214),
        .c(jinkela_wire_418)
    );

    or_bb _094_ (
        .b(jinkela_wire_171),
        .a(jinkela_wire_292),
        .c(jinkela_wire_398)
    );

    and_bb _095_ (
        .b(jinkela_wire_171),
        .a(jinkela_wire_292),
        .c(jinkela_wire_431)
    );

    or_bb _096_ (
        .b(jinkela_wire_297),
        .a(jinkela_wire_220),
        .c(jinkela_wire_409)
    );

    and_bb _097_ (
        .b(jinkela_wire_297),
        .a(jinkela_wire_220),
        .c(jinkela_wire_319)
    );

    or_bb _098_ (
        .b(jinkela_wire_273),
        .a(jinkela_wire_418),
        .c(jinkela_wire_306)
    );

    and_bb _099_ (
        .b(jinkela_wire_273),
        .a(jinkela_wire_418),
        .c(jinkela_wire_33)
    );

    or_bb _100_ (
        .b(jinkela_wire_361),
        .a(jinkela_wire_398),
        .c(jinkela_wire_129)
    );

    and_bb _101_ (
        .b(jinkela_wire_361),
        .a(jinkela_wire_398),
        .c(jinkela_wire_135)
    );

    or_bb _102_ (
        .b(jinkela_wire_302),
        .a(jinkela_wire_431),
        .c(jinkela_wire_5)
    );

    and_bb _103_ (
        .b(jinkela_wire_302),
        .a(jinkela_wire_431),
        .c(jinkela_wire_196)
    );

    or_bb _104_ (
        .b(jinkela_wire_206),
        .a(jinkela_wire_243),
        .c(jinkela_wire_86)
    );

    and_bb _105_ (
        .b(jinkela_wire_206),
        .a(jinkela_wire_243),
        .c(jinkela_wire_308)
    );

    or_bb _106_ (
        .b(jinkela_wire_445),
        .a(jinkela_wire_212),
        .c(jinkela_wire_336)
    );

    and_bb _107_ (
        .b(jinkela_wire_445),
        .a(jinkela_wire_212),
        .c(jinkela_wire_260)
    );

    or_bb _108_ (
        .b(jinkela_wire_190),
        .a(jinkela_wire_395),
        .c(jinkela_wire_102)
    );

    and_bb _109_ (
        .b(jinkela_wire_190),
        .a(jinkela_wire_395),
        .c(jinkela_wire_169)
    );

    or_bb _110_ (
        .b(jinkela_wire_381),
        .a(jinkela_wire_16),
        .c(jinkela_wire_303)
    );

    and_bb _111_ (
        .b(jinkela_wire_381),
        .a(jinkela_wire_16),
        .c(jinkela_wire_346)
    );

    or_bb _112_ (
        .b(jinkela_wire_86),
        .a(jinkela_wire_409),
        .c(jinkela_wire_239)
    );

    and_bb _113_ (
        .b(jinkela_wire_86),
        .a(jinkela_wire_409),
        .c(jinkela_wire_372)
    );

    or_bb _114_ (
        .b(jinkela_wire_336),
        .a(jinkela_wire_306),
        .c(jinkela_wire_394)
    );

    and_bb _115_ (
        .b(jinkela_wire_336),
        .a(jinkela_wire_306),
        .c(jinkela_wire_120)
    );

    or_bb _116_ (
        .b(jinkela_wire_102),
        .a(jinkela_wire_129),
        .c(jinkela_wire_406)
    );

    and_bb _117_ (
        .b(jinkela_wire_102),
        .a(jinkela_wire_129),
        .c(jinkela_wire_384)
    );

    or_bb _118_ (
        .b(jinkela_wire_303),
        .a(jinkela_wire_5),
        .c(jinkela_wire_128)
    );

    and_bb _119_ (
        .b(jinkela_wire_303),
        .a(jinkela_wire_5),
        .c(jinkela_wire_385)
    );

    or_bb _120_ (
        .b(jinkela_wire_385),
        .a(jinkela_wire_120),
        .c(jinkela_wire_316)
    );

    and_bb _121_ (
        .b(jinkela_wire_385),
        .a(jinkela_wire_120),
        .c(jinkela_wire_411)
    );

    or_bb _122_ (
        .b(jinkela_wire_384),
        .a(jinkela_wire_372),
        .c(jinkela_wire_417)
    );

    and_bb _123_ (
        .b(jinkela_wire_384),
        .a(jinkela_wire_372),
        .c(jinkela_wire_141)
    );

    or_bb _124_ (
        .b(jinkela_wire_316),
        .a(jinkela_wire_417),
        .c(jinkela_wire_338)
    );

    and_bb _125_ (
        .b(jinkela_wire_316),
        .a(jinkela_wire_417),
        .c(jinkela_wire_311)
    );

    or_bb _126_ (
        .b(jinkela_wire_411),
        .a(jinkela_wire_141),
        .c(jinkela_wire_386)
    );

    and_bb _127_ (
        .b(jinkela_wire_411),
        .a(jinkela_wire_141),
        .c(jinkela_wire_47)
    );

    or_bb _128_ (
        .b(jinkela_wire_128),
        .a(jinkela_wire_394),
        .c(jinkela_wire_81)
    );

    and_bb _129_ (
        .b(jinkela_wire_128),
        .a(jinkela_wire_394),
        .c(jinkela_wire_58)
    );

    or_bb _130_ (
        .b(jinkela_wire_406),
        .a(jinkela_wire_239),
        .c(jinkela_wire_46)
    );

    and_bb _131_ (
        .b(jinkela_wire_406),
        .a(jinkela_wire_239),
        .c(jinkela_wire_354)
    );

endmodule
