module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 );
  input G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 ;
  output G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 ;
  wire n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 ;
  assign n158 = G141 | G142 ;
  assign n159 = G139 | G140 ;
  assign n160 = n158 | n159 ;
  assign n161 = G121 | G2 ;
  assign n162 = G11 | n161 ;
  assign n163 = G115 & ~G74 ;
  assign n164 = G121 | G7 ;
  buffer buf_n165( .i (n164), .o (n165) );
  assign n166 = G119 | n165 ;
  assign n167 = G147 | n165 ;
  assign n168 = G53 & ~G96 ;
  assign n169 = G43 | G86 ;
  assign n170 = n168 & ~n169 ;
  buffer buf_n171( .i (n170), .o (n171) );
  assign n172 = ~G106 & G32 ;
  assign n173 = G64 | G76 ;
  assign n174 = n172 & ~n173 ;
  buffer buf_n175( .i (n174), .o (n175) );
  assign n176 = n171 | n175 ;
  buffer buf_n177( .i (n176), .o (n177) );
  assign n178 = G147 & ~n175 ;
  assign n179 = G119 & ~n171 ;
  assign n180 = n178 | n179 ;
  buffer buf_n181( .i (n180), .o (n181) );
  assign n182 = G145 | G146 ;
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n198 = G109 & ~n186 ;
  assign n199 = G79 & ~n186 ;
  assign n200 = n198 | n199 ;
  assign n201 = G89 & ~n186 ;
  buffer buf_n202( .i (n185), .o (n202) );
  assign n203 = G99 & ~n202 ;
  assign n204 = n201 | n203 ;
  assign n205 = n200 | n204 ;
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  assign n222 = G108 | n196 ;
  assign n223 = G98 & ~n196 ;
  assign n224 = n222 & ~n223 ;
  assign n225 = G88 & ~n196 ;
  buffer buf_n226( .i (n195), .o (n226) );
  assign n227 = G78 & ~n226 ;
  assign n228 = n225 | n227 ;
  assign n229 = n224 & ~n228 ;
  buffer buf_n230( .i (n229), .o (n230) );
  assign n233 = G80 | n202 ;
  assign n234 = G90 & ~n202 ;
  assign n235 = n233 & ~n234 ;
  assign n236 = G100 & ~n202 ;
  buffer buf_n237( .i (n185), .o (n237) );
  assign n238 = G110 & ~n237 ;
  assign n239 = n236 | n238 ;
  assign n240 = n235 & ~n239 ;
  buffer buf_n241( .i (n240), .o (n241) );
  assign n253 = G117 & ~G36 ;
  assign n254 = G117 & ~G68 ;
  assign n255 = G120 | n254 ;
  assign n256 = n253 & ~n255 ;
  assign n257 = G117 | G120 ;
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  assign n272 = G46 & ~n263 ;
  assign n273 = G57 & ~n263 ;
  assign n274 = n272 | n273 ;
  assign n275 = n256 & ~n274 ;
  buffer buf_n276( .i (n275), .o (n276) );
  assign n278 = G117 & ~G37 ;
  assign n279 = G117 & ~G69 ;
  assign n280 = G120 | n279 ;
  assign n281 = n278 & ~n280 ;
  assign n282 = G47 & ~n262 ;
  assign n283 = G58 & ~n262 ;
  assign n284 = n282 | n283 ;
  assign n285 = n281 & ~n284 ;
  buffer buf_n286( .i (n285), .o (n286) );
  assign n296 = G117 & ~G38 ;
  assign n297 = G117 & ~G70 ;
  assign n298 = G120 | n297 ;
  assign n299 = n296 & ~n298 ;
  assign n300 = G48 & ~n262 ;
  buffer buf_n301( .i (n261), .o (n301) );
  assign n302 = G59 & ~n301 ;
  assign n303 = n300 | n302 ;
  assign n304 = n299 & ~n303 ;
  buffer buf_n305( .i (n304), .o (n305) );
  assign n315 = G117 & ~G31 ;
  assign n316 = G117 & ~G63 ;
  assign n317 = G120 | n316 ;
  assign n318 = n315 & ~n317 ;
  assign n319 = G42 & ~n261 ;
  assign n320 = G52 & ~n261 ;
  assign n321 = n319 | n320 ;
  assign n322 = n318 & ~n321 ;
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  assign n336 = G122 | n335 ;
  assign n337 = G116 | G121 ;
  assign n338 = n181 | n337 ;
  buffer buf_n339( .i (n338), .o (n339) );
  assign n340 = G28 | n339 ;
  assign n341 = G1 & ~G3 ;
  assign n342 = n339 | n341 ;
  assign n343 = G117 | G39 ;
  assign n344 = G117 & ~G71 ;
  assign n345 = G120 | n344 ;
  assign n346 = n343 & ~n345 ;
  buffer buf_n347( .i (n260), .o (n347) );
  assign n348 = G49 & ~n347 ;
  assign n349 = G60 & ~n347 ;
  assign n350 = n348 | n349 ;
  assign n351 = n346 | n350 ;
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  assign n363 = G56 & ~n266 ;
  assign n364 = G117 | G35 ;
  assign n365 = G117 & ~G67 ;
  assign n366 = G120 | n365 ;
  assign n367 = n364 & ~n366 ;
  assign n368 = n363 & ~n367 ;
  buffer buf_n369( .i (n368), .o (n369) );
  assign n371 = G117 & ~G34 ;
  assign n372 = G117 & ~G66 ;
  assign n373 = G120 | n372 ;
  assign n374 = n371 & ~n373 ;
  assign n375 = G45 & ~n263 ;
  buffer buf_n376( .i (n301), .o (n376) );
  assign n377 = G55 & ~n376 ;
  assign n378 = n375 | n377 ;
  assign n379 = n374 & ~n378 ;
  buffer buf_n380( .i (n379), .o (n380) );
  assign n387 = G117 & ~G33 ;
  assign n388 = G117 & ~G65 ;
  assign n389 = G120 | n388 ;
  assign n390 = n387 & ~n389 ;
  assign n391 = G44 & ~n376 ;
  assign n392 = G54 & ~n376 ;
  assign n393 = n391 | n392 ;
  assign n394 = n390 & ~n393 ;
  buffer buf_n395( .i (n394), .o (n395) );
  assign n399 = G117 & ~G40 ;
  assign n400 = G117 & ~G72 ;
  assign n401 = G120 | n400 ;
  assign n402 = n399 & ~n401 ;
  assign n403 = G50 & ~n347 ;
  assign n404 = G61 & ~n347 ;
  assign n405 = n403 | n404 ;
  assign n406 = n402 & ~n405 ;
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  assign n420 = G123 | n417 ;
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  assign n421 = G123 & ~n314 ;
  assign n422 = n420 & ~n421 ;
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  assign n424 = G123 | n362 ;
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  assign n425 = ~G123 & n295 ;
  assign n426 = n424 & ~n425 ;
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  assign n428 = G118 & ~G122 ;
  assign n429 = n419 | n428 ;
  assign n430 = G123 & ~n333 ;
  assign n431 = G118 | G123 ;
  assign n432 = n417 & ~n431 ;
  assign n433 = n430 | n432 ;
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n197( .i (n196), .o (n197) );
  assign n435 = G77 & ~n197 ;
  assign n436 = G97 & ~n197 ;
  assign n437 = n435 & ~n436 ;
  assign n438 = G107 & ~n197 ;
  assign n439 = G87 & ~n197 ;
  assign n440 = n438 | n439 ;
  assign n441 = n437 & ~n440 ;
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  assign n450 = G143 | n449 ;
  assign n451 = G143 & ~n449 ;
  assign n452 = n450 & ~n451 ;
  assign n453 = G144 | n452 ;
  assign n454 = ~G19 & G23 ;
  buffer buf_n455( .i (n226), .o (n455) );
  assign n456 = G75 & ~n455 ;
  assign n457 = G85 & ~n455 ;
  assign n458 = n456 & ~n457 ;
  assign n459 = G95 & ~n455 ;
  assign n460 = G105 & ~n455 ;
  assign n461 = n459 | n460 ;
  assign n462 = n458 & ~n461 ;
  buffer buf_n463( .i (n462), .o (n463) );
  assign n465 = G23 & ~n463 ;
  assign n466 = n454 & ~n465 ;
  assign n467 = G135 & ~n466 ;
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  assign n471 = G12 & ~G13 ;
  assign n472 = G12 & ~n325 ;
  assign n473 = n471 & ~n472 ;
  assign n474 = G125 & ~n473 ;
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  assign n478 = G12 & ~G15 ;
  assign n479 = ~G12 & n287 ;
  assign n480 = n478 & ~n479 ;
  assign n481 = G130 & ~n480 ;
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  assign n485 = n477 | n484 ;
  assign n486 = n470 | n485 ;
  assign n487 = G12 & ~G5 ;
  assign n488 = G12 & ~n306 ;
  assign n489 = n487 & ~n488 ;
  assign n490 = G129 & ~n489 ;
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  assign n493 = ~G21 & G23 ;
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  assign n494 = G23 & ~n252 ;
  assign n495 = n493 & ~n494 ;
  assign n496 = G140 & ~n495 ;
  buffer buf_n497( .i (n496), .o (n497) );
  assign n498 = n492 | n497 ;
  assign n499 = G23 & ~G27 ;
  assign n500 = G23 & ~n230 ;
  assign n501 = n499 & ~n500 ;
  assign n502 = G142 & ~n501 ;
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  assign n505 = n468 | n504 ;
  assign n506 = n498 | n505 ;
  assign n507 = G12 & ~G14 ;
  assign n508 = ~G12 & n354 ;
  assign n509 = n507 & ~n508 ;
  assign n510 = G128 & ~n509 ;
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  assign n513 = G12 & ~G4 ;
  assign n514 = G12 & ~n409 ;
  assign n515 = n513 & ~n514 ;
  assign n516 = G126 & ~n515 ;
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  assign n519 = n512 | n518 ;
  assign n520 = G23 & ~G26 ;
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  assign n521 = G23 & ~n216 ;
  assign n522 = n520 & ~n521 ;
  assign n523 = G141 & ~n522 ;
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  assign n526 = n497 | n525 ;
  assign n527 = n519 | n526 ;
  assign n528 = n506 | n527 ;
  assign n529 = n486 | n528 ;
  assign n530 = G23 & ~G24 ;
  buffer buf_n531( .i (n226), .o (n531) );
  assign n532 = G93 & ~n531 ;
  assign n533 = G103 & ~n531 ;
  assign n534 = n532 & ~n533 ;
  assign n535 = G113 & ~n531 ;
  assign n536 = G83 & ~n531 ;
  assign n537 = n535 | n536 ;
  assign n538 = n534 & ~n537 ;
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  assign n541 = G23 & ~n540 ;
  assign n542 = n530 & ~n541 ;
  buffer buf_n543( .i (n542), .o (n543) );
  assign n544 = G136 | n543 ;
  assign n545 = G136 & ~n543 ;
  assign n546 = n544 & ~n545 ;
  assign n547 = G12 & ~G16 ;
  buffer buf_n277( .i (n276), .o (n277) );
  assign n548 = G12 & ~n277 ;
  assign n549 = n547 & ~n548 ;
  buffer buf_n550( .i (n549), .o (n550) );
  assign n551 = G131 | n550 ;
  assign n552 = G131 & ~n550 ;
  assign n553 = n551 & ~n552 ;
  assign n554 = ~G20 & G23 ;
  buffer buf_n555( .i (n226), .o (n555) );
  assign n556 = G82 & ~n555 ;
  assign n557 = G102 & ~n555 ;
  assign n558 = n556 & ~n557 ;
  assign n559 = G112 & ~n555 ;
  assign n560 = G92 & ~n555 ;
  assign n561 = n559 | n560 ;
  assign n562 = n558 & ~n561 ;
  buffer buf_n563( .i (n562), .o (n563) );
  assign n566 = G23 & ~n563 ;
  assign n567 = n554 & ~n566 ;
  buffer buf_n568( .i (n567), .o (n568) );
  assign n569 = G138 | n568 ;
  assign n570 = G138 & ~n568 ;
  assign n571 = n569 & ~n570 ;
  assign n572 = n553 | n571 ;
  assign n573 = n546 | n572 ;
  assign n574 = G23 & ~G25 ;
  buffer buf_n575( .i (n195), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  assign n577 = G81 & ~n576 ;
  assign n578 = G101 & ~n576 ;
  assign n579 = n577 & ~n578 ;
  assign n580 = G111 & ~n576 ;
  assign n581 = G91 & ~n576 ;
  assign n582 = n580 | n581 ;
  assign n583 = n579 & ~n582 ;
  assign n584 = G23 & ~n583 ;
  assign n585 = n574 & ~n584 ;
  assign n586 = G139 & ~n585 ;
  buffer buf_n587( .i (n586), .o (n587) );
  assign n588 = n482 | n587 ;
  assign n589 = G12 & ~G18 ;
  assign n590 = G12 & ~n395 ;
  assign n591 = n589 & ~n590 ;
  assign n592 = G134 & ~n591 ;
  buffer buf_n593( .i (n592), .o (n593) );
  assign n594 = n517 | n593 ;
  assign n595 = n588 | n594 ;
  assign n596 = G12 & ~G6 ;
  assign n597 = G12 & ~n380 ;
  assign n598 = n596 & ~n597 ;
  assign n599 = G133 & ~n598 ;
  buffer buf_n600( .i (n599), .o (n600) );
  assign n601 = G23 & ~n443 ;
  assign n602 = ~G22 & G23 ;
  assign n603 = G9 | n602 ;
  assign n604 = n601 | n603 ;
  assign n605 = n600 | n604 ;
  assign n606 = n503 | n600 ;
  assign n607 = n605 | n606 ;
  assign n608 = n595 | n607 ;
  assign n609 = n491 | n524 ;
  assign n610 = n475 | n511 ;
  assign n611 = n609 | n610 ;
  assign n612 = n587 | n593 ;
  assign n613 = G12 & ~G17 ;
  assign n614 = G12 & ~n369 ;
  assign n615 = n613 & ~n614 ;
  assign n616 = G132 & ~n615 ;
  assign n617 = n612 | n616 ;
  assign n618 = n611 | n617 ;
  assign n619 = n608 | n618 ;
  assign n620 = n573 | n619 ;
  assign n621 = n529 | n620 ;
  buffer buf_n622( .i (n621), .o (n622) );
  assign n623 = G117 & ~G41 ;
  assign n624 = G117 & ~G73 ;
  assign n625 = G120 | n624 ;
  assign n626 = n623 & ~n625 ;
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  assign n627 = G51 & ~n271 ;
  assign n628 = G62 & ~n271 ;
  assign n629 = n627 | n628 ;
  assign n630 = n626 & ~n629 ;
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  assign n633 = G122 & ~n632 ;
  assign n634 = G122 | n633 ;
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  assign n635 = n232 | n443 ;
  assign n636 = n232 & ~n443 ;
  assign n637 = n635 & ~n636 ;
  buffer buf_n638( .i (n637), .o (n638) );
  assign n639 = n221 | n638 ;
  assign n640 = ~n221 & n638 ;
  assign n641 = n639 & ~n640 ;
  assign n642 = G29 | n641 ;
  buffer buf_n643( .i (n642), .o (n643) );
  inverter inv_n789( .i (n643), .o (n789) );
  assign n644 = G123 & ~n631 ;
  assign n645 = G123 | n644 ;
  buffer buf_n646( .i (n645), .o (n646) );
  assign n647 = G127 | n241 ;
  buffer buf_n648( .i (n647), .o (n648) );
  assign n649 = G30 | n206 ;
  buffer buf_n650( .i (n649), .o (n650) );
  assign n651 = n648 | n650 ;
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  assign n657 = ~G8 & n654 ;
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  assign n668 = ~G133 & n667 ;
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  assign n669 = G8 | n654 ;
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  assign n679 = n386 | n678 ;
  assign n680 = ~G132 & n665 ;
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  assign n681 = G129 & n656 ;
  assign n682 = G140 & ~n656 ;
  assign n683 = n681 & ~n682 ;
  assign n684 = n306 & ~n683 ;
  buffer buf_n685( .i (n684), .o (n685) );
  assign n686 = ~G128 & n653 ;
  assign n687 = G139 & ~n653 ;
  assign n688 = n686 | n687 ;
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  assign n692 = ~n354 & n691 ;
  assign n693 = ~G126 & n653 ;
  buffer buf_n694( .i (n652), .o (n694) );
  assign n695 = G138 & ~n694 ;
  assign n696 = n693 | n695 ;
  buffer buf_n697( .i (n696), .o (n697) );
  assign n698 = n407 | n697 ;
  assign n699 = ~G125 & n654 ;
  buffer buf_n700( .i (n694), .o (n700) );
  assign n701 = G136 & ~n700 ;
  assign n702 = n699 | n701 ;
  assign n703 = ~n323 & n702 ;
  assign n704 = n698 & n703 ;
  assign n705 = n407 & n697 ;
  assign n706 = n352 & n689 ;
  assign n707 = n705 | n706 ;
  assign n708 = n704 | n707 ;
  assign n709 = ~n692 & n708 ;
  assign n710 = n685 | n709 ;
  assign n711 = G8 & ~n286 ;
  assign n712 = G130 & n658 ;
  assign n713 = G141 & ~n670 ;
  assign n714 = n712 & ~n713 ;
  assign n715 = n711 & ~n714 ;
  buffer buf_n716( .i (n715), .o (n716) );
  assign n718 = n685 | n716 ;
  assign n719 = n710 & ~n718 ;
  buffer buf_n717( .i (n716), .o (n717) );
  assign n720 = G8 & ~n276 ;
  assign n721 = G131 & n659 ;
  assign n722 = G142 & ~n671 ;
  assign n723 = n721 & ~n722 ;
  assign n724 = n720 & ~n723 ;
  buffer buf_n725( .i (n724), .o (n725) );
  assign n727 = n717 | n725 ;
  assign n728 = n719 | n727 ;
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n370( .i (n369), .o (n370) );
  assign n729 = n370 & ~n675 ;
  assign n730 = n726 | n729 ;
  assign n731 = n728 & ~n730 ;
  assign n732 = n680 | n731 ;
  assign n733 = n679 & n732 ;
  assign n734 = n668 | n733 ;
  assign n735 = n648 & ~n650 ;
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  assign n748 = G136 | n539 ;
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  assign n752 = n747 & ~n751 ;
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  assign n753 = G138 | n565 ;
  assign n754 = n746 & ~n753 ;
  buffer buf_n755( .i (n754), .o (n755) );
  assign n759 = n752 & ~n755 ;
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n464( .i (n463), .o (n464) );
  assign n761 = G135 | n464 ;
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  assign n765 = G134 & ~n398 ;
  assign n766 = n762 & ~n765 ;
  assign n767 = n747 & ~n766 ;
  assign n768 = n755 | n767 ;
  assign n769 = G135 & ~n464 ;
  assign n770 = n749 & ~n769 ;
  assign n771 = n746 & ~n770 ;
  buffer buf_n772( .i (n771), .o (n772) );
  assign n774 = G134 | n398 ;
  assign n775 = n746 & ~n774 ;
  buffer buf_n776( .i (n775), .o (n776) );
  assign n777 = n772 | n776 ;
  assign n778 = n768 | n777 ;
  assign n779 = n760 & ~n778 ;
  assign n780 = n734 & n779 ;
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  assign n781 = n764 & ~n776 ;
  assign n782 = n773 & ~n781 ;
  assign n783 = n760 & ~n782 ;
  assign n784 = n758 | n783 ;
  assign n785 = ~n780 & ~n784 ;
  assign n786 = G10 & ~n181 ;
  assign n787 = n643 & n786 ;
  inverter inv_n788( .i (n787), .o (n788) );
  assign G2531 = G115 ;
  assign G2532 = G115 ;
  assign G2533 = G115 ;
  assign G2534 = G124 ;
  assign G2535 = G124 ;
  assign G2536 = G137 ;
  assign G2537 = G137 ;
  assign G2538 = G137 ;
  assign G2539 = G32 ;
  assign G2540 = G106 ;
  assign G2541 = G64 ;
  assign G2542 = G76 ;
  assign G2543 = G53 ;
  assign G2544 = G96 ;
  assign G2545 = G43 ;
  assign G2546 = G86 ;
  assign G2547 = n160 ;
  assign G2548 = n162 ;
  assign G2549 = G115 ;
  assign G2550 = n163 ;
  assign G2551 = n165 ;
  assign G2552 = n166 ;
  assign G2553 = n167 ;
  assign G2554 = n177 ;
  assign G2555 = n177 ;
  assign G2556 = n181 ;
  assign G2557 = n206 ;
  assign G2558 = n230 ;
  assign G2559 = n241 ;
  assign G2560 = n276 ;
  assign G2561 = n286 ;
  assign G2562 = n305 ;
  assign G2563 = n336 ;
  assign G2564 = n340 ;
  assign G2565 = n342 ;
  assign G2566 = n352 ;
  assign G2567 = n305 ;
  assign G2568 = n286 ;
  assign G2569 = n276 ;
  assign G2570 = n369 ;
  assign G2571 = n380 ;
  assign G2572 = n395 ;
  assign G2573 = n423 ;
  assign G2574 = n423 ;
  assign G2575 = n427 ;
  assign G2576 = n427 ;
  assign G2577 = n429 ;
  assign G2578 = n434 ;
  assign G2579 = n434 ;
  assign G2580 = n453 ;
  assign G2581 = ~G10 ;
  assign G2582 = 1'b0 ;
  assign G2583 = 1'b0 ;
  assign G2584 = n622 ;
  assign G2585 = n622 ;
  assign G2586 = n634 ;
  assign G2587 = n789 ;
  assign G2588 = n646 ;
  assign G2589 = n646 ;
  assign G2590 = 1'b0 ;
  assign G2591 = n785 ;
  assign G2592 = 1'b0 ;
  assign G2593 = n788 ;
  assign G2594 = n788 ;
endmodule
