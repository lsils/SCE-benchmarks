module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 , y1 , y2 , y3 , y4 , y5 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 , y1 , y2 , y3 , y4 , y5 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 ;
  buffer buf_n10( .i (x0), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n34( .i (x1), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n103( .i (x4), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n149( .i (x6), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n126( .i (x5), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n172( .i (x7), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  assign n218 = n137 & n183 ;
  buffer buf_n219( .i (n218), .o (n219) );
  assign n220 = ( ~n116 & n162 ) | ( ~n116 & n219 ) | ( n162 & n219 ) ;
  assign n221 = n117 & n220 ;
  buffer buf_n59( .i (x2), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n81( .i (x3), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  assign n222 = n70 & n92 ;
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  assign n228 = ( n25 & n221 ) | ( n25 & n225 ) | ( n221 & n225 ) ;
  assign n229 = n50 & ~n228 ;
  assign n230 = ( n27 & n51 ) | ( n27 & ~n229 ) | ( n51 & ~n229 ) ;
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  assign n239 = ( n74 & ~n164 ) | ( n74 & n187 ) | ( ~n164 & n187 ) ;
  buffer buf_n240( .i (n239), .o (n240) );
  assign n241 = ( n98 & n189 ) | ( n98 & ~n240 ) | ( n189 & ~n240 ) ;
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  assign n242 = ( ~n76 & n98 ) | ( ~n76 & n240 ) | ( n98 & n240 ) ;
  assign n243 = n241 & ~n242 ;
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  assign n246 = n53 & n145 ;
  assign n247 = ( n123 & ~n244 ) | ( n123 & n246 ) | ( ~n244 & n246 ) ;
  assign n248 = n245 & n247 ;
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  assign n251 = n33 & n249 ;
  assign n252 = ~n16 & n65 ;
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  assign n267 = n45 & n256 ;
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  assign n278 = n139 & ~n162 ;
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  assign n285 = n123 & n284 ;
  assign n286 = ( n102 & ~n276 ) | ( n102 & n285 ) | ( ~n276 & n285 ) ;
  assign n287 = n277 & n286 ;
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  assign n288 = ~n17 & n41 ;
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  assign n299 = n44 & ~n91 ;
  buffer buf_n300( .i (n299), .o (n300) );
  assign n306 = ( n22 & n71 ) | ( n22 & n300 ) | ( n71 & n300 ) ;
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  assign n309 = ( ~n73 & n95 ) | ( ~n73 & n307 ) | ( n95 & n307 ) ;
  assign n310 = ( n49 & n308 ) | ( n49 & n309 ) | ( n308 & n309 ) ;
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  assign n313 = n73 & ~n117 ;
  buffer buf_n314( .i (n313), .o (n314) );
  assign n315 = n97 & n314 ;
  assign n316 = n311 | n315 ;
  assign n317 = ( n298 & n312 ) | ( n298 & n316 ) | ( n312 & n316 ) ;
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  assign n321 = ( n23 & n47 ) | ( n23 & n139 ) | ( n47 & n139 ) ;
  assign n322 = ( n48 & ~n95 ) | ( n48 & n321 ) | ( ~n95 & n321 ) ;
  buffer buf_n323( .i (n322), .o (n323) );
  assign n326 = n50 & ~n323 ;
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  assign n329 = n325 | n327 ;
  assign n330 = ( ~n53 & n328 ) | ( ~n53 & n329 ) | ( n328 & n329 ) ;
  assign n331 = ( n79 & n318 ) | ( n79 & n330 ) | ( n318 & n330 ) ;
  assign n332 = n124 & ~n331 ;
  assign n333 = ( n125 & n320 ) | ( n125 & ~n332 ) | ( n320 & ~n332 ) ;
  assign n334 = n287 | n333 ;
  assign n335 = ( n250 & ~n251 ) | ( n250 & n334 ) | ( ~n251 & n334 ) ;
  buffer buf_n336( .i (n335), .o (n336) );
  assign n337 = n160 | n183 ;
  buffer buf_n338( .i (n337), .o (n338) );
  assign n340 = n139 | n338 ;
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  assign n344 = n120 & ~n343 ;
  assign n345 = ( n28 & n77 ) | ( n28 & n344 ) | ( n77 & n344 ) ;
  assign n346 = ~n29 & n345 ;
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  assign n349 = n162 & n219 ;
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  assign n355 = n28 & ~n121 ;
  assign n356 = ( n78 & n354 ) | ( n78 & n355 ) | ( n354 & n355 ) ;
  assign n357 = ~n79 & n356 ;
  assign n358 = ~n347 & n357 ;
  buffer buf_n193( .i (x8), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n359 = ~n102 & n214 ;
  assign n360 = ( n348 & n358 ) | ( n348 & n359 ) | ( n358 & n359 ) ;
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  assign n363 = ~n58 & n361 ;
  assign n364 = ( n69 & ~n91 ) | ( n69 & n159 ) | ( ~n91 & n159 ) ;
  buffer buf_n365( .i (n364), .o (n365) );
  assign n370 = ( n46 & ~n161 ) | ( n46 & n365 ) | ( ~n161 & n365 ) ;
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  assign n375 = ( n73 & ~n95 ) | ( n73 & n371 ) | ( ~n95 & n371 ) ;
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  assign n378 = ~n369 & n376 ;
  assign n379 = ( ~n374 & n377 ) | ( ~n374 & n378 ) | ( n377 & n378 ) ;
  assign n380 = n121 & n379 ;
  assign n381 = n29 | n380 ;
  buffer buf_n382( .i (n72), .o (n382) );
  assign n383 = n48 | n382 ;
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n389( .i (n161), .o (n389) );
  assign n390 = ~n116 & n389 ;
  buffer buf_n391( .i (n390), .o (n391) );
  assign n394 = n96 & n391 ;
  assign n395 = ~n384 & n394 ;
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  assign n398 = n29 & ~n397 ;
  assign n399 = n381 & ~n398 ;
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  assign n402 = ~n148 & n400 ;
  assign n403 = ~n91 & n113 ;
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  assign n414 = ~n133 & n156 ;
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  assign n427 = n275 & n426 ;
  assign n428 = n413 & n427 ;
  assign n429 = ( n72 & n94 ) | ( n72 & ~n116 ) | ( n94 & ~n116 ) ;
  buffer buf_n430( .i (n429), .o (n430) );
  assign n434 = ( n25 & ~n96 ) | ( n25 & n430 ) | ( ~n96 & n430 ) ;
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  assign n438 = ( ~n76 & n98 ) | ( ~n76 & n435 ) | ( n98 & n435 ) ;
  assign n439 = n433 & ~n438 ;
  buffer buf_n440( .i (n28), .o (n440) );
  assign n441 = ( ~n437 & n439 ) | ( ~n437 & n440 ) | ( n439 & n440 ) ;
  buffer buf_n442( .i (n94), .o (n442) );
  assign n443 = ( n140 & ~n382 ) | ( n140 & n442 ) | ( ~n382 & n442 ) ;
  buffer buf_n444( .i (n443), .o (n444) );
  assign n446 = n65 & ~n132 ;
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  assign n455 = ( n49 & n96 ) | ( n49 & ~n454 ) | ( n96 & ~n454 ) ;
  assign n456 = ~n444 & n455 ;
  assign n457 = ( n27 & n120 ) | ( n27 & n456 ) | ( n120 & n456 ) ;
  assign n458 = n19 & ~n43 ;
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n467( .i (n442), .o (n467) );
  assign n468 = ( n454 & n463 ) | ( n454 & n467 ) | ( n463 & n467 ) ;
  assign n469 = ~n97 & n468 ;
  assign n470 = n120 & n469 ;
  buffer buf_n471( .i (n27), .o (n471) );
  assign n472 = ( n457 & n470 ) | ( n457 & ~n471 ) | ( n470 & ~n471 ) ;
  buffer buf_n473( .i (n472), .o (n473) );
  assign n474 = ( ~n54 & n441 ) | ( ~n54 & n473 ) | ( n441 & n473 ) ;
  assign n475 = ~n22 & n115 ;
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  assign n482 = ( n77 & n99 ) | ( n77 & n471 ) | ( n99 & n471 ) ;
  buffer buf_n483( .i (n26), .o (n483) );
  buffer buf_n484( .i (n119), .o (n484) );
  assign n485 = ( n76 & n483 ) | ( n76 & ~n484 ) | ( n483 & ~n484 ) ;
  assign n486 = n99 | n485 ;
  assign n487 = ( n481 & ~n482 ) | ( n481 & n486 ) | ( ~n482 & n486 ) ;
  assign n488 = ( n54 & n473 ) | ( n54 & ~n487 ) | ( n473 & ~n487 ) ;
  assign n489 = n474 | n488 ;
  assign n490 = n428 | n489 ;
  assign n491 = ( n401 & ~n402 ) | ( n401 & n490 ) | ( ~n402 & n490 ) ;
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  assign n492 = ~n161 & n184 ;
  buffer buf_n493( .i (n492), .o (n493) );
  assign n494 = ( n117 & n140 ) | ( n117 & n493 ) | ( n140 & n493 ) ;
  assign n495 = ~n118 & n494 ;
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n503( .i (n97), .o (n503) );
  assign n504 = n496 & n503 ;
  assign n505 = ( n77 & n466 ) | ( n77 & n504 ) | ( n466 & n504 ) ;
  assign n506 = ~n78 & n505 ;
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n90), .o (n510) );
  assign n511 = ( ~n136 & n182 ) | ( ~n136 & n510 ) | ( n182 & n510 ) ;
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n160), .o (n513) );
  assign n514 = ( n93 & n512 ) | ( n93 & ~n513 ) | ( n512 & ~n513 ) ;
  buffer buf_n515( .i (n514), .o (n515) );
  assign n518 = n442 & ~n515 ;
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  assign n521 = n517 | n519 ;
  assign n522 = ( ~n503 & n520 ) | ( ~n503 & n521 ) | ( n520 & n521 ) ;
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  assign n525 = ( n78 & n122 ) | ( n78 & ~n523 ) | ( n122 & ~n523 ) ;
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  assign n526 = n68 | n90 ;
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  assign n533 = n142 & ~n532 ;
  assign n534 = ( n166 & n189 ) | ( n166 & n533 ) | ( n189 & n533 ) ;
  assign n535 = ~n190 & n534 ;
  assign n536 = n122 & n535 ;
  assign n537 = ( n524 & n525 ) | ( n524 & n536 ) | ( n525 & n536 ) ;
  assign n538 = ( ~n31 & n507 ) | ( ~n31 & n537 ) | ( n507 & n537 ) ;
  assign n539 = n56 & ~n538 ;
  assign n540 = ( n57 & n509 ) | ( n57 & ~n539 ) | ( n509 & ~n539 ) ;
  assign n541 = n491 | n540 ;
  assign n542 = ( n362 & ~n363 ) | ( n362 & n541 ) | ( ~n363 & n541 ) ;
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  assign n543 = ( ~n70 & n92 ) | ( ~n70 & n114 ) | ( n92 & n114 ) ;
  assign n544 = ( ~n71 & n138 ) | ( ~n71 & n543 ) | ( n138 & n543 ) ;
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n115), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  assign n550 = ( n140 & ~n545 ) | ( n140 & n549 ) | ( ~n545 & n549 ) ;
  assign n551 = n467 & n550 ;
  assign n552 = ( n75 & n547 ) | ( n75 & ~n551 ) | ( n547 & ~n551 ) ;
  assign n553 = n483 & ~n552 ;
  assign n554 = n141 & n467 ;
  buffer buf_n555( .i (n467), .o (n555) );
  assign n556 = ( n314 & n554 ) | ( n314 & ~n555 ) | ( n554 & ~n555 ) ;
  assign n557 = n483 | n556 ;
  assign n558 = ( ~n471 & n553 ) | ( ~n471 & n557 ) | ( n553 & n557 ) ;
  assign n559 = n53 & ~n558 ;
  buffer buf_n560( .i (n138), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  assign n562 = ( n442 & n549 ) | ( n442 & n561 ) | ( n549 & n561 ) ;
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n94), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  assign n567 = ( n25 & ~n118 ) | ( n25 & n566 ) | ( ~n118 & n566 ) ;
  assign n568 = n563 | n567 ;
  assign n569 = ( ~n143 & n564 ) | ( ~n143 & n568 ) | ( n564 & n568 ) ;
  buffer buf_n570( .i (n75), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  assign n572 = ~n569 & n571 ;
  buffer buf_n573( .i (n52), .o (n573) );
  assign n574 = n572 | n573 ;
  assign n575 = ~n559 & n574 ;
  assign n576 = n115 & n138 ;
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  assign n581 = n555 & ~n579 ;
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n580( .i (n579), .o (n580) );
  assign n584 = ( n51 & n503 ) | ( n51 & ~n580 ) | ( n503 & ~n580 ) ;
  assign n585 = ~n582 & n584 ;
  assign n586 = ( n100 & ~n583 ) | ( n100 & n585 ) | ( ~n583 & n585 ) ;
  assign n587 = ( ~n30 & n79 ) | ( ~n30 & n586 ) | ( n79 & n586 ) ;
  assign n588 = ( ~n266 & n575 ) | ( ~n266 & n587 ) | ( n575 & n587 ) ;
  assign n589 = ~n45 & n70 ;
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n80( .i (n79), .o (n80) );
  assign n600 = ( n23 & n548 ) | ( n23 & n560 ) | ( n548 & n560 ) ;
  buffer buf_n601( .i (n600), .o (n601) );
  assign n606 = ( ~n141 & n566 ) | ( ~n141 & n601 ) | ( n566 & n601 ) ;
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  assign n611 = ( n483 & n484 ) | ( n483 & n607 ) | ( n484 & n607 ) ;
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  assign n614 = ~n605 & n612 ;
  assign n615 = ( ~n610 & n613 ) | ( ~n610 & n614 ) | ( n613 & n614 ) ;
  assign n616 = ( ~n55 & n80 ) | ( ~n55 & n615 ) | ( n80 & n615 ) ;
  assign n617 = ( n588 & ~n599 ) | ( n588 & n616 ) | ( ~n599 & n616 ) ;
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  assign n620 = n184 & n205 ;
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  assign n628 = ~n169 & n627 ;
  assign n629 = ( n124 & n147 ) | ( n124 & n628 ) | ( n147 & n628 ) ;
  assign n630 = ~n125 & n629 ;
  assign n631 = n157 | n201 ;
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  assign n634 = ( ~n137 & n183 ) | ( ~n137 & n633 ) | ( n183 & n633 ) ;
  buffer buf_n635( .i (n137), .o (n635) );
  assign n636 = n634 | n635 ;
  assign n637 = n548 & ~n636 ;
  assign n638 = ( ~n294 & n382 ) | ( ~n294 & n637 ) | ( n382 & n637 ) ;
  assign n639 = n295 & n638 ;
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  assign n643 = ~n157 & n201 ;
  assign n644 = ~n181 & n643 ;
  assign n645 = ~n136 & n644 ;
  buffer buf_n646( .i (n69), .o (n646) );
  assign n647 = ( n45 & n645 ) | ( n45 & n646 ) | ( n645 & n646 ) ;
  assign n648 = ~n46 & n647 ;
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  assign n652 = ~n71 & n635 ;
  assign n653 = n47 & n652 ;
  assign n654 = n177 & ~n198 ;
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  assign n666 = ( n649 & n653 ) | ( n649 & n662 ) | ( n653 & n662 ) ;
  assign n667 = n164 & ~n666 ;
  assign n668 = ( n165 & n651 ) | ( n165 & ~n667 ) | ( n651 & ~n667 ) ;
  assign n669 = ( ~n484 & n640 ) | ( ~n484 & n668 ) | ( n640 & n668 ) ;
  assign n670 = n471 & ~n669 ;
  assign n671 = ( n440 & n642 ) | ( n440 & ~n670 ) | ( n642 & ~n670 ) ;
  assign n672 = ~n101 & n671 ;
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  assign n675 = n20 | n44 ;
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  assign n685 = ~n69 & n510 ;
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  assign n695 = ~n684 & n694 ;
  buffer buf_n696( .i (n695), .o (n696) );
  assign n697 = n673 | n696 ;
  assign n698 = ( n630 & n674 ) | ( n630 & n697 ) | ( n674 & n697 ) ;
  assign n699 = ( ~n113 & n136 ) | ( ~n113 & n510 ) | ( n136 & n510 ) ;
  assign n700 = ( n92 & ~n160 ) | ( n92 & n699 ) | ( ~n160 & n699 ) ;
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n704( .i (n93), .o (n704) );
  assign n705 = ~n701 & n704 ;
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  assign n708 = n703 | n706 ;
  assign n709 = ( ~n555 & n707 ) | ( ~n555 & n708 ) | ( n707 & n708 ) ;
  assign n710 = n51 & ~n709 ;
  assign n711 = n118 & n421 ;
  assign n712 = ~n555 & n711 ;
  buffer buf_n713( .i (n50), .o (n713) );
  assign n714 = n712 | n713 ;
  assign n715 = ~n710 & n714 ;
  buffer buf_n716( .i (n571), .o (n716) );
  assign n717 = n715 | n716 ;
  buffer buf_n718( .i (n549), .o (n718) );
  assign n719 = ( n164 & ~n566 ) | ( n164 & n718 ) | ( ~n566 & n718 ) ;
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n566), .o (n721) );
  assign n722 = ( n119 & n142 ) | ( n119 & ~n721 ) | ( n142 & ~n721 ) ;
  assign n723 = n720 & ~n722 ;
  assign n724 = ~n52 & n723 ;
  assign n725 = n716 & ~n724 ;
  assign n726 = n717 & ~n725 ;
  assign n727 = n31 & ~n726 ;
  assign n728 = ( ~n503 & n570 ) | ( ~n503 & n713 ) | ( n570 & n713 ) ;
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  assign n729 = ( n166 & n305 ) | ( n166 & n570 ) | ( n305 & n570 ) ;
  assign n730 = n728 & ~n729 ;
  assign n731 = n121 | n396 ;
  assign n732 = ( n397 & n730 ) | ( n397 & n731 ) | ( n730 & n731 ) ;
  assign n733 = n146 & n732 ;
  assign n734 = n31 | n733 ;
  assign n735 = ~n727 & n734 ;
  assign n736 = ( ~n113 & n159 ) | ( ~n113 & n510 ) | ( n159 & n510 ) ;
  buffer buf_n737( .i (n736), .o (n737) );
  assign n738 = ( n46 & ~n513 ) | ( n46 & n737 ) | ( ~n513 & n737 ) ;
  buffer buf_n739( .i (n44), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  assign n741 = ( n93 & ~n737 ) | ( n93 & n740 ) | ( ~n737 & n740 ) ;
  assign n742 = n738 & ~n741 ;
  assign n743 = n24 & ~n742 ;
  assign n744 = ~n88 & n156 ;
  buffer buf_n745( .i (n744), .o (n745) );
  assign n748 = n112 & n745 ;
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  assign n752 = n47 & n751 ;
  assign n753 = n24 | n752 ;
  assign n754 = ~n743 & n753 ;
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  assign n757 = ( n189 & n570 ) | ( n189 & n755 ) | ( n570 & n755 ) ;
  assign n758 = n389 & n704 ;
  buffer buf_n759( .i (n758), .o (n759) );
  assign n762 = ( ~n270 & n718 ) | ( ~n270 & n759 ) | ( n718 & n759 ) ;
  assign n763 = n271 & n762 ;
  buffer buf_n764( .i (n188), .o (n764) );
  assign n765 = n763 & ~n764 ;
  assign n766 = ( n756 & ~n757 ) | ( n756 & n765 ) | ( ~n757 & n765 ) ;
  assign n767 = n145 & n766 ;
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  assign n770 = ( n119 & n188 ) | ( n119 & ~n721 ) | ( n188 & ~n721 ) ;
  assign n771 = ~n720 & n770 ;
  assign n772 = ~n144 & n771 ;
  assign n773 = ( n573 & n716 ) | ( n573 & n772 ) | ( n716 & n772 ) ;
  assign n774 = ~n54 & n773 ;
  assign n775 = n768 | n774 ;
  assign n776 = ( n32 & n769 ) | ( n32 & n775 ) | ( n769 & n775 ) ;
  assign n777 = n735 | n776 ;
  assign n778 = ( ~n618 & n698 ) | ( ~n618 & n777 ) | ( n698 & n777 ) ;
  assign n779 = n619 | n778 ;
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  assign n780 = ~n561 & n565 ;
  buffer buf_n781( .i (n780), .o (n781) );
  assign n783 = ~n188 & n781 ;
  assign n784 = n26 & n75 ;
  assign n785 = ( n713 & n783 ) | ( n713 & n784 ) | ( n783 & n784 ) ;
  assign n786 = ~n52 & n785 ;
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  assign n789 = ( n72 & n185 ) | ( n72 & ~n704 ) | ( n185 & ~n704 ) ;
  buffer buf_n790( .i (n789), .o (n790) );
  assign n791 = ( n141 & ~n187 ) | ( n141 & n790 ) | ( ~n187 & n790 ) ;
  buffer buf_n792( .i (n561), .o (n792) );
  assign n793 = ( n74 & ~n790 ) | ( n74 & n792 ) | ( ~n790 & n792 ) ;
  assign n794 = n791 & ~n793 ;
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n26), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n713), .o (n799) );
  assign n800 = ( n795 & n798 ) | ( n795 & ~n799 ) | ( n798 & ~n799 ) ;
  buffer buf_n801( .i (n565), .o (n801) );
  assign n802 = n187 & n801 ;
  assign n803 = n142 & n802 ;
  assign n804 = n594 & n803 ;
  assign n805 = ~n798 & n804 ;
  assign n806 = ( n796 & ~n800 ) | ( n796 & n805 ) | ( ~n800 & n805 ) ;
  assign n807 = n134 & ~n180 ;
  buffer buf_n808( .i (n807), .o (n808) );
  assign n816 = n90 & ~n181 ;
  assign n817 = ~n89 & n134 ;
  buffer buf_n818( .i (n817), .o (n818) );
  assign n821 = ( ~n808 & n816 ) | ( ~n808 & n818 ) | ( n816 & n818 ) ;
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n718), .o (n827) );
  assign n828 = n826 & n827 ;
  buffer buf_n829( .i (n24), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n74), .o (n831) );
  assign n832 = n830 & ~n831 ;
  buffer buf_n833( .i (n49), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  assign n835 = ( n828 & n832 ) | ( n828 & n834 ) | ( n832 & n834 ) ;
  assign n836 = ~n799 & n835 ;
  buffer buf_n837( .i (n836), .o (n837) );
  assign n838 = ( ~n787 & n806 ) | ( ~n787 & n837 ) | ( n806 & n837 ) ;
  assign n839 = n123 & ~n837 ;
  assign n840 = ( n788 & n838 ) | ( n788 & ~n839 ) | ( n838 & ~n839 ) ;
  assign n841 = n171 & n840 ;
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n842( .i (n721), .o (n842) );
  assign n843 = n815 & ~n842 ;
  buffer buf_n844( .i (n484), .o (n844) );
  assign n845 = n843 & ~n844 ;
  assign n846 = n440 & n845 ;
  assign n847 = ~n388 & n846 ;
  assign n848 = ( ~n186 & n382 ) | ( ~n186 & n561 ) | ( n382 & n561 ) ;
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n792), .o (n850) );
  assign n851 = ( n827 & ~n849 ) | ( n827 & n850 ) | ( ~n849 & n850 ) ;
  assign n852 = ( n827 & ~n831 ) | ( n827 & n849 ) | ( ~n831 & n849 ) ;
  assign n853 = n851 & ~n852 ;
  assign n854 = n99 & n853 ;
  assign n855 = ( n440 & n573 ) | ( n440 & n854 ) | ( n573 & n854 ) ;
  assign n856 = ~n30 & n855 ;
  assign n857 = n847 | n856 ;
  assign n858 = ~n171 & n857 ;
  assign n859 = n841 | n858 ;
  buffer buf_n860( .i (n182), .o (n860) );
  assign n861 = ~n646 & n860 ;
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n23), .o (n864) );
  buffer buf_n865( .i (n560), .o (n865) );
  assign n866 = ( n863 & n864 ) | ( n863 & ~n865 ) | ( n864 & ~n865 ) ;
  buffer buf_n867( .i (n646), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  assign n869 = ( n560 & n862 ) | ( n560 & n868 ) | ( n862 & n868 ) ;
  assign n870 = ( n186 & n864 ) | ( n186 & ~n869 ) | ( n864 & ~n869 ) ;
  assign n871 = ~n866 & n870 ;
  assign n872 = n827 | n871 ;
  buffer buf_n873( .i (n868), .o (n873) );
  assign n874 = n864 | n873 ;
  assign n875 = n813 & ~n874 ;
  buffer buf_n876( .i (n718), .o (n876) );
  assign n877 = ~n875 & n876 ;
  assign n878 = n872 & ~n877 ;
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  assign n881 = ( n100 & ~n168 ) | ( n100 & n879 ) | ( ~n168 & n879 ) ;
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  assign n882 = n814 & n876 ;
  assign n883 = ( n227 & n797 ) | ( n227 & n882 ) | ( n797 & n882 ) ;
  assign n884 = ~n798 & n883 ;
  assign n885 = n168 & n884 ;
  assign n886 = ( n880 & ~n881 ) | ( n880 & n885 ) | ( ~n881 & n885 ) ;
  assign n887 = n865 | n873 ;
  buffer buf_n888( .i (n48), .o (n888) );
  buffer buf_n889( .i (n549), .o (n889) );
  assign n890 = ( n887 & ~n888 ) | ( n887 & n889 ) | ( ~n888 & n889 ) ;
  assign n891 = n833 | n890 ;
  buffer buf_n892( .i (n43), .o (n892) );
  buffer buf_n893( .i (n135), .o (n893) );
  assign n894 = ~n892 & n893 ;
  assign n895 = ~n20 & n893 ;
  assign n896 = ( n291 & n894 ) | ( n291 & ~n895 ) | ( n894 & ~n895 ) ;
  buffer buf_n897( .i (n114), .o (n897) );
  assign n898 = ( n867 & ~n896 ) | ( n867 & n897 ) | ( ~n896 & n897 ) ;
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  assign n901 = n873 & ~n899 ;
  assign n902 = ( n889 & ~n900 ) | ( n889 & n901 ) | ( ~n900 & n901 ) ;
  assign n903 = n22 & n740 ;
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  assign n906 = n548 & ~n868 ;
  assign n907 = ( n476 & n904 ) | ( n476 & ~n906 ) | ( n904 & ~n906 ) ;
  assign n908 = ( ~n888 & n905 ) | ( ~n888 & n907 ) | ( n905 & n907 ) ;
  assign n909 = n902 | n908 ;
  assign n910 = n891 & ~n909 ;
  buffer buf_n911( .i (n68), .o (n911) );
  assign n912 = ( n290 & n818 ) | ( n290 & n911 ) | ( n818 & n911 ) ;
  assign n913 = ~n646 & n912 ;
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  assign n916 = n17 & ~n133 ;
  assign n917 = ( n253 & ~n447 ) | ( n253 & n916 ) | ( ~n447 & n916 ) ;
  buffer buf_n918( .i (n89), .o (n918) );
  assign n919 = ( n43 & n917 ) | ( n43 & ~n918 ) | ( n917 & ~n918 ) ;
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  assign n922 = ~n739 & n920 ;
  buffer buf_n923( .i (n918), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  assign n926 = ( n921 & n922 ) | ( n921 & n925 ) | ( n922 & n925 ) ;
  assign n927 = ( n86 & n131 ) | ( n86 & n154 ) | ( n131 & n154 ) ;
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  assign n930 = ~n133 & n928 ;
  assign n931 = ( ~n89 & n929 ) | ( ~n89 & n930 ) | ( n929 & n930 ) ;
  assign n932 = n68 & n931 ;
  assign n933 = ( n20 & n892 ) | ( n20 & n932 ) | ( n892 & n932 ) ;
  assign n934 = ~n21 & n933 ;
  buffer buf_n935( .i (n934), .o (n935) );
  assign n936 = ( ~n914 & n926 ) | ( ~n914 & n935 ) | ( n926 & n935 ) ;
  assign n937 = n389 & ~n935 ;
  assign n938 = ( n915 & n936 ) | ( n915 & ~n937 ) | ( n936 & ~n937 ) ;
  assign n939 = n889 & ~n938 ;
  assign n940 = ( ~n14 & n38 ) | ( ~n14 & n153 ) | ( n38 & n153 ) ;
  buffer buf_n941( .i (n940), .o (n941) );
  assign n946 = ( n16 & ~n87 ) | ( n16 & n941 ) | ( ~n87 & n941 ) ;
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  assign n951 = ( n42 & n157 ) | ( n42 & n947 ) | ( n157 & n947 ) ;
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  assign n954 = ~n945 & n952 ;
  assign n955 = ( ~n950 & n953 ) | ( ~n950 & n954 ) | ( n953 & n954 ) ;
  assign n956 = n867 | n955 ;
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  assign n957 = n459 & n747 ;
  assign n958 = n867 & ~n957 ;
  assign n959 = n956 & ~n958 ;
  assign n960 = n865 & n959 ;
  assign n961 = n889 | n960 ;
  assign n962 = ~n939 & n961 ;
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n842), .o (n964) );
  assign n965 = ( ~n910 & n963 ) | ( ~n910 & n964 ) | ( n963 & n964 ) ;
  buffer buf_n966( .i (n893), .o (n966) );
  assign n967 = ( n291 & ~n739 ) | ( n291 & n966 ) | ( ~n739 & n966 ) ;
  buffer buf_n968( .i (n911), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  assign n970 = ( n292 & n967 ) | ( n292 & n969 ) | ( n967 & n969 ) ;
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  assign n973 = ( n864 & ~n873 ) | ( n864 & n971 ) | ( ~n873 & n971 ) ;
  assign n974 = n972 | n973 ;
  assign n975 = n876 & ~n974 ;
  assign n976 = n892 & ~n911 ;
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n979( .i (n21), .o (n979) );
  assign n980 = ( n635 & n977 ) | ( n635 & n979 ) | ( n977 & n979 ) ;
  buffer buf_n981( .i (n980), .o (n981) );
  assign n982 = n865 | n981 ;
  buffer buf_n983( .i (n635), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  assign n985 = n981 & n984 ;
  assign n986 = n982 & ~n985 ;
  assign n987 = n876 | n986 ;
  buffer buf_n988( .i (n897), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  assign n993 = ( n975 & n987 ) | ( n975 & ~n992 ) | ( n987 & ~n992 ) ;
  assign n994 = ( n963 & ~n964 ) | ( n963 & n993 ) | ( ~n964 & n993 ) ;
  assign n995 = n965 | n994 ;
  buffer buf_n996( .i (n995), .o (n996) );
  assign n997 = ( n55 & n886 ) | ( n55 & n996 ) | ( n886 & n996 ) ;
  assign n998 = ( n135 & n181 ) | ( n135 & n918 ) | ( n181 & n918 ) ;
  assign n999 = ( ~n159 & n182 ) | ( ~n159 & n998 ) | ( n182 & n998 ) ;
  buffer buf_n1000( .i (n999), .o (n1000) );
  assign n1003 = n184 & ~n1000 ;
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  assign n1006 = n1002 | n1004 ;
  buffer buf_n1007( .i (n186), .o (n1007) );
  assign n1008 = ( n1005 & n1006 ) | ( n1005 & ~n1007 ) | ( n1006 & ~n1007 ) ;
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n831), .o (n1011) );
  assign n1012 = ( n992 & n1009 ) | ( n992 & n1011 ) | ( n1009 & n1011 ) ;
  buffer buf_n1013( .i (n180), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  assign n1015 = ~n893 & n1014 ;
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  assign n1019 = n163 & n1018 ;
  assign n1020 = ~n801 & n1019 ;
  assign n1021 = n831 & n1020 ;
  assign n1022 = ~n992 & n1021 ;
  assign n1023 = ( n1010 & ~n1012 ) | ( n1010 & n1022 ) | ( ~n1012 & n1022 ) ;
  buffer buf_n1024( .i (n798), .o (n1024) );
  assign n1025 = n1023 & ~n1024 ;
  assign n1026 = ( n66 & n110 ) | ( n66 & ~n156 ) | ( n110 & ~n156 ) ;
  buffer buf_n1027( .i (n1026), .o (n1027) );
  assign n1032 = ( n158 & n1013 ) | ( n158 & n1027 ) | ( n1013 & n1027 ) ;
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  assign n1037 = ( n114 & n968 ) | ( n114 & n1033 ) | ( n968 & n1033 ) ;
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  assign n1040 = ~n1031 & n1038 ;
  assign n1041 = ( ~n1036 & n1039 ) | ( ~n1036 & n1040 ) | ( n1039 & n1040 ) ;
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  assign n1044 = ( ~n721 & n850 ) | ( ~n721 & n1042 ) | ( n850 & n1042 ) ;
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n1045( .i (n966), .o (n1045) );
  assign n1046 = ~n897 & n1045 ;
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1056( .i (n868), .o (n1056) );
  assign n1057 = ( ~n339 & n1047 ) | ( ~n339 & n1056 ) | ( n1047 & n1056 ) ;
  buffer buf_n1058( .i (n1056), .o (n1058) );
  assign n1059 = n1057 & ~n1058 ;
  buffer buf_n1060( .i (n801), .o (n1060) );
  assign n1061 = n1059 & n1060 ;
  assign n1062 = ( n1043 & ~n1044 ) | ( n1043 & n1061 ) | ( ~n1044 & n1061 ) ;
  assign n1063 = n493 & n984 ;
  assign n1064 = ~n801 & n1063 ;
  buffer buf_n1065( .i (n1058), .o (n1065) );
  assign n1066 = ( ~n991 & n1064 ) | ( ~n991 & n1065 ) | ( n1064 & n1065 ) ;
  assign n1067 = ~n1011 & n1066 ;
  assign n1068 = n1062 | n1067 ;
  assign n1069 = n1024 & n1068 ;
  assign n1070 = n1025 | n1069 ;
  assign n1071 = ( ~n55 & n996 ) | ( ~n55 & n1070 ) | ( n996 & n1070 ) ;
  assign n1072 = n997 | n1071 ;
  buffer buf_n1073( .i (n1072), .o (n1073) );
  assign n1074 = ( n217 & n859 ) | ( n217 & n1073 ) | ( n859 & n1073 ) ;
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  assign n1075 = n268 & ~n338 ;
  assign n1076 = ( n984 & n989 ) | ( n984 & n1075 ) | ( n989 & n1075 ) ;
  assign n1077 = ~n792 & n1076 ;
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  assign n1081 = n739 & n968 ;
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1085( .i (n740), .o (n1085) );
  assign n1086 = ~n1082 & n1085 ;
  buffer buf_n1087( .i (n1086), .o (n1087) );
  assign n1088 = n350 & n1087 ;
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  assign n1089 = ( n341 & n1084 ) | ( n341 & ~n1087 ) | ( n1084 & ~n1087 ) ;
  assign n1090 = ( n1065 & n1088 ) | ( n1065 & ~n1089 ) | ( n1088 & ~n1089 ) ;
  assign n1091 = ( ~n992 & n1078 ) | ( ~n992 & n1090 ) | ( n1078 & n1090 ) ;
  buffer buf_n1092( .i (n797), .o (n1092) );
  assign n1093 = ~n1091 & n1092 ;
  assign n1094 = ( n1024 & n1080 ) | ( n1024 & ~n1093 ) | ( n1080 & ~n1093 ) ;
  assign n1095 = ~n101 & n1094 ;
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  assign n1098 = n696 | n1096 ;
  assign n1099 = ( n502 & n1097 ) | ( n502 & n1098 ) | ( n1097 & n1098 ) ;
  assign n1100 = ( ~n217 & n1073 ) | ( ~n217 & n1099 ) | ( n1073 & n1099 ) ;
  assign n1101 = n1074 | n1100 ;
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  assign n1102 = ~n740 & n925 ;
  assign n1103 = ( n590 & n687 ) | ( n590 & ~n1102 ) | ( n687 & ~n1102 ) ;
  buffer buf_n1104( .i (n979), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  assign n1106 = ~n1103 & n1105 ;
  assign n1107 = ~n205 & n686 ;
  assign n1108 = n1085 & n1107 ;
  assign n1109 = n1105 | n1108 ;
  assign n1110 = ~n1106 & n1109 ;
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  assign n1113 = ( n166 & ~n764 ) | ( n166 & n1111 ) | ( ~n764 & n1111 ) ;
  assign n1114 = ( n163 & ~n207 ) | ( n163 & n1056 ) | ( ~n207 & n1056 ) ;
  assign n1115 = ( ~n207 & n565 ) | ( ~n207 & n1056 ) | ( n565 & n1056 ) ;
  assign n1116 = n1114 & ~n1115 ;
  assign n1117 = n296 & n1116 ;
  assign n1118 = n764 & n1117 ;
  assign n1119 = ( n1112 & ~n1113 ) | ( n1112 & n1118 ) | ( ~n1113 & n1118 ) ;
  assign n1120 = ( ~n208 & n888 ) | ( ~n208 & n1007 ) | ( n888 & n1007 ) ;
  buffer buf_n1121( .i (n704), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  assign n1123 = ( n208 & n1007 ) | ( n208 & ~n1122 ) | ( n1007 & ~n1122 ) ;
  assign n1124 = n1120 | n1123 ;
  assign n1125 = ~n165 & n830 ;
  assign n1126 = ( n1011 & ~n1124 ) | ( n1011 & n1125 ) | ( ~n1124 & n1125 ) ;
  assign n1127 = ~n571 & n1126 ;
  assign n1128 = n1119 | n1127 ;
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n1131 = ( ~n124 & n147 ) | ( ~n124 & n1129 ) | ( n147 & n1129 ) ;
  assign n1132 = ( n1055 & n1130 ) | ( n1055 & ~n1131 ) | ( n1130 & ~n1131 ) ;
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  assign n1135 = n393 & n665 ;
  assign n1136 = ( ~n13 & n175 ) | ( ~n13 & n196 ) | ( n175 & n196 ) ;
  buffer buf_n1137( .i (n1136), .o (n1137) );
  assign n1142 = ( n15 & ~n154 ) | ( n15 & n1137 ) | ( ~n154 & n1137 ) ;
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  assign n1147 = ( n179 & n200 ) | ( n179 & n1143 ) | ( n200 & n1143 ) ;
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  assign n1150 = ~n1141 & n1148 ;
  assign n1151 = ( ~n1146 & n1149 ) | ( ~n1146 & n1150 ) | ( n1149 & n1150 ) ;
  buffer buf_n1152( .i (n892), .o (n1152) );
  assign n1153 = n1151 | n1152 ;
  assign n1154 = ( n155 & n178 ) | ( n155 & n199 ) | ( n178 & n199 ) ;
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n155), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  assign n1159 = ~n1155 & n1158 ;
  assign n1160 = ( n202 & ~n1156 ) | ( n202 & n1159 ) | ( ~n1156 & n1159 ) ;
  buffer buf_n1161( .i (n19), .o (n1161) );
  assign n1162 = n1160 & ~n1161 ;
  assign n1163 = n1152 & ~n1162 ;
  assign n1164 = n1153 & ~n1163 ;
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  assign n1167 = ( n989 & n1121 ) | ( n989 & ~n1165 ) | ( n1121 & ~n1165 ) ;
  assign n1168 = n291 & ~n924 ;
  buffer buf_n1169( .i (n1168), .o (n1169) );
  assign n1174 = ~n513 & n660 ;
  assign n1175 = n1169 & n1174 ;
  assign n1176 = n989 & n1175 ;
  assign n1177 = ( n1166 & n1167 ) | ( n1166 & n1176 ) | ( n1167 & n1176 ) ;
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  assign n1180 = n1173 | n1178 ;
  assign n1181 = ( n1135 & n1179 ) | ( n1135 & n1180 ) | ( n1179 & n1180 ) ;
  assign n1182 = ( ~n145 & n716 ) | ( ~n145 & n1181 ) | ( n716 & n1181 ) ;
  assign n1183 = ( n87 & ~n109 ) | ( n87 & n199 ) | ( ~n109 & n199 ) ;
  assign n1184 = ( n88 & ~n179 ) | ( n88 & n1183 ) | ( ~n179 & n1183 ) ;
  buffer buf_n1185( .i (n1184), .o (n1185) );
  assign n1188 = n918 & ~n1185 ;
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  assign n1191 = n1187 | n1189 ;
  assign n1192 = ( ~n925 & n1190 ) | ( ~n925 & n1191 ) | ( n1190 & n1191 ) ;
  assign n1193 = n1085 & ~n1192 ;
  buffer buf_n1194( .i (n112), .o (n1194) );
  assign n1195 = n203 | n1194 ;
  assign n1196 = n860 | n1195 ;
  assign n1197 = n925 | n1196 ;
  assign n1198 = ~n1085 & n1197 ;
  assign n1199 = n1193 | n1198 ;
  buffer buf_n1200( .i (n163), .o (n1200) );
  assign n1201 = n1199 & ~n1200 ;
  buffer buf_n1202( .i (n88), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  assign n1204 = ( n202 & ~n1013 ) | ( n202 & n1203 ) | ( ~n1013 & n1203 ) ;
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  assign n1207 = ( ~n205 & n897 ) | ( ~n205 & n1206 ) | ( n897 & n1206 ) ;
  buffer buf_n1208( .i (n924), .o (n1208) );
  buffer buf_n1209( .i (n1194), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  assign n1211 = ( ~n1206 & n1208 ) | ( ~n1206 & n1210 ) | ( n1208 & n1210 ) ;
  assign n1212 = n1207 & ~n1211 ;
  buffer buf_n1213( .i (n1152), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  assign n1216 = n1212 & ~n1215 ;
  assign n1217 = n1200 & ~n1216 ;
  assign n1218 = n1201 | n1217 ;
  assign n1219 = n797 & ~n1218 ;
  assign n1220 = n179 | n200 ;
  assign n1221 = ( ~n180 & n656 ) | ( ~n180 & n1220 ) | ( n656 & n1220 ) ;
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1234( .i (n42), .o (n1234) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n158), .o (n1236) );
  assign n1237 = ( n1222 & n1235 ) | ( n1222 & n1236 ) | ( n1235 & n1236 ) ;
  buffer buf_n1238( .i (n1237), .o (n1238) );
  assign n1239 = ( ~n513 & n1208 ) | ( ~n513 & n1238 ) | ( n1208 & n1238 ) ;
  assign n1240 = ( n1208 & n1213 ) | ( n1208 & ~n1238 ) | ( n1213 & ~n1238 ) ;
  assign n1241 = n1239 & ~n1240 ;
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  assign n1244 = ( n87 & n155 ) | ( n87 & ~n178 ) | ( n155 & ~n178 ) ;
  buffer buf_n1245( .i (n86), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  assign n1247 = ( ~n200 & n1244 ) | ( ~n200 & n1246 ) | ( n1244 & n1246 ) ;
  buffer buf_n1248( .i (n1247), .o (n1248) );
  assign n1251 = n1203 & ~n1248 ;
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  assign n1254 = n1250 | n1252 ;
  assign n1255 = ( ~n1208 & n1253 ) | ( ~n1208 & n1254 ) | ( n1253 & n1254 ) ;
  assign n1256 = n1214 & ~n1255 ;
  assign n1257 = n632 | n1014 ;
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n924), .o (n1259) );
  assign n1260 = n1258 | n1259 ;
  assign n1261 = ~n1214 & n1260 ;
  assign n1262 = n1256 | n1261 ;
  buffer buf_n1263( .i (n1236), .o (n1263) );
  assign n1264 = n659 & n1263 ;
  assign n1265 = ( n404 & n1213 ) | ( n404 & n1264 ) | ( n1213 & n1264 ) ;
  assign n1266 = ~n1214 & n1265 ;
  buffer buf_n1267( .i (n1266), .o (n1267) );
  assign n1268 = ( n1242 & n1262 ) | ( n1242 & ~n1267 ) | ( n1262 & ~n1267 ) ;
  assign n1269 = n990 & ~n1267 ;
  assign n1270 = ( ~n1243 & n1268 ) | ( ~n1243 & n1269 ) | ( n1268 & n1269 ) ;
  buffer buf_n1271( .i (n830), .o (n1271) );
  assign n1272 = n1270 & ~n1271 ;
  assign n1273 = ( n1092 & ~n1219 ) | ( n1092 & n1272 ) | ( ~n1219 & n1272 ) ;
  buffer buf_n1274( .i (n571), .o (n1274) );
  buffer buf_n1275( .i (n144), .o (n1275) );
  assign n1276 = ( ~n1273 & n1274 ) | ( ~n1273 & n1275 ) | ( n1274 & n1275 ) ;
  assign n1277 = n1182 & n1276 ;
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  assign n1280 = ( n67 & ~n1158 ) | ( n67 & n1202 ) | ( ~n1158 & n1202 ) ;
  buffer buf_n1281( .i (n1280), .o (n1281) );
  assign n1282 = ( ~n923 & n1194 ) | ( ~n923 & n1281 ) | ( n1194 & n1281 ) ;
  assign n1283 = ( n911 & n1194 ) | ( n911 & ~n1281 ) | ( n1194 & ~n1281 ) ;
  assign n1284 = n1282 & ~n1283 ;
  assign n1285 = n1213 & ~n1284 ;
  assign n1286 = n749 & n968 ;
  buffer buf_n1287( .i (n1152), .o (n1287) );
  assign n1288 = n1286 | n1287 ;
  assign n1289 = ~n1285 & n1288 ;
  assign n1290 = ~n984 & n1289 ;
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  assign n1293 = n112 & n158 ;
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n969), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n983), .o (n1300) );
  assign n1301 = ( n1297 & n1299 ) | ( n1297 & n1300 ) | ( n1299 & n1300 ) ;
  assign n1302 = ~n1058 & n1301 ;
  assign n1303 = n1291 | n1302 ;
  assign n1304 = ( ~n834 & n1292 ) | ( ~n834 & n1303 ) | ( n1292 & n1303 ) ;
  assign n1305 = ( n211 & n1092 ) | ( n211 & n1304 ) | ( n1092 & n1304 ) ;
  buffer buf_n1306( .i (n1305), .o (n1306) );
  assign n1307 = ( n192 & ~n213 ) | ( n192 & n1306 ) | ( ~n213 & n1306 ) ;
  assign n1308 = ( n30 & n192 ) | ( n30 & ~n1306 ) | ( n192 & ~n1306 ) ;
  assign n1309 = n1307 & ~n1308 ;
  buffer buf_n1310( .i (n178), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  assign n1312 = n201 & ~n1311 ;
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1317( .i (n135), .o (n1317) );
  assign n1318 = n1313 & n1317 ;
  buffer buf_n1319( .i (n1318), .o (n1319) );
  assign n1321 = n1210 & n1319 ;
  buffer buf_n1322( .i (n204), .o (n1322) );
  assign n1323 = n1210 & n1322 ;
  assign n1324 = ( n822 & n1210 ) | ( n822 & n1322 ) | ( n1210 & n1322 ) ;
  assign n1325 = ( n1321 & ~n1323 ) | ( n1321 & n1324 ) | ( ~n1323 & n1324 ) ;
  buffer buf_n1326( .i (n389), .o (n1326) );
  assign n1327 = ~n1325 & n1326 ;
  buffer buf_n1328( .i (n923), .o (n1328) );
  assign n1329 = ( n966 & n1205 ) | ( n966 & ~n1328 ) | ( n1205 & ~n1328 ) ;
  assign n1330 = ( n860 & ~n966 ) | ( n860 & n1205 ) | ( ~n966 & n1205 ) ;
  assign n1331 = n1329 & n1330 ;
  assign n1332 = n988 & n1331 ;
  assign n1333 = n1326 | n1332 ;
  assign n1334 = ~n1327 & n1333 ;
  assign n1335 = n830 & ~n1334 ;
  buffer buf_n1336( .i (n199), .o (n1336) );
  assign n1337 = ( n1157 & ~n1310 ) | ( n1157 & n1336 ) | ( ~n1310 & n1336 ) ;
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1158), .o (n1342) );
  assign n1343 = ~n1338 & n1342 ;
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  assign n1346 = ( n204 & n1328 ) | ( n204 & n1344 ) | ( n1328 & n1344 ) ;
  assign n1347 = ( ~n1341 & n1345 ) | ( ~n1341 & n1346 ) | ( n1345 & n1346 ) ;
  assign n1348 = n988 & ~n1347 ;
  assign n1349 = ~n1258 & n1259 ;
  assign n1350 = n988 | n1349 ;
  assign n1351 = ~n1348 & n1350 ;
  assign n1352 = n792 & n1351 ;
  buffer buf_n1353( .i (n829), .o (n1353) );
  assign n1354 = n1352 | n1353 ;
  assign n1355 = ~n1335 & n1354 ;
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  assign n1358 = ( n573 & n1274 ) | ( n573 & n1356 ) | ( n1274 & n1356 ) ;
  assign n1359 = n406 & n1215 ;
  assign n1360 = n829 & n1359 ;
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  assign n1363 = n165 & n623 ;
  assign n1364 = ( n143 & ~n1361 ) | ( n143 & n1363 ) | ( ~n1361 & n1363 ) ;
  assign n1365 = n1362 & n1364 ;
  assign n1366 = ~n1274 & n1365 ;
  assign n1367 = ( n1357 & ~n1358 ) | ( n1357 & n1366 ) | ( ~n1358 & n1366 ) ;
  buffer buf_n1368( .i (n860), .o (n1368) );
  assign n1369 = ( ~n1259 & n1295 ) | ( ~n1259 & n1368 ) | ( n1295 & n1368 ) ;
  assign n1370 = ( ~n1263 & n1294 ) | ( ~n1263 & n1328 ) | ( n1294 & n1328 ) ;
  buffer buf_n1371( .i (n1209), .o (n1371) );
  assign n1372 = ( n1368 & ~n1370 ) | ( n1368 & n1371 ) | ( ~n1370 & n1371 ) ;
  assign n1373 = ~n1369 & n1372 ;
  buffer buf_n1374( .i (n111), .o (n1374) );
  assign n1375 = n415 & ~n1374 ;
  buffer buf_n1376( .i (n1375), .o (n1376) );
  assign n1377 = n1328 & n1376 ;
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  assign n1380 = n983 | n1378 ;
  assign n1381 = ( n1373 & n1379 ) | ( n1373 & n1380 ) | ( n1379 & n1380 ) ;
  assign n1382 = n829 | n1381 ;
  buffer buf_n1383( .i (n1374), .o (n1383) );
  assign n1384 = ( n1236 & n1317 ) | ( n1236 & n1383 ) | ( n1317 & n1383 ) ;
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n1387( .i (n1317), .o (n1387) );
  buffer buf_n1388( .i (n1014), .o (n1388) );
  assign n1389 = ( ~n1209 & n1387 ) | ( ~n1209 & n1388 ) | ( n1387 & n1388 ) ;
  assign n1390 = ~n1385 & n1389 ;
  buffer buf_n1391( .i (n1263), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  assign n1393 = ( ~n1386 & n1390 ) | ( ~n1386 & n1392 ) | ( n1390 & n1392 ) ;
  assign n1394 = ~n1121 & n1393 ;
  buffer buf_n1395( .i (n1105), .o (n1395) );
  assign n1396 = ~n1394 & n1395 ;
  assign n1397 = n1382 & ~n1396 ;
  assign n1398 = n1011 & n1397 ;
  assign n1399 = ( n111 & ~n1158 ) | ( n111 & n1311 ) | ( ~n1158 & n1311 ) ;
  buffer buf_n1400( .i (n1399), .o (n1400) );
  assign n1404 = ( n1161 & n1236 ) | ( n1161 & n1400 ) | ( n1236 & n1400 ) ;
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  assign n1408 = ( n1371 & n1391 ) | ( n1371 & ~n1405 ) | ( n1391 & ~n1405 ) ;
  assign n1409 = n1403 | n1408 ;
  assign n1410 = ( n1105 & ~n1407 ) | ( n1105 & n1409 ) | ( ~n1407 & n1409 ) ;
  buffer buf_n1411( .i (n1300), .o (n1411) );
  assign n1412 = ~n1410 & n1411 ;
  assign n1413 = n1060 & n1412 ;
  buffer buf_n1414( .i (n1065), .o (n1414) );
  assign n1415 = n1413 | n1414 ;
  buffer buf_n1416( .i (n1414), .o (n1416) );
  assign n1417 = ( n1398 & n1415 ) | ( n1398 & ~n1416 ) | ( n1415 & ~n1416 ) ;
  buffer buf_n1418( .i (n1235), .o (n1418) );
  assign n1419 = ( ~n527 & n1376 ) | ( ~n527 & n1418 ) | ( n1376 & n1418 ) ;
  assign n1420 = ~n1287 & n1419 ;
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  assign n1424 = ( n85 & n107 ) | ( n85 & n153 ) | ( n107 & n153 ) ;
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1157), .o (n1428) );
  assign n1429 = ( ~n134 & n1427 ) | ( ~n134 & n1428 ) | ( n1427 & n1428 ) ;
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1433( .i (n1342), .o (n1433) );
  assign n1434 = ~n1430 & n1433 ;
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  assign n1437 = n1432 | n1435 ;
  assign n1438 = ( ~n1392 & n1436 ) | ( ~n1392 & n1437 ) | ( n1436 & n1437 ) ;
  assign n1439 = ( n1215 & n1421 ) | ( n1215 & n1438 ) | ( n1421 & n1438 ) ;
  assign n1440 = n1058 & ~n1439 ;
  assign n1441 = ( n1065 & n1423 ) | ( n1065 & ~n1440 ) | ( n1423 & ~n1440 ) ;
  assign n1442 = ( n109 & ~n132 ) | ( n109 & n1425 ) | ( ~n132 & n1425 ) ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  assign n1446 = n111 & ~n1443 ;
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  assign n1449 = n1445 | n1447 ;
  assign n1450 = ( ~n1209 & n1448 ) | ( ~n1209 & n1449 ) | ( n1448 & n1449 ) ;
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  assign n1453 = ~n1287 & n1368 ;
  assign n1454 = ( n1298 & n1451 ) | ( n1298 & ~n1453 ) | ( n1451 & ~n1453 ) ;
  assign n1455 = n1452 & ~n1454 ;
  buffer buf_n1456( .i (n1455), .o (n1456) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1007), .o (n1458) );
  assign n1459 = ~n1456 & n1458 ;
  assign n1460 = ( n1441 & n1457 ) | ( n1441 & ~n1459 ) | ( n1457 & ~n1459 ) ;
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n799), .o (n1462) );
  assign n1463 = ( n1417 & n1461 ) | ( n1417 & n1462 ) | ( n1461 & n1462 ) ;
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n1464( .i (n923), .o (n1464) );
  assign n1465 = n1388 & ~n1464 ;
  assign n1466 = ( n820 & n1016 ) | ( n820 & ~n1465 ) | ( n1016 & ~n1465 ) ;
  buffer buf_n1467( .i (n67), .o (n1467) );
  assign n1468 = n1374 & n1467 ;
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1472( .i (n1467), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  assign n1474 = ~n1469 & n1473 ;
  buffer buf_n1475( .i (n1474), .o (n1475) );
  assign n1476 = n1466 & n1475 ;
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  assign n1477 = ( n1017 & ~n1471 ) | ( n1017 & n1475 ) | ( ~n1471 & n1475 ) ;
  buffer buf_n1478( .i (n1371), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  assign n1480 = ( n1476 & n1477 ) | ( n1476 & n1479 ) | ( n1477 & n1479 ) ;
  assign n1481 = n1395 & n1480 ;
  assign n1482 = n1298 | n1478 ;
  assign n1483 = n969 & ~n1259 ;
  assign n1484 = n983 & ~n1483 ;
  assign n1485 = ( ~n577 & n1482 ) | ( ~n577 & n1484 ) | ( n1482 & n1484 ) ;
  assign n1486 = ~n1395 & n1485 ;
  assign n1487 = ( n1353 & ~n1481 ) | ( n1353 & n1486 ) | ( ~n1481 & n1486 ) ;
  buffer buf_n1488( .i (n1200), .o (n1488) );
  buffer buf_n1489( .i (n1488), .o (n1489) );
  assign n1490 = n1487 | n1489 ;
  buffer buf_n1491( .i (n110), .o (n1491) );
  buffer buf_n1492( .i (n132), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  assign n1494 = ( n1311 & n1491 ) | ( n1311 & ~n1493 ) | ( n1491 & ~n1493 ) ;
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  assign n1499 = n1383 & ~n1495 ;
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1464), .o (n1502) );
  assign n1503 = ( ~n1045 & n1500 ) | ( ~n1045 & n1502 ) | ( n1500 & n1502 ) ;
  assign n1504 = ( ~n1498 & n1501 ) | ( ~n1498 & n1503 ) | ( n1501 & n1503 ) ;
  buffer buf_n1505( .i (n1104), .o (n1505) );
  assign n1506 = ( ~n1299 & n1504 ) | ( ~n1299 & n1505 ) | ( n1504 & n1505 ) ;
  assign n1507 = ( n512 & n1371 ) | ( n512 & ~n1502 ) | ( n1371 & ~n1502 ) ;
  buffer buf_n1508( .i (n1383), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  assign n1510 = ( n512 & n1045 ) | ( n512 & ~n1509 ) | ( n1045 & ~n1509 ) ;
  assign n1511 = n1507 & n1510 ;
  assign n1512 = ( n1299 & n1505 ) | ( n1299 & ~n1511 ) | ( n1505 & ~n1511 ) ;
  assign n1513 = n1506 & ~n1512 ;
  assign n1514 = n1388 & n1508 ;
  assign n1515 = n1045 & n1514 ;
  assign n1516 = n1104 & n1515 ;
  assign n1517 = ( n1121 & n1299 ) | ( n1121 & n1516 ) | ( n1299 & n1516 ) ;
  assign n1518 = ~n1122 & n1517 ;
  assign n1519 = n1513 | n1518 ;
  assign n1520 = n1489 & n1519 ;
  assign n1521 = n1490 & ~n1520 ;
  assign n1522 = ( ~n1461 & n1462 ) | ( ~n1461 & n1521 ) | ( n1462 & n1521 ) ;
  assign n1523 = ~n1463 & n1522 ;
  assign n1524 = ~n1367 & n1523 ;
  assign n1525 = ( n1278 & ~n1309 ) | ( n1278 & n1524 ) | ( ~n1309 & n1524 ) ;
  assign n1526 = ~n1279 & n1525 ;
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  assign n1527 = ( n1263 & n1418 ) | ( n1263 & n1464 ) | ( n1418 & n1464 ) ;
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1533( .i (n1387), .o (n1533) );
  buffer buf_n1534( .i (n1533), .o (n1534) );
  assign n1535 = ( ~n1392 & n1528 ) | ( ~n1392 & n1534 ) | ( n1528 & n1534 ) ;
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  assign n1540 = ( n888 & n1122 ) | ( n888 & n1536 ) | ( n1122 & n1536 ) ;
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  assign n1543 = ~n1532 & n1541 ;
  assign n1544 = ( ~n1539 & n1542 ) | ( ~n1539 & n1543 ) | ( n1542 & n1543 ) ;
  assign n1545 = n1274 | n1544 ;
  buffer buf_n782( .i (n781), .o (n782) );
  assign n1546 = n1200 | n1411 ;
  assign n1547 = n1060 | n1546 ;
  assign n1548 = ( n782 & ~n842 ) | ( n782 & n1547 ) | ( ~n842 & n1547 ) ;
  assign n1549 = n799 | n1548 ;
  buffer buf_n1550( .i (n1416), .o (n1550) );
  assign n1551 = n1549 & n1550 ;
  assign n1552 = n1545 & ~n1551 ;
  buffer buf_n1553( .i (n1024), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  assign n1555 = ( n1233 & n1552 ) | ( n1233 & n1554 ) | ( n1552 & n1554 ) ;
  buffer buf_n445( .i (n444), .o (n445) );
  assign n1556 = ( n444 & n1060 ) | ( n444 & n1488 ) | ( n1060 & n1488 ) ;
  assign n1557 = n445 | n1556 ;
  assign n1558 = ~n692 & n1557 ;
  assign n1559 = n1462 & ~n1558 ;
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  assign n1560 = n143 & n761 ;
  assign n1561 = n1416 & n1560 ;
  assign n1562 = n1462 | n1561 ;
  assign n1563 = ~n1559 & n1562 ;
  assign n1564 = ( n1233 & ~n1554 ) | ( n1233 & n1563 ) | ( ~n1554 & n1563 ) ;
  assign n1565 = n1555 & n1564 ;
  assign n1566 = ~n1014 & n1235 ;
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  assign n1569 = ( ~n206 & n1104 ) | ( ~n206 & n1568 ) | ( n1104 & n1568 ) ;
  assign n1570 = ( n1322 & n1368 ) | ( n1322 & n1567 ) | ( n1368 & n1567 ) ;
  buffer buf_n1571( .i (n979), .o (n1571) );
  buffer buf_n1572( .i (n1287), .o (n1572) );
  assign n1573 = ( ~n1570 & n1571 ) | ( ~n1570 & n1572 ) | ( n1571 & n1572 ) ;
  assign n1574 = ~n1569 & n1573 ;
  assign n1575 = n1122 & ~n1574 ;
  assign n1576 = n621 & ~n678 ;
  buffer buf_n1577( .i (n1502), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  assign n1580 = n1576 | n1579 ;
  assign n1581 = ~n1575 & n1580 ;
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  assign n1584 = ( n144 & n167 ) | ( n144 & n1582 ) | ( n167 & n1582 ) ;
  assign n1585 = n1322 | n1533 ;
  assign n1586 = ( ~n219 & n661 ) | ( ~n219 & n1585 ) | ( n661 & n1585 ) ;
  assign n1587 = ( n1215 & n1578 ) | ( n1215 & ~n1586 ) | ( n1578 & ~n1586 ) ;
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1579), .o (n1589) );
  assign n1590 = ( n1353 & n1588 ) | ( n1353 & ~n1589 ) | ( n1588 & ~n1589 ) ;
  assign n1591 = ( n833 & n1353 ) | ( n833 & ~n1588 ) | ( n1353 & ~n1588 ) ;
  assign n1592 = n1590 & ~n1591 ;
  assign n1593 = ~n167 & n1592 ;
  assign n1594 = ( n1583 & ~n1584 ) | ( n1583 & n1593 ) | ( ~n1584 & n1593 ) ;
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  assign n1597 = ~n80 & n1595 ;
  buffer buf_n1598( .i (n185), .o (n1598) );
  assign n1599 = ( n1505 & n1578 ) | ( n1505 & ~n1598 ) | ( n1578 & ~n1598 ) ;
  assign n1600 = ( n1300 & ~n1505 ) | ( n1300 & n1598 ) | ( ~n1505 & n1598 ) ;
  assign n1601 = n1599 | n1600 ;
  buffer buf_n1602( .i (n1298), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  assign n1605 = ( n833 & ~n1601 ) | ( n833 & n1604 ) | ( ~n1601 & n1604 ) ;
  buffer buf_n1320( .i (n1319), .o (n1320) );
  assign n1606 = n1320 & n1577 ;
  buffer buf_n1607( .i (n1571), .o (n1607) );
  buffer buf_n1608( .i (n1572), .o (n1608) );
  assign n1609 = ( n1606 & n1607 ) | ( n1606 & n1608 ) | ( n1607 & n1608 ) ;
  assign n1610 = ~n1395 & n1609 ;
  assign n1611 = n1604 & n1610 ;
  assign n1612 = ( ~n834 & n1605 ) | ( ~n834 & n1611 ) | ( n1605 & n1611 ) ;
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n978( .i (n977), .o (n978) );
  assign n1615 = n676 & n1502 ;
  assign n1616 = ( n223 & n978 ) | ( n223 & ~n1615 ) | ( n978 & ~n1615 ) ;
  assign n1617 = ( n207 & n1300 ) | ( n207 & n1616 ) | ( n1300 & n1616 ) ;
  buffer buf_n1618( .i (n1617), .o (n1618) );
  assign n1619 = ( ~n209 & n1458 ) | ( ~n209 & n1618 ) | ( n1458 & n1618 ) ;
  assign n1620 = ( n850 & n1458 ) | ( n850 & ~n1618 ) | ( n1458 & ~n1618 ) ;
  assign n1621 = n1619 & ~n1620 ;
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  assign n1622 = ( n1316 & n1534 ) | ( n1316 & n1577 ) | ( n1534 & n1577 ) ;
  assign n1623 = ~n1578 & n1622 ;
  assign n1624 = ~n1603 & n1623 ;
  buffer buf_n1625( .i (n1607), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1608), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  assign n1629 = ( n1624 & n1626 ) | ( n1624 & n1628 ) | ( n1626 & n1628 ) ;
  assign n1630 = ~n1271 & n1629 ;
  assign n1631 = ( n167 & n1621 ) | ( n167 & n1630 ) | ( n1621 & n1630 ) ;
  assign n1632 = ~n1613 & n1631 ;
  assign n1633 = ( n169 & n1614 ) | ( n169 & n1632 ) | ( n1614 & n1632 ) ;
  assign n1634 = ( n1392 & n1534 ) | ( n1392 & n1572 ) | ( n1534 & n1572 ) ;
  assign n1635 = n1602 & n1634 ;
  assign n1636 = ( n1579 & ~n1625 ) | ( n1579 & n1635 ) | ( ~n1625 & n1635 ) ;
  assign n1637 = ( n42 & n67 ) | ( n42 & n1428 ) | ( n67 & n1428 ) ;
  buffer buf_n1638( .i (n1493), .o (n1638) );
  assign n1639 = ( n1467 & n1637 ) | ( n1467 & ~n1638 ) | ( n1637 & ~n1638 ) ;
  buffer buf_n1640( .i (n1639), .o (n1640) );
  assign n1643 = n1473 & ~n1640 ;
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  assign n1646 = n1642 | n1644 ;
  assign n1647 = ( ~n1602 & n1645 ) | ( ~n1602 & n1646 ) | ( n1645 & n1646 ) ;
  assign n1648 = ( n1579 & n1625 ) | ( n1579 & n1647 ) | ( n1625 & n1647 ) ;
  assign n1649 = n1636 & n1648 ;
  assign n1650 = ( n279 & n303 ) | ( n279 & n1603 ) | ( n303 & n1603 ) ;
  assign n1651 = ~n1604 & n1650 ;
  assign n1652 = n1649 | n1651 ;
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  assign n1655 = ( n191 & n212 ) | ( n191 & n1653 ) | ( n212 & n1653 ) ;
  assign n1656 = ( n627 & n1654 ) | ( n627 & ~n1655 ) | ( n1654 & ~n1655 ) ;
  assign n1657 = n1633 | n1656 ;
  assign n1658 = ( n1596 & ~n1597 ) | ( n1596 & n1657 ) | ( ~n1597 & n1657 ) ;
  assign n1659 = n1565 | n1658 ;
  assign n1660 = ( n1133 & n1526 ) | ( n1133 & ~n1659 ) | ( n1526 & ~n1659 ) ;
  assign n1661 = ~n1134 & n1660 ;
  assign y0 = n238 ;
  assign y1 = n336 ;
  assign y2 = n542 ;
  assign y3 = n779 ;
  assign y4 = n1101 ;
  assign y5 = ~n1661 ;
endmodule
