module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( in_18_ , in_1_ , in_7_ , in_109_ , in_13_ , in_106_ , in_54_ , in_118_ , in_101_ , in_3_ , in_0_ , in_113_ , in_56_ , in_30_ , in_89_ , in_35_ , in_70_ , in_38_ , in_100_ , in_105_ , in_28_ , in_10_ , in_9_ , in_78_ , in_29_ , in_60_ , in_94_ , in_108_ , in_117_ , in_103_ , in_67_ , in_44_ , in_57_ , in_76_ , in_47_ , in_20_ , in_84_ , in_17_ , in_72_ , in_116_ , in_16_ , in_120_ , in_104_ , in_64_ , in_125_ , in_58_ , in_42_ , in_40_ , in_81_ , in_115_ , in_88_ , in_24_ , in_33_ , in_123_ , in_61_ , in_79_ , in_31_ , in_36_ , in_82_ , in_111_ , in_68_ , in_2_ , in_87_ , in_74_ , in_114_ , in_53_ , in_83_ , in_86_ , in_65_ , in_102_ , in_6_ , in_75_ , in_4_ , in_93_ , in_45_ , in_90_ , in_80_ , in_73_ , in_46_ , in_25_ , in_107_ , in_37_ , in_85_ , in_49_ , in_39_ , in_63_ , in_12_ , in_112_ , in_32_ , in_119_ , in_77_ , in_34_ , in_41_ , in_122_ , in_124_ , in_48_ , in_92_ , in_15_ , in_55_ , in_50_ , in_5_ , in_127_ , in_96_ , in_22_ , in_43_ , in_52_ , in_51_ , in_21_ , in_95_ , in_59_ , in_69_ , in_121_ , in_97_ , in_11_ , in_98_ , in_126_ , in_14_ , in_91_ , in_26_ , in_99_ , in_27_ , in_71_ , in_8_ , in_23_ , in_110_ , in_62_ , in_66_ , in_19_ , out_3_ , out_2_ , out_5_ , out_1_ , out_0_ , out_7_ , out_4_ , out_6_ );
  input in_18_ , in_1_ , in_7_ , in_109_ , in_13_ , in_106_ , in_54_ , in_118_ , in_101_ , in_3_ , in_0_ , in_113_ , in_56_ , in_30_ , in_89_ , in_35_ , in_70_ , in_38_ , in_100_ , in_105_ , in_28_ , in_10_ , in_9_ , in_78_ , in_29_ , in_60_ , in_94_ , in_108_ , in_117_ , in_103_ , in_67_ , in_44_ , in_57_ , in_76_ , in_47_ , in_20_ , in_84_ , in_17_ , in_72_ , in_116_ , in_16_ , in_120_ , in_104_ , in_64_ , in_125_ , in_58_ , in_42_ , in_40_ , in_81_ , in_115_ , in_88_ , in_24_ , in_33_ , in_123_ , in_61_ , in_79_ , in_31_ , in_36_ , in_82_ , in_111_ , in_68_ , in_2_ , in_87_ , in_74_ , in_114_ , in_53_ , in_83_ , in_86_ , in_65_ , in_102_ , in_6_ , in_75_ , in_4_ , in_93_ , in_45_ , in_90_ , in_80_ , in_73_ , in_46_ , in_25_ , in_107_ , in_37_ , in_85_ , in_49_ , in_39_ , in_63_ , in_12_ , in_112_ , in_32_ , in_119_ , in_77_ , in_34_ , in_41_ , in_122_ , in_124_ , in_48_ , in_92_ , in_15_ , in_55_ , in_50_ , in_5_ , in_127_ , in_96_ , in_22_ , in_43_ , in_52_ , in_51_ , in_21_ , in_95_ , in_59_ , in_69_ , in_121_ , in_97_ , in_11_ , in_98_ , in_126_ , in_14_ , in_91_ , in_26_ , in_99_ , in_27_ , in_71_ , in_8_ , in_23_ , in_110_ , in_62_ , in_66_ , in_19_ ;
  output out_3_ , out_2_ , out_5_ , out_1_ , out_0_ , out_7_ , out_4_ , out_6_ ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 ;
  assign n129 = in_127_ & in_126_ ;
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  assign n140 = in_125_ | in_124_ ;
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  assign n149 = in_117_ | in_116_ ;
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  assign n153 = in_113_ | in_112_ ;
  buffer buf_n154( .i (n153), .o (n154) );
  assign n155 = in_115_ & in_114_ ;
  buffer buf_n156( .i (n155), .o (n156) );
  assign n157 = ( n150 & n154 ) | ( n150 & n156 ) | ( n154 & n156 ) ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n164 = ( ~n150 & n154 ) | ( ~n150 & n156 ) | ( n154 & n156 ) ;
  buffer buf_n165( .i (n164), .o (n165) );
  assign n166 = ( n152 & ~n158 ) | ( n152 & n165 ) | ( ~n158 & n165 ) ;
  buffer buf_n167( .i (n166), .o (n167) );
  assign n168 = in_123_ & in_122_ ;
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  assign n172 = in_118_ & in_119_ ;
  buffer buf_n173( .i (n172), .o (n173) );
  assign n174 = in_120_ | in_121_ ;
  buffer buf_n175( .i (n174), .o (n175) );
  assign n176 = ( n169 & n173 ) | ( n169 & n175 ) | ( n173 & n175 ) ;
  buffer buf_n177( .i (n176), .o (n177) );
  assign n183 = ( ~n169 & n173 ) | ( ~n169 & n175 ) | ( n173 & n175 ) ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n185 = ( n171 & ~n177 ) | ( n171 & n184 ) | ( ~n177 & n184 ) ;
  buffer buf_n186( .i (n185), .o (n186) );
  assign n187 = ( n145 & n167 ) | ( n145 & n186 ) | ( n167 & n186 ) ;
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  assign n192 = ( ~n145 & n167 ) | ( ~n145 & n186 ) | ( n167 & n186 ) ;
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  assign n195 = ( n148 & ~n189 ) | ( n148 & n194 ) | ( ~n189 & n194 ) ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n197 = n139 & n196 ;
  buffer buf_n198( .i (n197), .o (n198) );
  assign n199 = n139 | n196 ;
  buffer buf_n200( .i (n199), .o (n200) );
  assign n201 = ~n198 & n200 ;
  buffer buf_n202( .i (n201), .o (n202) );
  assign n203 = in_111_ & in_110_ ;
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  assign n214 = in_109_ | in_108_ ;
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  assign n223 = in_101_ | in_100_ ;
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  assign n227 = in_96_ | in_97_ ;
  buffer buf_n228( .i (n227), .o (n228) );
  assign n229 = in_98_ & in_99_ ;
  buffer buf_n230( .i (n229), .o (n230) );
  assign n231 = ( ~n224 & n228 ) | ( ~n224 & n230 ) | ( n228 & n230 ) ;
  buffer buf_n232( .i (n231), .o (n232) );
  assign n233 = ( n224 & n228 ) | ( n224 & n230 ) | ( n228 & n230 ) ;
  buffer buf_n234( .i (n233), .o (n234) );
  assign n240 = ( n226 & n232 ) | ( n226 & ~n234 ) | ( n232 & ~n234 ) ;
  buffer buf_n241( .i (n240), .o (n241) );
  assign n242 = in_106_ & in_107_ ;
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  assign n246 = in_103_ & in_102_ ;
  buffer buf_n247( .i (n246), .o (n247) );
  assign n248 = in_105_ | in_104_ ;
  buffer buf_n249( .i (n248), .o (n249) );
  assign n250 = ( n243 & n247 ) | ( n243 & n249 ) | ( n247 & n249 ) ;
  buffer buf_n251( .i (n250), .o (n251) );
  assign n257 = ( ~n243 & n247 ) | ( ~n243 & n249 ) | ( n247 & n249 ) ;
  buffer buf_n258( .i (n257), .o (n258) );
  assign n259 = ( n245 & ~n251 ) | ( n245 & n258 ) | ( ~n251 & n258 ) ;
  buffer buf_n260( .i (n259), .o (n260) );
  assign n261 = ( n219 & n241 ) | ( n219 & n260 ) | ( n241 & n260 ) ;
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  assign n266 = ( ~n219 & n241 ) | ( ~n219 & n260 ) | ( n241 & n260 ) ;
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  assign n269 = ( n222 & ~n263 ) | ( n222 & n268 ) | ( ~n263 & n268 ) ;
  buffer buf_n270( .i (n269), .o (n270) );
  assign n271 = n213 & n270 ;
  buffer buf_n272( .i (n271), .o (n272) );
  assign n273 = n213 | n270 ;
  buffer buf_n274( .i (n273), .o (n274) );
  assign n275 = ~n272 & n274 ;
  buffer buf_n276( .i (n275), .o (n276) );
  assign n277 = n202 & n276 ;
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  assign n282 = n202 | n276 ;
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  assign n285 = ~n279 & n284 ;
  buffer buf_n286( .i (n285), .o (n286) );
  assign n287 = in_94_ & in_95_ ;
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  assign n298 = in_93_ | in_92_ ;
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  assign n307 = in_84_ | in_85_ ;
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  assign n311 = in_81_ | in_80_ ;
  buffer buf_n312( .i (n311), .o (n312) );
  assign n313 = in_82_ & in_83_ ;
  buffer buf_n314( .i (n313), .o (n314) );
  assign n315 = ( n308 & n312 ) | ( n308 & n314 ) | ( n312 & n314 ) ;
  buffer buf_n316( .i (n315), .o (n316) );
  assign n322 = ( ~n308 & n312 ) | ( ~n308 & n314 ) | ( n312 & n314 ) ;
  buffer buf_n323( .i (n322), .o (n323) );
  assign n324 = ( n310 & ~n316 ) | ( n310 & n323 ) | ( ~n316 & n323 ) ;
  buffer buf_n325( .i (n324), .o (n325) );
  assign n326 = in_90_ & in_91_ ;
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  assign n330 = in_87_ & in_86_ ;
  buffer buf_n331( .i (n330), .o (n331) );
  assign n332 = in_89_ | in_88_ ;
  buffer buf_n333( .i (n332), .o (n333) );
  assign n334 = ( n327 & n331 ) | ( n327 & n333 ) | ( n331 & n333 ) ;
  buffer buf_n335( .i (n334), .o (n335) );
  assign n341 = ( ~n327 & n331 ) | ( ~n327 & n333 ) | ( n331 & n333 ) ;
  buffer buf_n342( .i (n341), .o (n342) );
  assign n343 = ( n329 & ~n335 ) | ( n329 & n342 ) | ( ~n335 & n342 ) ;
  buffer buf_n344( .i (n343), .o (n344) );
  assign n345 = ( n303 & n325 ) | ( n303 & n344 ) | ( n325 & n344 ) ;
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  assign n350 = ( ~n303 & n325 ) | ( ~n303 & n344 ) | ( n325 & n344 ) ;
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  assign n353 = ( n306 & ~n347 ) | ( n306 & n352 ) | ( ~n347 & n352 ) ;
  buffer buf_n354( .i (n353), .o (n354) );
  assign n355 = n297 & n354 ;
  buffer buf_n356( .i (n355), .o (n356) );
  assign n357 = n297 | n354 ;
  buffer buf_n358( .i (n357), .o (n358) );
  assign n359 = ~n356 & n358 ;
  buffer buf_n360( .i (n359), .o (n360) );
  assign n361 = in_78_ & in_79_ ;
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  assign n372 = in_76_ | in_77_ ;
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  assign n381 = in_68_ | in_69_ ;
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  assign n385 = in_64_ | in_65_ ;
  buffer buf_n386( .i (n385), .o (n386) );
  assign n387 = in_67_ & in_66_ ;
  buffer buf_n388( .i (n387), .o (n388) );
  assign n389 = ( n382 & n386 ) | ( n382 & n388 ) | ( n386 & n388 ) ;
  buffer buf_n390( .i (n389), .o (n390) );
  assign n396 = ( ~n382 & n386 ) | ( ~n382 & n388 ) | ( n386 & n388 ) ;
  buffer buf_n397( .i (n396), .o (n397) );
  assign n398 = ( n384 & ~n390 ) | ( n384 & n397 ) | ( ~n390 & n397 ) ;
  buffer buf_n399( .i (n398), .o (n399) );
  assign n400 = in_74_ & in_75_ ;
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  assign n404 = in_70_ & in_71_ ;
  buffer buf_n405( .i (n404), .o (n405) );
  assign n406 = in_72_ | in_73_ ;
  buffer buf_n407( .i (n406), .o (n407) );
  assign n408 = ( n401 & n405 ) | ( n401 & n407 ) | ( n405 & n407 ) ;
  buffer buf_n409( .i (n408), .o (n409) );
  assign n415 = ( ~n401 & n405 ) | ( ~n401 & n407 ) | ( n405 & n407 ) ;
  buffer buf_n416( .i (n415), .o (n416) );
  assign n417 = ( n403 & ~n409 ) | ( n403 & n416 ) | ( ~n409 & n416 ) ;
  buffer buf_n418( .i (n417), .o (n418) );
  assign n419 = ( n377 & n399 ) | ( n377 & n418 ) | ( n399 & n418 ) ;
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  assign n424 = ( ~n377 & n399 ) | ( ~n377 & n418 ) | ( n399 & n418 ) ;
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  assign n427 = ( n380 & ~n421 ) | ( n380 & n426 ) | ( ~n421 & n426 ) ;
  buffer buf_n428( .i (n427), .o (n428) );
  assign n429 = n371 & n428 ;
  buffer buf_n430( .i (n429), .o (n430) );
  assign n431 = n371 | n428 ;
  buffer buf_n432( .i (n431), .o (n432) );
  assign n433 = ~n430 & n432 ;
  buffer buf_n434( .i (n433), .o (n434) );
  assign n435 = n360 & n434 ;
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  assign n440 = n360 | n434 ;
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  assign n443 = ~n437 & n442 ;
  buffer buf_n444( .i (n443), .o (n444) );
  assign n445 = n286 & n444 ;
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  assign n451 = ( n163 & n182 ) | ( n163 & n189 ) | ( n182 & n189 ) ;
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n457( .i (n188), .o (n457) );
  assign n458 = ( n163 & n182 ) | ( n163 & ~n457 ) | ( n182 & ~n457 ) ;
  buffer buf_n459( .i (n458), .o (n459) );
  assign n460 = ( n191 & ~n452 ) | ( n191 & n459 ) | ( ~n452 & n459 ) ;
  buffer buf_n461( .i (n460), .o (n461) );
  assign n462 = n198 & n461 ;
  buffer buf_n463( .i (n462), .o (n463) );
  assign n464 = n198 | n461 ;
  buffer buf_n465( .i (n464), .o (n465) );
  assign n466 = ~n463 & n465 ;
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  assign n469 = ( n239 & n256 ) | ( n239 & n263 ) | ( n256 & n263 ) ;
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n475( .i (n262), .o (n475) );
  assign n476 = ( n239 & n256 ) | ( n239 & ~n475 ) | ( n256 & ~n475 ) ;
  buffer buf_n477( .i (n476), .o (n477) );
  assign n478 = ( n265 & ~n470 ) | ( n265 & n477 ) | ( ~n470 & n477 ) ;
  buffer buf_n479( .i (n478), .o (n479) );
  assign n480 = n272 & n479 ;
  buffer buf_n481( .i (n480), .o (n481) );
  assign n482 = n272 | n479 ;
  buffer buf_n483( .i (n482), .o (n483) );
  assign n484 = ~n481 & n483 ;
  buffer buf_n485( .i (n484), .o (n485) );
  assign n487 = n467 & n485 ;
  assign n488 = n467 | n485 ;
  assign n489 = ~n487 & n488 ;
  buffer buf_n490( .i (n489), .o (n490) );
  assign n491 = n281 & n490 ;
  assign n492 = n281 | n490 ;
  assign n493 = ~n491 & n492 ;
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  assign n495 = ( n321 & n340 ) | ( n321 & n347 ) | ( n340 & n347 ) ;
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n501( .i (n346), .o (n501) );
  assign n502 = ( n321 & n340 ) | ( n321 & ~n501 ) | ( n340 & ~n501 ) ;
  buffer buf_n503( .i (n502), .o (n503) );
  assign n504 = ( n349 & ~n496 ) | ( n349 & n503 ) | ( ~n496 & n503 ) ;
  buffer buf_n505( .i (n504), .o (n505) );
  assign n506 = n356 & n505 ;
  buffer buf_n507( .i (n506), .o (n507) );
  assign n508 = n356 | n505 ;
  buffer buf_n509( .i (n508), .o (n509) );
  assign n510 = ~n507 & n509 ;
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  assign n513 = ( n395 & n414 ) | ( n395 & n421 ) | ( n414 & n421 ) ;
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n519( .i (n420), .o (n519) );
  assign n520 = ( n395 & n414 ) | ( n395 & ~n519 ) | ( n414 & ~n519 ) ;
  buffer buf_n521( .i (n520), .o (n521) );
  assign n522 = ( n423 & ~n514 ) | ( n423 & n521 ) | ( ~n514 & n521 ) ;
  buffer buf_n523( .i (n522), .o (n523) );
  assign n524 = n430 & n523 ;
  buffer buf_n525( .i (n524), .o (n525) );
  assign n526 = n430 | n523 ;
  buffer buf_n527( .i (n526), .o (n527) );
  assign n528 = ~n525 & n527 ;
  buffer buf_n529( .i (n528), .o (n529) );
  assign n531 = n511 & n529 ;
  assign n532 = n511 | n529 ;
  assign n533 = ~n531 & n532 ;
  buffer buf_n534( .i (n533), .o (n534) );
  assign n535 = n439 & n534 ;
  assign n536 = n439 | n534 ;
  assign n537 = ~n535 & n536 ;
  buffer buf_n538( .i (n537), .o (n538) );
  assign n539 = n494 & n538 ;
  assign n540 = n494 | n538 ;
  assign n541 = ~n539 & n540 ;
  buffer buf_n542( .i (n541), .o (n542) );
  assign n543 = n450 & n542 ;
  assign n544 = n450 | n542 ;
  assign n545 = ~n543 & n544 ;
  buffer buf_n546( .i (n545), .o (n546) );
  assign n547 = n286 | n444 ;
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  assign n550 = ~n447 & n549 ;
  buffer buf_n551( .i (n550), .o (n551) );
  assign n552 = in_30_ & in_31_ ;
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  assign n563 = in_28_ | in_29_ ;
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  assign n572 = in_26_ & in_27_ ;
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  assign n576 = in_22_ & in_23_ ;
  buffer buf_n577( .i (n576), .o (n577) );
  assign n578 = in_24_ | in_25_ ;
  buffer buf_n579( .i (n578), .o (n579) );
  assign n580 = ( n573 & n577 ) | ( n573 & n579 ) | ( n577 & n579 ) ;
  buffer buf_n581( .i (n580), .o (n581) );
  assign n587 = ( ~n573 & n577 ) | ( ~n573 & n579 ) | ( n577 & n579 ) ;
  buffer buf_n588( .i (n587), .o (n588) );
  assign n589 = ( n575 & ~n581 ) | ( n575 & n588 ) | ( ~n581 & n588 ) ;
  buffer buf_n590( .i (n589), .o (n590) );
  assign n591 = in_20_ | in_21_ ;
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  assign n595 = in_17_ | in_16_ ;
  buffer buf_n596( .i (n595), .o (n596) );
  assign n597 = in_18_ & in_19_ ;
  buffer buf_n598( .i (n597), .o (n598) );
  assign n599 = ( n592 & n596 ) | ( n592 & n598 ) | ( n596 & n598 ) ;
  buffer buf_n600( .i (n599), .o (n600) );
  assign n606 = ( ~n592 & n596 ) | ( ~n592 & n598 ) | ( n596 & n598 ) ;
  buffer buf_n607( .i (n606), .o (n607) );
  assign n608 = ( n594 & ~n600 ) | ( n594 & n607 ) | ( ~n600 & n607 ) ;
  buffer buf_n609( .i (n608), .o (n609) );
  assign n610 = ( n568 & n590 ) | ( n568 & n609 ) | ( n590 & n609 ) ;
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  assign n615 = ( ~n568 & n590 ) | ( ~n568 & n609 ) | ( n590 & n609 ) ;
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  assign n618 = ( n571 & ~n612 ) | ( n571 & n617 ) | ( ~n612 & n617 ) ;
  buffer buf_n619( .i (n618), .o (n619) );
  assign n620 = n562 & n619 ;
  buffer buf_n621( .i (n620), .o (n621) );
  assign n622 = n562 | n619 ;
  buffer buf_n623( .i (n622), .o (n623) );
  assign n624 = ~n621 & n623 ;
  buffer buf_n625( .i (n624), .o (n625) );
  assign n626 = in_15_ & in_14_ ;
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  assign n637 = in_13_ | in_12_ ;
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  assign n646 = in_4_ | in_5_ ;
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  assign n650 = in_1_ | in_0_ ;
  buffer buf_n651( .i (n650), .o (n651) );
  assign n652 = in_3_ & in_2_ ;
  buffer buf_n653( .i (n652), .o (n653) );
  assign n654 = ( n647 & n651 ) | ( n647 & n653 ) | ( n651 & n653 ) ;
  buffer buf_n655( .i (n654), .o (n655) );
  assign n661 = ( ~n647 & n651 ) | ( ~n647 & n653 ) | ( n651 & n653 ) ;
  buffer buf_n662( .i (n661), .o (n662) );
  assign n663 = ( n649 & ~n655 ) | ( n649 & n662 ) | ( ~n655 & n662 ) ;
  buffer buf_n664( .i (n663), .o (n664) );
  assign n665 = in_10_ & in_11_ ;
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  assign n669 = in_7_ & in_6_ ;
  buffer buf_n670( .i (n669), .o (n670) );
  assign n671 = in_9_ | in_8_ ;
  buffer buf_n672( .i (n671), .o (n672) );
  assign n673 = ( n666 & n670 ) | ( n666 & n672 ) | ( n670 & n672 ) ;
  buffer buf_n674( .i (n673), .o (n674) );
  assign n680 = ( ~n666 & n670 ) | ( ~n666 & n672 ) | ( n670 & n672 ) ;
  buffer buf_n681( .i (n680), .o (n681) );
  assign n682 = ( n668 & ~n674 ) | ( n668 & n681 ) | ( ~n674 & n681 ) ;
  buffer buf_n683( .i (n682), .o (n683) );
  assign n684 = ( n642 & n664 ) | ( n642 & n683 ) | ( n664 & n683 ) ;
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  assign n689 = ( ~n642 & n664 ) | ( ~n642 & n683 ) | ( n664 & n683 ) ;
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  assign n692 = ( n645 & ~n686 ) | ( n645 & n691 ) | ( ~n686 & n691 ) ;
  buffer buf_n693( .i (n692), .o (n693) );
  assign n694 = n636 & n693 ;
  buffer buf_n695( .i (n694), .o (n695) );
  assign n696 = n636 | n693 ;
  buffer buf_n697( .i (n696), .o (n697) );
  assign n698 = ~n695 & n697 ;
  buffer buf_n699( .i (n698), .o (n699) );
  assign n700 = n625 & n699 ;
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  assign n705 = n625 | n699 ;
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  assign n708 = ~n702 & n707 ;
  buffer buf_n709( .i (n708), .o (n709) );
  assign n710 = in_47_ & in_46_ ;
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  assign n721 = in_44_ | in_45_ ;
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  assign n730 = in_36_ | in_37_ ;
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  assign n734 = in_33_ | in_32_ ;
  buffer buf_n735( .i (n734), .o (n735) );
  assign n736 = in_35_ & in_34_ ;
  buffer buf_n737( .i (n736), .o (n737) );
  assign n738 = ( n731 & n735 ) | ( n731 & n737 ) | ( n735 & n737 ) ;
  buffer buf_n739( .i (n738), .o (n739) );
  assign n745 = ( ~n731 & n735 ) | ( ~n731 & n737 ) | ( n735 & n737 ) ;
  buffer buf_n746( .i (n745), .o (n746) );
  assign n747 = ( n733 & ~n739 ) | ( n733 & n746 ) | ( ~n739 & n746 ) ;
  buffer buf_n748( .i (n747), .o (n748) );
  assign n749 = in_42_ & in_43_ ;
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  assign n753 = in_38_ & in_39_ ;
  buffer buf_n754( .i (n753), .o (n754) );
  assign n755 = in_40_ | in_41_ ;
  buffer buf_n756( .i (n755), .o (n756) );
  assign n757 = ( n750 & n754 ) | ( n750 & n756 ) | ( n754 & n756 ) ;
  buffer buf_n758( .i (n757), .o (n758) );
  assign n764 = ( ~n750 & n754 ) | ( ~n750 & n756 ) | ( n754 & n756 ) ;
  buffer buf_n765( .i (n764), .o (n765) );
  assign n766 = ( n752 & ~n758 ) | ( n752 & n765 ) | ( ~n758 & n765 ) ;
  buffer buf_n767( .i (n766), .o (n767) );
  assign n768 = ( n726 & n748 ) | ( n726 & n767 ) | ( n748 & n767 ) ;
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  assign n773 = ( ~n726 & n748 ) | ( ~n726 & n767 ) | ( n748 & n767 ) ;
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  assign n776 = ( n729 & ~n770 ) | ( n729 & n775 ) | ( ~n770 & n775 ) ;
  buffer buf_n777( .i (n776), .o (n777) );
  assign n778 = n720 & n777 ;
  buffer buf_n779( .i (n778), .o (n779) );
  assign n780 = n720 | n777 ;
  buffer buf_n781( .i (n780), .o (n781) );
  assign n782 = ~n779 & n781 ;
  buffer buf_n783( .i (n782), .o (n783) );
  assign n784 = in_63_ & in_62_ ;
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  assign n795 = in_60_ | in_61_ ;
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  assign n804 = in_58_ & in_59_ ;
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  assign n808 = in_54_ & in_55_ ;
  buffer buf_n809( .i (n808), .o (n809) );
  assign n810 = in_56_ | in_57_ ;
  buffer buf_n811( .i (n810), .o (n811) );
  assign n812 = ( n805 & n809 ) | ( n805 & n811 ) | ( n809 & n811 ) ;
  buffer buf_n813( .i (n812), .o (n813) );
  assign n819 = ( ~n805 & n809 ) | ( ~n805 & n811 ) | ( n809 & n811 ) ;
  buffer buf_n820( .i (n819), .o (n820) );
  assign n821 = ( n807 & ~n813 ) | ( n807 & n820 ) | ( ~n813 & n820 ) ;
  buffer buf_n822( .i (n821), .o (n822) );
  assign n823 = in_53_ | in_52_ ;
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  assign n827 = in_49_ | in_48_ ;
  buffer buf_n828( .i (n827), .o (n828) );
  assign n829 = in_50_ & in_51_ ;
  buffer buf_n830( .i (n829), .o (n830) );
  assign n831 = ( n824 & n828 ) | ( n824 & n830 ) | ( n828 & n830 ) ;
  buffer buf_n832( .i (n831), .o (n832) );
  assign n838 = ( ~n824 & n828 ) | ( ~n824 & n830 ) | ( n828 & n830 ) ;
  buffer buf_n839( .i (n838), .o (n839) );
  assign n840 = ( n826 & ~n832 ) | ( n826 & n839 ) | ( ~n832 & n839 ) ;
  buffer buf_n841( .i (n840), .o (n841) );
  assign n842 = ( n800 & n822 ) | ( n800 & n841 ) | ( n822 & n841 ) ;
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  assign n847 = ( ~n800 & n822 ) | ( ~n800 & n841 ) | ( n822 & n841 ) ;
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  assign n850 = ( n803 & ~n844 ) | ( n803 & n849 ) | ( ~n844 & n849 ) ;
  buffer buf_n851( .i (n850), .o (n851) );
  assign n852 = n794 & n851 ;
  buffer buf_n853( .i (n852), .o (n853) );
  assign n854 = n794 | n851 ;
  buffer buf_n855( .i (n854), .o (n855) );
  assign n856 = ~n853 & n855 ;
  buffer buf_n857( .i (n856), .o (n857) );
  assign n858 = n783 | n857 ;
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  assign n861 = n783 & n857 ;
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  assign n866 = n860 & ~n863 ;
  buffer buf_n867( .i (n866), .o (n867) );
  assign n868 = n709 & n867 ;
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  assign n874 = n709 | n867 ;
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  assign n877 = ~n870 & n876 ;
  buffer buf_n878( .i (n877), .o (n878) );
  assign n879 = n551 & n878 ;
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  assign n886 = ( n586 & n605 ) | ( n586 & n612 ) | ( n605 & n612 ) ;
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n892( .i (n611), .o (n892) );
  assign n893 = ( n586 & n605 ) | ( n586 & ~n892 ) | ( n605 & ~n892 ) ;
  buffer buf_n894( .i (n893), .o (n894) );
  assign n895 = ( n614 & ~n887 ) | ( n614 & n894 ) | ( ~n887 & n894 ) ;
  buffer buf_n896( .i (n895), .o (n896) );
  assign n897 = n621 | n896 ;
  buffer buf_n898( .i (n897), .o (n898) );
  assign n899 = n621 & n896 ;
  buffer buf_n900( .i (n899), .o (n900) );
  assign n901 = n898 & ~n900 ;
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  assign n904 = ( n660 & n679 ) | ( n660 & n686 ) | ( n679 & n686 ) ;
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n910( .i (n685), .o (n910) );
  assign n911 = ( n660 & n679 ) | ( n660 & ~n910 ) | ( n679 & ~n910 ) ;
  buffer buf_n912( .i (n911), .o (n912) );
  assign n913 = ( n688 & ~n905 ) | ( n688 & n912 ) | ( ~n905 & n912 ) ;
  buffer buf_n914( .i (n913), .o (n914) );
  assign n915 = n695 & n914 ;
  buffer buf_n916( .i (n915), .o (n916) );
  assign n917 = n695 | n914 ;
  buffer buf_n918( .i (n917), .o (n918) );
  assign n919 = ~n916 & n918 ;
  buffer buf_n920( .i (n919), .o (n920) );
  assign n922 = n902 & n920 ;
  assign n923 = n902 | n920 ;
  assign n924 = ~n922 & n923 ;
  buffer buf_n925( .i (n924), .o (n925) );
  assign n926 = n704 & n925 ;
  assign n927 = n704 | n925 ;
  assign n928 = ~n926 & n927 ;
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  assign n930 = ( n818 & n837 ) | ( n818 & n844 ) | ( n837 & n844 ) ;
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n936( .i (n843), .o (n936) );
  assign n937 = ( n818 & n837 ) | ( n818 & ~n936 ) | ( n837 & ~n936 ) ;
  buffer buf_n938( .i (n937), .o (n938) );
  assign n939 = ( n846 & ~n931 ) | ( n846 & n938 ) | ( ~n931 & n938 ) ;
  buffer buf_n940( .i (n939), .o (n940) );
  assign n941 = n853 & n940 ;
  buffer buf_n942( .i (n941), .o (n942) );
  assign n943 = n853 | n940 ;
  buffer buf_n944( .i (n943), .o (n944) );
  assign n945 = ~n942 & n944 ;
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  assign n948 = ( n744 & n763 ) | ( n744 & n770 ) | ( n763 & n770 ) ;
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n954( .i (n769), .o (n954) );
  assign n955 = ( n744 & n763 ) | ( n744 & ~n954 ) | ( n763 & ~n954 ) ;
  buffer buf_n956( .i (n955), .o (n956) );
  assign n957 = ( n772 & ~n949 ) | ( n772 & n956 ) | ( ~n949 & n956 ) ;
  buffer buf_n958( .i (n957), .o (n958) );
  assign n959 = n779 & n958 ;
  buffer buf_n960( .i (n959), .o (n960) );
  assign n961 = n779 | n958 ;
  buffer buf_n962( .i (n961), .o (n962) );
  assign n963 = ~n960 & n962 ;
  buffer buf_n964( .i (n963), .o (n964) );
  assign n966 = n946 & n964 ;
  assign n967 = n946 | n964 ;
  assign n968 = ~n966 & n967 ;
  buffer buf_n969( .i (n968), .o (n969) );
  assign n970 = n865 & n969 ;
  assign n971 = n865 | n969 ;
  assign n972 = ~n970 & n971 ;
  buffer buf_n973( .i (n972), .o (n973) );
  assign n974 = n929 & n973 ;
  assign n975 = n929 | n973 ;
  assign n976 = ~n974 & n975 ;
  buffer buf_n977( .i (n976), .o (n977) );
  assign n978 = n873 & n977 ;
  assign n979 = n873 | n977 ;
  assign n980 = ~n978 & n979 ;
  buffer buf_n981( .i (n980), .o (n981) );
  assign n982 = ( n546 & n882 ) | ( n546 & n981 ) | ( n882 & n981 ) ;
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  assign n988 = ( n870 & n929 ) | ( n870 & n973 ) | ( n929 & n973 ) ;
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n921( .i (n920), .o (n921) );
  assign n994 = ( n702 & n903 ) | ( n702 & n921 ) | ( n903 & n921 ) ;
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  assign n999 = n891 & n900 ;
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  assign n1006 = n891 | n900 ;
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  assign n1009 = ~n1001 & n1008 ;
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  assign n1011 = n909 & n916 ;
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  assign n1018 = n909 | n916 ;
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  assign n1021 = ~n1013 & n1020 ;
  buffer buf_n1022( .i (n1021), .o (n1022) );
  assign n1023 = n1010 & n1022 ;
  assign n1024 = n1010 | n1022 ;
  assign n1025 = ~n1023 & n1024 ;
  buffer buf_n1026( .i (n1025), .o (n1026) );
  assign n1027 = n998 & n1026 ;
  assign n1028 = n998 | n1026 ;
  assign n1029 = ~n1027 & n1028 ;
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  assign n1031 = n953 & n960 ;
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  assign n1038 = n953 | n960 ;
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  assign n1041 = ~n1033 & n1040 ;
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  assign n1043 = n935 & n942 ;
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  assign n1050 = n935 | n942 ;
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  assign n1053 = ~n1045 & n1052 ;
  buffer buf_n1054( .i (n1053), .o (n1054) );
  assign n1055 = n1042 & n1054 ;
  assign n1056 = n1042 | n1054 ;
  assign n1057 = ~n1055 & n1056 ;
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n965( .i (n964), .o (n965) );
  assign n1059 = ( n863 & n947 ) | ( n863 & n965 ) | ( n947 & n965 ) ;
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  assign n1064 = n1058 & n1063 ;
  assign n1065 = n1058 | n1063 ;
  assign n1066 = ~n1064 & n1065 ;
  buffer buf_n1067( .i (n1066), .o (n1067) );
  assign n1068 = n1030 & n1067 ;
  assign n1069 = n1030 | n1067 ;
  assign n1070 = ~n1068 & n1069 ;
  buffer buf_n1071( .i (n1070), .o (n1071) );
  assign n1072 = n993 & n1071 ;
  assign n1073 = n993 | n1071 ;
  assign n1074 = ~n1072 & n1073 ;
  buffer buf_n1075( .i (n1074), .o (n1075) );
  assign n1076 = ( n447 & n494 ) | ( n447 & n538 ) | ( n494 & n538 ) ;
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n486( .i (n485), .o (n486) );
  assign n1082 = ( n279 & n468 ) | ( n279 & n486 ) | ( n468 & n486 ) ;
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  assign n1087 = n456 & n463 ;
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  assign n1094 = n456 | n463 ;
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  assign n1097 = ~n1089 & n1096 ;
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  assign n1099 = n474 & n481 ;
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  assign n1106 = n474 | n481 ;
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  assign n1109 = ~n1101 & n1108 ;
  buffer buf_n1110( .i (n1109), .o (n1110) );
  assign n1111 = n1098 & n1110 ;
  assign n1112 = n1098 | n1110 ;
  assign n1113 = ~n1111 & n1112 ;
  buffer buf_n1114( .i (n1113), .o (n1114) );
  assign n1115 = n1086 & n1114 ;
  assign n1116 = n1086 | n1114 ;
  assign n1117 = ~n1115 & n1116 ;
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n530( .i (n529), .o (n530) );
  assign n1119 = ( n437 & n512 ) | ( n437 & n530 ) | ( n512 & n530 ) ;
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  assign n1124 = n500 & n507 ;
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  assign n1131 = n500 | n507 ;
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  assign n1134 = ~n1126 & n1133 ;
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  assign n1136 = n518 & n525 ;
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  assign n1143 = n518 | n525 ;
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  assign n1146 = ~n1138 & n1145 ;
  buffer buf_n1147( .i (n1146), .o (n1147) );
  assign n1148 = n1135 & n1147 ;
  assign n1149 = n1135 | n1147 ;
  assign n1150 = ~n1148 & n1149 ;
  buffer buf_n1151( .i (n1150), .o (n1151) );
  assign n1152 = n1123 & n1151 ;
  assign n1153 = n1123 | n1151 ;
  assign n1154 = ~n1152 & n1153 ;
  buffer buf_n1155( .i (n1154), .o (n1155) );
  assign n1156 = n1118 & n1155 ;
  assign n1157 = n1118 | n1155 ;
  assign n1158 = ~n1156 & n1157 ;
  buffer buf_n1159( .i (n1158), .o (n1159) );
  assign n1160 = n1081 & n1159 ;
  assign n1161 = n1081 | n1159 ;
  assign n1162 = ~n1160 & n1161 ;
  buffer buf_n1163( .i (n1162), .o (n1163) );
  assign n1164 = n1075 & n1163 ;
  assign n1165 = n1075 | n1163 ;
  assign n1166 = ~n1164 & n1165 ;
  buffer buf_n1167( .i (n1166), .o (n1167) );
  assign n1168 = n987 & n1167 ;
  assign n1169 = n987 | n1167 ;
  assign n1170 = ~n1168 & n1169 ;
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  assign n1174 = n546 & n981 ;
  assign n1175 = n546 | n981 ;
  assign n1176 = ~n1174 & n1175 ;
  buffer buf_n1177( .i (n1176), .o (n1177) );
  assign n1178 = n885 & n1177 ;
  assign n1179 = n885 | n1177 ;
  assign n1180 = ~n1178 & n1179 ;
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  assign n1187 = ( n990 & n1030 ) | ( n990 & n1067 ) | ( n1030 & n1067 ) ;
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  assign n1189 = n1002 & n1014 ;
  assign n1190 = n1002 | n1014 ;
  assign n1191 = ~n1189 & n1190 ;
  buffer buf_n1192( .i (n1191), .o (n1192) );
  assign n1193 = ( n995 & n1010 ) | ( n995 & n1022 ) | ( n1010 & n1022 ) ;
  buffer buf_n1194( .i (n1193), .o (n1194) );
  assign n1195 = n1192 & n1194 ;
  assign n1196 = n1192 | n1194 ;
  assign n1197 = ~n1195 & n1196 ;
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  assign n1202 = n1034 & n1046 ;
  assign n1203 = n1034 | n1046 ;
  assign n1204 = ~n1202 & n1203 ;
  buffer buf_n1205( .i (n1204), .o (n1205) );
  assign n1206 = ( n1042 & n1054 ) | ( n1042 & n1060 ) | ( n1054 & n1060 ) ;
  buffer buf_n1207( .i (n1206), .o (n1207) );
  assign n1208 = n1205 & n1207 ;
  assign n1209 = n1205 | n1207 ;
  assign n1210 = ~n1208 & n1209 ;
  buffer buf_n1211( .i (n1210), .o (n1211) );
  assign n1215 = n1198 & n1211 ;
  assign n1216 = n1198 | n1211 ;
  assign n1217 = ~n1215 & n1216 ;
  buffer buf_n1218( .i (n1217), .o (n1218) );
  assign n1219 = n1188 & n1218 ;
  assign n1220 = n1188 | n1218 ;
  assign n1221 = ~n1219 & n1220 ;
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  assign n1226 = ( n984 & n1075 ) | ( n984 & n1163 ) | ( n1075 & n1163 ) ;
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  assign n1228 = n1090 & n1102 ;
  assign n1229 = n1090 | n1102 ;
  assign n1230 = ~n1228 & n1229 ;
  buffer buf_n1231( .i (n1230), .o (n1231) );
  assign n1232 = ( n1083 & n1098 ) | ( n1083 & n1110 ) | ( n1098 & n1110 ) ;
  buffer buf_n1233( .i (n1232), .o (n1233) );
  assign n1234 = n1231 & n1233 ;
  assign n1235 = n1231 | n1233 ;
  assign n1236 = ~n1234 & n1235 ;
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  assign n1241 = n1127 & n1139 ;
  assign n1242 = n1127 | n1139 ;
  assign n1243 = ~n1241 & n1242 ;
  buffer buf_n1244( .i (n1243), .o (n1244) );
  assign n1245 = ( n1120 & n1135 ) | ( n1120 & n1147 ) | ( n1135 & n1147 ) ;
  buffer buf_n1246( .i (n1245), .o (n1246) );
  assign n1247 = n1244 & n1246 ;
  assign n1248 = n1244 | n1246 ;
  assign n1249 = ~n1247 & n1248 ;
  buffer buf_n1250( .i (n1249), .o (n1250) );
  assign n1254 = n1237 & n1250 ;
  assign n1255 = n1237 | n1250 ;
  assign n1256 = ~n1254 & n1255 ;
  buffer buf_n1257( .i (n1256), .o (n1257) );
  assign n1258 = ( n1078 & n1118 ) | ( n1078 & n1155 ) | ( n1118 & n1155 ) ;
  buffer buf_n1259( .i (n1258), .o (n1259) );
  assign n1260 = n1257 & n1259 ;
  assign n1261 = n1257 | n1259 ;
  assign n1262 = ~n1260 & n1261 ;
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  assign n1267 = ( n1225 & n1227 ) | ( n1225 & n1266 ) | ( n1227 & n1266 ) ;
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  assign n1269 = ( n1188 & n1201 ) | ( n1188 & n1214 ) | ( n1201 & n1214 ) ;
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  assign n1271 = ( n1005 & n1017 ) | ( n1005 & n1194 ) | ( n1017 & n1194 ) ;
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  assign n1279 = ( n1037 & n1049 ) | ( n1037 & n1207 ) | ( n1049 & n1207 ) ;
  buffer buf_n1280( .i (n1279), .o (n1280) );
  assign n1287 = n1272 & n1280 ;
  assign n1288 = n1272 | n1280 ;
  assign n1289 = ~n1287 & n1288 ;
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  assign n1294 = n1270 & n1293 ;
  assign n1295 = n1270 | n1293 ;
  assign n1296 = ~n1294 & n1295 ;
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  assign n1301 = ( n1093 & n1105 ) | ( n1093 & n1233 ) | ( n1105 & n1233 ) ;
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  assign n1309 = ( n1130 & n1142 ) | ( n1130 & n1246 ) | ( n1142 & n1246 ) ;
  buffer buf_n1310( .i (n1309), .o (n1310) );
  assign n1317 = n1302 & n1310 ;
  assign n1318 = n1302 | n1310 ;
  assign n1319 = ~n1317 & n1318 ;
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  assign n1324 = ( n1240 & n1253 ) | ( n1240 & n1259 ) | ( n1253 & n1259 ) ;
  buffer buf_n1325( .i (n1324), .o (n1325) );
  assign n1326 = n1323 & n1325 ;
  assign n1327 = n1323 | n1325 ;
  assign n1328 = ~n1326 & n1327 ;
  buffer buf_n1329( .i (n1328), .o (n1329) );
  assign n1333 = n1297 & n1329 ;
  assign n1334 = n1297 | n1329 ;
  assign n1335 = ~n1333 & n1334 ;
  buffer buf_n1336( .i (n1335), .o (n1336) );
  assign n1337 = n1268 & n1336 ;
  assign n1338 = n1268 | n1336 ;
  assign n1339 = ~n1337 & n1338 ;
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  assign n1342 = n551 | n878 ;
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  assign n1345 = ~n881 & n1344 ;
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  assign n1357 = ( n1270 & n1278 ) | ( n1270 & n1286 ) | ( n1278 & n1286 ) ;
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  assign n1365 = ( n1268 & n1300 ) | ( n1268 & n1332 ) | ( n1300 & n1332 ) ;
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  assign n1367 = ( n1308 & n1316 ) | ( n1308 & n1325 ) | ( n1316 & n1325 ) ;
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  assign n1375 = ( n1364 & n1366 ) | ( n1364 & n1374 ) | ( n1366 & n1374 ) ;
  buffer buf_n1376( .i (n1375), .o (n1376) );
  assign n1377 = n1222 & n1263 ;
  assign n1378 = n1222 | n1263 ;
  assign n1379 = ~n1377 & n1378 ;
  buffer buf_n1380( .i (n1379), .o (n1380) );
  assign n1381 = n1227 & n1380 ;
  assign n1382 = n1227 | n1380 ;
  assign n1383 = ~n1381 & n1382 ;
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  assign n1388 = n1358 & n1368 ;
  assign n1389 = n1358 | n1368 ;
  assign n1390 = ~n1388 & n1389 ;
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  assign n1395 = n1366 & n1394 ;
  assign n1396 = n1366 | n1394 ;
  assign n1397 = ~n1395 & n1396 ;
  assign out_3_ = n1173 ;
  assign out_2_ = n1186 ;
  assign out_5_ = n1341 ;
  assign out_1_ = n1356 ;
  assign out_0_ = 1'b0 ;
  assign out_7_ = n1376 ;
  assign out_4_ = n1387 ;
  assign out_6_ = n1397 ;
endmodule
