module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 ;
  buffer buf_n347( .i (x10), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n315( .i (x9), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n380( .i (x11), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  assign n482 = ~n322 & n387 ;
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  assign n498 = n362 | n489 ;
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n247( .i (x7), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n413( .i (x12), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n447( .i (x13), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  assign n518 = ~n419 & n453 ;
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n79( .i (x2), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n282( .i (x8), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  assign n538 = n292 & n390 ;
  buffer buf_n539( .i (n538), .o (n539) );
  assign n559 = n327 & n539 ;
  buffer buf_n560( .i (n559), .o (n560) );
  assign n572 = n361 & ~n560 ;
  buffer buf_n328( .i (n327), .o (n328) );
  assign n573 = n328 | n360 ;
  buffer buf_n574( .i (n573), .o (n574) );
  assign n585 = ( ~n362 & n572 ) | ( ~n362 & n574 ) | ( n572 & n574 ) ;
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n112( .i (x3), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n178( .i (x5), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n599 = n120 & n186 ;
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  assign n620 = ( n100 & n590 ) | ( n100 & n611 ) | ( n590 & n611 ) ;
  buffer buf_n145( .i (x4), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  assign n621 = n152 & ~n185 ;
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  assign n642 = ( ~n100 & n590 ) | ( ~n100 & n634 ) | ( n590 & n634 ) ;
  assign n643 = n620 & n642 ;
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n212( .i (x6), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  assign n646 = n98 & ~n197 ;
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  assign n647 = ( n97 & n163 ) | ( n97 & n196 ) | ( n163 & n196 ) ;
  buffer buf_n648( .i (n647), .o (n648) );
  assign n653 = ( n232 & n646 ) | ( n232 & n648 ) | ( n646 & n648 ) ;
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n591( .i (n590), .o (n591) );
  assign n656 = ( n134 & ~n591 ) | ( n134 & n654 ) | ( ~n591 & n654 ) ;
  assign n657 = n129 | n229 ;
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  assign n661 = ~n157 & n190 ;
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  assign n674 = ( n133 & ~n660 ) | ( n133 & n669 ) | ( ~n660 & n669 ) ;
  assign n675 = n591 & n674 ;
  assign n676 = ( n655 & ~n656 ) | ( n655 & n675 ) | ( ~n656 & n675 ) ;
  assign n677 = ~n644 & n676 ;
  assign n678 = ( n536 & n645 ) | ( n536 & n677 ) | ( n645 & n677 ) ;
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n48( .i (x1), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  assign n681 = ( n75 & n274 ) | ( n75 & ~n679 ) | ( n274 & ~n679 ) ;
  assign n682 = ~n290 & n388 ;
  buffer buf_n683( .i (n682), .o (n683) );
  assign n689 = n323 | n388 ;
  buffer buf_n690( .i (n689), .o (n690) );
  assign n705 = ( ~n390 & n683 ) | ( ~n390 & n690 ) | ( n683 & n690 ) ;
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  assign n716 = ( n298 & n363 ) | ( n298 & ~n396 ) | ( n363 & ~n396 ) ;
  assign n717 = n332 & ~n716 ;
  buffer buf_n397( .i (n396), .o (n397) );
  assign n718 = ( ~n286 & n319 ) | ( ~n286 & n384 ) | ( n319 & n384 ) ;
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  assign n727 = n360 & ~n726 ;
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  assign n743 = ( ~n262 & n297 ) | ( ~n262 & n728 ) | ( n297 & n728 ) ;
  assign n744 = n396 & ~n743 ;
  assign n745 = ( n397 & n730 ) | ( n397 & ~n744 ) | ( n730 & ~n744 ) ;
  assign n746 = n717 | n745 ;
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  assign n757 = n267 | n747 ;
  assign n758 = ( n715 & n748 ) | ( n715 & n757 ) | ( n748 & n757 ) ;
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  assign n767 = n266 & ~n399 ;
  assign n768 = n367 & n767 ;
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  assign n771 = n234 | n769 ;
  assign n772 = ( n759 & n770 ) | ( n759 & n771 ) | ( n770 & n771 ) ;
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n15( .i (x0), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  assign n775 = n37 | n167 ;
  assign n776 = n124 | n190 ;
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  assign n786 = ( n37 & ~n167 ) | ( n37 & n785 ) | ( ~n167 & n785 ) ;
  assign n787 = n122 & ~n155 ;
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n198( .i (n197), .o (n198) );
  assign n801 = n99 | n198 ;
  assign n802 = n130 | n163 ;
  buffer buf_n803( .i (n802), .o (n803) );
  assign n806 = ( ~n132 & n796 ) | ( ~n132 & n803 ) | ( n796 & n803 ) ;
  assign n807 = ( n797 & n801 ) | ( n797 & n806 ) | ( n801 & n806 ) ;
  assign n808 = n37 & n807 ;
  assign n809 = ( n775 & ~n786 ) | ( n775 & n808 ) | ( ~n786 & n808 ) ;
  assign n810 = n437 & n809 ;
  assign n811 = ( n472 & n773 ) | ( n472 & ~n810 ) | ( n773 & ~n810 ) ;
  assign n812 = n774 & ~n811 ;
  assign n813 = n75 & n812 ;
  assign n814 = ( n680 & n681 ) | ( n680 & n813 ) | ( n681 & n813 ) ;
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  assign n818 = ( n136 & n202 ) | ( n136 & n800 ) | ( n202 & n800 ) ;
  assign n819 = ( ~n136 & n202 ) | ( ~n136 & n800 ) | ( n202 & n800 ) ;
  assign n820 = ( n137 & ~n818 ) | ( n137 & n819 ) | ( ~n818 & n819 ) ;
  buffer buf_n821( .i (n820), .o (n821) );
  assign n825 = ~n474 & n821 ;
  assign n826 = ( n441 & n597 ) | ( n441 & ~n825 ) | ( n597 & ~n825 ) ;
  assign n827 = n598 & ~n826 ;
  assign n828 = ( n109 & n815 ) | ( n109 & n827 ) | ( n815 & n827 ) ;
  assign n829 = n278 & ~n828 ;
  assign n830 = ( n279 & n817 ) | ( n279 & ~n829 ) | ( n817 & ~n829 ) ;
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  assign n833 = n306 & ~n437 ;
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  assign n838 = ( n476 & n823 ) | ( n476 & ~n837 ) | ( n823 & ~n837 ) ;
  assign n839 = n824 & ~n838 ;
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n76( .i (n75), .o (n76) );
  assign n842 = ( ~n120 & n153 ) | ( ~n120 & n220 ) | ( n153 & n220 ) ;
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  assign n857 = ~n165 & n853 ;
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  assign n860 = ( ~n201 & n856 ) | ( ~n201 & n859 ) | ( n856 & n859 ) ;
  assign n861 = n129 & ~n793 ;
  assign n862 = n97 & n861 ;
  assign n863 = ( n164 & n795 ) | ( n164 & ~n862 ) | ( n795 & ~n862 ) ;
  assign n864 = ( n232 & n796 ) | ( n232 & n863 ) | ( n796 & n863 ) ;
  assign n865 = n199 & n864 ;
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  assign n868 = n102 | n866 ;
  assign n869 = ( n860 & n867 ) | ( n860 & n868 ) | ( n867 & n868 ) ;
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n537( .i (n536), .o (n537) );
  assign n872 = ( n308 & n537 ) | ( n308 & ~n870 ) | ( n537 & ~n870 ) ;
  assign n873 = n871 & n872 ;
  assign n874 = ( n76 & n275 ) | ( n76 & n873 ) | ( n275 & n873 ) ;
  assign n875 = n32 & n129 ;
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  assign n882 = n258 & ~n458 ;
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  assign n890 = ( n432 & n876 ) | ( n432 & n889 ) | ( n876 & n889 ) ;
  assign n891 = ~n877 & n890 ;
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  assign n895 = n299 & n528 ;
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  assign n900 = n185 | n254 ;
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  assign n920 = ( n892 & n899 ) | ( n892 & ~n914 ) | ( n899 & ~n914 ) ;
  assign n921 = n102 & ~n920 ;
  assign n922 = ( n103 & n894 ) | ( n103 & ~n921 ) | ( n894 & ~n921 ) ;
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  assign n925 = ( ~n171 & n238 ) | ( ~n171 & n923 ) | ( n238 & n923 ) ;
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  assign n926 = n426 & n883 ;
  assign n927 = ~n159 & n926 ;
  buffer buf_n928( .i (n927), .o (n928) );
  assign n936 = n31 & n928 ;
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  assign n940 = ( n196 & ~n265 ) | ( n196 & n937 ) | ( ~n265 & n937 ) ;
  assign n941 = n896 & ~n940 ;
  assign n942 = ( n897 & n939 ) | ( n897 & ~n941 ) | ( n939 & ~n941 ) ;
  assign n943 = ~n100 & n942 ;
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  assign n946 = n935 | n944 ;
  assign n947 = ( n39 & n945 ) | ( n39 & n946 ) | ( n945 & n946 ) ;
  assign n948 = ~n267 & n897 ;
  assign n949 = ( n166 & n199 ) | ( n166 & n948 ) | ( n199 & n948 ) ;
  assign n950 = ~n167 & n949 ;
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  assign n953 = n136 | n951 ;
  assign n954 = ( n947 & n952 ) | ( n947 & n953 ) | ( n952 & n953 ) ;
  assign n955 = ~n238 & n954 ;
  assign n956 = ( n924 & ~n925 ) | ( n924 & n955 ) | ( ~n925 & n955 ) ;
  assign n957 = n76 & n956 ;
  assign n958 = ( ~n276 & n874 ) | ( ~n276 & n957 ) | ( n874 & n957 ) ;
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n110( .i (n109), .o (n110) );
  assign n962 = ( n110 & ~n278 ) | ( n110 & n959 ) | ( ~n278 & n959 ) ;
  assign n963 = n840 & ~n962 ;
  assign n964 = ( n841 & n961 ) | ( n841 & ~n963 ) | ( n961 & ~n963 ) ;
  assign n965 = n831 | n964 ;
  assign n966 = ( n517 & n832 ) | ( n517 & n965 ) | ( n832 & n965 ) ;
  assign n967 = n127 & n160 ;
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  assign n979 = n673 & ~n976 ;
  assign n980 = n438 & ~n472 ;
  assign n981 = ( n977 & n979 ) | ( n977 & n980 ) | ( n979 & n980 ) ;
  assign n982 = ~n238 & n273 ;
  assign n983 = ( n75 & n981 ) | ( n75 & n982 ) | ( n981 & n982 ) ;
  assign n984 = ~n76 & n983 ;
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  assign n987 = ( n45 & n109 ) | ( n45 & ~n985 ) | ( n109 & ~n985 ) ;
  assign n988 = n58 | n188 ;
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  assign n999 = n163 | n230 ;
  buffer buf_n1000( .i (n999), .o (n1000) );
  assign n1005 = ( n68 & ~n198 ) | ( n68 & n1000 ) | ( ~n198 & n1000 ) ;
  assign n1006 = n156 | n189 ;
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  assign n1019 = ( ~n162 & n630 ) | ( ~n162 & n1011 ) | ( n630 & n1011 ) ;
  buffer buf_n1020( .i (n1019), .o (n1020) );
  assign n1026 = ( n632 & n658 ) | ( n632 & n1020 ) | ( n658 & n1020 ) ;
  assign n1027 = n68 & n1026 ;
  assign n1028 = ( n998 & ~n1005 ) | ( n998 & n1027 ) | ( ~n1005 & n1027 ) ;
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  assign n1032 = n472 & ~n1031 ;
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1033( .i (n135), .o (n1033) );
  assign n1034 = n1025 & n1033 ;
  buffer buf_n1035( .i (n471), .o (n1035) );
  assign n1036 = n1034 | n1035 ;
  assign n1037 = ~n1032 & n1036 ;
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  assign n1040 = ~n261 & n296 ;
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  assign n1055 = ( n441 & n1038 ) | ( n441 & ~n1053 ) | ( n1038 & ~n1053 ) ;
  assign n1056 = n1039 & ~n1055 ;
  assign n1057 = n109 & n1056 ;
  assign n1058 = ( n986 & n987 ) | ( n986 & n1057 ) | ( n987 & n1057 ) ;
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1061 = ~n91 & n190 ;
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  assign n1079 = ~n60 & n91 ;
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  assign n1091 = ( n169 & ~n1072 ) | ( n169 & n1090 ) | ( ~n1072 & n1090 ) ;
  assign n1092 = n40 & ~n1091 ;
  assign n1093 = n60 & n157 ;
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  assign n1109 = n40 | n1105 ;
  assign n1110 = ( ~n41 & n1092 ) | ( ~n41 & n1109 ) | ( n1092 & n1109 ) ;
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  assign n1113 = ~n232 & n433 ;
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  assign n1121 = ( n275 & ~n1111 ) | ( n275 & n1120 ) | ( ~n1111 & n1120 ) ;
  assign n1122 = n1112 & n1121 ;
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  assign n1125 = ~n435 & n1047 ;
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  assign n1133 = n1078 & n1132 ;
  assign n1134 = ~n1123 & n1133 ;
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  assign n1135 = n143 & ~n478 ;
  assign n1136 = ( n1124 & n1134 ) | ( n1124 & n1135 ) | ( n1134 & n1135 ) ;
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  assign n1137 = ( ~n63 & n94 ) | ( ~n63 & n160 ) | ( n94 & n160 ) ;
  assign n1138 = n159 & n192 ;
  assign n1139 = ( n94 & n160 ) | ( n94 & n1138 ) | ( n160 & n1138 ) ;
  assign n1140 = ( n1096 & n1137 ) | ( n1096 & ~n1139 ) | ( n1137 & ~n1139 ) ;
  assign n1141 = n662 & n1080 ;
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  assign n1144 = n128 | n1142 ;
  assign n1145 = ( ~n1140 & n1143 ) | ( ~n1140 & n1144 ) | ( n1143 & n1144 ) ;
  assign n1146 = n33 & ~n1145 ;
  assign n1147 = n65 & n968 ;
  assign n1148 = n33 | n1147 ;
  assign n1149 = ~n1146 & n1148 ;
  buffer buf_n1150( .i (n1149), .o (n1150) );
  assign n1159 = n224 & n706 ;
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  assign n1162 = n361 | n1160 ;
  assign n1163 = ( ~n395 & n1161 ) | ( ~n395 & n1162 ) | ( n1161 & n1162 ) ;
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  assign n1170 = n1150 & n1168 ;
  assign n1171 = n435 & ~n1170 ;
  assign n1172 = ( n96 & n162 ) | ( n96 & ~n586 ) | ( n162 & ~n586 ) ;
  buffer buf_n1173( .i (n1172), .o (n1173) );
  assign n1174 = ~n197 & n1173 ;
  assign n1175 = ( ~n197 & n588 ) | ( ~n197 & n1173 ) | ( n588 & n1173 ) ;
  assign n1176 = ( n589 & n1174 ) | ( n589 & ~n1175 ) | ( n1174 & ~n1175 ) ;
  assign n1177 = n133 & n1176 ;
  assign n1178 = n435 | n1177 ;
  assign n1179 = ~n1171 & n1178 ;
  assign n1180 = ~n471 & n1179 ;
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  assign n1183 = n470 & n1029 ;
  assign n1184 = ( n437 & n593 ) | ( n437 & ~n1183 ) | ( n593 & ~n1183 ) ;
  assign n1185 = n594 & ~n1184 ;
  assign n1186 = n1181 | n1185 ;
  assign n1187 = ( n106 & n1182 ) | ( n106 & n1186 ) | ( n1182 & n1186 ) ;
  assign n1188 = n275 & n1187 ;
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  assign n1191 = n440 & n754 ;
  assign n1192 = ( n475 & n1157 ) | ( n475 & ~n1191 ) | ( n1157 & ~n1191 ) ;
  assign n1193 = n1158 & ~n1192 ;
  assign n1194 = n1189 | n1193 ;
  assign n1195 = ( n243 & n1190 ) | ( n243 & n1194 ) | ( n1190 & n1194 ) ;
  buffer buf_n1196( .i (n1195), .o (n1196) );
  assign n1197 = ( ~n1059 & n1136 ) | ( ~n1059 & n1196 ) | ( n1136 & n1196 ) ;
  assign n1198 = n515 | n1196 ;
  assign n1199 = ( n1060 & n1197 ) | ( n1060 & n1198 ) | ( n1197 & n1198 ) ;
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  assign n1201 = n132 & ~n1100 ;
  assign n1202 = n36 & n1201 ;
  assign n1203 = n28 & ~n92 ;
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  assign n1210 = n67 & ~n131 ;
  assign n1211 = ( ~n35 & n1209 ) | ( ~n35 & n1210 ) | ( n1209 & n1210 ) ;
  assign n1212 = n1168 & n1211 ;
  assign n1213 = ( n1169 & n1202 ) | ( n1169 & n1212 ) | ( n1202 & n1212 ) ;
  assign n1214 = n92 | n125 ;
  buffer buf_n1215( .i (n1214), .o (n1215) );
  assign n1231 = n92 & ~n125 ;
  buffer buf_n1232( .i (n1231), .o (n1232) );
  assign n1233 = ( ~n94 & n1215 ) | ( ~n94 & n1232 ) | ( n1215 & n1232 ) ;
  buffer buf_n1234( .i (n1233), .o (n1234) );
  assign n1240 = n586 & n1234 ;
  assign n1241 = n431 | n1240 ;
  assign n1242 = n30 | n63 ;
  assign n1243 = n30 & ~n1232 ;
  assign n1244 = n1242 & ~n1243 ;
  assign n1245 = n1164 & n1244 ;
  assign n1246 = n431 & ~n1245 ;
  assign n1247 = n1241 & ~n1246 ;
  assign n1248 = n165 & n1247 ;
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n434), .o (n1251) );
  assign n1252 = n1249 | n1251 ;
  assign n1253 = ( n1213 & n1250 ) | ( n1213 & n1252 ) | ( n1250 & n1252 ) ;
  assign n1254 = ~n471 & n1253 ;
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  assign n1257 = n68 | n99 ;
  assign n1258 = ~n85 & n118 ;
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1278( .i (n67), .o (n1278) );
  assign n1279 = n1271 & n1278 ;
  assign n1280 = ( ~n69 & n1257 ) | ( ~n69 & n1279 ) | ( n1257 & n1279 ) ;
  buffer buf_n1281( .i (n1280), .o (n1281) );
  assign n1285 = n470 & n1281 ;
  buffer buf_n1286( .i (n436), .o (n1286) );
  assign n1287 = ( n593 & ~n1285 ) | ( n593 & n1286 ) | ( ~n1285 & n1286 ) ;
  assign n1288 = n594 & ~n1287 ;
  assign n1289 = n1255 | n1288 ;
  assign n1290 = ( n172 & n1256 ) | ( n172 & n1289 ) | ( n1256 & n1289 ) ;
  buffer buf_n1291( .i (n274), .o (n1291) );
  assign n1292 = n1290 & n1291 ;
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n1295( .i (n159), .o (n1295) );
  assign n1296 = ( n63 & ~n127 ) | ( n63 & n1295 ) | ( ~n127 & n1295 ) ;
  assign n1297 = n128 & ~n1296 ;
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n128), .o (n1300) );
  assign n1301 = n162 & ~n1300 ;
  assign n1302 = ( n97 & n1298 ) | ( n97 & n1301 ) | ( n1298 & n1301 ) ;
  assign n1303 = n1299 | n1302 ;
  assign n1304 = n30 & ~n1215 ;
  buffer buf_n1305( .i (n29), .o (n1305) );
  assign n1306 = n791 & ~n1305 ;
  assign n1307 = ( n31 & ~n1304 ) | ( n31 & n1306 ) | ( ~n1304 & n1306 ) ;
  assign n1308 = n65 & ~n1307 ;
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  assign n1311 = n34 | n1309 ;
  assign n1312 = ( n1303 & n1310 ) | ( n1303 & n1311 ) | ( n1310 & n1311 ) ;
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  assign n1319 = n440 & n1318 ;
  assign n1320 = ( n475 & n755 ) | ( n475 & ~n1319 ) | ( n755 & ~n1319 ) ;
  assign n1321 = n756 & ~n1320 ;
  assign n1322 = n1293 | n1321 ;
  assign n1323 = ( n243 & n1294 ) | ( n243 & n1322 ) | ( n1294 & n1322 ) ;
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  assign n1326 = ~n211 & n1324 ;
  buffer buf_n1327( .i (n158), .o (n1327) );
  assign n1328 = ~n461 & n1327 ;
  buffer buf_n1329( .i (n93), .o (n1329) );
  assign n1330 = ( n193 & n1328 ) | ( n193 & n1329 ) | ( n1328 & n1329 ) ;
  assign n1331 = ~n194 & n1330 ;
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  assign n1342 = ~n134 & n234 ;
  assign n1343 = ( n201 & n1274 ) | ( n201 & ~n1342 ) | ( n1274 & ~n1342 ) ;
  assign n1344 = ~n185 & n219 ;
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  assign n1362 = n1272 & n1357 ;
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  assign n1365 = n168 | n1363 ;
  assign n1366 = ( ~n1343 & n1364 ) | ( ~n1343 & n1365 ) | ( n1364 & n1365 ) ;
  assign n1367 = ( n73 & n1339 ) | ( n73 & n1366 ) | ( n1339 & n1366 ) ;
  assign n1368 = n473 & ~n1367 ;
  assign n1369 = ( n474 & n1341 ) | ( n474 & ~n1368 ) | ( n1341 & ~n1368 ) ;
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  assign n1374 = n272 & n594 ;
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n1378( .i (n1377), .o (n1378) );
  buffer buf_n1379( .i (n1378), .o (n1379) );
  assign n1380 = ( n444 & n1372 ) | ( n444 & ~n1379 ) | ( n1372 & ~n1379 ) ;
  assign n1381 = n1373 & ~n1380 ;
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  assign n1382 = ( n307 & n536 ) | ( n307 & ~n1283 ) | ( n536 & ~n1283 ) ;
  assign n1383 = n1284 & n1382 ;
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  assign n1386 = ( n434 & ~n1046 ) | ( n434 & n1238 ) | ( ~n1046 & n1238 ) ;
  assign n1387 = n1239 & ~n1386 ;
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n470), .o (n1390) );
  assign n1391 = ( ~n169 & n1388 ) | ( ~n169 & n1390 ) | ( n1388 & n1390 ) ;
  assign n1392 = ( n269 & n1114 ) | ( n269 & ~n1313 ) | ( n1114 & ~n1313 ) ;
  assign n1393 = n1314 & n1392 ;
  assign n1394 = ~n1390 & n1393 ;
  assign n1395 = ( n1389 & ~n1391 ) | ( n1389 & n1394 ) | ( ~n1391 & n1394 ) ;
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  assign n1399 = ( n172 & ~n274 ) | ( n172 & n1396 ) | ( ~n274 & n1396 ) ;
  assign n1400 = n1384 & ~n1399 ;
  assign n1401 = ( n1385 & n1398 ) | ( n1385 & ~n1400 ) | ( n1398 & ~n1400 ) ;
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  assign n1404 = ( n209 & n513 ) | ( n209 & ~n1402 ) | ( n513 & ~n1402 ) ;
  buffer buf_n1054( .i (n1053), .o (n1054) );
  assign n1405 = ( n442 & ~n1054 ) | ( n442 & n1370 ) | ( ~n1054 & n1370 ) ;
  assign n1406 = n1371 & ~n1405 ;
  assign n1407 = n513 & n1406 ;
  assign n1408 = ( n1403 & n1404 ) | ( n1403 & n1407 ) | ( n1404 & n1407 ) ;
  assign n1409 = n1381 | n1408 ;
  assign n1410 = ( n1325 & ~n1326 ) | ( n1325 & n1409 ) | ( ~n1326 & n1409 ) ;
  buffer buf_n1411( .i (n1410), .o (n1411) );
  assign n1412 = ( n166 & n199 ) | ( n166 & ~n468 ) | ( n199 & ~n468 ) ;
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1415( .i (n166), .o (n1415) );
  assign n1416 = ( n134 & n469 ) | ( n134 & n1415 ) | ( n469 & n1415 ) ;
  assign n1417 = n1413 & ~n1416 ;
  assign n1418 = ( ~n202 & n1414 ) | ( ~n202 & n1417 ) | ( n1414 & n1417 ) ;
  assign n1419 = n89 & ~n155 ;
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n96), .o (n1428) );
  assign n1429 = ( n196 & n1426 ) | ( n196 & n1428 ) | ( n1426 & n1428 ) ;
  buffer buf_n1430( .i (n161), .o (n1430) );
  assign n1431 = ( n195 & n1300 ) | ( n195 & n1430 ) | ( n1300 & n1430 ) ;
  assign n1432 = ( ~n1300 & n1425 ) | ( ~n1300 & n1430 ) | ( n1425 & n1430 ) ;
  assign n1433 = n1431 | n1432 ;
  assign n1434 = ( n1427 & ~n1429 ) | ( n1427 & n1433 ) | ( ~n1429 & n1433 ) ;
  assign n1435 = n467 & n1434 ;
  buffer buf_n1436( .i (n1435), .o (n1436) );
  assign n1438 = n70 & n1436 ;
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  assign n1441 = n103 | n1439 ;
  assign n1442 = ( n1418 & n1440 ) | ( n1418 & n1441 ) | ( n1440 & n1441 ) ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  assign n1445 = ( n440 & ~n1375 ) | ( n440 & n1443 ) | ( ~n1375 & n1443 ) ;
  assign n1446 = n1444 & ~n1445 ;
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  assign n1449 = ~n242 & n1447 ;
  assign n1450 = ( n64 & n95 ) | ( n64 & n194 ) | ( n95 & n194 ) ;
  assign n1451 = n194 & n792 ;
  assign n1452 = ( ~n65 & n1450 ) | ( ~n65 & n1451 ) | ( n1450 & n1451 ) ;
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  assign n1455 = ( ~n85 & n118 ) | ( ~n85 & n184 ) | ( n118 & n184 ) ;
  buffer buf_n1456( .i (n1455), .o (n1456) );
  assign n1477 = n153 & ~n1456 ;
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  assign n1488 = ( ~n21 & n85 ) | ( ~n21 & n184 ) | ( n85 & n184 ) ;
  assign n1489 = ( n21 & n118 ) | ( n21 & n184 ) | ( n118 & n184 ) ;
  assign n1490 = ~n1488 & n1489 ;
  assign n1491 = ( ~n20 & n117 ) | ( ~n20 & n183 ) | ( n117 & n183 ) ;
  assign n1492 = ~n19 & n149 ;
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1504( .i (n117), .o (n1504) );
  assign n1505 = ( n1491 & n1493 ) | ( n1491 & ~n1504 ) | ( n1493 & ~n1504 ) ;
  buffer buf_n1506( .i (n1505), .o (n1506) );
  assign n1517 = ( n56 & n1490 ) | ( n56 & n1506 ) | ( n1490 & n1506 ) ;
  assign n1518 = ~n622 & n1517 ;
  assign n1519 = ( n58 & n623 ) | ( n58 & n1518 ) | ( n623 & n1518 ) ;
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n1522( .i (n1521), .o (n1522) );
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  assign n1528 = ( ~n1453 & n1487 ) | ( ~n1453 & n1527 ) | ( n1487 & n1527 ) ;
  assign n1529 = n27 | n1520 ;
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  buffer buf_n1534( .i (n1533), .o (n1534) );
  buffer buf_n1535( .i (n1534), .o (n1535) );
  buffer buf_n1536( .i (n1535), .o (n1536) );
  assign n1537 = ( n1454 & n1528 ) | ( n1454 & n1536 ) | ( n1528 & n1536 ) ;
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  assign n1543 = ( ~n259 & n359 ) | ( ~n259 & n392 ) | ( n359 & n392 ) ;
  buffer buf_n1544( .i (n1543), .o (n1544) );
  assign n1548 = ( n261 & ~n329 ) | ( n261 & n1544 ) | ( ~n329 & n1544 ) ;
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  assign n1554 = ( n263 & n363 ) | ( n263 & ~n1549 ) | ( n363 & ~n1549 ) ;
  assign n1555 = n1547 | n1554 ;
  buffer buf_n1556( .i (n1555), .o (n1556) );
  buffer buf_n1557( .i (n1556), .o (n1557) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  assign n1558 = ~n334 & n1556 ;
  assign n1559 = ( ~n1553 & n1557 ) | ( ~n1553 & n1558 ) | ( n1557 & n1558 ) ;
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  assign n1563 = n1286 & n1562 ;
  assign n1564 = ( n1035 & n1541 ) | ( n1035 & ~n1563 ) | ( n1541 & ~n1563 ) ;
  assign n1565 = n1542 & ~n1564 ;
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  assign n1568 = ( n240 & n310 ) | ( n240 & ~n1566 ) | ( n310 & ~n1566 ) ;
  buffer buf_n1437( .i (n1436), .o (n1437) );
  assign n1569 = n231 & ~n432 ;
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  assign n1573 = ( n270 & n1437 ) | ( n270 & n1572 ) | ( n1437 & n1572 ) ;
  assign n1574 = ~n271 & n1573 ;
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  assign n1577 = ( n74 & n508 ) | ( n74 & ~n1575 ) | ( n508 & ~n1575 ) ;
  assign n1578 = ( n195 & ~n430 ) | ( n195 & n1430 ) | ( ~n430 & n1430 ) ;
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1430), .o (n1581) );
  assign n1582 = ( n130 & n431 ) | ( n130 & n1581 ) | ( n431 & n1581 ) ;
  assign n1583 = n1579 & ~n1582 ;
  assign n1584 = ( ~n198 & n1580 ) | ( ~n198 & n1583 ) | ( n1580 & n1583 ) ;
  assign n1585 = ~n268 & n1584 ;
  assign n1586 = n234 & n1585 ;
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  assign n1589 = ( ~n103 & n1390 ) | ( ~n103 & n1587 ) | ( n1390 & n1587 ) ;
  assign n1590 = ( n269 & n1114 ) | ( n269 & ~n1538 ) | ( n1114 & ~n1538 ) ;
  assign n1591 = n1539 & n1590 ;
  assign n1592 = ~n1390 & n1591 ;
  assign n1593 = ( n1588 & ~n1589 ) | ( n1588 & n1592 ) | ( ~n1589 & n1592 ) ;
  assign n1594 = n508 & n1593 ;
  assign n1595 = ( n1576 & n1577 ) | ( n1576 & n1594 ) | ( n1577 & n1594 ) ;
  assign n1596 = n310 & n1595 ;
  assign n1597 = ( n1567 & n1568 ) | ( n1567 & n1596 ) | ( n1568 & n1596 ) ;
  buffer buf_n1598( .i (n91), .o (n1598) );
  assign n1599 = ~n460 & n1598 ;
  buffer buf_n1600( .i (n1599), .o (n1600) );
  assign n1603 = n1329 & ~n1600 ;
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n1605( .i (n64), .o (n1605) );
  assign n1606 = n1604 & ~n1605 ;
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  assign n1607 = ( n1300 & ~n1602 ) | ( n1300 & n1604 ) | ( ~n1602 & n1604 ) ;
  assign n1608 = ( ~n465 & n1606 ) | ( ~n465 & n1607 ) | ( n1606 & n1607 ) ;
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n1613( .i (n1612), .o (n1613) );
  assign n1614 = n271 & n1613 ;
  buffer buf_n1615( .i (n593), .o (n1615) );
  assign n1616 = ( n438 & ~n1614 ) | ( n438 & n1615 ) | ( ~n1614 & n1615 ) ;
  assign n1617 = n595 & ~n1616 ;
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  assign n1620 = ( ~n240 & n641 ) | ( ~n240 & n1618 ) | ( n641 & n1618 ) ;
  assign n1621 = n228 & ~n263 ;
  assign n1622 = n263 & n429 ;
  assign n1623 = ~n227 & n1305 ;
  assign n1624 = n429 & ~n1623 ;
  assign n1625 = ( n1621 & n1622 ) | ( n1621 & ~n1624 ) | ( n1622 & ~n1624 ) ;
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  assign n1628 = ( n466 & ~n1270 ) | ( n466 & n1626 ) | ( ~n1270 & n1626 ) ;
  assign n1629 = n1627 & ~n1628 ;
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n1633( .i (n231), .o (n1633) );
  assign n1634 = ~n1278 & n1633 ;
  buffer buf_n1635( .i (n99), .o (n1635) );
  assign n1636 = n1634 & n1635 ;
  assign n1637 = ( ~n269 & n1630 ) | ( ~n269 & n1636 ) | ( n1630 & n1636 ) ;
  assign n1638 = n534 & ~n1637 ;
  assign n1639 = ( n535 & n1632 ) | ( n535 & ~n1638 ) | ( n1632 & ~n1638 ) ;
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  assign n1642 = ( n308 & n508 ) | ( n308 & ~n1640 ) | ( n508 & ~n1640 ) ;
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  assign n1643 = n233 & ~n468 ;
  assign n1644 = ( n1251 & ~n1560 ) | ( n1251 & n1643 ) | ( ~n1560 & n1643 ) ;
  assign n1645 = n1561 & n1644 ;
  buffer buf_n1646( .i (n102), .o (n1646) );
  assign n1647 = ( n881 & n1645 ) | ( n881 & n1646 ) | ( n1645 & n1646 ) ;
  assign n1648 = ~n104 & n1647 ;
  assign n1649 = n308 & n1648 ;
  assign n1650 = ( n1641 & n1642 ) | ( n1641 & n1649 ) | ( n1642 & n1649 ) ;
  assign n1651 = ~n641 & n1650 ;
  assign n1652 = ( n1619 & ~n1620 ) | ( n1619 & n1651 ) | ( ~n1620 & n1651 ) ;
  assign n1653 = n1597 | n1652 ;
  assign n1654 = ( n1448 & ~n1449 ) | ( n1448 & n1653 ) | ( ~n1449 & n1653 ) ;
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  buffer buf_n1658( .i (n1657), .o (n1658) );
  assign n1659 = n188 & n457 ;
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1663( .i (n189), .o (n1663) );
  assign n1664 = ~n1660 & n1663 ;
  buffer buf_n1665( .i (n1664), .o (n1665) );
  assign n1666 = n93 & n1665 ;
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  assign n1667 = ( n1094 & ~n1662 ) | ( n1094 & n1665 ) | ( ~n1662 & n1665 ) ;
  assign n1668 = ( n462 & n1666 ) | ( n462 & n1667 ) | ( n1666 & n1667 ) ;
  assign n1669 = ~n455 & n1259 ;
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  assign n1673 = ( n58 & ~n843 ) | ( n58 & n1670 ) | ( ~n843 & n1670 ) ;
  assign n1674 = n458 & ~n1673 ;
  assign n1675 = ( n459 & n1672 ) | ( n459 & ~n1674 ) | ( n1672 & ~n1674 ) ;
  assign n1676 = ( n55 & n219 ) | ( n55 & ~n454 ) | ( n219 & ~n454 ) ;
  assign n1677 = ( n152 & n219 ) | ( n152 & n454 ) | ( n219 & n454 ) ;
  assign n1678 = n1676 & n1677 ;
  assign n1679 = n182 & ~n451 ;
  assign n1680 = n51 & ~n215 ;
  assign n1681 = n451 & ~n1680 ;
  assign n1682 = n1679 | n1681 ;
  assign n1683 = n151 & ~n1682 ;
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  assign n1686 = n186 | n1684 ;
  assign n1687 = ( ~n1678 & n1685 ) | ( ~n1678 & n1686 ) | ( n1685 & n1686 ) ;
  assign n1688 = n89 & n1687 ;
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  assign n1691 = n1663 | n1689 ;
  assign n1692 = ( n1675 & n1690 ) | ( n1675 & n1691 ) | ( n1690 & n1691 ) ;
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  assign n1695 = n127 & ~n1693 ;
  assign n1696 = ( n1668 & n1694 ) | ( n1668 & ~n1695 ) | ( n1694 & ~n1695 ) ;
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  assign n1707 = n298 & ~n331 ;
  buffer buf_n1708( .i (n1707), .o (n1708) );
  assign n1709 = ( n300 & n365 ) | ( n300 & n1708 ) | ( n365 & n1708 ) ;
  assign n1710 = ( ~n300 & n365 ) | ( ~n300 & n1708 ) | ( n365 & n1708 ) ;
  assign n1711 = ( n301 & ~n1709 ) | ( n301 & n1710 ) | ( ~n1709 & n1710 ) ;
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  assign n1719 = n1706 & n1718 ;
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  assign n1722 = n157 | n1263 ;
  assign n1723 = ( ~n603 & n1264 ) | ( ~n603 & n1722 ) | ( n1264 & n1722 ) ;
  buffer buf_n1724( .i (n57), .o (n1724) );
  assign n1725 = ( ~n89 & n122 ) | ( ~n89 & n1724 ) | ( n122 & n1724 ) ;
  buffer buf_n1726( .i (n88), .o (n1726) );
  assign n1727 = ( ~n155 & n1724 ) | ( ~n155 & n1726 ) | ( n1724 & n1726 ) ;
  assign n1728 = ~n1725 & n1727 ;
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  assign n1731 = n61 | n1729 ;
  assign n1732 = ( n1723 & n1730 ) | ( n1723 & n1731 ) | ( n1730 & n1731 ) ;
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  assign n1741 = n468 & n1712 ;
  assign n1742 = ( n1251 & n1739 ) | ( n1251 & ~n1741 ) | ( n1739 & ~n1741 ) ;
  assign n1743 = n1740 & ~n1742 ;
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  assign n1746 = ( n237 & n272 ) | ( n237 & ~n1744 ) | ( n272 & ~n1744 ) ;
  assign n1747 = n88 & n187 ;
  buffer buf_n1748( .i (n1747), .o (n1748) );
  assign n1762 = ~n1478 & n1724 ;
  assign n1763 = ( n1479 & n1748 ) | ( n1479 & ~n1762 ) | ( n1748 & ~n1762 ) ;
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  assign n1772 = n320 & ~n385 ;
  assign n1773 = ~n250 & n318 ;
  buffer buf_n1774( .i (n1773), .o (n1774) );
  assign n1793 = ( ~n287 & n320 ) | ( ~n287 & n1774 ) | ( n320 & n1774 ) ;
  assign n1794 = ( n719 & n1772 ) | ( n719 & ~n1793 ) | ( n1772 & ~n1793 ) ;
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  assign n1807 = ( ~n34 & n1770 ) | ( ~n34 & n1806 ) | ( n1770 & n1806 ) ;
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  assign n1808 = n193 & ~n1204 ;
  assign n1809 = n1010 & ~n1808 ;
  assign n1810 = n1605 & n1809 ;
  assign n1811 = ( n66 & n1516 ) | ( n66 & n1810 ) | ( n1516 & n1810 ) ;
  assign n1812 = ~n1806 & n1811 ;
  assign n1813 = ( n1771 & ~n1807 ) | ( n1771 & n1812 ) | ( ~n1807 & n1812 ) ;
  assign n1814 = n421 & ~n1795 ;
  buffer buf_n1815( .i (n1814), .o (n1815) );
  assign n1817 = n188 & n1815 ;
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n90), .o (n1820) );
  assign n1821 = ( ~n27 & n1818 ) | ( ~n27 & n1820 ) | ( n1818 & n1820 ) ;
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1822( .i (n154), .o (n1822) );
  assign n1823 = ( ~n25 & n1815 ) | ( ~n25 & n1822 ) | ( n1815 & n1822 ) ;
  assign n1824 = n288 & n321 ;
  buffer buf_n1825( .i (n1824), .o (n1825) );
  assign n1843 = n255 & ~n1825 ;
  assign n1844 = ~n422 & n1843 ;
  assign n1845 = ~n1822 & n1844 ;
  assign n1846 = ( n1816 & ~n1823 ) | ( n1816 & n1845 ) | ( ~n1823 & n1845 ) ;
  assign n1847 = ~n1820 & n1846 ;
  assign n1848 = ( n1819 & ~n1821 ) | ( n1819 & n1847 ) | ( ~n1821 & n1847 ) ;
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  assign n1852 = ( n61 & n191 ) | ( n61 & ~n1800 ) | ( n191 & ~n1800 ) ;
  assign n1853 = ( n158 & n191 ) | ( n158 & n1800 ) | ( n191 & n1800 ) ;
  assign n1854 = n1852 & ~n1853 ;
  assign n1855 = ( n1305 & n1849 ) | ( n1305 & n1854 ) | ( n1849 & n1854 ) ;
  assign n1856 = n429 & ~n1855 ;
  assign n1857 = ( n430 & n1851 ) | ( n430 & ~n1856 ) | ( n1851 & ~n1856 ) ;
  assign n1858 = n130 & n1857 ;
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1860( .i (n1859), .o (n1860) );
  assign n1861 = n433 | n1859 ;
  assign n1862 = ( n1813 & n1860 ) | ( n1813 & n1861 ) | ( n1860 & n1861 ) ;
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n1865( .i (n469), .o (n1865) );
  assign n1866 = ( ~n370 & n1863 ) | ( ~n370 & n1865 ) | ( n1863 & n1865 ) ;
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n1867( .i (n187), .o (n1867) );
  assign n1868 = ( n1726 & n1822 ) | ( n1726 & ~n1867 ) | ( n1822 & ~n1867 ) ;
  assign n1869 = n123 & ~n1868 ;
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  assign n1872 = ( n1521 & n1764 ) | ( n1521 & ~n1870 ) | ( n1764 & ~n1870 ) ;
  assign n1873 = ( n1530 & n1871 ) | ( n1530 & n1872 ) | ( n1871 & n1872 ) ;
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n1876( .i (n1875), .o (n1876) );
  assign n1887 = ( n300 & n492 ) | ( n300 & n1876 ) | ( n492 & n1876 ) ;
  assign n1888 = n328 & ~n360 ;
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  assign n1902 = n1876 & n1892 ;
  assign n1903 = ( ~n301 & n1887 ) | ( ~n301 & n1902 ) | ( n1887 & n1902 ) ;
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  assign n1906 = ( n268 & n434 ) | ( n268 & ~n1904 ) | ( n434 & ~n1904 ) ;
  assign n1907 = n789 & ~n1598 ;
  buffer buf_n1908( .i (n1907), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  buffer buf_n1915( .i (n430), .o (n1915) );
  assign n1916 = n1835 & ~n1915 ;
  assign n1917 = ( n366 & n1912 ) | ( n366 & n1916 ) | ( n1912 & n1916 ) ;
  assign n1918 = ~n367 & n1917 ;
  assign n1919 = n268 & n1918 ;
  assign n1920 = ( n1905 & n1906 ) | ( n1905 & n1919 ) | ( n1906 & n1919 ) ;
  assign n1921 = ~n1865 & n1920 ;
  assign n1922 = ( n1864 & ~n1866 ) | ( n1864 & n1921 ) | ( ~n1866 & n1921 ) ;
  assign n1923 = n237 & n1922 ;
  assign n1924 = ( n1745 & n1746 ) | ( n1745 & n1923 ) | ( n1746 & n1923 ) ;
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  assign n1928 = ( ~n441 & n1291 ) | ( ~n441 & n1925 ) | ( n1291 & n1925 ) ;
  assign n1929 = n1720 & ~n1928 ;
  assign n1930 = ( n1721 & n1927 ) | ( n1721 & ~n1929 ) | ( n1927 & ~n1929 ) ;
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n1934( .i (n1933), .o (n1934) );
  buffer buf_n1935( .i (n1934), .o (n1935) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n1936( .i (n156), .o (n1936) );
  assign n1937 = n224 & ~n1936 ;
  buffer buf_n1938( .i (n1937), .o (n1938) );
  assign n1945 = n192 | n1938 ;
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  assign n1952 = ( n433 & ~n1609 ) | ( n433 & n1950 ) | ( ~n1609 & n1950 ) ;
  assign n1953 = ( n124 & n224 ) | ( n124 & ~n1820 ) | ( n224 & ~n1820 ) ;
  buffer buf_n1954( .i (n223), .o (n1954) );
  assign n1955 = ( n1820 & n1936 ) | ( n1820 & n1954 ) | ( n1936 & n1954 ) ;
  assign n1956 = ~n1953 & n1955 ;
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  assign n1959 = ( n123 & n189 ) | ( n123 & ~n223 ) | ( n189 & ~n223 ) ;
  assign n1960 = n1936 & ~n1959 ;
  buffer buf_n1961( .i (n1960), .o (n1961) );
  assign n1971 = ~n90 & n223 ;
  assign n1972 = n124 & n1971 ;
  buffer buf_n1973( .i (n1972), .o (n1973) );
  assign n1983 = ( n461 & n1961 ) | ( n461 & n1973 ) | ( n1961 & n1973 ) ;
  assign n1984 = ~n1957 & n1983 ;
  assign n1985 = ( n463 & n1958 ) | ( n463 & n1984 ) | ( n1958 & n1984 ) ;
  buffer buf_n1986( .i (n1985), .o (n1986) );
  buffer buf_n1987( .i (n1986), .o (n1987) );
  assign n1988 = ~n66 & n1986 ;
  assign n1989 = n457 | n1726 ;
  assign n1990 = n57 & n121 ;
  assign n1991 = n457 & ~n1990 ;
  assign n1992 = n1989 & ~n1991 ;
  buffer buf_n1993( .i (n1992), .o (n1993) );
  buffer buf_n1994( .i (n1993), .o (n1994) );
  assign n1995 = ~n225 & n1993 ;
  assign n1996 = ( ~n1327 & n1994 ) | ( ~n1327 & n1995 ) | ( n1994 & n1995 ) ;
  buffer buf_n1997( .i (n1996), .o (n1997) );
  buffer buf_n1998( .i (n1997), .o (n1998) );
  assign n1999 = ( n225 & n460 ) | ( n225 & ~n1598 ) | ( n460 & ~n1598 ) ;
  assign n2000 = ( ~n125 & n460 ) | ( ~n125 & n1598 ) | ( n460 & n1598 ) ;
  assign n2001 = ~n1999 & n2000 ;
  assign n2002 = n459 & ~n1954 ;
  assign n2003 = ( n61 & n158 ) | ( n61 & n2002 ) | ( n158 & n2002 ) ;
  assign n2004 = ~n1327 & n2003 ;
  assign n2005 = ( n193 & n2001 ) | ( n193 & n2004 ) | ( n2001 & n2004 ) ;
  assign n2006 = ~n1997 & n2005 ;
  assign n2007 = ( n195 & n1998 ) | ( n195 & n2006 ) | ( n1998 & n2006 ) ;
  assign n2008 = n1332 | n2007 ;
  assign n2009 = ( n1987 & ~n1988 ) | ( n1987 & n2008 ) | ( ~n1988 & n2008 ) ;
  buffer buf_n2010( .i (n432), .o (n2010) );
  assign n2011 = n2009 & ~n2010 ;
  assign n2012 = ( n1951 & ~n1952 ) | ( n1951 & n2011 ) | ( ~n1952 & n2011 ) ;
  buffer buf_n2013( .i (n2012), .o (n2013) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  assign n2015 = n323 & n355 ;
  buffer buf_n2016( .i (n2015), .o (n2016) );
  buffer buf_n2017( .i (n2016), .o (n2017) );
  buffer buf_n2018( .i (n2017), .o (n2018) );
  buffer buf_n2019( .i (n2018), .o (n2019) );
  buffer buf_n2020( .i (n2019), .o (n2020) );
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  assign n2031 = n336 & ~n2027 ;
  buffer buf_n2032( .i (n2031), .o (n2032) );
  assign n2033 = n2013 & n2032 ;
  buffer buf_n2028( .i (n2027), .o (n2028) );
  buffer buf_n2029( .i (n2028), .o (n2029) );
  assign n2034 = ~n161 & n1267 ;
  buffer buf_n2035( .i (n428), .o (n2035) );
  buffer buf_n2036( .i (n2035), .o (n2036) );
  assign n2037 = n2034 & ~n2036 ;
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  assign n2040 = n1874 & n2035 ;
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  assign n2050 = n463 & n1733 ;
  assign n2051 = ~n2036 & n2050 ;
  buffer buf_n2052( .i (n2051), .o (n2052) );
  assign n2055 = ( ~n2038 & n2042 ) | ( ~n2038 & n2052 ) | ( n2042 & n2052 ) ;
  assign n2056 = n466 & ~n2052 ;
  assign n2057 = ( n2039 & n2055 ) | ( n2039 & ~n2056 ) | ( n2055 & ~n2056 ) ;
  assign n2058 = n1697 & ~n1915 ;
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  assign n2065 = n1633 | n2059 ;
  assign n2066 = ( n2057 & n2060 ) | ( n2057 & n2065 ) | ( n2060 & n2065 ) ;
  buffer buf_n2067( .i (n2066), .o (n2067) );
  assign n2068 = ( ~n2029 & n2032 ) | ( ~n2029 & n2067 ) | ( n2032 & n2067 ) ;
  assign n2069 = ( n371 & n2033 ) | ( n371 & n2068 ) | ( n2033 & n2068 ) ;
  assign n2070 = n272 & ~n2069 ;
  buffer buf_n2014( .i (n2013), .o (n2014) );
  assign n2071 = n371 & n2014 ;
  buffer buf_n2072( .i (n271), .o (n2072) );
  assign n2073 = n2071 | n2072 ;
  assign n2074 = ~n2070 & n2073 ;
  assign n2075 = n309 & n2074 ;
  buffer buf_n2076( .i (n2075), .o (n2076) );
  buffer buf_n2077( .i (n2076), .o (n2077) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  buffer buf_n1879( .i (n1878), .o (n1879) );
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  buffer buf_n1886( .i (n1885), .o (n1886) );
  assign n2078 = n236 | n371 ;
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n2079( .i (n370), .o (n2079) );
  assign n2080 = ( n236 & n704 ) | ( n236 & ~n2079 ) | ( n704 & ~n2079 ) ;
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1897( .i (n1896), .o (n1897) );
  assign n2081 = n301 | n399 ;
  assign n2082 = ( n302 & n367 ) | ( n302 & ~n2081 ) | ( n367 & ~n2081 ) ;
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n337( .i (n336), .o (n337) );
  assign n2085 = ( ~n337 & n369 ) | ( ~n337 & n2083 ) | ( n369 & n2083 ) ;
  assign n2086 = ( n1897 & ~n2084 ) | ( n1897 & n2085 ) | ( ~n2084 & n2085 ) ;
  assign n2087 = n236 & n2086 ;
  assign n2088 = ( n2078 & ~n2080 ) | ( n2078 & n2087 ) | ( ~n2080 & n2087 ) ;
  assign n2089 = n439 & n2088 ;
  assign n2090 = ( n474 & n1885 ) | ( n474 & ~n2089 ) | ( n1885 & ~n2089 ) ;
  assign n2091 = n1886 & ~n2090 ;
  assign n2092 = n2076 | n2091 ;
  assign n2093 = ( n277 & n2077 ) | ( n277 & n2092 ) | ( n2077 & n2092 ) ;
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2099( .i (n1865), .o (n2099) );
  assign n2100 = n2047 & ~n2099 ;
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n2102( .i (n2101), .o (n2102) );
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  assign n2107 = ( n378 & n558 ) | ( n378 & n2106 ) | ( n558 & n2106 ) ;
  assign n2108 = ~n379 & n2107 ;
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  assign n2111 = ( n270 & n370 ) | ( n270 & n2067 ) | ( n370 & n2067 ) ;
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  assign n2116 = ~n372 & n2112 ;
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  buffer buf_n2119( .i (n273), .o (n2119) );
  assign n2120 = ( n309 & n2117 ) | ( n309 & ~n2119 ) | ( n2117 & ~n2119 ) ;
  assign n2121 = ( n2115 & n2118 ) | ( n2115 & n2120 ) | ( n2118 & n2120 ) ;
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n359), .o (n2124) );
  assign n2125 = n393 & n2124 ;
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  buffer buf_n2129( .i (n2128), .o (n2129) );
  buffer buf_n2130( .i (n2129), .o (n2130) );
  buffer buf_n2131( .i (n2130), .o (n2131) );
  buffer buf_n2132( .i (n2131), .o (n2132) );
  buffer buf_n2133( .i (n2132), .o (n2133) );
  assign n2134 = ( ~n369 & n2045 ) | ( ~n369 & n2133 ) | ( n2045 & n2133 ) ;
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n2137( .i (n267), .o (n2137) );
  assign n2138 = n1914 & n2137 ;
  assign n2139 = ( n369 & n1251 ) | ( n369 & n2138 ) | ( n1251 & n2138 ) ;
  assign n2140 = ~n436 & n2139 ;
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  assign n2141 = n368 & n2054 ;
  buffer buf_n2142( .i (n2137), .o (n2142) );
  assign n2143 = n2141 & n2142 ;
  buffer buf_n2144( .i (n2143), .o (n2144) );
  assign n2145 = ( ~n2135 & n2140 ) | ( ~n2135 & n2144 ) | ( n2140 & n2144 ) ;
  assign n2146 = n2099 & ~n2144 ;
  assign n2147 = ( n2136 & n2145 ) | ( n2136 & ~n2146 ) | ( n2145 & ~n2146 ) ;
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  assign n2150 = ( ~n239 & n309 ) | ( ~n239 & n2148 ) | ( n309 & n2148 ) ;
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  buffer buf_n2064( .i (n2063), .o (n2064) );
  assign n2151 = n372 & n2064 ;
  assign n2152 = n273 & n2151 ;
  buffer buf_n2153( .i (n307), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  assign n2155 = n2152 & ~n2154 ;
  assign n2156 = ( n2149 & ~n2150 ) | ( n2149 & n2155 ) | ( ~n2150 & n2155 ) ;
  assign n2157 = n373 & n2101 ;
  assign n2158 = ( n239 & n2119 ) | ( n239 & n2157 ) | ( n2119 & n2157 ) ;
  assign n2159 = ~n240 & n2158 ;
  assign n2160 = ( n344 & n2156 ) | ( n344 & n2159 ) | ( n2156 & n2159 ) ;
  assign n2161 = ~n2122 & n2160 ;
  assign n2162 = ( n346 & n2123 ) | ( n346 & n2161 ) | ( n2123 & n2161 ) ;
  buffer buf_n2163( .i (n2162), .o (n2163) );
  buffer buf_n2164( .i (n2163), .o (n2164) );
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n280( .i (n279), .o (n280) );
  assign n2166 = ( n245 & ~n280 ) | ( n245 & n2163 ) | ( ~n280 & n2163 ) ;
  assign n2167 = n2109 & ~n2166 ;
  assign n2168 = ( n2110 & n2165 ) | ( n2110 & ~n2167 ) | ( n2165 & ~n2167 ) ;
  assign n2169 = ( n230 & n333 ) | ( n230 & n2041 ) | ( n333 & n2041 ) ;
  assign n2170 = n330 & n1908 ;
  assign n2171 = ( n363 & n2035 ) | ( n363 & n2170 ) | ( n2035 & n2170 ) ;
  assign n2172 = ~n2036 & n2171 ;
  assign n2173 = n230 & n2172 ;
  assign n2174 = ( ~n334 & n2169 ) | ( ~n334 & n2173 ) | ( n2169 & n2173 ) ;
  buffer buf_n2175( .i (n2174), .o (n2175) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n1915), .o (n2178) );
  assign n2179 = ( n98 & n609 ) | ( n98 & ~n2178 ) | ( n609 & ~n2178 ) ;
  buffer buf_n2180( .i (n123), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  assign n2182 = n225 & n2181 ;
  assign n2183 = n1327 & n2182 ;
  buffer buf_n2184( .i (n2183), .o (n2184) );
  buffer buf_n2192( .i (n192), .o (n2192) );
  buffer buf_n2193( .i (n2192), .o (n2193) );
  assign n2194 = ~n2184 & n2193 ;
  buffer buf_n2195( .i (n2193), .o (n2195) );
  assign n2196 = ( n1011 & n2194 ) | ( n1011 & ~n2195 ) | ( n2194 & ~n2195 ) ;
  buffer buf_n2197( .i (n2196), .o (n2197) );
  assign n2199 = ( n98 & n2178 ) | ( n98 & ~n2197 ) | ( n2178 & ~n2197 ) ;
  assign n2200 = n2179 & ~n2199 ;
  assign n2201 = ( n336 & n2175 ) | ( n336 & n2200 ) | ( n2175 & n2200 ) ;
  buffer buf_n2202( .i (n368), .o (n2202) );
  assign n2203 = ~n2201 & n2202 ;
  buffer buf_n2204( .i (n2202), .o (n2204) );
  assign n2205 = ( n2177 & ~n2203 ) | ( n2177 & n2204 ) | ( ~n2203 & n2204 ) ;
  assign n2206 = ~n306 & n2205 ;
  buffer buf_n2207( .i (n2206), .o (n2207) );
  buffer buf_n2208( .i (n2207), .o (n2208) );
  buffer buf_n2198( .i (n2197), .o (n2198) );
  buffer buf_n2209( .i (n1428), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  assign n2211 = ~n2198 & n2210 ;
  buffer buf_n2212( .i (n126), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  buffer buf_n2214( .i (n2213), .o (n2214) );
  assign n2215 = n1947 & n2214 ;
  buffer buf_n2216( .i (n2215), .o (n2216) );
  assign n2223 = ~n2209 & n2216 ;
  buffer buf_n2224( .i (n2223), .o (n2224) );
  assign n2230 = ( n1635 & ~n2211 ) | ( n1635 & n2224 ) | ( ~n2211 & n2224 ) ;
  assign n2231 = ( n337 & n2202 ) | ( n337 & ~n2230 ) | ( n2202 & ~n2230 ) ;
  buffer buf_n2232( .i (n2231), .o (n2232) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  assign n2234 = n339 & ~n2232 ;
  assign n2235 = ( n372 & ~n2233 ) | ( n372 & n2234 ) | ( ~n2233 & n2234 ) ;
  assign n2236 = n2207 | n2235 ;
  buffer buf_n2237( .i (n439), .o (n2237) );
  assign n2238 = ( n2208 & n2236 ) | ( n2208 & ~n2237 ) | ( n2236 & ~n2237 ) ;
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  assign n2241 = ~n276 & n2239 ;
  assign n2242 = ( ~n336 & n368 ) | ( ~n336 & n2137 ) | ( n368 & n2137 ) ;
  assign n2243 = n337 & ~n2242 ;
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  assign n2246 = ~n338 & n2204 ;
  assign n2247 = ( n306 & n2244 ) | ( n306 & n2246 ) | ( n2244 & n2246 ) ;
  assign n2248 = n2245 | n2247 ;
  assign n2249 = n439 & n2248 ;
  assign n2250 = ( n239 & ~n1885 ) | ( n239 & n2249 ) | ( ~n1885 & n2249 ) ;
  assign n2251 = n1886 & n2250 ;
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n2225( .i (n2224), .o (n2225) );
  buffer buf_n2226( .i (n2225), .o (n2226) );
  buffer buf_n2227( .i (n2226), .o (n2227) );
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n2252( .i (n133), .o (n2252) );
  assign n2253 = ( ~n101 & n1415 ) | ( ~n101 & n2252 ) | ( n1415 & n2252 ) ;
  assign n2254 = n651 & ~n2253 ;
  buffer buf_n2255( .i (n201), .o (n2255) );
  assign n2256 = ( n652 & n2254 ) | ( n652 & ~n2255 ) | ( n2254 & ~n2255 ) ;
  assign n2257 = ~n2228 & n2256 ;
  assign n2258 = ( n834 & n2229 ) | ( n834 & n2257 ) | ( n2229 & n2257 ) ;
  assign n2259 = ( ~n1901 & n2119 ) | ( ~n1901 & n2258 ) | ( n2119 & n2258 ) ;
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  assign n2260 = ( n237 & n2048 ) | ( n237 & ~n2072 ) | ( n2048 & ~n2072 ) ;
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  assign n2261 = n1126 & n1761 ;
  buffer buf_n2262( .i (n235), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  assign n2264 = n2261 & ~n2263 ;
  assign n2265 = ( n2049 & ~n2260 ) | ( n2049 & n2264 ) | ( ~n2260 & n2264 ) ;
  assign n2266 = ~n1901 & n2265 ;
  assign n2267 = ( ~n1291 & n2259 ) | ( ~n1291 & n2266 ) | ( n2259 & n2266 ) ;
  assign n2268 = n2251 | n2267 ;
  assign n2269 = ( n2240 & ~n2241 ) | ( n2240 & n2268 ) | ( ~n2241 & n2268 ) ;
  buffer buf_n2270( .i (n2269), .o (n2270) );
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n479( .i (n478), .o (n479) );
  assign n2272 = ( ~n412 & n479 ) | ( ~n412 & n2270 ) | ( n479 & n2270 ) ;
  assign n2273 = ( ~n72 & n1033 ) | ( ~n72 & n2262 ) | ( n1033 & n2262 ) ;
  assign n2274 = ( n60 & n1936 ) | ( n60 & n1954 ) | ( n1936 & n1954 ) ;
  buffer buf_n2275( .i (n2274), .o (n2275) );
  buffer buf_n2276( .i (n2275), .o (n2276) );
  buffer buf_n2277( .i (n2276), .o (n2277) );
  buffer buf_n2278( .i (n2277), .o (n2278) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  buffer buf_n2280( .i (n2279), .o (n2280) );
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  assign n2287 = ~n2273 & n2286 ;
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n2289( .i (n2288), .o (n2289) );
  buffer buf_n2290( .i (n1867), .o (n2290) );
  buffer buf_n2291( .i (n222), .o (n2291) );
  assign n2292 = n2290 & ~n2291 ;
  buffer buf_n2293( .i (n2292), .o (n2293) );
  buffer buf_n2294( .i (n2293), .o (n2294) );
  buffer buf_n2295( .i (n2294), .o (n2295) );
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n2297( .i (n2296), .o (n2297) );
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  assign n2307 = ( ~n170 & n203 ) | ( ~n170 & n2263 ) | ( n203 & n2263 ) ;
  assign n2308 = n72 & n2262 ;
  buffer buf_n2309( .i (n2308), .o (n2309) );
  assign n2310 = ( n2306 & n2307 ) | ( n2306 & ~n2309 ) | ( n2307 & ~n2309 ) ;
  assign n2311 = n200 & ~n855 ;
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n1967( .i (n1966), .o (n1967) );
  buffer buf_n1968( .i (n1967), .o (n1968) );
  buffer buf_n1969( .i (n1968), .o (n1969) );
  buffer buf_n1970( .i (n1969), .o (n1970) );
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  assign n2314 = ( n71 & n1970 ) | ( n71 & n1982 ) | ( n1970 & n1982 ) ;
  assign n2315 = ~n2312 & n2314 ;
  assign n2316 = ( n73 & n2313 ) | ( n73 & n2315 ) | ( n2313 & n2315 ) ;
  buffer buf_n2317( .i (n2316), .o (n2317) );
  assign n2318 = ( ~n2288 & n2310 ) | ( ~n2288 & n2317 ) | ( n2310 & n2317 ) ;
  assign n2319 = n106 | n2317 ;
  assign n2320 = ( n2289 & n2318 ) | ( n2289 & n2319 ) | ( n2318 & n2319 ) ;
  buffer buf_n2321( .i (n2320), .o (n2321) );
  buffer buf_n2322( .i (n2321), .o (n2322) );
  assign n2323 = ( n342 & n374 ) | ( n342 & n2119 ) | ( n374 & n2119 ) ;
  buffer buf_n2324( .i (n2072), .o (n2324) );
  assign n2325 = ( n373 & n2153 ) | ( n373 & ~n2324 ) | ( n2153 & ~n2324 ) ;
  assign n2326 = n342 & n2325 ;
  assign n2327 = ( n1053 & n2323 ) | ( n1053 & ~n2326 ) | ( n2323 & ~n2326 ) ;
  assign n2328 = n476 & n2327 ;
  assign n2329 = ( n443 & n2321 ) | ( n443 & ~n2328 ) | ( n2321 & ~n2328 ) ;
  assign n2330 = n2322 & ~n2329 ;
  assign n2331 = n412 & n2330 ;
  assign n2332 = ( n2271 & ~n2272 ) | ( n2271 & n2331 ) | ( ~n2272 & n2331 ) ;
  buffer buf_n2333( .i (n2332), .o (n2333) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n111( .i (n110), .o (n111) );
  assign n2335 = ( n259 & n294 ) | ( n259 & n359 ) | ( n294 & n359 ) ;
  assign n2336 = ( ~n328 & n2124 ) | ( ~n328 & n2335 ) | ( n2124 & n2335 ) ;
  buffer buf_n2337( .i (n2336), .o (n2337) );
  assign n2340 = n362 & ~n2337 ;
  buffer buf_n2341( .i (n2340), .o (n2341) );
  buffer buf_n2342( .i (n2341), .o (n2342) );
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  assign n2343 = n2339 | n2341 ;
  assign n2344 = ( ~n365 & n2342 ) | ( ~n365 & n2343 ) | ( n2342 & n2343 ) ;
  buffer buf_n2345( .i (n2344), .o (n2345) );
  buffer buf_n2346( .i (n2345), .o (n2346) );
  assign n2350 = ( ~n1068 & n2010 ) | ( ~n1068 & n2345 ) | ( n2010 & n2345 ) ;
  assign n2351 = n2346 & ~n2350 ;
  buffer buf_n2352( .i (n2351), .o (n2352) );
  buffer buf_n2353( .i (n2352), .o (n2353) );
  assign n2354 = ( n259 & ~n294 ) | ( n259 & n327 ) | ( ~n294 & n327 ) ;
  buffer buf_n2355( .i (n2354), .o (n2355) );
  buffer buf_n2356( .i (n2355), .o (n2356) );
  assign n2357 = ( n296 & n361 ) | ( n296 & ~n2355 ) | ( n361 & ~n2355 ) ;
  assign n2358 = n2356 & ~n2357 ;
  assign n2359 = n1041 | n2358 ;
  buffer buf_n2360( .i (n2359), .o (n2360) );
  buffer buf_n2361( .i (n2360), .o (n2361) );
  buffer buf_n2362( .i (n2361), .o (n2362) );
  buffer buf_n2363( .i (n2362), .o (n2363) );
  buffer buf_n2364( .i (n2363), .o (n2364) );
  assign n2368 = n35 & n2010 ;
  assign n2369 = ( n1635 & ~n2363 ) | ( n1635 & n2368 ) | ( ~n2363 & n2368 ) ;
  assign n2370 = n2364 & n2369 ;
  assign n2371 = ( n33 & n66 ) | ( n33 & n2360 ) | ( n66 & n2360 ) ;
  buffer buf_n2372( .i (n32), .o (n2372) );
  buffer buf_n2373( .i (n2195), .o (n2373) );
  assign n2374 = ( ~n2360 & n2372 ) | ( ~n2360 & n2373 ) | ( n2372 & n2373 ) ;
  assign n2375 = n2371 & ~n2374 ;
  assign n2376 = n2010 & n2375 ;
  assign n2377 = n1635 & n2376 ;
  buffer buf_n2378( .i (n2377), .o (n2378) );
  assign n2379 = ( ~n2352 & n2370 ) | ( ~n2352 & n2378 ) | ( n2370 & n2378 ) ;
  assign n2380 = n135 & ~n2378 ;
  assign n2381 = ( n2353 & n2379 ) | ( n2353 & ~n2380 ) | ( n2379 & ~n2380 ) ;
  assign n2382 = n170 & n2381 ;
  buffer buf_n2383( .i (n2382), .o (n2383) );
  buffer buf_n2384( .i (n2383), .o (n2384) );
  assign n2385 = n70 | n798 ;
  buffer buf_n2386( .i (n36), .o (n2386) );
  assign n2387 = n200 & n2386 ;
  assign n2388 = ( n799 & ~n2385 ) | ( n799 & n2387 ) | ( ~n2385 & n2387 ) ;
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2391( .i (n2373), .o (n2391) );
  buffer buf_n2392( .i (n2391), .o (n2392) );
  buffer buf_n2393( .i (n2392), .o (n2393) );
  assign n2394 = ( n36 & ~n69 ) | ( n36 & n2393 ) | ( ~n69 & n2393 ) ;
  buffer buf_n2395( .i (n2394), .o (n2395) );
  buffer buf_n2396( .i (n200), .o (n2396) );
  assign n2397 = ( n135 & ~n2395 ) | ( n135 & n2396 ) | ( ~n2395 & n2396 ) ;
  buffer buf_n2398( .i (n2252), .o (n2398) );
  assign n2399 = ( ~n38 & n2395 ) | ( ~n38 & n2398 ) | ( n2395 & n2398 ) ;
  assign n2400 = n2397 & ~n2399 ;
  assign n2401 = ~n2389 & n2400 ;
  buffer buf_n2365( .i (n2364), .o (n2365) );
  buffer buf_n2366( .i (n2365), .o (n2366) );
  buffer buf_n2367( .i (n2366), .o (n2367) );
  assign n2402 = n438 & n2367 ;
  assign n2403 = ( n2390 & n2401 ) | ( n2390 & n2402 ) | ( n2401 & n2402 ) ;
  assign n2404 = n2383 | n2403 ;
  assign n2405 = ( n107 & n2384 ) | ( n107 & n2404 ) | ( n2384 & n2404 ) ;
  assign n2406 = n409 & n2405 ;
  buffer buf_n2407( .i (n2406), .o (n2407) );
  buffer buf_n2408( .i (n2407), .o (n2408) );
  assign n2409 = ( n341 & n406 ) | ( n341 & n2324 ) | ( n406 & n2324 ) ;
  buffer buf_n2410( .i (n305), .o (n2410) );
  assign n2411 = n2079 | n2410 ;
  buffer buf_n2412( .i (n2411), .o (n2412) );
  assign n2419 = n341 & ~n2412 ;
  assign n2420 = ( ~n407 & n2409 ) | ( ~n407 & n2419 ) | ( n2409 & n2419 ) ;
  buffer buf_n2421( .i (n2420), .o (n2421) );
  buffer buf_n2422( .i (n2421), .o (n2422) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  assign n2423 = n742 & ~n2421 ;
  assign n2424 = n164 & ~n609 ;
  buffer buf_n2425( .i (n1605), .o (n2425) );
  assign n2426 = n2373 & ~n2425 ;
  assign n2427 = ( ~n164 & n609 ) | ( ~n164 & n2426 ) | ( n609 & n2426 ) ;
  assign n2428 = n2424 | n2427 ;
  assign n2429 = ( n28 & n191 ) | ( n28 & ~n2181 ) | ( n191 & ~n2181 ) ;
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  assign n2432 = n31 & n2431 ;
  assign n2433 = ( n1295 & n1305 ) | ( n1295 & ~n2430 ) | ( n1305 & ~n2430 ) ;
  assign n2434 = n2431 | n2433 ;
  assign n2435 = ~n2432 & n2434 ;
  assign n2436 = n2425 & n2435 ;
  buffer buf_n2437( .i (n2436), .o (n2437) );
  buffer buf_n2438( .i (n2437), .o (n2438) );
  assign n2439 = n35 | n2437 ;
  assign n2440 = ( n2428 & n2438 ) | ( n2428 & n2439 ) | ( n2438 & n2439 ) ;
  buffer buf_n2441( .i (n2440), .o (n2441) );
  assign n2449 = n436 & n2441 ;
  buffer buf_n2450( .i (n2449), .o (n2450) );
  buffer buf_n2451( .i (n2450), .o (n2451) );
  buffer buf_n2452( .i (n2451), .o (n2452) );
  buffer buf_n2453( .i (n2452), .o (n2453) );
  buffer buf_n2454( .i (n2453), .o (n2454) );
  buffer buf_n2455( .i (n2454), .o (n2455) );
  assign n2456 = ( n2422 & n2423 ) | ( n2422 & n2455 ) | ( n2423 & n2455 ) ;
  assign n2457 = n2407 | n2456 ;
  assign n2458 = ( n111 & n2408 ) | ( n111 & n2457 ) | ( n2408 & n2457 ) ;
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n2460( .i (n2459), .o (n2460) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  assign n2461 = ( ~n246 & n481 ) | ( ~n246 & n2459 ) | ( n481 & n2459 ) ;
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  assign n2462 = n918 | n1226 ;
  buffer buf_n2463( .i (n2462), .o (n2463) );
  buffer buf_n2464( .i (n2463), .o (n2464) );
  assign n2465 = n406 | n2412 ;
  assign n2466 = n2237 | n2465 ;
  buffer buf_n2467( .i (n2263), .o (n2467) );
  buffer buf_n2468( .i (n2467), .o (n2468) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  assign n2470 = ( ~n2463 & n2466 ) | ( ~n2463 & n2469 ) | ( n2466 & n2469 ) ;
  assign n2471 = ( n104 & ~n507 ) | ( n104 & n2450 ) | ( ~n507 & n2450 ) ;
  buffer buf_n2472( .i (n507), .o (n2472) );
  assign n2473 = n2471 & n2472 ;
  assign n2474 = n303 & ~n2393 ;
  assign n2475 = ~n1222 & n2474 ;
  assign n2476 = n2029 & n2475 ;
  assign n2477 = ( n404 & n1286 ) | ( n404 & n2476 ) | ( n1286 & n2476 ) ;
  buffer buf_n2478( .i (n1286), .o (n2478) );
  assign n2479 = n2477 & ~n2478 ;
  assign n2480 = n2324 & n2479 ;
  buffer buf_n2481( .i (n2324), .o (n2481) );
  assign n2482 = ( n2473 & n2480 ) | ( n2473 & n2481 ) | ( n2480 & n2481 ) ;
  assign n2483 = ~n2469 & n2482 ;
  assign n2484 = ( n2464 & n2470 ) | ( n2464 & ~n2483 ) | ( n2470 & ~n2483 ) ;
  buffer buf_n2485( .i (n2484), .o (n2485) );
  buffer buf_n2486( .i (n2485), .o (n2486) );
  buffer buf_n2487( .i (n2486), .o (n2487) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  buffer buf_n2443( .i (n2442), .o (n2443) );
  buffer buf_n2444( .i (n2443), .o (n2444) );
  buffer buf_n2445( .i (n2444), .o (n2445) );
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n2448( .i (n2447), .o (n2448) );
  assign n2488 = ~n405 & n2478 ;
  buffer buf_n2489( .i (n2488), .o (n2489) );
  buffer buf_n2490( .i (n2489), .o (n2490) );
  buffer buf_n2491( .i (n2490), .o (n2491) );
  assign n2492 = ( n376 & ~n2447 ) | ( n376 & n2491 ) | ( ~n2447 & n2491 ) ;
  assign n2493 = n2448 & n2492 ;
  assign n2494 = ( n110 & ~n2485 ) | ( n110 & n2493 ) | ( ~n2485 & n2493 ) ;
  assign n2495 = n279 & ~n2494 ;
  assign n2496 = ( ~n280 & n2487 ) | ( ~n280 & n2495 ) | ( n2487 & n2495 ) ;
  assign n2497 = n481 | n2496 ;
  assign n2498 = ( ~n2460 & n2461 ) | ( ~n2460 & n2497 ) | ( n2461 & n2497 ) ;
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n2499( .i (n165), .o (n2499) );
  assign n2500 = n2137 & n2499 ;
  buffer buf_n2501( .i (n2500), .o (n2501) );
  buffer buf_n2502( .i (n2501), .o (n2502) );
  buffer buf_n2503( .i (n2502), .o (n2503) );
  buffer buf_n2504( .i (n2503), .o (n2504) );
  buffer buf_n2505( .i (n2504), .o (n2505) );
  buffer buf_n2506( .i (n2505), .o (n2506) );
  assign n2507 = ( n206 & n1228 ) | ( n206 & n2506 ) | ( n1228 & n2506 ) ;
  assign n2508 = ~n1229 & n2507 ;
  buffer buf_n2509( .i (n2508), .o (n2509) );
  buffer buf_n2510( .i (n2509), .o (n2510) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  assign n2511 = ~n374 & n407 ;
  buffer buf_n2512( .i (n2237), .o (n2512) );
  assign n2513 = n2511 & ~n2512 ;
  assign n2514 = ~n344 & n2513 ;
  assign n2515 = n312 & n2514 ;
  assign n2516 = ( n478 & n2509 ) | ( n478 & ~n2515 ) | ( n2509 & ~n2515 ) ;
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  assign n2517 = ( n126 & n1062 ) | ( n126 & ~n1080 ) | ( n1062 & ~n1080 ) ;
  assign n2518 = ~n121 & n187 ;
  buffer buf_n2519( .i (n2518), .o (n2519) );
  assign n2528 = ( n59 & n90 ) | ( n59 & n2519 ) | ( n90 & n2519 ) ;
  buffer buf_n2529( .i (n1726), .o (n2529) );
  buffer buf_n2530( .i (n2529), .o (n2530) );
  assign n2531 = n2528 & ~n2530 ;
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n2532), .o (n2533) );
  buffer buf_n2534( .i (n156), .o (n2534) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  buffer buf_n2536( .i (n2535), .o (n2536) );
  assign n2537 = n2532 | n2536 ;
  assign n2538 = ( ~n2517 & n2533 ) | ( ~n2517 & n2537 ) | ( n2533 & n2537 ) ;
  buffer buf_n2539( .i (n2538), .o (n2539) );
  assign n2551 = n2036 & n2539 ;
  buffer buf_n2552( .i (n2551), .o (n2552) );
  buffer buf_n2553( .i (n2552), .o (n2553) );
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2555( .i (n2554), .o (n2555) );
  buffer buf_n2556( .i (n2555), .o (n2556) );
  buffer buf_n2557( .i (n2556), .o (n2557) );
  buffer buf_n2558( .i (n2557), .o (n2558) );
  buffer buf_n2559( .i (n2558), .o (n2559) );
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  assign n2563 = ( n44 & ~n765 ) | ( n44 & n2562 ) | ( ~n765 & n2562 ) ;
  assign n2564 = n766 & n2563 ;
  assign n2565 = ~n478 & n2564 ;
  assign n2566 = ( n2510 & ~n2516 ) | ( n2510 & n2565 ) | ( ~n2516 & n2565 ) ;
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n2568( .i (n2567), .o (n2568) );
  assign n2569 = n62 | n2536 ;
  assign n2570 = ~n1062 & n2536 ;
  assign n2571 = n2569 & ~n2570 ;
  buffer buf_n2572( .i (n2571), .o (n2572) );
  buffer buf_n2573( .i (n2572), .o (n2573) );
  buffer buf_n2574( .i (n2573), .o (n2574) );
  buffer buf_n2575( .i (n2574), .o (n2575) );
  buffer buf_n2576( .i (n2575), .o (n2576) );
  buffer buf_n2577( .i (n2576), .o (n2577) );
  buffer buf_n2578( .i (n2577), .o (n2578) );
  buffer buf_n2579( .i (n2578), .o (n2579) );
  buffer buf_n2580( .i (n2579), .o (n2580) );
  buffer buf_n2581( .i (n2580), .o (n2581) );
  buffer buf_n2582( .i (n2581), .o (n2582) );
  buffer buf_n2583( .i (n2582), .o (n2583) );
  assign n2584 = n2512 & n2583 ;
  assign n2585 = ( n476 & n765 ) | ( n476 & ~n2584 ) | ( n765 & ~n2584 ) ;
  assign n2586 = n766 & ~n2585 ;
  buffer buf_n2587( .i (n2586), .o (n2587) );
  buffer buf_n2588( .i (n2587), .o (n2588) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n144( .i (n143), .o (n144) );
  assign n2589 = ( n47 & n144 ) | ( n47 & ~n2587 ) | ( n144 & ~n2587 ) ;
  buffer buf_n2590( .i (n266), .o (n2590) );
  buffer buf_n2591( .i (n2590), .o (n2591) );
  assign n2592 = ~n590 & n2591 ;
  assign n2593 = n302 & n502 ;
  assign n2594 = n2591 | n2593 ;
  assign n2595 = ~n2592 & n2594 ;
  buffer buf_n2596( .i (n2595), .o (n2596) );
  assign n2597 = n169 | n2596 ;
  assign n2598 = ~n292 & n325 ;
  buffer buf_n2599( .i (n2598), .o (n2599) );
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  buffer buf_n2602( .i (n2601), .o (n2602) );
  buffer buf_n2603( .i (n2602), .o (n2603) );
  buffer buf_n2604( .i (n2603), .o (n2604) );
  buffer buf_n2605( .i (n2604), .o (n2605) );
  buffer buf_n2606( .i (n2605), .o (n2606) );
  buffer buf_n2607( .i (n2606), .o (n2607) );
  buffer buf_n2608( .i (n2607), .o (n2608) );
  buffer buf_n2609( .i (n2608), .o (n2609) );
  assign n2617 = n2133 & n2609 ;
  assign n2618 = ~n915 & n2617 ;
  buffer buf_n2619( .i (n168), .o (n2619) );
  assign n2620 = ~n2618 & n2619 ;
  assign n2621 = n2597 & ~n2620 ;
  buffer buf_n2622( .i (n2621), .o (n2622) );
  buffer buf_n2623( .i (n2622), .o (n2623) );
  assign n2624 = n358 | n391 ;
  buffer buf_n2625( .i (n2624), .o (n2625) );
  buffer buf_n2626( .i (n2625), .o (n2626) );
  buffer buf_n2627( .i (n2626), .o (n2627) );
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  buffer buf_n2631( .i (n2630), .o (n2631) );
  buffer buf_n2632( .i (n2631), .o (n2632) );
  buffer buf_n2633( .i (n2632), .o (n2633) );
  buffer buf_n2634( .i (n2633), .o (n2634) );
  buffer buf_n2635( .i (n2634), .o (n2635) );
  buffer buf_n2636( .i (n2635), .o (n2636) );
  buffer buf_n2637( .i (n2636), .o (n2637) );
  buffer buf_n2638( .i (n2637), .o (n2638) );
  buffer buf_n2347( .i (n2346), .o (n2347) );
  buffer buf_n2642( .i (n1581), .o (n2642) );
  assign n2643 = n399 & ~n2642 ;
  buffer buf_n2644( .i (n2643), .o (n2644) );
  assign n2648 = ( n2346 & n2393 ) | ( n2346 & ~n2644 ) | ( n2393 & ~n2644 ) ;
  assign n2649 = n2347 & ~n2648 ;
  buffer buf_n2650( .i (n2649), .o (n2650) );
  buffer buf_n2651( .i (n2650), .o (n2651) );
  buffer buf_n2652( .i (n2651), .o (n2652) );
  buffer buf_n2610( .i (n2609), .o (n2610) );
  buffer buf_n2611( .i (n2610), .o (n2611) );
  assign n2653 = ~n261 & n2536 ;
  buffer buf_n2654( .i (n2653), .o (n2654) );
  buffer buf_n2655( .i (n2654), .o (n2655) );
  buffer buf_n2656( .i (n2655), .o (n2656) );
  buffer buf_n2657( .i (n2656), .o (n2657) );
  buffer buf_n2658( .i (n2657), .o (n2658) );
  buffer buf_n2659( .i (n2658), .o (n2659) );
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2393), .o (n2661) );
  assign n2662 = n2660 & n2661 ;
  buffer buf_n2663( .i (n2662), .o (n2663) );
  assign n2665 = ( n2611 & n2650 ) | ( n2611 & n2663 ) | ( n2650 & n2663 ) ;
  assign n2666 = n2637 | n2665 ;
  assign n2667 = ( ~n2638 & n2652 ) | ( ~n2638 & n2666 ) | ( n2652 & n2666 ) ;
  assign n2668 = n73 & n1035 ;
  buffer buf_n2669( .i (n2668), .o (n2669) );
  buffer buf_n2670( .i (n473), .o (n2670) );
  assign n2671 = ( n2667 & ~n2669 ) | ( n2667 & n2670 ) | ( ~n2669 & n2670 ) ;
  assign n2672 = ( n2622 & ~n2669 ) | ( n2622 & n2670 ) | ( ~n2669 & n2670 ) ;
  assign n2673 = ( n2623 & n2671 ) | ( n2623 & ~n2672 ) | ( n2671 & ~n2672 ) ;
  buffer buf_n2674( .i (n2673), .o (n2674) );
  buffer buf_n2675( .i (n2674), .o (n2675) );
  buffer buf_n2676( .i (n108), .o (n2676) );
  assign n2677 = ( n443 & n2674 ) | ( n443 & ~n2676 ) | ( n2674 & ~n2676 ) ;
  buffer buf_n2612( .i (n2611), .o (n2612) );
  buffer buf_n2613( .i (n2612), .o (n2613) );
  assign n2678 = n373 & n2613 ;
  assign n2679 = ( n407 & n2670 ) | ( n407 & n2678 ) | ( n2670 & n2678 ) ;
  assign n2680 = ~n475 & n2679 ;
  assign n2681 = n637 | n1646 ;
  assign n2682 = n2099 & n2596 ;
  assign n2683 = ( n638 & ~n2681 ) | ( n638 & n2682 ) | ( ~n2681 & n2682 ) ;
  assign n2684 = n74 & n2683 ;
  buffer buf_n2685( .i (n2684), .o (n2685) );
  buffer buf_n2686( .i (n2685), .o (n2686) );
  buffer buf_n919( .i (n918), .o (n919) );
  assign n2687 = ~n105 & n171 ;
  assign n2688 = ~n919 & n2687 ;
  assign n2689 = n2685 | n2688 ;
  assign n2690 = ( n2680 & n2686 ) | ( n2680 & n2689 ) | ( n2686 & n2689 ) ;
  assign n2691 = ~n443 & n2690 ;
  assign n2692 = ( n2675 & ~n2677 ) | ( n2675 & n2691 ) | ( ~n2677 & n2691 ) ;
  assign n2693 = n144 & n2692 ;
  assign n2694 = ( n2588 & n2589 ) | ( n2588 & n2693 ) | ( n2589 & n2693 ) ;
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  assign n2695 = ( n34 & ~n501 ) | ( n34 & n2552 ) | ( ~n501 & n2552 ) ;
  assign n2696 = n502 & n2695 ;
  buffer buf_n2697( .i (n2696), .o (n2697) );
  buffer buf_n2698( .i (n2697), .o (n2698) );
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  assign n2700 = n366 & n1836 ;
  buffer buf_n2701( .i (n2178), .o (n2701) );
  assign n2702 = ( n400 & n2700 ) | ( n400 & n2701 ) | ( n2700 & n2701 ) ;
  buffer buf_n2703( .i (n2701), .o (n2703) );
  assign n2704 = n2702 & ~n2703 ;
  assign n2705 = ( ~n1222 & n2697 ) | ( ~n1222 & n2704 ) | ( n2697 & n2704 ) ;
  assign n2706 = n1017 | n2705 ;
  assign n2707 = ( ~n1018 & n2699 ) | ( ~n1018 & n2706 ) | ( n2699 & n2706 ) ;
  buffer buf_n2708( .i (n2707), .o (n2708) );
  buffer buf_n2709( .i (n2708), .o (n2709) );
  buffer buf_n2710( .i (n2072), .o (n2710) );
  assign n2711 = ( n2467 & n2708 ) | ( n2467 & ~n2710 ) | ( n2708 & ~n2710 ) ;
  assign n2712 = n262 | n297 ;
  buffer buf_n2713( .i (n2712), .o (n2713) );
  buffer buf_n2714( .i (n2713), .o (n2714) );
  buffer buf_n2715( .i (n2714), .o (n2715) );
  buffer buf_n2716( .i (n2715), .o (n2716) );
  buffer buf_n2717( .i (n2716), .o (n2717) );
  assign n2722 = n401 | n2717 ;
  buffer buf_n2723( .i (n2703), .o (n2723) );
  assign n2724 = ( ~n2202 & n2722 ) | ( ~n2202 & n2723 ) | ( n2722 & n2723 ) ;
  assign n2725 = n2204 | n2724 ;
  assign n2726 = n1018 | n2725 ;
  assign n2727 = n1225 | n2726 ;
  assign n2728 = n2467 | n2727 ;
  assign n2729 = ( ~n2709 & n2711 ) | ( ~n2709 & n2728 ) | ( n2711 & n2728 ) ;
  buffer buf_n2730( .i (n2729), .o (n2730) );
  buffer buf_n2731( .i (n2730), .o (n2731) );
  buffer buf_n2732( .i (n2731), .o (n2732) );
  buffer buf_n2540( .i (n2539), .o (n2540) );
  buffer buf_n2541( .i (n2540), .o (n2541) );
  buffer buf_n2542( .i (n2541), .o (n2542) );
  buffer buf_n2543( .i (n2542), .o (n2543) );
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  assign n2733 = ( n374 & n2489 ) | ( n374 & ~n2549 ) | ( n2489 & ~n2549 ) ;
  assign n2734 = n2550 & n2733 ;
  assign n2735 = ( n44 & ~n2730 ) | ( n44 & n2734 ) | ( ~n2730 & n2734 ) ;
  assign n2736 = n277 & ~n2735 ;
  assign n2737 = ( ~n278 & n2732 ) | ( ~n278 & n2736 ) | ( n2732 & n2736 ) ;
  assign n2738 = n32 & ~n464 ;
  assign n2739 = ( n1915 & ~n2573 ) | ( n1915 & n2738 ) | ( ~n2573 & n2738 ) ;
  assign n2740 = n2574 & n2739 ;
  buffer buf_n2741( .i (n2740), .o (n2741) );
  buffer buf_n2742( .i (n2741), .o (n2742) );
  assign n2743 = n154 & ~n221 ;
  buffer buf_n2744( .i (n2743), .o (n2744) );
  assign n2757 = n59 & ~n2744 ;
  assign n2758 = n989 & ~n2757 ;
  buffer buf_n2759( .i (n2530), .o (n2759) );
  assign n2760 = n2758 & n2759 ;
  buffer buf_n2761( .i (n2760), .o (n2761) );
  buffer buf_n2762( .i (n2761), .o (n2762) );
  buffer buf_n2763( .i (n1663), .o (n2763) );
  assign n2764 = ( n2293 & ~n2535 ) | ( n2293 & n2763 ) | ( ~n2535 & n2763 ) ;
  buffer buf_n2765( .i (n2764), .o (n2765) );
  assign n2769 = n2761 | n2765 ;
  assign n2770 = ( n64 & n2762 ) | ( n64 & n2769 ) | ( n2762 & n2769 ) ;
  buffer buf_n2771( .i (n2770), .o (n2771) );
  assign n2773 = n465 & n2771 ;
  assign n2774 = ~n2178 & n2773 ;
  buffer buf_n2775( .i (n2774), .o (n2775) );
  buffer buf_n2772( .i (n2771), .o (n2772) );
  assign n2779 = n464 & ~n1834 ;
  buffer buf_n2780( .i (n2035), .o (n2780) );
  buffer buf_n2781( .i (n2780), .o (n2781) );
  assign n2782 = ( n2771 & ~n2779 ) | ( n2771 & n2781 ) | ( ~n2779 & n2781 ) ;
  assign n2783 = n2772 & ~n2782 ;
  buffer buf_n2784( .i (n2783), .o (n2784) );
  assign n2785 = ( ~n2741 & n2775 ) | ( ~n2741 & n2784 ) | ( n2775 & n2784 ) ;
  assign n2786 = n401 & ~n2784 ;
  assign n2787 = ( n2742 & n2785 ) | ( n2742 & ~n2786 ) | ( n2785 & ~n2786 ) ;
  assign n2788 = n2204 & ~n2787 ;
  buffer buf_n2776( .i (n2775), .o (n2776) );
  buffer buf_n2789( .i (n335), .o (n2789) );
  buffer buf_n2790( .i (n2789), .o (n2790) );
  assign n2791 = n2776 & n2790 ;
  buffer buf_n2792( .i (n366), .o (n2792) );
  buffer buf_n2793( .i (n2792), .o (n2793) );
  buffer buf_n2794( .i (n2793), .o (n2794) );
  buffer buf_n2795( .i (n2794), .o (n2795) );
  assign n2796 = n2791 | n2795 ;
  assign n2797 = ~n2788 & n2796 ;
  buffer buf_n2798( .i (n270), .o (n2798) );
  buffer buf_n2799( .i (n2798), .o (n2799) );
  assign n2800 = n2797 & n2799 ;
  buffer buf_n2801( .i (n2800), .o (n2801) );
  buffer buf_n2802( .i (n2801), .o (n2802) );
  buffer buf_n2803( .i (n2781), .o (n2803) );
  assign n2804 = ( n889 & ~n2574 ) | ( n889 & n2803 ) | ( ~n2574 & n2803 ) ;
  assign n2805 = n2575 & n2804 ;
  assign n2806 = ~n233 & n2805 ;
  assign n2807 = n2386 & n2806 ;
  buffer buf_n2808( .i (n2807), .o (n2808) );
  buffer buf_n2809( .i (n2808), .o (n2809) );
  buffer buf_n2810( .i (n2809), .o (n2810) );
  buffer buf_n2777( .i (n2776), .o (n2777) );
  buffer buf_n2778( .i (n2777), .o (n2778) );
  assign n2811 = ( n2778 & ~n2798 ) | ( n2778 & n2808 ) | ( ~n2798 & n2808 ) ;
  assign n2812 = n307 & ~n2811 ;
  assign n2813 = ( n2153 & n2810 ) | ( n2153 & ~n2812 ) | ( n2810 & ~n2812 ) ;
  assign n2814 = n2801 | n2813 ;
  assign n2815 = ( n510 & n2802 ) | ( n510 & n2814 ) | ( n2802 & n2814 ) ;
  assign n2816 = n141 & n2815 ;
  buffer buf_n2817( .i (n2816), .o (n2817) );
  buffer buf_n2818( .i (n2817), .o (n2818) );
  buffer buf_n2819( .i (n477), .o (n2819) );
  assign n2820 = ~n2817 & n2819 ;
  assign n2821 = ( n2737 & ~n2818 ) | ( n2737 & n2820 ) | ( ~n2818 & n2820 ) ;
  buffer buf_n2822( .i (n2821), .o (n2822) );
  assign n2823 = ( n2567 & ~n2694 ) | ( n2567 & n2822 ) | ( ~n2694 & n2822 ) ;
  assign n2824 = ~n246 & n2822 ;
  assign n2825 = ( ~n2568 & n2823 ) | ( ~n2568 & n2824 ) | ( n2823 & n2824 ) ;
  assign n2826 = n410 | n477 ;
  assign n2827 = n444 | n2826 ;
  buffer buf_n2828( .i (n2827), .o (n2828) );
  assign n2829 = n297 | n574 ;
  buffer buf_n2830( .i (n2829), .o (n2830) );
  buffer buf_n2831( .i (n2830), .o (n2831) );
  buffer buf_n2832( .i (n2831), .o (n2832) );
  buffer buf_n2833( .i (n2832), .o (n2833) );
  buffer buf_n2834( .i (n2833), .o (n2834) );
  buffer buf_n2835( .i (n2834), .o (n2835) );
  buffer buf_n2836( .i (n2835), .o (n2836) );
  buffer buf_n2837( .i (n2836), .o (n2837) );
  buffer buf_n2838( .i (n2837), .o (n2838) );
  buffer buf_n2839( .i (n2838), .o (n2839) );
  buffer buf_n2840( .i (n2839), .o (n2840) );
  buffer buf_n2841( .i (n2840), .o (n2841) );
  buffer buf_n2842( .i (n2841), .o (n2842) );
  buffer buf_n2843( .i (n2842), .o (n2843) );
  buffer buf_n2844( .i (n2843), .o (n2844) );
  buffer buf_n2845( .i (n2844), .o (n2845) );
  buffer buf_n2846( .i (n2845), .o (n2846) );
  assign n2847 = n2828 | n2846 ;
  assign n2848 = ~n323 & n519 ;
  assign n2849 = n1345 & n2848 ;
  buffer buf_n2850( .i (n2849), .o (n2850) );
  buffer buf_n2851( .i (n2850), .o (n2851) );
  buffer buf_n2852( .i (n2851), .o (n2852) );
  assign n2853 = ( n221 & n324 ) | ( n221 & ~n422 ) | ( n324 & ~n422 ) ;
  assign n2854 = ( n221 & n324 ) | ( n221 & ~n456 ) | ( n324 & ~n456 ) ;
  assign n2855 = ~n2853 & n2854 ;
  assign n2856 = ( ~n26 & n2850 ) | ( ~n26 & n2855 ) | ( n2850 & n2855 ) ;
  assign n2857 = n1663 & ~n2856 ;
  assign n2858 = ( n2763 & n2852 ) | ( n2763 & ~n2857 ) | ( n2852 & ~n2857 ) ;
  buffer buf_n2859( .i (n2858), .o (n2859) );
  buffer buf_n2860( .i (n2859), .o (n2860) );
  buffer buf_n2861( .i (n258), .o (n2861) );
  buffer buf_n2862( .i (n358), .o (n2862) );
  assign n2863 = n2861 & ~n2862 ;
  buffer buf_n2864( .i (n2863), .o (n2864) );
  buffer buf_n2865( .i (n2864), .o (n2865) );
  buffer buf_n2868( .i (n296), .o (n2868) );
  assign n2869 = ( ~n2859 & n2865 ) | ( ~n2859 & n2868 ) | ( n2865 & n2868 ) ;
  assign n2870 = n2860 & n2869 ;
  buffer buf_n2871( .i (n2870), .o (n2871) );
  buffer buf_n2872( .i (n2871), .o (n2872) );
  buffer buf_n2873( .i (n2872), .o (n2873) );
  assign n2874 = n1353 & ~n2713 ;
  assign n2875 = ( n529 & n2871 ) | ( n529 & n2874 ) | ( n2871 & n2874 ) ;
  assign n2876 = n2025 & ~n2875 ;
  assign n2877 = ( n2026 & n2873 ) | ( n2026 & ~n2876 ) | ( n2873 & ~n2876 ) ;
  assign n2878 = n69 & n2877 ;
  buffer buf_n2879( .i (n2878), .o (n2879) );
  buffer buf_n2880( .i (n2879), .o (n2880) );
  buffer buf_n2881( .i (n467), .o (n2881) );
  assign n2882 = ( ~n1570 & n2346 ) | ( ~n1570 & n2881 ) | ( n2346 & n2881 ) ;
  assign n2883 = n2347 & ~n2882 ;
  assign n2884 = n2879 | n2883 ;
  assign n2885 = ( ~n2255 & n2880 ) | ( ~n2255 & n2884 ) | ( n2880 & n2884 ) ;
  assign n2886 = n170 | n2885 ;
  buffer buf_n2887( .i (n327), .o (n2887) );
  assign n2888 = n260 & ~n2887 ;
  buffer buf_n2889( .i (n2888), .o (n2889) );
  buffer buf_n2890( .i (n326), .o (n2890) );
  assign n2891 = n2861 | n2890 ;
  buffer buf_n2892( .i (n2891), .o (n2892) );
  buffer buf_n2893( .i (n2892), .o (n2893) );
  assign n2894 = ( ~n262 & n2889 ) | ( ~n262 & n2893 ) | ( n2889 & n2893 ) ;
  buffer buf_n2895( .i (n2894), .o (n2895) );
  buffer buf_n2896( .i (n2895), .o (n2896) );
  buffer buf_n2897( .i (n2896), .o (n2897) );
  buffer buf_n2898( .i (n2897), .o (n2898) );
  buffer buf_n2903( .i (n364), .o (n2903) );
  assign n2904 = n465 & ~n2903 ;
  assign n2905 = ( n2803 & n2897 ) | ( n2803 & ~n2904 ) | ( n2897 & ~n2904 ) ;
  assign n2906 = n2898 & ~n2905 ;
  assign n2907 = n303 & n2906 ;
  buffer buf_n2908( .i (n233), .o (n2908) );
  assign n2909 = ( n2661 & n2907 ) | ( n2661 & n2908 ) | ( n2907 & n2908 ) ;
  assign n2910 = ~n2396 & n2909 ;
  assign n2911 = ~n72 & n2910 ;
  buffer buf_n2912( .i (n2619), .o (n2912) );
  assign n2913 = ~n2911 & n2912 ;
  assign n2914 = n2886 & ~n2913 ;
  assign n2915 = n106 & ~n2914 ;
  buffer buf_n2899( .i (n2898), .o (n2899) );
  buffer buf_n2900( .i (n2899), .o (n2900) );
  assign n2916 = n467 | n2792 ;
  assign n2917 = ( n2703 & n2899 ) | ( n2703 & n2916 ) | ( n2899 & n2916 ) ;
  assign n2918 = n2900 & ~n2917 ;
  assign n2919 = n305 & n2918 ;
  assign n2920 = ( n2255 & n2262 ) | ( n2255 & n2919 ) | ( n2262 & n2919 ) ;
  assign n2921 = ~n203 & n2920 ;
  assign n2922 = n171 & n2921 ;
  buffer buf_n2923( .i (n105), .o (n2923) );
  assign n2924 = n2922 | n2923 ;
  assign n2925 = ~n2915 & n2924 ;
  assign n2926 = n141 & ~n2925 ;
  assign n2927 = n254 & n289 ;
  buffer buf_n2928( .i (n2927), .o (n2928) );
  buffer buf_n2929( .i (n2928), .o (n2929) );
  buffer buf_n2930( .i (n2929), .o (n2930) );
  buffer buf_n2931( .i (n2930), .o (n2931) );
  buffer buf_n2932( .i (n2931), .o (n2932) );
  buffer buf_n2933( .i (n2932), .o (n2933) );
  buffer buf_n2934( .i (n2933), .o (n2934) );
  buffer buf_n2935( .i (n2934), .o (n2935) );
  buffer buf_n2936( .i (n2935), .o (n2936) );
  buffer buf_n2937( .i (n2936), .o (n2937) );
  buffer buf_n2938( .i (n2937), .o (n2938) );
  buffer buf_n2939( .i (n2938), .o (n2939) );
  assign n2946 = ~n1633 & n2939 ;
  buffer buf_n2947( .i (n2946), .o (n2947) );
  buffer buf_n2948( .i (n2947), .o (n2948) );
  buffer buf_n2949( .i (n2948), .o (n2949) );
  assign n2950 = ( n1017 & n1865 ) | ( n1017 & n2948 ) | ( n1865 & n2948 ) ;
  buffer buf_n2718( .i (n2717), .o (n2718) );
  assign n2951 = n161 & n228 ;
  buffer buf_n2952( .i (n2951), .o (n2952) );
  buffer buf_n2953( .i (n2952), .o (n2953) );
  buffer buf_n2954( .i (n2953), .o (n2954) );
  buffer buf_n2955( .i (n2954), .o (n2955) );
  buffer buf_n2960( .i (n2392), .o (n2960) );
  assign n2961 = ( n2717 & n2955 ) | ( n2717 & n2960 ) | ( n2955 & n2960 ) ;
  assign n2962 = ~n2718 & n2961 ;
  buffer buf_n2963( .i (n469), .o (n2963) );
  assign n2964 = n2962 & ~n2963 ;
  assign n2965 = ( n2949 & ~n2950 ) | ( n2949 & n2964 ) | ( ~n2950 & n2964 ) ;
  assign n2966 = n340 & n2965 ;
  buffer buf_n2967( .i (n2079), .o (n2967) );
  buffer buf_n2968( .i (n2967), .o (n2968) );
  buffer buf_n2969( .i (n2478), .o (n2969) );
  assign n2970 = ( n2966 & n2968 ) | ( n2966 & n2969 ) | ( n2968 & n2969 ) ;
  assign n2971 = ~n2237 & n2970 ;
  assign n2972 = ~n107 & n2971 ;
  assign n2973 = n141 | n2972 ;
  assign n2974 = ~n2926 & n2973 ;
  assign n2975 = n411 & n2974 ;
  buffer buf_n2976( .i (n2975), .o (n2976) );
  buffer buf_n2977( .i (n2976), .o (n2977) );
  buffer buf_n2978( .i (n235), .o (n2978) );
  assign n2979 = n1224 | n2978 ;
  buffer buf_n2980( .i (n2979), .o (n2980) );
  buffer buf_n2981( .i (n2980), .o (n2981) );
  buffer buf_n2982( .i (n2981), .o (n2982) );
  buffer buf_n2983( .i (n2982), .o (n2983) );
  buffer buf_n2984( .i (n2983), .o (n2984) );
  buffer buf_n2985( .i (n2984), .o (n2985) );
  buffer buf_n2986( .i (n277), .o (n2986) );
  assign n2987 = ( ~n209 & n2985 ) | ( ~n209 & n2986 ) | ( n2985 & n2986 ) ;
  assign n2988 = n210 | n2987 ;
  assign n2989 = ~n2976 & n2988 ;
  assign n2990 = ( n2847 & ~n2977 ) | ( n2847 & n2989 ) | ( ~n2977 & n2989 ) ;
  buffer buf_n2991( .i (n2990), .o (n2991) );
  buffer buf_n2413( .i (n2412), .o (n2413) );
  buffer buf_n2414( .i (n2413), .o (n2414) );
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n2416( .i (n2415), .o (n2416) );
  buffer buf_n2417( .i (n2416), .o (n2417) );
  buffer buf_n2418( .i (n2417), .o (n2418) );
  assign n2992 = n279 | n2418 ;
  assign n2993 = n2828 | n2992 ;
  buffer buf_n2664( .i (n2663), .o (n2664) );
  assign n2994 = ~n2723 & n2794 ;
  assign n2995 = ~n2963 & n2994 ;
  buffer buf_n2996( .i (n2995), .o (n2996) );
  assign n2998 = n2664 & n2996 ;
  assign n2999 = ( n1226 & n2613 ) | ( n1226 & n2998 ) | ( n2613 & n2998 ) ;
  assign n3000 = ~n1227 & n2999 ;
  buffer buf_n3001( .i (n3000), .o (n3001) );
  buffer buf_n3002( .i (n3001), .o (n3002) );
  assign n3003 = ( n28 & ~n2124 ) | ( n28 & n2887 ) | ( ~n2124 & n2887 ) ;
  buffer buf_n3004( .i (n2535), .o (n3004) );
  buffer buf_n3005( .i (n2124), .o (n3005) );
  assign n3006 = ( n3003 & n3004 ) | ( n3003 & ~n3005 ) | ( n3004 & ~n3005 ) ;
  buffer buf_n3007( .i (n3006), .o (n3007) );
  buffer buf_n3010( .i (n3005), .o (n3010) );
  buffer buf_n3011( .i (n3010), .o (n3011) );
  assign n3012 = n3007 & n3011 ;
  buffer buf_n3013( .i (n3012), .o (n3013) );
  buffer buf_n3014( .i (n3013), .o (n3014) );
  buffer buf_n3008( .i (n3007), .o (n3008) );
  buffer buf_n3009( .i (n3008), .o (n3009) );
  assign n3015 = n3009 & ~n3013 ;
  buffer buf_n3016( .i (n2903), .o (n3016) );
  assign n3017 = ( ~n3014 & n3015 ) | ( ~n3014 & n3016 ) | ( n3015 & n3016 ) ;
  buffer buf_n3018( .i (n3017), .o (n3018) );
  buffer buf_n3019( .i (n3018), .o (n3019) );
  buffer buf_n3020( .i (n466), .o (n3020) );
  assign n3021 = n302 & ~n3020 ;
  assign n3022 = ( n2703 & n3018 ) | ( n2703 & n3021 ) | ( n3018 & n3021 ) ;
  assign n3023 = ~n3019 & n3022 ;
  buffer buf_n3024( .i (n3023), .o (n3024) );
  buffer buf_n3025( .i (n3024), .o (n3025) );
  buffer buf_n3026( .i (n101), .o (n3026) );
  buffer buf_n3027( .i (n2142), .o (n3027) );
  assign n3028 = n3026 & n3027 ;
  assign n3029 = ( n2255 & ~n3024 ) | ( n2255 & n3028 ) | ( ~n3024 & n3028 ) ;
  assign n3030 = n3025 & n3029 ;
  buffer buf_n3031( .i (n3030), .o (n3031) );
  buffer buf_n3032( .i (n3031), .o (n3032) );
  buffer buf_n3033( .i (n74), .o (n3033) );
  assign n3034 = ( n139 & ~n3031 ) | ( n139 & n3033 ) | ( ~n3031 & n3033 ) ;
  buffer buf_n2348( .i (n2347), .o (n2348) );
  buffer buf_n2349( .i (n2348), .o (n2349) );
  assign n3035 = ( ~n636 & n2348 ) | ( ~n636 & n2963 ) | ( n2348 & n2963 ) ;
  assign n3036 = n2349 & ~n3035 ;
  assign n3037 = ( n104 & ~n2478 ) | ( n104 & n3036 ) | ( ~n2478 & n3036 ) ;
  assign n3038 = n464 & n2604 ;
  assign n3039 = n2903 & n3038 ;
  assign n3040 = ~n57 & n154 ;
  buffer buf_n3041( .i (n3040), .o (n3041) );
  buffer buf_n3042( .i (n3041), .o (n3042) );
  buffer buf_n3043( .i (n3042), .o (n3043) );
  buffer buf_n3044( .i (n3043), .o (n3044) );
  buffer buf_n3045( .i (n3044), .o (n3045) );
  buffer buf_n3046( .i (n3045), .o (n3046) );
  buffer buf_n3047( .i (n3046), .o (n3047) );
  buffer buf_n3048( .i (n3047), .o (n3048) );
  buffer buf_n3049( .i (n3048), .o (n3049) );
  assign n3053 = n3039 & n3049 ;
  assign n3054 = ~n912 & n3053 ;
  buffer buf_n3055( .i (n3054), .o (n3055) );
  buffer buf_n3056( .i (n3055), .o (n3056) );
  buffer buf_n3057( .i (n3056), .o (n3057) );
  buffer buf_n3058( .i (n456), .o (n3058) );
  assign n3059 = ~n325 & n3058 ;
  assign n3060 = ~n358 & n3059 ;
  buffer buf_n3061( .i (n3060), .o (n3061) );
  buffer buf_n3062( .i (n3061), .o (n3062) );
  buffer buf_n3063( .i (n3062), .o (n3063) );
  buffer buf_n3064( .i (n3063), .o (n3064) );
  buffer buf_n3065( .i (n3064), .o (n3065) );
  buffer buf_n3066( .i (n3065), .o (n3066) );
  assign n3067 = n630 & ~n1605 ;
  assign n3068 = n3066 & n3067 ;
  buffer buf_n3069( .i (n3068), .o (n3069) );
  assign n3070 = ( n1278 & n3020 ) | ( n1278 & ~n3069 ) | ( n3020 & ~n3069 ) ;
  buffer buf_n3071( .i (n2862), .o (n3071) );
  assign n3072 = ( n2535 & n2887 ) | ( n2535 & ~n3071 ) | ( n2887 & ~n3071 ) ;
  buffer buf_n3073( .i (n2763), .o (n3073) );
  assign n3074 = ( ~n3005 & n3072 ) | ( ~n3005 & n3073 ) | ( n3072 & n3073 ) ;
  buffer buf_n3075( .i (n3074), .o (n3075) );
  assign n3078 = n3011 & n3075 ;
  buffer buf_n3079( .i (n3078), .o (n3079) );
  buffer buf_n3080( .i (n3079), .o (n3080) );
  buffer buf_n3076( .i (n3075), .o (n3076) );
  buffer buf_n3077( .i (n3076), .o (n3077) );
  assign n3081 = n3077 & ~n3079 ;
  assign n3082 = ( n3016 & ~n3080 ) | ( n3016 & n3081 ) | ( ~n3080 & n3081 ) ;
  assign n3083 = ~n3069 & n3082 ;
  buffer buf_n3084( .i (n1278), .o (n3084) );
  assign n3085 = ( n3070 & n3083 ) | ( n3070 & ~n3084 ) | ( n3083 & ~n3084 ) ;
  assign n3086 = ( n2142 & n3055 ) | ( n2142 & ~n3085 ) | ( n3055 & ~n3085 ) ;
  assign n3087 = n305 & ~n3086 ;
  assign n3088 = ( n2410 & n3057 ) | ( n2410 & ~n3087 ) | ( n3057 & ~n3087 ) ;
  buffer buf_n3089( .i (n1646), .o (n3089) );
  buffer buf_n3090( .i (n2723), .o (n3090) );
  buffer buf_n3091( .i (n3090), .o (n3091) );
  buffer buf_n3092( .i (n3091), .o (n3092) );
  assign n3093 = ( ~n3088 & n3089 ) | ( ~n3088 & n3092 ) | ( n3089 & n3092 ) ;
  assign n3094 = n3037 & ~n3093 ;
  assign n3095 = n139 & n3094 ;
  assign n3096 = ( n3032 & n3034 ) | ( n3032 & n3095 ) | ( n3034 & n3095 ) ;
  buffer buf_n2745( .i (n2744), .o (n2745) );
  buffer buf_n2746( .i (n2745), .o (n2746) );
  buffer buf_n2747( .i (n2746), .o (n2747) );
  buffer buf_n2748( .i (n2747), .o (n2748) );
  buffer buf_n2749( .i (n2748), .o (n2749) );
  buffer buf_n2750( .i (n2749), .o (n2750) );
  buffer buf_n2751( .i (n2750), .o (n2751) );
  buffer buf_n2752( .i (n2751), .o (n2752) );
  buffer buf_n2753( .i (n2752), .o (n2753) );
  buffer buf_n2754( .i (n2753), .o (n2754) );
  buffer buf_n2755( .i (n2754), .o (n2755) );
  buffer buf_n2756( .i (n2755), .o (n2756) );
  assign n3097 = ( ~n1223 & n2396 ) | ( ~n1223 & n2756 ) | ( n2396 & n2756 ) ;
  buffer buf_n3098( .i (n2396), .o (n3098) );
  assign n3099 = n3097 & ~n3098 ;
  buffer buf_n3100( .i (n3099), .o (n3100) );
  buffer buf_n3101( .i (n3100), .o (n3101) );
  buffer buf_n2997( .i (n2996), .o (n2997) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  assign n3102 = n1842 & n2799 ;
  assign n3103 = ( n2997 & ~n3100 ) | ( n2997 & n3102 ) | ( ~n3100 & n3102 ) ;
  assign n3104 = n3101 & n3103 ;
  buffer buf_n3105( .i (n3104), .o (n3105) );
  assign n3106 = ( ~n3001 & n3096 ) | ( ~n3001 & n3105 ) | ( n3096 & n3105 ) ;
  assign n3107 = n241 | n3105 ;
  assign n3108 = ( n3002 & n3106 ) | ( n3002 & n3107 ) | ( n3106 & n3107 ) ;
  assign n3109 = n411 & n3108 ;
  buffer buf_n3110( .i (n3109), .o (n3110) );
  buffer buf_n3111( .i (n3110), .o (n3111) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  assign n3112 = n208 | n1230 ;
  assign n3113 = ( ~n176 & n243 ) | ( ~n176 & n3112 ) | ( n243 & n3112 ) ;
  assign n3114 = n177 | n3113 ;
  assign n3115 = ~n3110 & n3114 ;
  assign n3116 = ( n2993 & ~n3111 ) | ( n2993 & n3115 ) | ( ~n3111 & n3115 ) ;
  buffer buf_n3117( .i (n3116), .o (n3117) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n3118( .i (n299), .o (n3118) );
  assign n3119 = n2024 & n3118 ;
  buffer buf_n3120( .i (n3119), .o (n3120) );
  buffer buf_n3121( .i (n3120), .o (n3121) );
  buffer buf_n3122( .i (n3121), .o (n3122) );
  buffer buf_n3123( .i (n3122), .o (n3123) );
  buffer buf_n3124( .i (n3123), .o (n3124) );
  buffer buf_n3125( .i (n3124), .o (n3125) );
  buffer buf_n3126( .i (n3125), .o (n3126) );
  buffer buf_n3127( .i (n2661), .o (n3127) );
  assign n3128 = n3027 & ~n3127 ;
  assign n3129 = ~n2978 & n3128 ;
  assign n3130 = ( n3092 & n3125 ) | ( n3092 & ~n3129 ) | ( n3125 & ~n3129 ) ;
  buffer buf_n2956( .i (n2955), .o (n2956) );
  buffer buf_n2957( .i (n2956), .o (n2957) );
  assign n3131 = ( ~n2348 & n2957 ) | ( ~n2348 & n3127 ) | ( n2957 & n3127 ) ;
  assign n3132 = n2349 & n3131 ;
  assign n3133 = ~n3092 & n3132 ;
  assign n3134 = ( n3126 & ~n3130 ) | ( n3126 & n3133 ) | ( ~n3130 & n3133 ) ;
  assign n3135 = ( ~n2670 & n2923 ) | ( ~n2670 & n3134 ) | ( n2923 & n3134 ) ;
  buffer buf_n3136( .i (n2210), .o (n3136) );
  assign n3137 = ~n1015 & n3136 ;
  assign n3138 = ( n70 & n2386 ) | ( n70 & n3137 ) | ( n2386 & n3137 ) ;
  assign n3139 = ~n38 & n3138 ;
  buffer buf_n3140( .i (n3139), .o (n3140) );
  buffer buf_n3141( .i (n3140), .o (n3141) );
  assign n3142 = ~n338 & n3090 ;
  assign n3143 = n2079 & n3142 ;
  buffer buf_n2719( .i (n2718), .o (n2719) );
  buffer buf_n2720( .i (n2719), .o (n2720) );
  assign n3144 = ~n2720 & n2978 ;
  assign n3145 = ( ~n3140 & n3143 ) | ( ~n3140 & n3144 ) | ( n3143 & n3144 ) ;
  assign n3146 = n3141 & n3145 ;
  buffer buf_n3147( .i (n473), .o (n3147) );
  assign n3148 = n3146 & ~n3147 ;
  assign n3149 = ( ~n107 & n3135 ) | ( ~n107 & n3148 ) | ( n3135 & n3148 ) ;
  buffer buf_n3150( .i (n140), .o (n3150) );
  assign n3151 = n3149 & ~n3150 ;
  buffer buf_n3152( .i (n62), .o (n3152) );
  buffer buf_n3153( .i (n3152), .o (n3153) );
  buffer buf_n3154( .i (n3153), .o (n3154) );
  buffer buf_n3155( .i (n463), .o (n3155) );
  assign n3156 = n3154 & ~n3155 ;
  assign n3157 = n364 | n2780 ;
  assign n3158 = ( n2425 & ~n3156 ) | ( n2425 & n3157 ) | ( ~n3156 & n3157 ) ;
  buffer buf_n3159( .i (n3118), .o (n3159) );
  assign n3160 = n3158 | n3159 ;
  assign n3161 = ( n335 & ~n1633 ) | ( n335 & n3160 ) | ( ~n1633 & n3160 ) ;
  buffer buf_n3162( .i (n231), .o (n3162) );
  buffer buf_n3163( .i (n3162), .o (n3163) );
  assign n3164 = n3161 | n3163 ;
  buffer buf_n3165( .i (n3164), .o (n3165) );
  buffer buf_n3166( .i (n3165), .o (n3166) );
  buffer buf_n3167( .i (n183), .o (n3167) );
  buffer buf_n3168( .i (n3167), .o (n3168) );
  assign n3169 = n322 & n3168 ;
  buffer buf_n3170( .i (n3169), .o (n3170) );
  assign n3176 = ( n356 & n456 ) | ( n356 & n3170 ) | ( n456 & n3170 ) ;
  assign n3177 = ~n3058 & n3176 ;
  buffer buf_n3178( .i (n3177), .o (n3178) );
  buffer buf_n3179( .i (n3178), .o (n3179) );
  buffer buf_n3180( .i (n3179), .o (n3180) );
  buffer buf_n3181( .i (n59), .o (n3181) );
  buffer buf_n3182( .i (n2290), .o (n3182) );
  assign n3183 = ( ~n3178 & n3181 ) | ( ~n3178 & n3182 ) | ( n3181 & n3182 ) ;
  assign n3184 = n3061 & n3183 ;
  assign n3185 = ( n3062 & n3180 ) | ( n3062 & ~n3184 ) | ( n3180 & ~n3184 ) ;
  buffer buf_n3186( .i (n3185), .o (n3186) );
  buffer buf_n3187( .i (n3186), .o (n3187) );
  buffer buf_n3188( .i (n1295), .o (n3188) );
  buffer buf_n3189( .i (n428), .o (n3189) );
  assign n3190 = ( n3186 & ~n3188 ) | ( n3186 & n3189 ) | ( ~n3188 & n3189 ) ;
  assign n3191 = n1007 | n3071 ;
  assign n3192 = ( ~n329 & n461 ) | ( ~n329 & n3191 ) | ( n461 & n3191 ) ;
  assign n3193 = n330 | n3192 ;
  assign n3194 = n3189 | n3193 ;
  assign n3195 = ( ~n3187 & n3190 ) | ( ~n3187 & n3194 ) | ( n3190 & n3194 ) ;
  buffer buf_n3196( .i (n3195), .o (n3196) );
  buffer buf_n3197( .i (n3196), .o (n3197) );
  buffer buf_n3198( .i (n229), .o (n3198) );
  buffer buf_n3199( .i (n3198), .o (n3199) );
  assign n3200 = ( n3159 & n3196 ) | ( n3159 & n3199 ) | ( n3196 & n3199 ) ;
  buffer buf_n3201( .i (n218), .o (n3201) );
  assign n3202 = n322 & n3201 ;
  buffer buf_n3203( .i (n3202), .o (n3203) );
  assign n3218 = n356 & n3203 ;
  assign n3219 = ( ~n521 & n1822 ) | ( ~n521 & n3218 ) | ( n1822 & n3218 ) ;
  assign n3220 = n522 & n3219 ;
  buffer buf_n3221( .i (n3220), .o (n3221) );
  buffer buf_n3222( .i (n3221), .o (n3222) );
  buffer buf_n3223( .i (n3222), .o (n3223) );
  assign n3224 = n222 & n2016 ;
  assign n3225 = n22 & ~n152 ;
  buffer buf_n3226( .i (n3225), .o (n3226) );
  assign n3229 = n24 & ~n3226 ;
  buffer buf_n3230( .i (n3229), .o (n3230) );
  assign n3231 = n3224 & n3230 ;
  buffer buf_n3227( .i (n3226), .o (n3227) );
  buffer buf_n3228( .i (n3227), .o (n3228) );
  buffer buf_n3232( .i (n321), .o (n3232) );
  assign n3233 = ( n354 & n3201 ) | ( n354 & n3232 ) | ( n3201 & n3232 ) ;
  buffer buf_n3234( .i (n3233), .o (n3234) );
  buffer buf_n3235( .i (n3234), .o (n3235) );
  buffer buf_n3236( .i (n220), .o (n3236) );
  assign n3237 = ~n3234 & n3236 ;
  assign n3238 = ( n325 & ~n3235 ) | ( n325 & n3237 ) | ( ~n3235 & n3237 ) ;
  assign n3239 = ( ~n3228 & n3230 ) | ( ~n3228 & n3238 ) | ( n3230 & n3238 ) ;
  assign n3240 = ( ~n2534 & n3231 ) | ( ~n2534 & n3239 ) | ( n3231 & n3239 ) ;
  buffer buf_n3241( .i (n459), .o (n3241) );
  assign n3242 = ( n3221 & n3240 ) | ( n3221 & ~n3241 ) | ( n3240 & ~n3241 ) ;
  assign n3243 = n427 & ~n3242 ;
  assign n3244 = ( n428 & n3223 ) | ( n428 & ~n3243 ) | ( n3223 & ~n3243 ) ;
  buffer buf_n3245( .i (n3244), .o (n3245) );
  buffer buf_n3246( .i (n3245), .o (n3246) );
  assign n3247 = ( n2195 & n3154 ) | ( n2195 & ~n3245 ) | ( n3154 & ~n3245 ) ;
  assign n3248 = n525 & n1350 ;
  assign n3249 = ( ~n574 & n1295 ) | ( ~n574 & n3248 ) | ( n1295 & n3248 ) ;
  assign n3250 = ~n3188 & n3249 ;
  assign n3251 = n3154 & n3250 ;
  assign n3252 = ( n3246 & n3247 ) | ( n3246 & n3251 ) | ( n3247 & n3251 ) ;
  assign n3253 = n3159 & n3252 ;
  assign n3254 = ( ~n3197 & n3200 ) | ( ~n3197 & n3253 ) | ( n3200 & n3253 ) ;
  buffer buf_n3255( .i (n3254), .o (n3255) );
  buffer buf_n3256( .i (n3255), .o (n3256) );
  buffer buf_n3257( .i (n3256), .o (n3257) );
  assign n3258 = ( n1415 & n2661 ) | ( n1415 & ~n3255 ) | ( n2661 & ~n3255 ) ;
  assign n3259 = ~n3165 & n3258 ;
  assign n3260 = ( n3166 & ~n3257 ) | ( n3166 & n3259 ) | ( ~n3257 & n3259 ) ;
  buffer buf_n3261( .i (n3260), .o (n3261) );
  buffer buf_n3262( .i (n3261), .o (n3262) );
  assign n3263 = ( n105 & n2710 ) | ( n105 & n3261 ) | ( n2710 & n3261 ) ;
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  assign n3264 = ( n1098 & n2903 ) | ( n1098 & n3118 ) | ( n2903 & n3118 ) ;
  assign n3265 = ( n299 & ~n1097 ) | ( n299 & n3154 ) | ( ~n1097 & n3154 ) ;
  buffer buf_n3266( .i (n364), .o (n3266) );
  assign n3267 = ( n1581 & n3265 ) | ( n1581 & n3266 ) | ( n3265 & n3266 ) ;
  assign n3268 = ~n3264 & n3267 ;
  assign n3269 = n3020 & ~n3268 ;
  buffer buf_n3270( .i (n2534), .o (n3270) );
  assign n3271 = n295 | n3270 ;
  buffer buf_n3272( .i (n3271), .o (n3272) );
  buffer buf_n3273( .i (n3272), .o (n3273) );
  buffer buf_n3274( .i (n3273), .o (n3274) );
  buffer buf_n3275( .i (n3274), .o (n3275) );
  buffer buf_n3276( .i (n3275), .o (n3276) );
  assign n3277 = n3016 & ~n3276 ;
  assign n3278 = n3020 | n3277 ;
  assign n3279 = ~n3269 & n3278 ;
  buffer buf_n3280( .i (n3279), .o (n3280) );
  buffer buf_n3281( .i (n3280), .o (n3281) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  assign n3282 = ( ~n1792 & n3090 ) | ( ~n1792 & n3280 ) | ( n3090 & n3280 ) ;
  assign n3283 = n3281 & ~n3282 ;
  assign n3284 = n1361 & n3283 ;
  buffer buf_n3285( .i (n3089), .o (n3285) );
  assign n3286 = n3284 & n3285 ;
  assign n3287 = ( ~n3262 & n3263 ) | ( ~n3262 & n3286 ) | ( n3263 & n3286 ) ;
  assign n3288 = n256 & n324 ;
  buffer buf_n3289( .i (n3288), .o (n3289) );
  buffer buf_n3290( .i (n3289), .o (n3290) );
  buffer buf_n3291( .i (n3290), .o (n3291) );
  buffer buf_n3292( .i (n3291), .o (n3292) );
  buffer buf_n3293( .i (n3292), .o (n3293) );
  buffer buf_n3294( .i (n3293), .o (n3294) );
  buffer buf_n3295( .i (n3294), .o (n3295) );
  buffer buf_n3296( .i (n3295), .o (n3296) );
  buffer buf_n3297( .i (n3296), .o (n3297) );
  buffer buf_n3298( .i (n3297), .o (n3298) );
  buffer buf_n3299( .i (n3159), .o (n3299) );
  assign n3300 = ( n2792 & ~n3298 ) | ( n2792 & n3299 ) | ( ~n3298 & n3299 ) ;
  buffer buf_n3301( .i (n3118), .o (n3301) );
  assign n3302 = ( ~n266 & n3297 ) | ( ~n266 & n3301 ) | ( n3297 & n3301 ) ;
  assign n3303 = ( ~n335 & n2792 ) | ( ~n335 & n3302 ) | ( n2792 & n3302 ) ;
  assign n3304 = n3300 & ~n3303 ;
  buffer buf_n3305( .i (n3304), .o (n3305) );
  buffer buf_n3306( .i (n3305), .o (n3306) );
  assign n3307 = ( ~n1572 & n2963 ) | ( ~n1572 & n3305 ) | ( n2963 & n3305 ) ;
  assign n3308 = n3306 & ~n3307 ;
  assign n3309 = ~n203 & n3308 ;
  buffer buf_n3310( .i (n2912), .o (n3310) );
  assign n3311 = ( n3285 & n3309 ) | ( n3285 & n3310 ) | ( n3309 & n3310 ) ;
  assign n3312 = ~n2923 & n3311 ;
  assign n3313 = n3287 | n3312 ;
  assign n3314 = n3150 & n3313 ;
  assign n3315 = n3151 | n3314 ;
  assign n3316 = n411 & n3315 ;
  buffer buf_n3317( .i (n3316), .o (n3317) );
  buffer buf_n3318( .i (n3317), .o (n3318) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n3204( .i (n3203), .o (n3204) );
  buffer buf_n3205( .i (n3204), .o (n3205) );
  buffer buf_n3206( .i (n3205), .o (n3206) );
  buffer buf_n3207( .i (n3206), .o (n3207) );
  buffer buf_n3208( .i (n3207), .o (n3208) );
  buffer buf_n3209( .i (n3208), .o (n3209) );
  buffer buf_n3210( .i (n3209), .o (n3210) );
  buffer buf_n3211( .i (n3210), .o (n3211) );
  buffer buf_n3212( .i (n3211), .o (n3212) );
  buffer buf_n3213( .i (n3212), .o (n3213) );
  buffer buf_n3214( .i (n3213), .o (n3214) );
  buffer buf_n3215( .i (n3214), .o (n3215) );
  buffer buf_n3216( .i (n3215), .o (n3216) );
  buffer buf_n3217( .i (n3216), .o (n3217) );
  buffer buf_n3319( .i (n3084), .o (n3319) );
  buffer buf_n3320( .i (n2881), .o (n3320) );
  assign n3321 = n3319 | n3320 ;
  assign n3322 = ( n71 & n3217 ) | ( n71 & ~n3321 ) | ( n3217 & ~n3321 ) ;
  buffer buf_n3323( .i (n3322), .o (n3323) );
  buffer buf_n3324( .i (n3323), .o (n3324) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  assign n3325 = ( n615 & n2912 ) | ( n615 & ~n3323 ) | ( n2912 & ~n3323 ) ;
  assign n3326 = n3324 & n3325 ;
  buffer buf_n3327( .i (n3326), .o (n3327) );
  buffer buf_n3328( .i (n3327), .o (n3328) );
  buffer buf_n3329( .i (n2923), .o (n3329) );
  assign n3330 = ( n2512 & n3327 ) | ( n2512 & ~n3329 ) | ( n3327 & ~n3329 ) ;
  buffer buf_n3331( .i (n1035), .o (n3331) );
  assign n3332 = ( ~n204 & n2980 ) | ( ~n204 & n3331 ) | ( n2980 & n3331 ) ;
  assign n3333 = n205 | n3332 ;
  assign n3334 = n2512 | n3333 ;
  assign n3335 = ( ~n3328 & n3330 ) | ( ~n3328 & n3334 ) | ( n3330 & n3334 ) ;
  assign n3336 = n377 | n3335 ;
  buffer buf_n3337( .i (n410), .o (n3337) );
  assign n3338 = ( ~n313 & n3336 ) | ( ~n313 & n3337 ) | ( n3336 & n3337 ) ;
  assign n3339 = n314 | n3338 ;
  assign n3340 = ~n3317 & n3339 ;
  assign n3341 = ( n281 & ~n3318 ) | ( n281 & n3340 ) | ( ~n3318 & n3340 ) ;
  buffer buf_n3342( .i (n3341), .o (n3342) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  assign n3343 = ~n137 & n1473 ;
  buffer buf_n3344( .i (n3343), .o (n3344) );
  buffer buf_n3345( .i (n3344), .o (n3345) );
  assign n3346 = ( n172 & ~n205 ) | ( n172 & n3344 ) | ( ~n205 & n3344 ) ;
  assign n3347 = ( n1476 & n3345 ) | ( n1476 & n3346 ) | ( n3345 & n3346 ) ;
  buffer buf_n3348( .i (n3347), .o (n3348) );
  buffer buf_n3349( .i (n3348), .o (n3349) );
  buffer buf_n2940( .i (n2939), .o (n2940) );
  buffer buf_n2941( .i (n2940), .o (n2941) );
  buffer buf_n2942( .i (n2941), .o (n2942) );
  buffer buf_n2943( .i (n2942), .o (n2943) );
  buffer buf_n2944( .i (n2943), .o (n2944) );
  buffer buf_n2945( .i (n2944), .o (n2945) );
  assign n3350 = n330 & n2126 ;
  buffer buf_n3351( .i (n3350), .o (n3351) );
  buffer buf_n3352( .i (n3351), .o (n3352) );
  buffer buf_n3353( .i (n3352), .o (n3353) );
  buffer buf_n3354( .i (n3353), .o (n3354) );
  buffer buf_n3355( .i (n3354), .o (n3355) );
  buffer buf_n3356( .i (n3355), .o (n3356) );
  buffer buf_n3357( .i (n3356), .o (n3357) );
  buffer buf_n3358( .i (n3357), .o (n3358) );
  buffer buf_n3359( .i (n3358), .o (n3359) );
  buffer buf_n3360( .i (n3359), .o (n3360) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  assign n3361 = n584 | n3359 ;
  assign n3362 = ( n2945 & n3360 ) | ( n2945 & ~n3361 ) | ( n3360 & ~n3361 ) ;
  buffer buf_n3363( .i (n3362), .o (n3363) );
  buffer buf_n3364( .i (n3363), .o (n3364) );
  assign n3365 = ~n2469 & n3363 ;
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  assign n3366 = n204 | n1277 ;
  buffer buf_n3367( .i (n3310), .o (n3367) );
  assign n3368 = n3366 | n3367 ;
  assign n3369 = n492 & ~n2714 ;
  buffer buf_n3370( .i (n3369), .o (n3370) );
  buffer buf_n3371( .i (n3370), .o (n3371) );
  buffer buf_n3372( .i (n3371), .o (n3372) );
  buffer buf_n3373( .i (n3372), .o (n3373) );
  buffer buf_n3374( .i (n3373), .o (n3374) );
  buffer buf_n3375( .i (n3374), .o (n3375) );
  buffer buf_n3376( .i (n3375), .o (n3376) );
  buffer buf_n3377( .i (n3376), .o (n3377) );
  buffer buf_n3378( .i (n1954), .o (n3378) );
  assign n3379 = n260 | n3378 ;
  buffer buf_n3380( .i (n3379), .o (n3380) );
  buffer buf_n3381( .i (n3380), .o (n3381) );
  buffer buf_n3382( .i (n3381), .o (n3382) );
  buffer buf_n3383( .i (n3382), .o (n3383) );
  buffer buf_n3384( .i (n3383), .o (n3384) );
  buffer buf_n3385( .i (n3384), .o (n3385) );
  buffer buf_n3386( .i (n3385), .o (n3386) );
  buffer buf_n3387( .i (n3386), .o (n3387) );
  buffer buf_n3388( .i (n3387), .o (n3388) );
  buffer buf_n3389( .i (n3388), .o (n3389) );
  buffer buf_n3390( .i (n3389), .o (n3390) );
  assign n3391 = ( ~n1899 & n2263 ) | ( ~n1899 & n3390 ) | ( n2263 & n3390 ) ;
  assign n3392 = n41 & n3391 ;
  assign n3393 = ~n3377 & n3392 ;
  assign n3394 = n3368 & n3393 ;
  assign n3395 = ( ~n3364 & n3365 ) | ( ~n3364 & n3394 ) | ( n3365 & n3394 ) ;
  assign n3396 = n2634 & n2908 ;
  assign n3397 = ( n2635 & n3127 ) | ( n2635 & n3396 ) | ( n3127 & n3396 ) ;
  assign n3398 = ~n2798 & n3397 ;
  assign n3399 = ~n395 & n2192 ;
  assign n3400 = ( n331 & ~n2193 ) | ( n331 & n3399 ) | ( ~n2193 & n3399 ) ;
  buffer buf_n3401( .i (n3400), .o (n3401) );
  buffer buf_n3402( .i (n3401), .o (n3402) );
  assign n3403 = ( n333 & n3266 ) | ( n333 & n3401 ) | ( n3266 & n3401 ) ;
  assign n3404 = ( n578 & n3402 ) | ( n578 & ~n3403 ) | ( n3402 & ~n3403 ) ;
  buffer buf_n3405( .i (n3404), .o (n3405) );
  buffer buf_n3406( .i (n3405), .o (n3406) );
  buffer buf_n3407( .i (n132), .o (n3407) );
  assign n3408 = ~n3405 & n3407 ;
  assign n3409 = n578 | n1756 ;
  assign n3410 = ( n1757 & ~n3354 ) | ( n1757 & n3409 ) | ( ~n3354 & n3409 ) ;
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n3411( .i (n29), .o (n3411) );
  buffer buf_n3412( .i (n3411), .o (n3412) );
  assign n3413 = ( ~n575 & n1503 ) | ( ~n575 & n3412 ) | ( n1503 & n3412 ) ;
  buffer buf_n3414( .i (n3413), .o (n3414) );
  buffer buf_n3415( .i (n3414), .o (n3415) );
  buffer buf_n3416( .i (n3415), .o (n3416) );
  assign n3417 = ( ~n2372 & n3352 ) | ( ~n2372 & n3414 ) | ( n3352 & n3414 ) ;
  assign n3418 = n2391 & ~n3417 ;
  assign n3419 = ( n2392 & n3416 ) | ( n2392 & ~n3418 ) | ( n3416 & ~n3418 ) ;
  assign n3420 = n3410 & ~n3419 ;
  assign n3421 = ( n3406 & n3408 ) | ( n3406 & n3420 ) | ( n3408 & n3420 ) ;
  assign n3422 = n235 & ~n3421 ;
  assign n3423 = n2798 & ~n3422 ;
  assign n3424 = n3398 | n3423 ;
  buffer buf_n3425( .i (n3424), .o (n3425) );
  buffer buf_n3426( .i (n3425), .o (n3426) );
  assign n3427 = n2154 | n3425 ;
  assign n3428 = ( n2373 & ~n3198 ) | ( n2373 & n3266 ) | ( ~n3198 & n3266 ) ;
  assign n3429 = n131 & n3428 ;
  buffer buf_n3430( .i (n131), .o (n3430) );
  assign n3431 = ( n2392 & n3429 ) | ( n2392 & ~n3430 ) | ( n3429 & ~n3430 ) ;
  buffer buf_n3432( .i (n3431), .o (n3432) );
  buffer buf_n3433( .i (n3432), .o (n3433) );
  assign n3434 = n2386 & ~n3432 ;
  buffer buf_n3435( .i (n265), .o (n3435) );
  assign n3436 = n2391 & n3435 ;
  assign n3437 = n3162 & n3436 ;
  assign n3438 = n2131 & n3299 ;
  assign n3439 = n3437 & n3438 ;
  assign n3440 = n785 & ~n3439 ;
  assign n3441 = ( n3433 & n3434 ) | ( n3433 & n3440 ) | ( n3434 & n3440 ) ;
  buffer buf_n3442( .i (n3441), .o (n3442) );
  buffer buf_n3443( .i (n3442), .o (n3443) );
  assign n3444 = ( n340 & ~n2912 ) | ( n340 & n3442 ) | ( ~n2912 & n3442 ) ;
  assign n3445 = n227 | n1889 ;
  buffer buf_n3446( .i (n3445), .o (n3446) );
  buffer buf_n3447( .i (n3446), .o (n3447) );
  buffer buf_n3449( .i (n295), .o (n3449) );
  assign n3450 = n93 & ~n3449 ;
  buffer buf_n3451( .i (n260), .o (n3451) );
  buffer buf_n3452( .i (n3451), .o (n3452) );
  assign n3453 = ( n2126 & n3450 ) | ( n2126 & n3452 ) | ( n3450 & n3452 ) ;
  buffer buf_n3454( .i (n3452), .o (n3454) );
  assign n3455 = n3453 & ~n3454 ;
  assign n3456 = n3446 & ~n3455 ;
  assign n3457 = ( n2372 & n3447 ) | ( n2372 & ~n3456 ) | ( n3447 & ~n3456 ) ;
  buffer buf_n3458( .i (n3457), .o (n3458) );
  buffer buf_n3459( .i (n3458), .o (n3459) );
  buffer buf_n3460( .i (n2372), .o (n3460) );
  buffer buf_n3461( .i (n3460), .o (n3461) );
  assign n3462 = ( n3430 & n3458 ) | ( n3430 & n3461 ) | ( n3458 & n3461 ) ;
  assign n3463 = ( n878 & n3459 ) | ( n878 & ~n3462 ) | ( n3459 & ~n3462 ) ;
  buffer buf_n3464( .i (n3463), .o (n3464) );
  buffer buf_n3465( .i (n3464), .o (n3465) );
  assign n3466 = n3127 & ~n3464 ;
  buffer buf_n3467( .i (n1724), .o (n3467) );
  assign n3468 = n26 & n3467 ;
  assign n3469 = ( n2180 & n2530 ) | ( n2180 & n3468 ) | ( n2530 & n3468 ) ;
  assign n3470 = ~n2181 & n3469 ;
  buffer buf_n3471( .i (n3470), .o (n3471) );
  buffer buf_n3472( .i (n3471), .o (n3472) );
  buffer buf_n3473( .i (n3472), .o (n3473) );
  buffer buf_n3474( .i (n3473), .o (n3474) );
  buffer buf_n3475( .i (n3474), .o (n3475) );
  buffer buf_n3476( .i (n3412), .o (n3476) );
  assign n3477 = ( n2936 & ~n3473 ) | ( n2936 & n3476 ) | ( ~n3473 & n3476 ) ;
  buffer buf_n3478( .i (n2214), .o (n3478) );
  assign n3479 = n3477 & n3478 ;
  buffer buf_n3480( .i (n3478), .o (n3480) );
  assign n3481 = ( n3475 & ~n3479 ) | ( n3475 & n3480 ) | ( ~n3479 & n3480 ) ;
  buffer buf_n3482( .i (n3481), .o (n3482) );
  buffer buf_n3483( .i (n3482), .o (n3483) );
  assign n3484 = ~n2793 & n3482 ;
  buffer buf_n3485( .i (n2960), .o (n3485) );
  assign n3486 = ( n3483 & n3484 ) | ( n3483 & n3485 ) | ( n3484 & n3485 ) ;
  buffer buf_n3487( .i (n2391), .o (n3487) );
  buffer buf_n3488( .i (n3016), .o (n3488) );
  assign n3489 = ( n3430 & ~n3487 ) | ( n3430 & n3488 ) | ( ~n3487 & n3488 ) ;
  assign n3490 = ( n1272 & n2960 ) | ( n1272 & n3489 ) | ( n2960 & n3489 ) ;
  buffer buf_n3448( .i (n3447), .o (n3448) );
  assign n3491 = n2212 | n3471 ;
  assign n3492 = ( ~n3412 & n3472 ) | ( ~n3412 & n3491 ) | ( n3472 & n3491 ) ;
  buffer buf_n3493( .i (n3492), .o (n3493) );
  buffer buf_n3494( .i (n3493), .o (n3494) );
  assign n3495 = ~n398 & n3493 ;
  assign n3496 = ( ~n3448 & n3494 ) | ( ~n3448 & n3495 ) | ( n3494 & n3495 ) ;
  buffer buf_n3497( .i (n3496), .o (n3497) );
  buffer buf_n3498( .i (n3497), .o (n3498) );
  buffer buf_n3499( .i (n3461), .o (n3499) );
  assign n3500 = ~n3497 & n3499 ;
  assign n3501 = ( n3490 & n3498 ) | ( n3490 & ~n3500 ) | ( n3498 & ~n3500 ) ;
  assign n3502 = n3486 | n3501 ;
  assign n3503 = ( n3465 & n3466 ) | ( n3465 & ~n3502 ) | ( n3466 & ~n3502 ) ;
  buffer buf_n3504( .i (n2619), .o (n3504) );
  assign n3505 = n3503 | n3504 ;
  assign n3506 = ( n3443 & ~n3444 ) | ( n3443 & n3505 ) | ( ~n3444 & n3505 ) ;
  buffer buf_n3507( .i (n56), .o (n3507) );
  assign n3508 = n88 & n3507 ;
  buffer buf_n3509( .i (n3508), .o (n3509) );
  buffer buf_n3510( .i (n3509), .o (n3510) );
  buffer buf_n3511( .i (n3510), .o (n3511) );
  buffer buf_n3512( .i (n3511), .o (n3512) );
  buffer buf_n3513( .i (n3512), .o (n3513) );
  assign n3523 = n3411 & n3513 ;
  buffer buf_n3524( .i (n3523), .o (n3524) );
  assign n3526 = n968 & n3524 ;
  buffer buf_n3527( .i (n2195), .o (n3527) );
  assign n3528 = ( n333 & n3526 ) | ( n333 & n3527 ) | ( n3526 & n3527 ) ;
  assign n3529 = ~n334 & n3528 ;
  buffer buf_n3530( .i (n3529), .o (n3530) );
  buffer buf_n3531( .i (n3530), .o (n3531) );
  buffer buf_n3532( .i (n3531), .o (n3532) );
  assign n3533 = ( ~n401 & n2789 ) | ( ~n401 & n3530 ) | ( n2789 & n3530 ) ;
  assign n3534 = n2718 | n3533 ;
  assign n3535 = ( ~n2719 & n3532 ) | ( ~n2719 & n3534 ) | ( n3532 & n3534 ) ;
  buffer buf_n3536( .i (n3535), .o (n3536) );
  buffer buf_n3537( .i (n3536), .o (n3537) );
  assign n3538 = ~n2967 & n3536 ;
  assign n3539 = ( ~n2181 & n2600 ) | ( ~n2181 & n2887 ) | ( n2600 & n2887 ) ;
  assign n3540 = n3451 & ~n3539 ;
  assign n3541 = n777 & ~n3451 ;
  assign n3542 = ( n3010 & n3540 ) | ( n3010 & ~n3541 ) | ( n3540 & ~n3541 ) ;
  buffer buf_n3543( .i (n3542), .o (n3543) );
  buffer buf_n3544( .i (n3011), .o (n3544) );
  assign n3545 = ( ~n264 & n3543 ) | ( ~n264 & n3544 ) | ( n3543 & n3544 ) ;
  assign n3546 = ( n396 & n490 ) | ( n396 & n2193 ) | ( n490 & n2193 ) ;
  assign n3547 = n3543 & n3546 ;
  assign n3548 = ( n265 & n3545 ) | ( n265 & n3547 ) | ( n3545 & n3547 ) ;
  buffer buf_n3549( .i (n3548), .o (n3549) );
  assign n3550 = ( n1894 & n2590 ) | ( n1894 & n3549 ) | ( n2590 & n3549 ) ;
  assign n3551 = n2210 & n3549 ;
  assign n3552 = ( ~n1895 & n3550 ) | ( ~n1895 & n3551 ) | ( n3550 & n3551 ) ;
  buffer buf_n3553( .i (n3552), .o (n3553) );
  buffer buf_n3554( .i (n3553), .o (n3554) );
  assign n3555 = n910 & ~n1892 ;
  buffer buf_n3556( .i (n3555), .o (n3556) );
  buffer buf_n3557( .i (n3556), .o (n3557) );
  buffer buf_n3558( .i (n2642), .o (n3558) );
  assign n3559 = ~n3556 & n3558 ;
  assign n3560 = ( n3499 & ~n3557 ) | ( n3499 & n3559 ) | ( ~n3557 & n3559 ) ;
  buffer buf_n3525( .i (n3524), .o (n3525) );
  buffer buf_n3561( .i (n3188), .o (n3561) );
  assign n3562 = ( n607 & ~n3524 ) | ( n607 & n3561 ) | ( ~n3524 & n3561 ) ;
  assign n3563 = n3525 & n3562 ;
  buffer buf_n3564( .i (n3563), .o (n3564) );
  buffer buf_n3565( .i (n3564), .o (n3565) );
  assign n3569 = n1894 | n2590 ;
  assign n3570 = ( n1895 & ~n3565 ) | ( n1895 & n3569 ) | ( ~n3565 & n3569 ) ;
  assign n3571 = ( n2908 & ~n3560 ) | ( n2908 & n3570 ) | ( ~n3560 & n3570 ) ;
  assign n3572 = n3553 & ~n3571 ;
  assign n3573 = ( n2978 & n3554 ) | ( n2978 & ~n3572 ) | ( n3554 & ~n3572 ) ;
  buffer buf_n3566( .i (n3565), .o (n3566) );
  buffer buf_n3567( .i (n3566), .o (n3567) );
  buffer buf_n3568( .i (n3567), .o (n3568) );
  assign n3574 = ~n291 & n483 ;
  assign n3575 = ~n902 & n3574 ;
  buffer buf_n3576( .i (n3575), .o (n3576) );
  buffer buf_n3577( .i (n3576), .o (n3577) );
  buffer buf_n3578( .i (n3577), .o (n3578) );
  buffer buf_n3579( .i (n153), .o (n3579) );
  buffer buf_n3580( .i (n3579), .o (n3580) );
  assign n3581 = ( n600 & n2929 ) | ( n600 & n3580 ) | ( n2929 & n3580 ) ;
  assign n3582 = ~n2930 & n3581 ;
  assign n3583 = ( n3181 & n3576 ) | ( n3181 & n3582 ) | ( n3576 & n3582 ) ;
  assign n3584 = n2759 & ~n3583 ;
  buffer buf_n3585( .i (n2759), .o (n3585) );
  assign n3586 = ( n3578 & ~n3584 ) | ( n3578 & n3585 ) | ( ~n3584 & n3585 ) ;
  assign n3587 = n3411 & n3586 ;
  buffer buf_n3588( .i (n3587), .o (n3588) );
  buffer buf_n3589( .i (n3588), .o (n3589) );
  assign n3590 = ( n1420 & n2180 ) | ( n1420 & ~n3182 ) | ( n2180 & ~n3182 ) ;
  buffer buf_n3591( .i (n2180), .o (n3591) );
  assign n3592 = n3590 & ~n3591 ;
  buffer buf_n3593( .i (n3592), .o (n3593) );
  buffer buf_n3594( .i (n3593), .o (n3594) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n3595( .i (n329), .o (n3595) );
  assign n3596 = ( n688 & n3593 ) | ( n688 & ~n3595 ) | ( n3593 & ~n3595 ) ;
  assign n3597 = ~n3594 & n3596 ;
  assign n3598 = n3588 | n3597 ;
  buffer buf_n3599( .i (n264), .o (n3599) );
  assign n3600 = ( n3589 & n3598 ) | ( n3589 & ~n3599 ) | ( n3598 & ~n3599 ) ;
  buffer buf_n3601( .i (n3600), .o (n3601) );
  assign n3602 = ( n3370 & ~n3564 ) | ( n3370 & n3601 ) | ( ~n3564 & n3601 ) ;
  assign n3603 = n3488 & ~n3601 ;
  assign n3604 = ( n3565 & n3602 ) | ( n3565 & ~n3603 ) | ( n3602 & ~n3603 ) ;
  buffer buf_n3605( .i (n3604), .o (n3605) );
  assign n3606 = ( n582 & n3567 ) | ( n582 & ~n3605 ) | ( n3567 & ~n3605 ) ;
  assign n3607 = n403 & ~n3605 ;
  assign n3608 = ( ~n3568 & n3606 ) | ( ~n3568 & n3607 ) | ( n3606 & n3607 ) ;
  assign n3609 = n3573 & n3608 ;
  assign n3610 = ( ~n3537 & n3538 ) | ( ~n3537 & n3609 ) | ( n3538 & n3609 ) ;
  assign n3611 = n3506 & n3610 ;
  assign n3612 = ( n3426 & ~n3427 ) | ( n3426 & n3611 ) | ( ~n3427 & n3611 ) ;
  buffer buf_n3613( .i (n3612), .o (n3613) );
  assign n3614 = ( n3348 & n3395 ) | ( n3348 & n3613 ) | ( n3395 & n3613 ) ;
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  assign n3615 = n78 & n3613 ;
  assign n3616 = ( ~n3349 & n3614 ) | ( ~n3349 & n3615 ) | ( n3614 & n3615 ) ;
  assign n3617 = n445 & ~n3616 ;
  assign n3618 = ~n295 & n3378 ;
  buffer buf_n3619( .i (n3618), .o (n3619) );
  buffer buf_n3620( .i (n3619), .o (n3620) );
  buffer buf_n3621( .i (n3620), .o (n3621) );
  buffer buf_n3622( .i (n3621), .o (n3622) );
  buffer buf_n3623( .i (n3622), .o (n3623) );
  buffer buf_n3624( .i (n3623), .o (n3624) );
  buffer buf_n3625( .i (n3624), .o (n3625) );
  buffer buf_n3626( .i (n3625), .o (n3626) );
  buffer buf_n3627( .i (n3626), .o (n3627) );
  assign n3628 = ( n1415 & n1759 ) | ( n1415 & ~n3626 ) | ( n1759 & ~n3626 ) ;
  assign n3629 = n3627 & n3628 ;
  buffer buf_n3630( .i (n3629), .o (n3630) );
  buffer buf_n3631( .i (n3630), .o (n3631) );
  buffer buf_n3632( .i (n3631), .o (n3632) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n3633( .i (n2908), .o (n3633) );
  buffer buf_n3634( .i (n3633), .o (n3634) );
  buffer buf_n3635( .i (n3634), .o (n3635) );
  assign n3636 = ( n571 & n3630 ) | ( n571 & ~n3635 ) | ( n3630 & ~n3635 ) ;
  assign n3637 = n2710 & ~n3636 ;
  assign n3638 = ( n2481 & n3632 ) | ( n2481 & ~n3637 ) | ( n3632 & ~n3637 ) ;
  buffer buf_n3639( .i (n3638), .o (n3639) );
  buffer buf_n3640( .i (n3639), .o (n3640) );
  assign n3641 = ( n376 & n3150 ) | ( n376 & ~n3639 ) | ( n3150 & ~n3639 ) ;
  assign n3642 = n3162 | n3487 ;
  buffer buf_n3643( .i (n3642), .o (n3643) );
  buffer buf_n3644( .i (n3643), .o (n3644) );
  buffer buf_n3645( .i (n3644), .o (n3645) );
  buffer buf_n3646( .i (n3645), .o (n3646) );
  buffer buf_n3647( .i (n3646), .o (n3647) );
  buffer buf_n2721( .i (n2720), .o (n2721) );
  buffer buf_n3648( .i (n3098), .o (n3648) );
  assign n3649 = n2721 & n3648 ;
  assign n3650 = ( ~n204 & n3647 ) | ( ~n204 & n3649 ) | ( n3647 & n3649 ) ;
  buffer buf_n3651( .i (n332), .o (n3651) );
  buffer buf_n3652( .i (n3651), .o (n3652) );
  buffer buf_n3653( .i (n3652), .o (n3653) );
  assign n3654 = ( n2590 & n3162 ) | ( n2590 & n3653 ) | ( n3162 & n3653 ) ;
  buffer buf_n3655( .i (n3654), .o (n3655) );
  buffer buf_n3656( .i (n3655), .o (n3656) );
  buffer buf_n3657( .i (n400), .o (n3657) );
  assign n3658 = ( ~n2591 & n3163 ) | ( ~n2591 & n3657 ) | ( n3163 & n3657 ) ;
  assign n3659 = n3655 | n3658 ;
  assign n3660 = ( ~n338 & n3656 ) | ( ~n338 & n3659 ) | ( n3656 & n3659 ) ;
  buffer buf_n3661( .i (n2795), .o (n3661) );
  assign n3662 = ( ~n1646 & n3660 ) | ( ~n1646 & n3661 ) | ( n3660 & n3661 ) ;
  assign n3663 = n3211 & n3561 ;
  assign n3664 = n1428 & n3663 ;
  buffer buf_n3665( .i (n3664), .o (n3665) );
  buffer buf_n3666( .i (n3665), .o (n3666) );
  assign n3667 = n3653 & ~n3665 ;
  assign n3668 = ( n2591 & n3666 ) | ( n2591 & ~n3667 ) | ( n3666 & ~n3667 ) ;
  assign n3669 = n304 & n3668 ;
  buffer buf_n3670( .i (n3485), .o (n3670) );
  assign n3671 = n3669 & n3670 ;
  assign n3672 = ~n3661 & n3671 ;
  assign n3673 = ( n3089 & n3662 ) | ( n3089 & ~n3672 ) | ( n3662 & ~n3672 ) ;
  buffer buf_n3674( .i (n3673), .o (n3674) );
  buffer buf_n3675( .i (n3285), .o (n3675) );
  assign n3676 = ( n3650 & n3674 ) | ( n3650 & n3675 ) | ( n3674 & n3675 ) ;
  assign n3677 = ( ~n392 & n2861 ) | ( ~n392 & n2890 ) | ( n2861 & n2890 ) ;
  buffer buf_n3678( .i (n3677), .o (n3678) );
  buffer buf_n3679( .i (n3678), .o (n3679) );
  buffer buf_n3680( .i (n3679), .o (n3680) );
  buffer buf_n3681( .i (n3680), .o (n3681) );
  buffer buf_n3682( .i (n3681), .o (n3682) );
  buffer buf_n3683( .i (n3682), .o (n3683) );
  buffer buf_n3684( .i (n3683), .o (n3684) );
  buffer buf_n3685( .i (n3684), .o (n3685) );
  buffer buf_n3686( .i (n3685), .o (n3686) );
  assign n3687 = ( n304 & ~n2142 ) | ( n304 & n3686 ) | ( ~n2142 & n3686 ) ;
  assign n3688 = ( ~n304 & n402 ) | ( ~n304 & n3686 ) | ( n402 & n3686 ) ;
  assign n3689 = n3687 & n3688 ;
  buffer buf_n3690( .i (n3689), .o (n3690) );
  buffer buf_n3691( .i (n3690), .o (n3691) );
  buffer buf_n2958( .i (n2957), .o (n2958) );
  buffer buf_n2959( .i (n2958), .o (n2959) );
  assign n3692 = ( n2959 & n3648 ) | ( n2959 & n3690 ) | ( n3648 & n3690 ) ;
  assign n3693 = ~n3691 & n3692 ;
  assign n3694 = ( ~n3674 & n3675 ) | ( ~n3674 & n3693 ) | ( n3675 & n3693 ) ;
  assign n3695 = n3676 & ~n3694 ;
  assign n3696 = n3150 & ~n3695 ;
  assign n3697 = ( n3640 & n3641 ) | ( n3640 & n3696 ) | ( n3641 & n3696 ) ;
  assign n3698 = n3358 & n3634 ;
  assign n3699 = n2944 & n3698 ;
  buffer buf_n3700( .i (n3699), .o (n3700) );
  buffer buf_n3701( .i (n3700), .o (n3701) );
  buffer buf_n3702( .i (n3701), .o (n3702) );
  buffer buf_n3703( .i (n2410), .o (n3703) );
  assign n3704 = n2637 & ~n3703 ;
  buffer buf_n3705( .i (n3435), .o (n3705) );
  buffer buf_n3706( .i (n3705), .o (n3706) );
  buffer buf_n3707( .i (n3706), .o (n3707) );
  assign n3708 = n2028 & n3707 ;
  buffer buf_n3709( .i (n3708), .o (n3709) );
  buffer buf_n3710( .i (n3709), .o (n3710) );
  assign n3711 = n3703 & ~n3710 ;
  assign n3712 = n3704 | n3711 ;
  assign n3713 = ( ~n3675 & n3700 ) | ( ~n3675 & n3712 ) | ( n3700 & n3712 ) ;
  assign n3714 = n2469 | n3713 ;
  assign n3715 = ( ~n241 & n3702 ) | ( ~n241 & n3714 ) | ( n3702 & n3714 ) ;
  assign n3716 = ~n400 & n3430 ;
  assign n3717 = ( ~n2960 & n3407 ) | ( ~n2960 & n3716 ) | ( n3407 & n3716 ) ;
  assign n3718 = n580 & n3706 ;
  buffer buf_n3719( .i (n3266), .o (n3719) );
  assign n3720 = n3199 & ~n3719 ;
  buffer buf_n3721( .i (n3199), .o (n3721) );
  assign n3722 = ( ~n3487 & n3720 ) | ( ~n3487 & n3721 ) | ( n3720 & n3721 ) ;
  assign n3723 = n3706 | n3722 ;
  assign n3724 = ( n3717 & n3718 ) | ( n3717 & n3723 ) | ( n3718 & n3723 ) ;
  buffer buf_n3725( .i (n3724), .o (n3725) );
  buffer buf_n3726( .i (n3725), .o (n3726) );
  assign n3727 = n2410 & ~n3725 ;
  buffer buf_n3728( .i (n357), .o (n3728) );
  assign n3729 = n293 & ~n3728 ;
  buffer buf_n3730( .i (n3729), .o (n3730) );
  buffer buf_n3731( .i (n3730), .o (n3731) );
  assign n3732 = ( n2600 & ~n3291 ) | ( n2600 & n3730 ) | ( ~n3291 & n3730 ) ;
  assign n3733 = ( n3005 & n3731 ) | ( n3005 & n3732 ) | ( n3731 & n3732 ) ;
  buffer buf_n3734( .i (n3733), .o (n3734) );
  buffer buf_n3735( .i (n3734), .o (n3735) );
  assign n3736 = n228 | n3734 ;
  buffer buf_n3737( .i (n2890), .o (n3737) );
  buffer buf_n3738( .i (n3737), .o (n3738) );
  assign n3739 = ( n3449 & ~n3451 ) | ( n3449 & n3738 ) | ( ~n3451 & n3738 ) ;
  assign n3740 = ( n3380 & n3595 ) | ( n3380 & ~n3739 ) | ( n3595 & ~n3739 ) ;
  assign n3741 = ( ~n354 & n387 ) | ( ~n354 & n3232 ) | ( n387 & n3232 ) ;
  assign n3742 = n290 & n3741 ;
  assign n3743 = ( ~n291 & n389 ) | ( ~n291 & n3742 ) | ( n389 & n3742 ) ;
  buffer buf_n3744( .i (n3743), .o (n3744) );
  assign n3745 = ( n293 & ~n3728 ) | ( n293 & n3744 ) | ( ~n3728 & n3744 ) ;
  assign n3746 = n2291 & n3744 ;
  assign n3747 = ( ~n294 & n3745 ) | ( ~n294 & n3746 ) | ( n3745 & n3746 ) ;
  buffer buf_n3748( .i (n3747), .o (n3748) );
  buffer buf_n3749( .i (n3748), .o (n3749) );
  assign n3750 = ~n3738 & n3748 ;
  assign n3751 = ( n3619 & n3749 ) | ( n3619 & n3750 ) | ( n3749 & n3750 ) ;
  assign n3752 = n3740 & n3751 ;
  assign n3753 = ( n3735 & ~n3736 ) | ( n3735 & n3752 ) | ( ~n3736 & n3752 ) ;
  buffer buf_n3754( .i (n3753), .o (n3754) );
  assign n3755 = ( ~n3301 & n3652 ) | ( ~n3301 & n3754 ) | ( n3652 & n3754 ) ;
  assign n3756 = n3480 & n3754 ;
  assign n3757 = ( n3299 & n3755 ) | ( n3299 & n3756 ) | ( n3755 & n3756 ) ;
  buffer buf_n3758( .i (n3757), .o (n3758) );
  buffer buf_n3759( .i (n3758), .o (n3759) );
  buffer buf_n3760( .i (n2499), .o (n3760) );
  assign n3761 = ( n3485 & ~n3758 ) | ( n3485 & n3760 ) | ( ~n3758 & n3760 ) ;
  assign n3762 = ( ~n1836 & n2631 ) | ( ~n1836 & n3719 ) | ( n2631 & n3719 ) ;
  buffer buf_n3763( .i (n298), .o (n3763) );
  assign n3764 = ( ~n264 & n397 ) | ( ~n264 & n3763 ) | ( n397 & n3763 ) ;
  assign n3765 = ( ~n575 & n2654 ) | ( ~n575 & n3188 ) | ( n2654 & n3188 ) ;
  assign n3766 = ~n3763 & n3765 ;
  assign n3767 = ( n3599 & n3764 ) | ( n3599 & ~n3766 ) | ( n3764 & ~n3766 ) ;
  buffer buf_n3768( .i (n3767), .o (n3768) );
  assign n3769 = ( n3705 & n3762 ) | ( n3705 & n3768 ) | ( n3762 & n3768 ) ;
  assign n3770 = n398 & ~n1835 ;
  assign n3771 = ( n578 & ~n2130 ) | ( n578 & n3770 ) | ( ~n2130 & n3770 ) ;
  assign n3772 = ( ~n3705 & n3768 ) | ( ~n3705 & n3771 ) | ( n3768 & n3771 ) ;
  assign n3773 = n3769 & n3772 ;
  assign n3774 = n3485 | n3773 ;
  assign n3775 = ( n3759 & n3761 ) | ( n3759 & n3774 ) | ( n3761 & n3774 ) ;
  buffer buf_n3776( .i (n3004), .o (n3776) );
  buffer buf_n3777( .i (n3776), .o (n3777) );
  assign n3778 = ( ~n331 & n3620 ) | ( ~n331 & n3777 ) | ( n3620 & n3777 ) ;
  assign n3779 = n186 & n290 ;
  buffer buf_n3780( .i (n3779), .o (n3780) );
  buffer buf_n3781( .i (n3780), .o (n3781) );
  buffer buf_n3782( .i (n3781), .o (n3782) );
  buffer buf_n3783( .i (n3782), .o (n3783) );
  buffer buf_n3784( .i (n3783), .o (n3784) );
  buffer buf_n3785( .i (n3784), .o (n3785) );
  assign n3786 = n394 & ~n3784 ;
  assign n3787 = ( n227 & ~n3785 ) | ( n227 & n3786 ) | ( ~n3785 & n3786 ) ;
  buffer buf_n3788( .i (n3595), .o (n3788) );
  assign n3789 = n3787 | n3788 ;
  assign n3790 = ( n3621 & ~n3778 ) | ( n3621 & n3789 ) | ( ~n3778 & n3789 ) ;
  assign n3791 = n3599 & n3790 ;
  assign n3792 = n229 | n491 ;
  assign n3793 = ~n3599 & n3792 ;
  assign n3794 = n3791 | n3793 ;
  assign n3795 = n3488 | n3794 ;
  buffer buf_n3796( .i (n3795), .o (n3796) );
  buffer buf_n3797( .i (n3796), .o (n3797) );
  assign n3798 = ~n2947 & n3796 ;
  assign n3799 = ( ~n3357 & n3797 ) | ( ~n3357 & n3798 ) | ( n3797 & n3798 ) ;
  assign n3800 = n3775 & n3799 ;
  assign n3801 = ( n3726 & n3727 ) | ( n3726 & n3800 ) | ( n3727 & n3800 ) ;
  buffer buf_n3802( .i (n226), .o (n3802) );
  buffer buf_n3803( .i (n3802), .o (n3803) );
  buffer buf_n3804( .i (n3803), .o (n3804) );
  assign n3805 = ( ~n397 & n3561 ) | ( ~n397 & n3804 ) | ( n3561 & n3804 ) ;
  buffer buf_n3806( .i (n2192), .o (n3806) );
  buffer buf_n3807( .i (n3806), .o (n3807) );
  buffer buf_n3808( .i (n395), .o (n3808) );
  buffer buf_n3809( .i (n3808), .o (n3809) );
  assign n3810 = ( n3804 & n3807 ) | ( n3804 & n3809 ) | ( n3807 & n3809 ) ;
  assign n3811 = ~n3805 & n3810 ;
  buffer buf_n3812( .i (n3811), .o (n3812) );
  buffer buf_n3813( .i (n3812), .o (n3813) );
  assign n3814 = n3435 & n3719 ;
  assign n3815 = ( n3653 & ~n3812 ) | ( n3653 & n3814 ) | ( ~n3812 & n3814 ) ;
  assign n3816 = n3813 & n3815 ;
  buffer buf_n3817( .i (n3816), .o (n3817) );
  buffer buf_n3818( .i (n3817), .o (n3818) );
  assign n3819 = ~n3294 & n3788 ;
  buffer buf_n3820( .i (n3819), .o (n3820) );
  assign n3821 = n3198 & n3820 ;
  assign n3822 = ( n3296 & n3527 ) | ( n3296 & ~n3820 ) | ( n3527 & ~n3820 ) ;
  assign n3823 = ( n3435 & n3821 ) | ( n3435 & ~n3822 ) | ( n3821 & ~n3822 ) ;
  buffer buf_n3824( .i (n3823), .o (n3824) );
  buffer buf_n3825( .i (n3824), .o (n3825) );
  assign n3826 = ( n2793 & n3407 ) | ( n2793 & n3824 ) | ( n3407 & n3824 ) ;
  assign n3827 = ( n1946 & n3788 ) | ( n1946 & ~n3808 ) | ( n3788 & ~n3808 ) ;
  assign n3828 = ( n697 & n3295 ) | ( n697 & ~n3827 ) | ( n3295 & ~n3827 ) ;
  buffer buf_n3829( .i (n3828), .o (n3829) );
  buffer buf_n3830( .i (n3829), .o (n3830) );
  assign n3831 = n3199 & n3829 ;
  assign n3832 = ( ~n2898 & n3830 ) | ( ~n2898 & n3831 ) | ( n3830 & n3831 ) ;
  assign n3833 = n2793 | n3832 ;
  assign n3834 = ( ~n3825 & n3826 ) | ( ~n3825 & n3833 ) | ( n3826 & n3833 ) ;
  assign n3835 = ( n2626 & n3004 ) | ( n2626 & ~n3738 ) | ( n3004 & ~n3738 ) ;
  assign n3836 = ( n3272 & n3595 ) | ( n3272 & n3835 ) | ( n3595 & n3835 ) ;
  buffer buf_n3837( .i (n3836), .o (n3837) );
  assign n3838 = ( ~n499 & n3763 ) | ( ~n499 & n3837 ) | ( n3763 & n3837 ) ;
  assign n3839 = n3804 & n3837 ;
  assign n3840 = ( n500 & n3838 ) | ( n500 & n3839 ) | ( n3838 & n3839 ) ;
  assign n3841 = ( ~n2868 & n3010 ) | ( ~n2868 & n3802 ) | ( n3010 & n3802 ) ;
  buffer buf_n3171( .i (n3170), .o (n3171) );
  buffer buf_n3172( .i (n3171), .o (n3172) );
  buffer buf_n3173( .i (n3172), .o (n3173) );
  buffer buf_n3174( .i (n3173), .o (n3174) );
  buffer buf_n3175( .i (n3174), .o (n3175) );
  assign n3842 = ( n3071 & ~n3591 ) | ( n3071 & n3737 ) | ( ~n3591 & n3737 ) ;
  assign n3843 = ( n126 & n3175 ) | ( n126 & n3842 ) | ( n3175 & n3842 ) ;
  assign n3844 = ( n2868 & n3802 ) | ( n2868 & n3843 ) | ( n3802 & n3843 ) ;
  assign n3845 = n3841 & ~n3844 ;
  buffer buf_n3846( .i (n3845), .o (n3846) );
  buffer buf_n3847( .i (n3846), .o (n3847) );
  assign n3848 = n3527 | n3846 ;
  assign n3849 = ( ~n3840 & n3847 ) | ( ~n3840 & n3848 ) | ( n3847 & n3848 ) ;
  assign n3850 = n3705 | n3849 ;
  buffer buf_n2766( .i (n2765), .o (n2766) );
  buffer buf_n2767( .i (n2766), .o (n2767) );
  buffer buf_n2768( .i (n2767), .o (n2768) );
  assign n3851 = ~n3544 & n3621 ;
  buffer buf_n3852( .i (n3544), .o (n3852) );
  assign n3853 = ( n2768 & n3851 ) | ( n2768 & ~n3852 ) | ( n3851 & ~n3852 ) ;
  assign n3854 = ~n3652 & n3853 ;
  buffer buf_n3855( .i (n3454), .o (n3855) );
  buffer buf_n3856( .i (n3855), .o (n3856) );
  buffer buf_n3857( .i (n3856), .o (n3857) );
  buffer buf_n3858( .i (n3857), .o (n3858) );
  assign n3859 = ~n3854 & n3858 ;
  assign n3860 = n3850 & ~n3859 ;
  buffer buf_n3861( .i (n3860), .o (n3861) );
  assign n3862 = ( n3817 & n3834 ) | ( n3817 & ~n3861 ) | ( n3834 & ~n3861 ) ;
  buffer buf_n3863( .i (n303), .o (n3863) );
  buffer buf_n3864( .i (n3863), .o (n3864) );
  assign n3865 = n3861 | n3864 ;
  assign n3866 = ( n3818 & ~n3862 ) | ( n3818 & n3865 ) | ( ~n3862 & n3865 ) ;
  buffer buf_n3867( .i (n3866), .o (n3867) );
  assign n3868 = ( n3285 & ~n3801 ) | ( n3285 & n3867 ) | ( ~n3801 & n3867 ) ;
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n2221( .i (n2220), .o (n2221) );
  buffer buf_n2222( .i (n2221), .o (n2222) );
  assign n3869 = n3707 & ~n3863 ;
  assign n3870 = ( ~n550 & n3864 ) | ( ~n550 & n3869 ) | ( n3864 & n3869 ) ;
  assign n3871 = n2221 | n3870 ;
  buffer buf_n3872( .i (n3163), .o (n3872) );
  assign n3873 = ( n402 & ~n2718 ) | ( n402 & n3872 ) | ( ~n2718 & n3872 ) ;
  assign n3874 = n3120 & n3858 ;
  buffer buf_n3875( .i (n3487), .o (n3875) );
  assign n3876 = n3874 & n3875 ;
  assign n3877 = n402 & n3876 ;
  assign n3878 = ( ~n3633 & n3873 ) | ( ~n3633 & n3877 ) | ( n3873 & n3877 ) ;
  assign n3879 = n2022 | n2213 ;
  assign n3880 = ( ~n630 & n2023 ) | ( ~n630 & n3879 ) | ( n2023 & n3879 ) ;
  buffer buf_n3881( .i (n3880), .o (n3881) );
  buffer buf_n3882( .i (n3881), .o (n3882) );
  assign n3883 = ( n778 & n2212 ) | ( n778 & n3776 ) | ( n2212 & n3776 ) ;
  buffer buf_n3884( .i (n3883), .o (n3884) );
  assign n3885 = ( n2128 & ~n3561 ) | ( n2128 & n3884 ) | ( ~n3561 & n3884 ) ;
  assign n3886 = n3855 & n3884 ;
  assign n3887 = ( n1581 & n3885 ) | ( n1581 & n3886 ) | ( n3885 & n3886 ) ;
  assign n3888 = n2862 | n3290 ;
  buffer buf_n3889( .i (n293), .o (n3889) );
  buffer buf_n3890( .i (n3889), .o (n3890) );
  assign n3891 = ( n3291 & n3888 ) | ( n3291 & n3890 ) | ( n3888 & n3890 ) ;
  assign n3892 = ~n393 & n3270 ;
  assign n3893 = ( ~n790 & n3891 ) | ( ~n790 & n3892 ) | ( n3891 & n3892 ) ;
  buffer buf_n3894( .i (n3893), .o (n3894) );
  buffer buf_n3895( .i (n3894), .o (n3895) );
  assign n3896 = n3806 & n3894 ;
  assign n3897 = ( n2627 & ~n2889 ) | ( n2627 & n3452 ) | ( ~n2889 & n3452 ) ;
  buffer buf_n3898( .i (n3591), .o (n3898) );
  assign n3899 = n394 | n3898 ;
  assign n3900 = ( ~n1832 & n2212 ) | ( ~n1832 & n3899 ) | ( n2212 & n3899 ) ;
  assign n3901 = n3897 & n3900 ;
  assign n3902 = ( ~n3895 & n3896 ) | ( ~n3895 & n3901 ) | ( n3896 & n3901 ) ;
  buffer buf_n3903( .i (n3902), .o (n3903) );
  assign n3904 = ( ~n3881 & n3887 ) | ( ~n3881 & n3903 ) | ( n3887 & n3903 ) ;
  assign n3905 = n3301 & n3903 ;
  assign n3906 = ( n3882 & n3904 ) | ( n3882 & n3905 ) | ( n3904 & n3905 ) ;
  buffer buf_n3907( .i (n3906), .o (n3907) );
  buffer buf_n3908( .i (n3907), .o (n3908) );
  assign n3909 = n3872 | n3907 ;
  assign n3910 = n2864 & ~n3004 ;
  buffer buf_n3911( .i (n3910), .o (n3911) );
  buffer buf_n3912( .i (n3911), .o (n3912) );
  buffer buf_n3913( .i (n3912), .o (n3913) );
  buffer buf_n2866( .i (n2865), .o (n2866) );
  buffer buf_n2867( .i (n2866), .o (n2867) );
  assign n3914 = ( n3777 & ~n3806 ) | ( n3777 & n3911 ) | ( ~n3806 & n3911 ) ;
  assign n3915 = ( n2214 & n2867 ) | ( n2214 & ~n3914 ) | ( n2867 & ~n3914 ) ;
  assign n3916 = ~n3913 & n3915 ;
  buffer buf_n3917( .i (n3916), .o (n3917) );
  buffer buf_n3918( .i (n3917), .o (n3918) );
  assign n3919 = ( n3299 & ~n3653 ) | ( n3299 & n3917 ) | ( ~n3653 & n3917 ) ;
  buffer buf_n2520( .i (n2519), .o (n2520) );
  buffer buf_n2521( .i (n2520), .o (n2521) );
  buffer buf_n2522( .i (n2521), .o (n2522) );
  buffer buf_n2523( .i (n2522), .o (n2523) );
  buffer buf_n2524( .i (n2523), .o (n2524) );
  buffer buf_n2525( .i (n2524), .o (n2525) );
  buffer buf_n2526( .i (n2525), .o (n2526) );
  buffer buf_n2527( .i (n2526), .o (n2527) );
  assign n3920 = ( n2527 & n3297 ) | ( n2527 & ~n3857 ) | ( n3297 & ~n3857 ) ;
  buffer buf_n3921( .i (n3301), .o (n3921) );
  assign n3922 = n3920 & n3921 ;
  assign n3923 = ( ~n3918 & n3919 ) | ( ~n3918 & n3922 ) | ( n3919 & n3922 ) ;
  assign n3924 = ~n2830 & n3855 ;
  buffer buf_n3925( .i (n3924), .o (n3925) );
  buffer buf_n3926( .i (n3925), .o (n3926) );
  buffer buf_n3927( .i (n3926), .o (n3927) );
  assign n3928 = ( n1835 & n2952 ) | ( n1835 & n3198 ) | ( n2952 & n3198 ) ;
  assign n3929 = ( n3480 & ~n3925 ) | ( n3480 & n3928 ) | ( ~n3925 & n3928 ) ;
  buffer buf_n3930( .i (n3527), .o (n3930) );
  buffer buf_n3931( .i (n3930), .o (n3931) );
  assign n3932 = n3929 & n3931 ;
  assign n3933 = ( n3875 & n3927 ) | ( n3875 & ~n3932 ) | ( n3927 & ~n3932 ) ;
  assign n3934 = n3923 | n3933 ;
  assign n3935 = ( ~n3908 & n3909 ) | ( ~n3908 & n3934 ) | ( n3909 & n3934 ) ;
  assign n3936 = n3878 | n3935 ;
  assign n3937 = ( ~n2222 & n3871 ) | ( ~n2222 & n3936 ) | ( n3871 & n3936 ) ;
  buffer buf_n3938( .i (n3089), .o (n3938) );
  assign n3939 = ( n3867 & n3937 ) | ( n3867 & ~n3938 ) | ( n3937 & ~n3938 ) ;
  assign n3940 = n3868 | n3939 ;
  buffer buf_n3941( .i (n3940), .o (n3941) );
  buffer buf_n3942( .i (n3941), .o (n3942) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  assign n3943 = n619 & ~n3941 ;
  assign n3944 = ( n3715 & n3942 ) | ( n3715 & ~n3943 ) | ( n3942 & ~n3943 ) ;
  assign n3945 = n3697 | n3944 ;
  assign n3946 = ~n445 & n3945 ;
  assign n3947 = n3617 | n3946 ;
  assign n3948 = n481 | n3947 ;
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  assign n3949 = ~n1105 & n2799 ;
  buffer buf_n3514( .i (n3513), .o (n3514) );
  buffer buf_n3515( .i (n3514), .o (n3515) );
  buffer buf_n3516( .i (n3515), .o (n3516) );
  buffer buf_n3517( .i (n3516), .o (n3517) );
  buffer buf_n3518( .i (n3517), .o (n3518) );
  buffer buf_n3519( .i (n3518), .o (n3519) );
  buffer buf_n3520( .i (n3519), .o (n3520) );
  buffer buf_n3521( .i (n3520), .o (n3521) );
  buffer buf_n3522( .i (n3521), .o (n3522) );
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  buffer buf_n2187( .i (n2186), .o (n2187) );
  buffer buf_n2188( .i (n2187), .o (n2188) );
  buffer buf_n2189( .i (n2188), .o (n2189) );
  buffer buf_n2190( .i (n2189), .o (n2190) );
  buffer buf_n2191( .i (n2190), .o (n2191) );
  assign n3950 = ( n2191 & n2635 ) | ( n2191 & ~n3521 ) | ( n2635 & ~n3521 ) ;
  assign n3951 = n2634 & ~n3707 ;
  buffer buf_n3952( .i (n3951), .o (n3952) );
  assign n3954 = ( n3522 & n3950 ) | ( n3522 & n3952 ) | ( n3950 & n3952 ) ;
  assign n3955 = n2501 & n3633 ;
  assign n3956 = n84 & n117 ;
  buffer buf_n3957( .i (n3956), .o (n3957) );
  buffer buf_n3958( .i (n3957), .o (n3958) );
  buffer buf_n3959( .i (n3958), .o (n3959) );
  buffer buf_n3960( .i (n3959), .o (n3960) );
  buffer buf_n3961( .i (n3960), .o (n3961) );
  buffer buf_n3962( .i (n3961), .o (n3962) );
  buffer buf_n3963( .i (n3962), .o (n3963) );
  buffer buf_n3964( .i (n3963), .o (n3964) );
  buffer buf_n3965( .i (n3964), .o (n3965) );
  buffer buf_n3966( .i (n3965), .o (n3966) );
  buffer buf_n3967( .i (n3966), .o (n3967) );
  buffer buf_n3968( .i (n3967), .o (n3968) );
  buffer buf_n3969( .i (n3968), .o (n3969) );
  buffer buf_n3970( .i (n3969), .o (n3970) );
  buffer buf_n3971( .i (n3970), .o (n3971) );
  buffer buf_n3972( .i (n3971), .o (n3972) );
  buffer buf_n3973( .i (n3972), .o (n3973) );
  assign n3974 = n71 & n3973 ;
  assign n3975 = n3955 & n3974 ;
  assign n3976 = n3954 | n3975 ;
  assign n3977 = ( n1106 & n3949 ) | ( n1106 & ~n3976 ) | ( n3949 & ~n3976 ) ;
  buffer buf_n3978( .i (n3977), .o (n3978) );
  buffer buf_n3979( .i (n3978), .o (n3979) );
  assign n3980 = ( n206 & ~n310 ) | ( n206 & n3978 ) | ( ~n310 & n3978 ) ;
  buffer buf_n2645( .i (n2644), .o (n2645) );
  buffer buf_n2646( .i (n2645), .o (n2646) );
  buffer buf_n2647( .i (n2646), .o (n2647) );
  buffer buf_n3981( .i (n3319), .o (n3981) );
  assign n3982 = ( n403 & n2795 ) | ( n403 & n3981 ) | ( n2795 & n3981 ) ;
  buffer buf_n3983( .i (n3981), .o (n3983) );
  assign n3984 = ( n2647 & n3982 ) | ( n2647 & ~n3983 ) | ( n3982 & ~n3983 ) ;
  assign n3985 = ( n398 & ~n2425 ) | ( n398 & n3852 ) | ( ~n2425 & n3852 ) ;
  buffer buf_n3986( .i (n3804), .o (n3986) );
  buffer buf_n3987( .i (n3809), .o (n3987) );
  assign n3988 = ~n3986 & n3987 ;
  assign n3989 = ( n67 & n3985 ) | ( n67 & n3988 ) | ( n3985 & n3988 ) ;
  buffer buf_n3990( .i (n3989), .o (n3990) );
  buffer buf_n3991( .i (n3990), .o (n3991) );
  assign n3992 = n2499 & ~n3990 ;
  assign n3993 = n3215 & n3971 ;
  assign n3994 = ( n3991 & n3992 ) | ( n3991 & n3993 ) | ( n3992 & n3993 ) ;
  buffer buf_n3995( .i (n3994), .o (n3995) );
  buffer buf_n3996( .i (n3995), .o (n3996) );
  assign n3997 = n3098 & n3995 ;
  assign n3998 = ( n3984 & n3996 ) | ( n3984 & n3997 ) | ( n3996 & n3997 ) ;
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n3050( .i (n3049), .o (n3050) );
  buffer buf_n3051( .i (n3050), .o (n3051) );
  buffer buf_n3052( .i (n3051), .o (n3052) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  assign n3999 = ( n1944 & n3050 ) | ( n1944 & n3518 ) | ( n3050 & n3518 ) ;
  assign n4000 = n3407 & ~n3999 ;
  assign n4001 = ( n2252 & n3052 ) | ( n2252 & ~n4000 ) | ( n3052 & ~n4000 ) ;
  assign n4002 = ~n3670 & n4001 ;
  assign n4003 = ( ~n2030 & n3709 ) | ( ~n2030 & n4002 ) | ( n3709 & n4002 ) ;
  buffer buf_n4004( .i (n4003), .o (n4004) );
  assign n4005 = ( n2710 & n3998 ) | ( n2710 & ~n4004 ) | ( n3998 & ~n4004 ) ;
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  assign n4006 = n1004 & ~n3661 ;
  assign n4007 = ~n340 & n4006 ;
  buffer buf_n4008( .i (n2799), .o (n4008) );
  assign n4009 = ( n4004 & n4007 ) | ( n4004 & n4008 ) | ( n4007 & n4008 ) ;
  assign n4010 = n4005 & ~n4009 ;
  buffer buf_n4011( .i (n2154), .o (n4011) );
  assign n4012 = n4010 | n4011 ;
  assign n4013 = ( n3979 & ~n3980 ) | ( n3979 & n4012 ) | ( ~n3980 & n4012 ) ;
  buffer buf_n4014( .i (n4013), .o (n4014) );
  buffer buf_n4015( .i (n4014), .o (n4015) );
  buffer buf_n2614( .i (n2613), .o (n2614) );
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  buffer buf_n2639( .i (n2638), .o (n2639) );
  buffer buf_n2640( .i (n2639), .o (n2640) );
  buffer buf_n2641( .i (n2640), .o (n2641) );
  assign n4016 = ( ~n276 & n2616 ) | ( ~n276 & n2641 ) | ( n2616 & n2641 ) ;
  assign n4017 = n3041 | n3509 ;
  assign n4018 = ( n788 & n3042 ) | ( n788 & n4017 ) | ( n3042 & n4017 ) ;
  buffer buf_n4019( .i (n4018), .o (n4019) );
  buffer buf_n4020( .i (n4019), .o (n4020) );
  buffer buf_n4021( .i (n4020), .o (n4021) );
  buffer buf_n4022( .i (n4021), .o (n4022) );
  buffer buf_n4023( .i (n4022), .o (n4023) );
  buffer buf_n4024( .i (n4023), .o (n4024) );
  buffer buf_n4025( .i (n4024), .o (n4025) );
  buffer buf_n4026( .i (n4025), .o (n4026) );
  buffer buf_n4027( .i (n4026), .o (n4027) );
  buffer buf_n4028( .i (n4027), .o (n4028) );
  buffer buf_n4029( .i (n4028), .o (n4029) );
  buffer buf_n4030( .i (n4029), .o (n4030) );
  buffer buf_n4031( .i (n4030), .o (n4031) );
  buffer buf_n4032( .i (n4031), .o (n4032) );
  buffer buf_n4033( .i (n2968), .o (n4033) );
  assign n4034 = n4032 & n4033 ;
  assign n4035 = ~n206 & n4034 ;
  assign n4036 = ~n2616 & n4035 ;
  buffer buf_n4037( .i (n1291), .o (n4037) );
  buffer buf_n4038( .i (n4037), .o (n4038) );
  assign n4039 = ( n4016 & ~n4036 ) | ( n4016 & n4038 ) | ( ~n4036 & n4038 ) ;
  buffer buf_n3953( .i (n3952), .o (n3953) );
  assign n4040 = n3357 & n3864 ;
  buffer buf_n4041( .i (n3027), .o (n4041) );
  assign n4042 = ~n4040 & n4041 ;
  assign n4043 = n3953 | n4042 ;
  buffer buf_n4044( .i (n4043), .o (n4044) );
  buffer buf_n4045( .i (n4044), .o (n4045) );
  buffer buf_n4046( .i (n4045), .o (n4046) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n4047( .i (n3648), .o (n4047) );
  assign n4048 = n2309 & n4047 ;
  assign n4049 = ( n978 & n4044 ) | ( n978 & n4048 ) | ( n4044 & n4048 ) ;
  assign n4050 = n3329 & ~n4049 ;
  assign n4051 = ( n108 & n4046 ) | ( n108 & ~n4050 ) | ( n4046 & ~n4050 ) ;
  assign n4052 = ( n3027 & n3633 ) | ( n3027 & ~n3670 ) | ( n3633 & ~n3670 ) ;
  buffer buf_n4053( .i (n3707), .o (n4053) );
  assign n4054 = ( ~n1897 & n3670 ) | ( ~n1897 & n4053 ) | ( n3670 & n4053 ) ;
  assign n4055 = n4052 | n4054 ;
  buffer buf_n4056( .i (n4055), .o (n4056) );
  buffer buf_n4057( .i (n4056), .o (n4057) );
  buffer buf_n4058( .i (n4057), .o (n4058) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  assign n4059 = n497 & ~n2795 ;
  buffer buf_n4060( .i (n3864), .o (n4060) );
  assign n4061 = n4059 & ~n4060 ;
  assign n4062 = n137 & n4061 ;
  assign n4063 = ( n4047 & n4056 ) | ( n4047 & n4062 ) | ( n4056 & n4062 ) ;
  assign n4064 = ~n2468 & n4063 ;
  buffer buf_n4065( .i (n2468), .o (n4065) );
  assign n4066 = ( n4058 & n4064 ) | ( n4058 & n4065 ) | ( n4064 & n4065 ) ;
  buffer buf_n4067( .i (n3875), .o (n4067) );
  assign n4068 = ( n858 & ~n3872 ) | ( n858 & n4067 ) | ( ~n3872 & n4067 ) ;
  assign n4069 = ( n856 & n859 ) | ( n856 & n4068 ) | ( n859 & n4068 ) ;
  buffer buf_n4070( .i (n4069), .o (n4070) );
  buffer buf_n4071( .i (n4070), .o (n4071) );
  buffer buf_n2901( .i (n2900), .o (n2901) );
  buffer buf_n2902( .i (n2901), .o (n2902) );
  buffer buf_n4072( .i (n2794), .o (n4072) );
  assign n4073 = n2901 & n4072 ;
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  assign n4074 = ( n805 & ~n2252 ) | ( n805 & n3643 ) | ( ~n2252 & n3643 ) ;
  assign n4075 = n3981 & n4074 ;
  assign n4076 = ( ~n2902 & n4073 ) | ( ~n2902 & n4075 ) | ( n4073 & n4075 ) ;
  buffer buf_n4077( .i (n3153), .o (n4077) );
  buffer buf_n4078( .i (n4077), .o (n4078) );
  buffer buf_n4079( .i (n4078), .o (n4079) );
  assign n4080 = ( n1943 & n2897 ) | ( n1943 & n4079 ) | ( n2897 & n4079 ) ;
  assign n4081 = n2897 & ~n3480 ;
  buffer buf_n4082( .i (n4079), .o (n4082) );
  assign n4083 = ( n4080 & n4081 ) | ( n4080 & ~n4082 ) | ( n4081 & ~n4082 ) ;
  buffer buf_n4084( .i (n4083), .o (n4084) );
  buffer buf_n4085( .i (n4084), .o (n4085) );
  buffer buf_n4086( .i (n3763), .o (n4086) );
  assign n4087 = ( n631 & n3651 ) | ( n631 & n4086 ) | ( n3651 & n4086 ) ;
  assign n4088 = n3651 & ~n3986 ;
  assign n4089 = ( ~n632 & n4087 ) | ( ~n632 & n4088 ) | ( n4087 & n4088 ) ;
  assign n4090 = ( n222 & n3780 ) | ( n222 & ~n3960 ) | ( n3780 & ~n3960 ) ;
  assign n4091 = n3961 & n4090 ;
  buffer buf_n4092( .i (n4091), .o (n4092) );
  buffer buf_n4093( .i (n4092), .o (n4093) );
  buffer buf_n4094( .i (n4093), .o (n4094) );
  buffer buf_n4095( .i (n2861), .o (n4095) );
  assign n4096 = ( n2763 & ~n4092 ) | ( n2763 & n4095 ) | ( ~n4092 & n4095 ) ;
  assign n4097 = n3738 & n4096 ;
  buffer buf_n4098( .i (n3737), .o (n4098) );
  buffer buf_n4099( .i (n4098), .o (n4099) );
  assign n4100 = ( n4094 & ~n4097 ) | ( n4094 & n4099 ) | ( ~n4097 & n4099 ) ;
  buffer buf_n4101( .i (n4100), .o (n4101) );
  buffer buf_n4102( .i (n4101), .o (n4102) );
  buffer buf_n4103( .i (n3777), .o (n4103) );
  assign n4104 = ( n4077 & ~n4101 ) | ( n4077 & n4103 ) | ( ~n4101 & n4103 ) ;
  assign n4105 = ~n908 & n1833 ;
  assign n4106 = n4077 & n4105 ;
  assign n4107 = ( n4102 & n4104 ) | ( n4102 & n4106 ) | ( n4104 & n4106 ) ;
  buffer buf_n4108( .i (n4107), .o (n4108) );
  assign n4109 = ( ~n3858 & n4089 ) | ( ~n3858 & n4108 ) | ( n4089 & n4108 ) ;
  assign n4110 = ( n1942 & ~n3651 ) | ( n1942 & n4078 ) | ( ~n3651 & n4078 ) ;
  assign n4111 = n3273 & n3803 ;
  buffer buf_n4112( .i (n3270), .o (n4112) );
  assign n4113 = ( n62 & n3449 ) | ( n62 & ~n4112 ) | ( n3449 & ~n4112 ) ;
  assign n4114 = n394 | n4112 ;
  assign n4115 = ( n3152 & ~n4113 ) | ( n3152 & n4114 ) | ( ~n4113 & n4114 ) ;
  buffer buf_n4116( .i (n393), .o (n4116) );
  buffer buf_n4117( .i (n4116), .o (n4117) );
  assign n4118 = ~n2192 & n4117 ;
  assign n4119 = n4115 & n4118 ;
  assign n4120 = ( ~n3274 & n4111 ) | ( ~n3274 & n4119 ) | ( n4111 & n4119 ) ;
  buffer buf_n4121( .i (n332), .o (n4121) );
  assign n4122 = n4120 | n4121 ;
  assign n4123 = ( n1943 & ~n4110 ) | ( n1943 & n4122 ) | ( ~n4110 & n4122 ) ;
  assign n4124 = ( n3858 & n4108 ) | ( n3858 & ~n4123 ) | ( n4108 & ~n4123 ) ;
  assign n4125 = n4109 | n4124 ;
  buffer buf_n4126( .i (n3181), .o (n4126) );
  buffer buf_n4127( .i (n4126), .o (n4127) );
  assign n4128 = ~n2275 & n4127 ;
  assign n4129 = ( ~n2276 & n3776 ) | ( ~n2276 & n4128 ) | ( n3776 & n4128 ) ;
  assign n4130 = ( ~n2892 & n3678 ) | ( ~n2892 & n4019 ) | ( n3678 & n4019 ) ;
  assign n4131 = n1825 & n3958 ;
  assign n4132 = ( n3507 & n3579 ) | ( n3507 & n4131 ) | ( n3579 & n4131 ) ;
  assign n4133 = ~n3580 & n4132 ;
  buffer buf_n4134( .i (n4133), .o (n4134) );
  buffer buf_n4135( .i (n4134), .o (n4135) );
  buffer buf_n4136( .i (n4135), .o (n4136) );
  buffer buf_n4137( .i (n122), .o (n4137) );
  buffer buf_n4138( .i (n4137), .o (n4138) );
  assign n4139 = ( n3181 & ~n4134 ) | ( n3181 & n4138 ) | ( ~n4134 & n4138 ) ;
  assign n4140 = n3270 & n4139 ;
  assign n4141 = ( n4112 & n4136 ) | ( n4112 & ~n4140 ) | ( n4136 & ~n4140 ) ;
  assign n4142 = n4130 | n4141 ;
  assign n4143 = n4129 | n4142 ;
  assign n4144 = ~n3807 & n4143 ;
  buffer buf_n4145( .i (n4144), .o (n4145) );
  buffer buf_n4146( .i (n4145), .o (n4146) );
  buffer buf_n4147( .i (n258), .o (n4147) );
  assign n4148 = ( n392 & n2890 ) | ( n392 & ~n4147 ) | ( n2890 & ~n4147 ) ;
  assign n4149 = ( n2600 & n4095 ) | ( n2600 & n4148 ) | ( n4095 & n4148 ) ;
  assign n4150 = n226 & ~n4149 ;
  buffer buf_n4151( .i (n3073), .o (n4151) );
  assign n4152 = n4150 & n4151 ;
  buffer buf_n4153( .i (n4152), .o (n4153) );
  buffer buf_n4154( .i (n4153), .o (n4154) );
  assign n4155 = n95 & n3777 ;
  assign n4156 = ( n2214 & ~n4153 ) | ( n2214 & n4155 ) | ( ~n4153 & n4155 ) ;
  assign n4157 = n4154 & n4156 ;
  assign n4158 = n4145 | n4157 ;
  assign n4159 = ( n4082 & n4146 ) | ( n4082 & n4158 ) | ( n4146 & n4158 ) ;
  buffer buf_n4160( .i (n4159), .o (n4160) );
  assign n4161 = ( ~n4084 & n4125 ) | ( ~n4084 & n4160 ) | ( n4125 & n4160 ) ;
  assign n4162 = n2794 & ~n4160 ;
  assign n4163 = ( n4085 & n4161 ) | ( n4085 & ~n4162 ) | ( n4161 & ~n4162 ) ;
  buffer buf_n4164( .i (n4163), .o (n4164) );
  assign n4165 = ( n4070 & n4076 ) | ( n4070 & ~n4164 ) | ( n4076 & ~n4164 ) ;
  buffer buf_n4166( .i (n3026), .o (n4166) );
  buffer buf_n4167( .i (n4166), .o (n4167) );
  assign n4168 = ~n4164 & n4167 ;
  assign n4169 = ( ~n4071 & n4165 ) | ( ~n4071 & n4168 ) | ( n4165 & n4168 ) ;
  buffer buf_n4170( .i (n4169), .o (n4170) );
  buffer buf_n4171( .i (n4170), .o (n4171) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  assign n4172 = n1108 & n4170 ;
  assign n4173 = ( n4066 & n4171 ) | ( n4066 & n4172 ) | ( n4171 & n4172 ) ;
  assign n4174 = n4051 & n4173 ;
  assign n4175 = ( ~n4014 & n4039 ) | ( ~n4014 & n4174 ) | ( n4039 & n4174 ) ;
  assign n4176 = n4015 & n4175 ;
  assign n4177 = n446 | n4176 ;
  assign n4178 = n481 & n4177 ;
  assign n4179 = n3948 & ~n4178 ;
  assign y0 = n966 ;
  assign y1 = n1200 ;
  assign y2 = n1411 ;
  assign y3 = n1658 ;
  assign y4 = n1935 ;
  assign y5 = n2098 ;
  assign y6 = n2168 ;
  assign y7 = n2334 ;
  assign y8 = ~n2498 ;
  assign y9 = ~n2825 ;
  assign y10 = ~n2991 ;
  assign y11 = ~n3117 ;
  assign y12 = ~n3342 ;
  assign y13 = n4179 ;
endmodule
