module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , y0 , y1 , y2 , y3 , y4 , y5 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 ;
  output y0 , y1 , y2 , y3 , y4 , y5 ;
  wire n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 ;
  buffer buf_n56( .i (x2), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n43( .i (x1), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n70( .i (x3), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  assign n240 = ( n53 & n66 ) | ( n53 & n80 ) | ( n66 & n80 ) ;
  buffer buf_n81( .i (x4), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  assign n241 = n53 & ~n91 ;
  assign n242 = ( ~n67 & n240 ) | ( ~n67 & n241 ) | ( n240 & n241 ) ;
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n28( .i (x0), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  assign n245 = ( ~n52 & n65 ) | ( ~n52 & n79 ) | ( n65 & n79 ) ;
  assign n246 = ~n52 & n90 ;
  assign n247 = ( ~n80 & n245 ) | ( ~n80 & n246 ) | ( n245 & n246 ) ;
  buffer buf_n116( .i (x8), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n112( .i (x7), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  assign n248 = n115 & ~n119 ;
  buffer buf_n99( .i (x6), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  assign n249 = ~n101 & n114 ;
  assign n250 = n119 & n249 ;
  assign n251 = ( n120 & n248 ) | ( n120 & ~n250 ) | ( n248 & ~n250 ) ;
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n92( .i (x5), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  assign n260 = n98 | n252 ;
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n140( .i (x11), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n121( .i (x9), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n128( .i (x10), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  assign n261 = n124 & ~n131 ;
  assign n262 = ( n103 & ~n144 ) | ( n103 & n261 ) | ( ~n144 & n261 ) ;
  assign n263 = ~n104 & n262 ;
  buffer buf_n151( .i (x12), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  assign n264 = n114 | n118 ;
  buffer buf_n265( .i (n264), .o (n265) );
  assign n272 = n155 & n265 ;
  assign n273 = n104 & n272 ;
  assign n274 = n263 | n273 ;
  assign n275 = ( ~n253 & n260 ) | ( ~n253 & n274 ) | ( n260 & n274 ) ;
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  assign n279 = n38 & n277 ;
  assign n280 = ( n247 & n278 ) | ( n247 & n279 ) | ( n278 & n279 ) ;
  buffer buf_n281( .i (n280), .o (n281) );
  assign n282 = ( n41 & n243 ) | ( n41 & ~n281 ) | ( n243 & ~n281 ) ;
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n158( .i (x13), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (x14), .o (n164) );
  assign n283 = ~n128 & n164 ;
  assign n284 = ~n141 & n283 ;
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  assign n288 = ( n115 & n119 ) | ( n115 & n285 ) | ( n119 & n285 ) ;
  assign n289 = n162 & ~n288 ;
  assign n290 = ( n163 & n287 ) | ( n163 & ~n289 ) | ( n287 & ~n289 ) ;
  assign n291 = ~n113 & n159 ;
  assign n292 = ~n118 & n291 ;
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = ( ~n105 & n290 ) | ( ~n105 & n295 ) | ( n290 & n295 ) ;
  buffer buf_n169( .i (x15), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  assign n297 = n173 & n265 ;
  assign n298 = ( n104 & n294 ) | ( n104 & n297 ) | ( n294 & n297 ) ;
  buffer buf_n299( .i (n298), .o (n299) );
  assign n300 = n296 | n299 ;
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  assign n306 = n281 | n305 ;
  assign n307 = ( n244 & ~n282 ) | ( n244 & n306 ) | ( ~n282 & n306 ) ;
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n182( .i (x17), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n174( .i (x16), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n198( .i (x22), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n192( .i (x20), .o (n192) );
  buffer buf_n194( .i (x21), .o (n194) );
  assign n311 = ( ~n192 & n194 ) | ( ~n192 & n198 ) | ( n194 & n198 ) ;
  buffer buf_n189( .i (x19), .o (n189) );
  assign n312 = n189 & ~n192 ;
  assign n313 = ( ~n199 & n311 ) | ( ~n199 & n312 ) | ( n311 & n312 ) ;
  assign n314 = ( n176 & ~n184 ) | ( n176 & n313 ) | ( ~n184 & n313 ) ;
  buffer buf_n187( .i (x18), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  assign n315 = ~n175 & n188 ;
  buffer buf_n316( .i (n315), .o (n316) );
  assign n317 = ( n185 & n314 ) | ( n185 & ~n316 ) | ( n314 & ~n316 ) ;
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  assign n324 = n277 & n323 ;
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n193( .i (n192), .o (n193) );
  assign n327 = ( n193 & n195 ) | ( n193 & n199 ) | ( n195 & n199 ) ;
  buffer buf_n190( .i (n189), .o (n190) );
  assign n328 = ~n190 & n193 ;
  assign n329 = ( ~n196 & n327 ) | ( ~n196 & n328 ) | ( n327 & n328 ) ;
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n332 = ( n178 & n186 ) | ( n178 & n330 ) | ( n186 & n330 ) ;
  assign n333 = n175 & ~n188 ;
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  assign n337 = ( ~n331 & n332 ) | ( ~n331 & n336 ) | ( n332 & n336 ) ;
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  assign n344 = ~n325 & n343 ;
  assign n345 = ( n305 & n326 ) | ( n305 & ~n344 ) | ( n326 & ~n344 ) ;
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  assign n350 = n44 & n71 ;
  assign n351 = ( ~n30 & n58 ) | ( ~n30 & n350 ) | ( n58 & n350 ) ;
  assign n352 = n31 & n351 ;
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n200( .i (x23), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  assign n356 = n176 & n202 ;
  buffer buf_n357( .i (n356), .o (n357) );
  assign n358 = n162 & n357 ;
  assign n359 = ( n86 & ~n353 ) | ( n86 & n358 ) | ( ~n353 & n358 ) ;
  assign n360 = n354 & n359 ;
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  assign n368 = n44 | n71 ;
  assign n369 = ( ~n30 & n58 ) | ( ~n30 & n368 ) | ( n58 & n368 ) ;
  assign n370 = n31 | n369 ;
  buffer buf_n371( .i (n370), .o (n371) );
  assign n372 = n176 | n202 ;
  buffer buf_n373( .i (n372), .o (n373) );
  assign n374 = n96 & ~n373 ;
  assign n375 = ( n86 & ~n371 ) | ( n86 & n374 ) | ( ~n371 & n374 ) ;
  assign n376 = ~n87 & n375 ;
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  assign n383 = n173 & n357 ;
  assign n384 = n86 & n383 ;
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n355( .i (n354), .o (n355) );
  assign n387 = ( n268 & n355 ) | ( n268 & ~n385 ) | ( n355 & ~n385 ) ;
  assign n388 = n155 & ~n373 ;
  buffer buf_n389( .i (n85), .o (n389) );
  assign n390 = ( ~n371 & n388 ) | ( ~n371 & n389 ) | ( n388 & n389 ) ;
  assign n391 = ~n87 & n390 ;
  assign n392 = n268 & n391 ;
  assign n393 = ( n386 & n387 ) | ( n386 & n392 ) | ( n387 & n392 ) ;
  assign n394 = n108 & ~n393 ;
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  assign n396 = n168 & n357 ;
  assign n397 = n389 & n396 ;
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  assign n400 = ( n147 & ~n355 ) | ( n147 & n398 ) | ( ~n355 & n398 ) ;
  buffer buf_n125( .i (n124), .o (n125) );
  assign n401 = n125 & ~n373 ;
  assign n402 = ( ~n371 & n389 ) | ( ~n371 & n401 ) | ( n389 & n401 ) ;
  assign n403 = ~n87 & n402 ;
  assign n404 = ~n147 & n403 ;
  assign n405 = ( n399 & ~n400 ) | ( n399 & n404 ) | ( ~n400 & n404 ) ;
  assign n406 = ~n137 & n405 ;
  assign n407 = n109 | n406 ;
  assign n408 = ~n395 & n407 ;
  buffer buf_n409( .i (n408), .o (n409) );
  assign n410 = ( ~n366 & n382 ) | ( ~n366 & n409 ) | ( n382 & n409 ) ;
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  assign n411 = n259 & ~n409 ;
  assign n412 = ( n367 & n410 ) | ( n367 & ~n411 ) | ( n410 & ~n411 ) ;
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  assign n416 = n71 & n201 ;
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  assign n424 = ( n90 & ~n301 ) | ( n90 & n423 ) | ( ~n301 & n423 ) ;
  assign n425 = n302 & n424 ;
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  assign n428 = n28 & n56 ;
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  assign n440 = ( n55 & ~n426 ) | ( n55 & n439 ) | ( ~n426 & n439 ) ;
  assign n441 = n427 & n440 ;
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n446( .i (n70), .o (n446) );
  assign n447 = n201 | n446 ;
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  assign n456 = ( n91 & n277 ) | ( n91 & n455 ) | ( n277 & n455 ) ;
  assign n457 = n278 & ~n456 ;
  assign n458 = ~n55 & n457 ;
  assign n459 = ( n41 & ~n69 ) | ( n41 & n458 ) | ( ~n69 & n458 ) ;
  assign n460 = ~n42 & n459 ;
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n203( .i (x24), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  assign n464 = n45 & n429 ;
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  assign n467 = n82 & n446 ;
  buffer buf_n468( .i (n175), .o (n468) );
  assign n469 = n467 & n468 ;
  buffer buf_n470( .i (n469), .o (n470) );
  assign n471 = ( n162 & ~n465 ) | ( n162 & n470 ) | ( ~n465 & n470 ) ;
  assign n472 = n466 & n471 ;
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n191( .i (n190), .o (n191) );
  assign n475 = n188 & n193 ;
  assign n476 = ( ~n184 & n191 ) | ( ~n184 & n475 ) | ( n191 & n475 ) ;
  assign n477 = n185 & n476 ;
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n238( .i (x26), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  assign n478 = n199 & n239 ;
  assign n479 = ( ~n196 & n202 ) | ( ~n196 & n478 ) | ( n202 & n478 ) ;
  assign n480 = n197 & n479 ;
  assign n481 = n477 & n480 ;
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  assign n484 = ( n253 & n473 ) | ( n253 & ~n483 ) | ( n473 & ~n483 ) ;
  assign n485 = n188 | n193 ;
  assign n486 = ( ~n184 & n191 ) | ( ~n184 & n485 ) | ( n191 & n485 ) ;
  assign n487 = n185 | n486 ;
  assign n488 = n199 | n239 ;
  assign n489 = ( ~n196 & n202 ) | ( ~n196 & n488 ) | ( n202 & n488 ) ;
  assign n490 = n197 | n489 ;
  assign n491 = n487 | n490 ;
  buffer buf_n492( .i (n491), .o (n492) );
  assign n496 = n82 | n446 ;
  buffer buf_n497( .i (n496), .o (n497) );
  assign n499 = n177 | n497 ;
  assign n500 = n96 & ~n499 ;
  assign n501 = n29 | n57 ;
  assign n502 = n45 | n501 ;
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  assign n505 = n500 & ~n504 ;
  assign n506 = ~n492 & n505 ;
  assign n507 = ~n253 & n506 ;
  assign n508 = ( n474 & ~n484 ) | ( n474 & n507 ) | ( ~n484 & n507 ) ;
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  assign n514 = ( n168 & ~n465 ) | ( n168 & n470 ) | ( ~n465 & n470 ) ;
  assign n515 = n466 & n514 ;
  assign n516 = n482 & n515 ;
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n498( .i (n497), .o (n498) );
  assign n519 = n498 | n503 ;
  buffer buf_n520( .i (n519), .o (n520) );
  assign n521 = ( n127 & n180 ) | ( n127 & ~n520 ) | ( n180 & ~n520 ) ;
  assign n522 = ~n181 & n521 ;
  assign n523 = n517 | n522 ;
  assign n524 = ( ~n495 & n518 ) | ( ~n495 & n523 ) | ( n518 & n523 ) ;
  assign n525 = ~n150 & n524 ;
  assign n526 = ~n139 & n525 ;
  assign n527 = n111 | n526 ;
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  assign n528 = ( n173 & ~n465 ) | ( n173 & n470 ) | ( ~n465 & n470 ) ;
  assign n529 = n466 & n528 ;
  assign n530 = n482 & n529 ;
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  assign n533 = ( n157 & n180 ) | ( n157 & ~n520 ) | ( n180 & ~n520 ) ;
  assign n534 = ~n181 & n533 ;
  assign n535 = n531 | n534 ;
  assign n536 = ( ~n495 & n532 ) | ( ~n495 & n535 ) | ( n532 & n535 ) ;
  assign n537 = n271 & n536 ;
  assign n538 = n110 & ~n537 ;
  buffer buf_n539( .i (n538), .o (n539) );
  assign n540 = n527 & ~n539 ;
  assign n541 = n513 | n540 ;
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n221( .i (x25), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  assign n544 = ~n237 & n542 ;
  assign n545 = ( ~n220 & n543 ) | ( ~n220 & n544 ) | ( n543 & n544 ) ;
  assign y0 = n310 ;
  assign y1 = n349 ;
  assign y2 = n415 ;
  assign y3 = n445 ;
  assign y4 = n463 ;
  assign y5 = n545 ;
endmodule
