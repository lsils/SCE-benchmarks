module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 ;
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n26( .i (x2), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n35( .i (x3), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  assign n76 = n27 | n36 ;
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n15( .i (x1), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  assign n81 = n3 | n16 ;
  buffer buf_n82( .i (n81), .o (n82) );
  assign n83 = n77 | n82 ;
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n43( .i (x4), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n52( .i (x5), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n60( .i (x6), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  assign n88 = n54 & n62 ;
  buffer buf_n89( .i (n88), .o (n89) );
  assign n94 = n47 & n89 ;
  buffer buf_n95( .i (n94), .o (n95) );
  assign n96 = n85 | n95 ;
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  assign n98 = ~n29 & n46 ;
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n68( .i (x7), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  assign n101 = n62 & n70 ;
  buffer buf_n102( .i (n101), .o (n102) );
  assign n103 = n56 | n102 ;
  buffer buf_n104( .i (n103), .o (n104) );
  assign n105 = n100 & n104 ;
  buffer buf_n106( .i (n105), .o (n106) );
  assign n107 = n97 | n106 ;
  assign n108 = ~n11 & n107 ;
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n37( .i (n36), .o (n37) );
  assign n110 = n28 & ~n37 ;
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  assign n115 = n60 | n68 ;
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  assign n120 = n44 | n53 ;
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  assign n124 = ( n47 & n118 ) | ( n47 & n122 ) | ( n118 & n122 ) ;
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  assign n128 = n114 & ~n126 ;
  buffer buf_n129( .i (n128), .o (n129) );
  assign n130 = ~n27 & n36 ;
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  assign n137 = n106 | n136 ;
  assign n138 = n129 | n137 ;
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  assign n139 = ~n11 & n24 ;
  assign n140 = ( n12 & n138 ) | ( n12 & ~n139 ) | ( n138 & ~n139 ) ;
  buffer buf_n63( .i (n62), .o (n63) );
  assign n141 = n55 | n63 ;
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  assign n145 = ~n8 & n143 ;
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  assign n148 = n49 | n80 ;
  buffer buf_n149( .i (n148), .o (n149) );
  assign n150 = n37 & n45 ;
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  assign n156 = n149 & ~n155 ;
  assign n157 = n147 & ~n156 ;
  assign n158 = n100 & ~n104 ;
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  assign n160 = n91 & n134 ;
  assign n161 = n22 | n160 ;
  assign n162 = n159 | n161 ;
  assign n163 = n129 | n162 ;
  assign n164 = ( ~n12 & n157 ) | ( ~n12 & n163 ) | ( n157 & n163 ) ;
  assign n165 = n44 & n53 ;
  buffer buf_n166( .i (n165), .o (n166) );
  assign n169 = n117 & n166 ;
  buffer buf_n170( .i (n169), .o (n170) );
  assign n172 = n18 & ~n77 ;
  buffer buf_n173( .i (n172), .o (n173) );
  assign n175 = ~n170 & n173 ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n177 = n9 | n176 ;
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  assign n180 = n55 & n117 ;
  buffer buf_n181( .i (n180), .o (n181) );
  assign n184 = n29 & ~n46 ;
  buffer buf_n185( .i (n184), .o (n185) );
  assign n186 = ~n181 & n185 ;
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n38( .i (n37), .o (n38) );
  assign n188 = n38 & ~n46 ;
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n30( .i (n29), .o (n30) );
  assign n191 = ~n30 & n89 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = n190 & ~n192 ;
  assign n194 = n187 | n193 ;
  buffer buf_n195( .i (n194), .o (n195) );
  assign n196 = ~n178 & n195 ;
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  assign n197 = ( n31 & ~n40 ) | ( n31 & n142 ) | ( ~n40 & n142 ) ;
  assign n198 = ( ~n31 & n40 ) | ( ~n31 & n142 ) | ( n40 & n142 ) ;
  assign n199 = ( ~n171 & n197 ) | ( ~n171 & n198 ) | ( n197 & n198 ) ;
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  assign n202 = ~n80 & n91 ;
  assign n203 = ~n43 & n68 ;
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  assign n210 = n202 & n209 ;
  assign n211 = n62 & ~n70 ;
  buffer buf_n212( .i (n211), .o (n212) );
  assign n213 = n19 | n212 ;
  buffer buf_n214( .i (n45), .o (n214) );
  assign n215 = ~n55 & n214 ;
  assign n216 = ~n78 & n215 ;
  assign n217 = ( n20 & n213 ) | ( n20 & n216 ) | ( n213 & n216 ) ;
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  assign n221 = n210 | n219 ;
  assign n222 = n201 & ~n221 ;
  assign n223 = ( n179 & ~n196 ) | ( n179 & n222 ) | ( ~n196 & n222 ) ;
  assign n224 = ~n38 & n214 ;
  buffer buf_n225( .i (n224), .o (n225) );
  assign n227 = ~n7 & n225 ;
  assign n228 = n17 & ~n28 ;
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  assign n233 = ~n90 & n230 ;
  assign n234 = ( n8 & ~n227 ) | ( n8 & n233 ) | ( ~n227 & n233 ) ;
  buffer buf_n235( .i (n234), .o (n235) );
  assign n236 = ~n146 & n235 ;
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  assign n237 = ~n176 & n232 ;
  assign n238 = n200 & n237 ;
  assign n239 = n236 | n238 ;
  buffer buf_n41( .i (n40), .o (n41) );
  assign n240 = n102 | n122 ;
  assign n241 = n30 | n118 ;
  assign n242 = n240 & n241 ;
  assign n243 = n41 & ~n242 ;
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  assign n244 = ( n57 & n112 ) | ( n57 & n168 ) | ( n112 & n168 ) ;
  buffer buf_n119( .i (n118), .o (n119) );
  assign n245 = ~n119 & n225 ;
  assign n246 = n244 | n245 ;
  assign n247 = n243 | n246 ;
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  assign n248 = n31 & n152 ;
  assign n249 = ( n66 & ~n80 ) | ( n66 & n248 ) | ( ~n80 & n248 ) ;
  assign n250 = ~n61 & n69 ;
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  assign n254 = ~n28 & n54 ;
  buffer buf_n255( .i (n254), .o (n255) );
  assign n256 = ~n252 & n255 ;
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  assign n259 = n249 | n258 ;
  assign n260 = n247 | n259 ;
  assign n261 = n111 | n132 ;
  assign n262 = n56 & ~n118 ;
  assign n263 = n261 & n262 ;
  assign n264 = n77 | n205 ;
  assign n265 = n89 & ~n264 ;
  buffer buf_n266( .i (n265), .o (n266) );
  assign n269 = n263 | n266 ;
  buffer buf_n270( .i (n269), .o (n270) );
  assign n271 = n219 | n270 ;
  assign n272 = n260 & ~n271 ;
  assign n273 = n239 | n272 ;
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n123( .i (n122), .o (n123) );
  assign n274 = n119 | n123 ;
  buffer buf_n275( .i (n274), .o (n275) );
  assign n276 = n86 | n275 ;
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n127( .i (n126), .o (n127) );
  assign n280 = n87 | n127 ;
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n144( .i (n143), .o (n144) );
  assign n283 = ~n126 & n144 ;
  assign n284 = n97 | n283 ;
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n30), .o (n287) );
  assign n288 = n20 | n287 ;
  assign n289 = n8 | n288 ;
  buffer buf_n226( .i (n225), .o (n226) );
  assign n290 = ~n91 & n226 ;
  assign n291 = n289 | n290 ;
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  assign n292 = ~n154 & n183 ;
  assign n293 = n54 | n116 ;
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n298( .i (n61), .o (n298) );
  assign n299 = ~n204 & n298 ;
  buffer buf_n300( .i (n299), .o (n300) );
  assign n302 = n294 & ~n300 ;
  assign n303 = ~n84 & n302 ;
  buffer buf_n304( .i (n303), .o (n304) );
  assign n305 = n183 | n304 ;
  assign n306 = ( n291 & ~n292 ) | ( n291 & n305 ) | ( ~n292 & n305 ) ;
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  assign n309 = n27 & n36 ;
  buffer buf_n310( .i (n309), .o (n310) );
  assign n311 = n82 | n310 ;
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n58( .i (n57), .o (n58) );
  assign n315 = n58 & n190 ;
  assign n316 = n314 | n315 ;
  buffer buf_n50( .i (n49), .o (n50) );
  assign n317 = ~n50 & n258 ;
  assign n318 = n316 | n317 ;
  buffer buf_n301( .i (n300), .o (n301) );
  assign n319 = ~n84 & n301 ;
  buffer buf_n320( .i (n319), .o (n320) );
  assign n321 = ~n218 & n320 ;
  assign n322 = ~n270 & n321 ;
  assign n323 = n318 | n322 ;
  buffer buf_n324( .i (n53), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  assign n326 = ~n5 & n325 ;
  assign n327 = ( n6 & n132 ) | ( n6 & ~n326 ) | ( n132 & ~n326 ) ;
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n29), .o (n329) );
  assign n330 = n151 & ~n329 ;
  assign n331 = ~n119 & n330 ;
  assign n332 = n328 | n331 ;
  assign n333 = n304 | n332 ;
  buffer buf_n334( .i (n333), .o (n334) );
  assign n335 = n99 | n152 ;
  assign n336 = ( n104 & n153 ) | ( n104 & n335 ) | ( n153 & n335 ) ;
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  assign n339 = n113 & n125 ;
  buffer buf_n340( .i (n339), .o (n340) );
  assign n342 = n337 & n340 ;
  assign n343 = ( n334 & n338 ) | ( n334 & n342 ) | ( n338 & n342 ) ;
  assign n344 = n323 | n343 ;
  buffer buf_n341( .i (n340), .o (n341) );
  assign n345 = n334 | n341 ;
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  assign n346 = n93 | n149 ;
  assign n347 = n220 & n346 ;
  assign n348 = n345 | n347 ;
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  assign n349 = ~n192 & n296 ;
  assign n350 = n50 & ~n349 ;
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n297( .i (n296), .o (n297) );
  assign n351 = n32 & n190 ;
  assign n352 = ( n33 & ~n297 ) | ( n33 & n351 ) | ( ~n297 & n351 ) ;
  assign n353 = n350 | n352 ;
  assign n354 = n39 | n47 ;
  assign n355 = ( n40 & n142 ) | ( n40 & n354 ) | ( n142 & n354 ) ;
  assign n356 = n257 | n355 ;
  assign n357 = n187 | n356 ;
  assign n358 = n23 | n357 ;
  assign n359 = ( n24 & ~n353 ) | ( n24 & n358 ) | ( ~n353 & n358 ) ;
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n174( .i (n173), .o (n174) );
  assign n360 = n48 | n90 ;
  assign n361 = n174 & n360 ;
  assign n362 = ~n45 & n324 ;
  assign n363 = ( ~n63 & n251 ) | ( ~n63 & n362 ) | ( n251 & n362 ) ;
  buffer buf_n364( .i (n363), .o (n364) );
  assign n365 = n133 & n364 ;
  buffer buf_n366( .i (n365), .o (n366) );
  assign n367 = n361 | n366 ;
  assign n368 = n268 | n367 ;
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  assign n369 = n72 & n167 ;
  assign n370 = n18 & n131 ;
  buffer buf_n371( .i (n370), .o (n371) );
  assign n372 = ~n369 & n371 ;
  buffer buf_n373( .i (n372), .o (n373) );
  assign n375 = ~n71 & n166 ;
  assign n376 = ~n78 & n375 ;
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  assign n379 = n373 | n378 ;
  assign n380 = ~n10 & n379 ;
  assign n381 = ( ~n11 & n368 ) | ( ~n11 & n380 ) | ( n368 & n380 ) ;
  assign n382 = ( n12 & n359 ) | ( n12 & ~n381 ) | ( n359 & ~n381 ) ;
  assign n383 = n132 & n212 ;
  assign n384 = ~n121 & n310 ;
  assign n385 = n19 | n384 ;
  assign n386 = n383 | n385 ;
  assign n387 = n377 | n386 ;
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  assign n390 = ~n72 & n329 ;
  assign n391 = ( n225 & n287 ) | ( n225 & n390 ) | ( n287 & n390 ) ;
  buffer buf_n253( .i (n252), .o (n253) );
  assign n392 = ( n65 & n168 ) | ( n65 & ~n253 ) | ( n168 & ~n253 ) ;
  assign n393 = n391 & ~n392 ;
  assign n394 = n131 & ~n325 ;
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  assign n397 = n48 & n364 ;
  assign n398 = n396 & n397 ;
  assign n399 = n393 | n398 ;
  assign n400 = ~n388 & n399 ;
  assign n401 = n56 & n72 ;
  assign n402 = n189 & n401 ;
  assign n403 = n39 | n102 ;
  assign n404 = n185 & n403 ;
  assign n405 = n402 | n404 ;
  buffer buf_n406( .i (n71), .o (n406) );
  assign n407 = n122 & n406 ;
  assign n408 = n64 & ~n329 ;
  assign n409 = ~n407 & n408 ;
  assign n410 = n95 | n409 ;
  assign n411 = n405 | n410 ;
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  assign n412 = n100 & ~n396 ;
  assign n413 = ~n123 & n133 ;
  buffer buf_n414( .i (n413), .o (n414) );
  assign n415 = ( ~n75 & n412 ) | ( ~n75 & n414 ) | ( n412 & n414 ) ;
  assign n416 = n411 | n415 ;
  assign n417 = ( ~n389 & n400 ) | ( ~n389 & n416 ) | ( n400 & n416 ) ;
  buffer buf_n374( .i (n373), .o (n374) );
  assign n418 = n235 | n374 ;
  buffer buf_n419( .i (n418), .o (n419) );
  assign n420 = n417 | n419 ;
  assign y0 = ~n13 ;
  assign y1 = ~n13 ;
  assign y2 = ~n13 ;
  assign y3 = n109 ;
  assign y4 = ~n140 ;
  assign y5 = n164 ;
  assign y6 = ~n223 ;
  assign y7 = ~n273 ;
  assign y8 = ~n279 ;
  assign y9 = ~n282 ;
  assign y10 = ~n286 ;
  assign y11 = ~n308 ;
  assign y12 = ~n344 ;
  assign y13 = ~n348 ;
  assign y14 = ~n382 ;
  assign y15 = ~n420 ;
endmodule
