module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 ;
  buffer buf_n351( .i (x10), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n319( .i (x9), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n384( .i (x11), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  assign n486 = ~n326 & n391 ;
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  assign n502 = n366 | n493 ;
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n249( .i (x7), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n417( .i (x12), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n451( .i (x13), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  assign n522 = ~n424 & n458 ;
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n79( .i (x2), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n285( .i (x8), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  assign n541 = n296 & n395 ;
  buffer buf_n542( .i (n541), .o (n542) );
  assign n561 = n332 & n542 ;
  buffer buf_n562( .i (n561), .o (n562) );
  assign n573 = n366 & ~n562 ;
  assign n574 = n332 | n364 ;
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  assign n586 = ( ~n367 & n573 ) | ( ~n367 & n576 ) | ( n573 & n576 ) ;
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n112( .i (x3), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n179( .i (x5), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n599 = n119 & n186 ;
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  assign n621 = ( n100 & n590 ) | ( n100 & n612 ) | ( n590 & n612 ) ;
  buffer buf_n145( .i (x4), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  assign n622 = n152 & ~n186 ;
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  assign n644 = ( ~n100 & n590 ) | ( ~n100 & n635 ) | ( n590 & n635 ) ;
  assign n645 = n621 & n644 ;
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n214( .i (x6), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  assign n648 = n98 & ~n198 ;
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  assign n649 = ( n97 & n163 ) | ( n97 & n197 ) | ( n163 & n197 ) ;
  buffer buf_n650( .i (n649), .o (n650) );
  assign n655 = ( n234 & n648 ) | ( n234 & n650 ) | ( n648 & n650 ) ;
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n591( .i (n590), .o (n591) );
  assign n658 = ( n134 & ~n591 ) | ( n134 & n656 ) | ( ~n591 & n656 ) ;
  assign n659 = n130 | n232 ;
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  assign n662 = ~n158 & n192 ;
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  assign n675 = ( n133 & ~n661 ) | ( n133 & n669 ) | ( ~n661 & n669 ) ;
  assign n676 = n591 & n675 ;
  assign n677 = ( n657 & ~n658 ) | ( n657 & n676 ) | ( ~n658 & n676 ) ;
  assign n678 = ~n646 & n677 ;
  assign n679 = ( n539 & n647 ) | ( n539 & n678 ) | ( n647 & n678 ) ;
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n48( .i (x1), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  assign n682 = ( n75 & n276 ) | ( n75 & ~n680 ) | ( n276 & ~n680 ) ;
  assign n683 = ~n294 & n393 ;
  buffer buf_n684( .i (n683), .o (n684) );
  assign n689 = n328 | n393 ;
  buffer buf_n690( .i (n689), .o (n690) );
  assign n704 = ( ~n395 & n684 ) | ( ~n395 & n690 ) | ( n684 & n690 ) ;
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  assign n714 = ( n301 & n367 ) | ( n301 & ~n400 ) | ( n367 & ~n400 ) ;
  assign n715 = n336 & ~n714 ;
  buffer buf_n401( .i (n400), .o (n401) );
  assign n716 = ( ~n288 & n322 ) | ( ~n288 & n387 ) | ( n322 & n387 ) ;
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  assign n726 = n364 & ~n725 ;
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  assign n742 = ( ~n264 & n300 ) | ( ~n264 & n727 ) | ( n300 & n727 ) ;
  assign n743 = n400 & ~n742 ;
  assign n744 = ( n401 & n729 ) | ( n401 & ~n743 ) | ( n729 & ~n743 ) ;
  assign n745 = n715 | n744 ;
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  assign n757 = n269 | n746 ;
  assign n758 = ( n713 & n747 ) | ( n713 & n757 ) | ( n747 & n757 ) ;
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  assign n767 = n268 & ~n403 ;
  assign n768 = n371 & n767 ;
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  assign n771 = n236 | n769 ;
  assign n772 = ( n759 & n770 ) | ( n759 & n771 ) | ( n770 & n771 ) ;
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n15( .i (x0), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  assign n775 = n37 | n167 ;
  assign n776 = n124 | n191 ;
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  assign n786 = ( n37 & ~n167 ) | ( n37 & n785 ) | ( ~n167 & n785 ) ;
  assign n787 = n122 & ~n155 ;
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n199( .i (n198), .o (n199) );
  assign n801 = n99 | n199 ;
  assign n802 = n130 | n163 ;
  buffer buf_n803( .i (n802), .o (n803) );
  assign n806 = ( ~n132 & n796 ) | ( ~n132 & n803 ) | ( n796 & n803 ) ;
  assign n807 = ( n797 & n801 ) | ( n797 & n806 ) | ( n801 & n806 ) ;
  assign n808 = n37 & n807 ;
  assign n809 = ( n775 & ~n786 ) | ( n775 & n808 ) | ( ~n786 & n808 ) ;
  assign n810 = n441 & n809 ;
  assign n811 = ( n476 & n773 ) | ( n476 & ~n810 ) | ( n773 & ~n810 ) ;
  assign n812 = n774 & ~n811 ;
  assign n813 = n75 & n812 ;
  assign n814 = ( n681 & n682 ) | ( n681 & n813 ) | ( n682 & n813 ) ;
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  assign n818 = ( n136 & n203 ) | ( n136 & n800 ) | ( n203 & n800 ) ;
  assign n819 = ( ~n136 & n203 ) | ( ~n136 & n800 ) | ( n203 & n800 ) ;
  assign n820 = ( n137 & ~n818 ) | ( n137 & n819 ) | ( ~n818 & n819 ) ;
  buffer buf_n821( .i (n820), .o (n821) );
  assign n825 = ~n478 & n821 ;
  assign n826 = ( n445 & n597 ) | ( n445 & ~n825 ) | ( n597 & ~n825 ) ;
  assign n827 = n598 & ~n826 ;
  assign n828 = ( n109 & n815 ) | ( n109 & n827 ) | ( n815 & n827 ) ;
  assign n829 = n280 & ~n828 ;
  assign n830 = ( n281 & n817 ) | ( n281 & ~n829 ) | ( n817 & ~n829 ) ;
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  assign n833 = n309 & ~n441 ;
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  assign n838 = ( n480 & n823 ) | ( n480 & ~n837 ) | ( n823 & ~n837 ) ;
  assign n839 = n824 & ~n838 ;
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n76( .i (n75), .o (n76) );
  assign n842 = ( ~n120 & n153 ) | ( ~n120 & n222 ) | ( n153 & n222 ) ;
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  assign n857 = ~n165 & n853 ;
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  assign n860 = ( ~n202 & n856 ) | ( ~n202 & n859 ) | ( n856 & n859 ) ;
  assign n861 = n129 & ~n793 ;
  assign n862 = n97 & n861 ;
  assign n863 = ( n164 & n795 ) | ( n164 & ~n862 ) | ( n795 & ~n862 ) ;
  assign n864 = ( n234 & n796 ) | ( n234 & n863 ) | ( n796 & n863 ) ;
  assign n865 = n200 & n864 ;
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  assign n868 = n102 | n866 ;
  assign n869 = ( n860 & n867 ) | ( n860 & n868 ) | ( n867 & n868 ) ;
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n540( .i (n539), .o (n540) );
  assign n872 = ( n311 & n540 ) | ( n311 & ~n870 ) | ( n540 & ~n870 ) ;
  assign n873 = n871 & n872 ;
  assign n874 = ( n76 & n277 ) | ( n76 & n873 ) | ( n277 & n873 ) ;
  assign n875 = n32 & n129 ;
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  assign n883 = n260 & ~n462 ;
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  assign n891 = ( n436 & n876 ) | ( n436 & n890 ) | ( n876 & n890 ) ;
  assign n892 = ~n877 & n891 ;
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  assign n896 = n302 & n531 ;
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  assign n901 = n186 | n256 ;
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  assign n921 = ( n893 & n900 ) | ( n893 & ~n915 ) | ( n900 & ~n915 ) ;
  assign n922 = n102 & ~n921 ;
  assign n923 = ( n103 & n895 ) | ( n103 & ~n922 ) | ( n895 & ~n922 ) ;
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  assign n926 = ( ~n171 & n240 ) | ( ~n171 & n924 ) | ( n240 & n924 ) ;
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  assign n927 = n430 & n884 ;
  assign n928 = ~n159 & n927 ;
  buffer buf_n929( .i (n928), .o (n929) );
  assign n937 = n31 & n929 ;
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  assign n941 = ( n197 & ~n267 ) | ( n197 & n938 ) | ( ~n267 & n938 ) ;
  assign n942 = n897 & ~n941 ;
  assign n943 = ( n898 & n940 ) | ( n898 & ~n942 ) | ( n940 & ~n942 ) ;
  assign n944 = ~n100 & n943 ;
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  assign n947 = n936 | n945 ;
  assign n948 = ( n39 & n946 ) | ( n39 & n947 ) | ( n946 & n947 ) ;
  assign n949 = ~n269 & n898 ;
  assign n950 = ( n166 & n200 ) | ( n166 & n949 ) | ( n200 & n949 ) ;
  assign n951 = ~n167 & n950 ;
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  assign n954 = n136 | n952 ;
  assign n955 = ( n948 & n953 ) | ( n948 & n954 ) | ( n953 & n954 ) ;
  assign n956 = ~n240 & n955 ;
  assign n957 = ( n925 & ~n926 ) | ( n925 & n956 ) | ( ~n926 & n956 ) ;
  assign n958 = n76 & n957 ;
  assign n959 = ( ~n278 & n874 ) | ( ~n278 & n958 ) | ( n874 & n958 ) ;
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n110( .i (n109), .o (n110) );
  assign n963 = ( n110 & ~n280 ) | ( n110 & n960 ) | ( ~n280 & n960 ) ;
  assign n964 = n840 & ~n963 ;
  assign n965 = ( n841 & n962 ) | ( n841 & ~n964 ) | ( n962 & ~n964 ) ;
  assign n966 = n831 | n965 ;
  assign n967 = ( n521 & n832 ) | ( n521 & n966 ) | ( n832 & n966 ) ;
  buffer buf_n77( .i (n76), .o (n77) );
  assign n968 = n127 & n160 ;
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  assign n980 = n674 & ~n978 ;
  assign n981 = n443 & ~n477 ;
  assign n982 = ( n979 & n980 ) | ( n979 & n981 ) | ( n980 & n981 ) ;
  buffer buf_n241( .i (n240), .o (n241) );
  assign n983 = ~n241 & n276 ;
  assign n984 = ( n76 & n982 ) | ( n76 & n983 ) | ( n982 & n983 ) ;
  assign n985 = ~n77 & n984 ;
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  assign n988 = ( n46 & n110 ) | ( n46 & ~n986 ) | ( n110 & ~n986 ) ;
  assign n989 = n58 | n189 ;
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  assign n1001 = n164 | n233 ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  assign n1006 = ( n69 & ~n200 ) | ( n69 & n1002 ) | ( ~n200 & n1002 ) ;
  assign n1007 = n157 | n191 ;
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  assign n1019 = ( ~n163 & n632 ) | ( ~n163 & n1012 ) | ( n632 & n1012 ) ;
  buffer buf_n1020( .i (n1019), .o (n1020) );
  assign n1026 = ( n634 & n660 ) | ( n634 & n1020 ) | ( n660 & n1020 ) ;
  assign n1027 = n69 & n1026 ;
  assign n1028 = ( n1000 & ~n1006 ) | ( n1000 & n1027 ) | ( ~n1006 & n1027 ) ;
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  assign n1032 = n477 & ~n1031 ;
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  assign n1033 = n137 & n1025 ;
  assign n1034 = n477 | n1033 ;
  assign n1035 = ~n1032 & n1034 ;
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n446( .i (n445), .o (n446) );
  assign n1038 = ~n263 & n299 ;
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  assign n1054 = ( n446 & n1036 ) | ( n446 & ~n1052 ) | ( n1036 & ~n1052 ) ;
  assign n1055 = n1037 & ~n1054 ;
  assign n1056 = n110 & n1055 ;
  assign n1057 = ( n987 & n988 ) | ( n987 & n1056 ) | ( n988 & n1056 ) ;
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  assign n1060 = ~n91 & n191 ;
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  assign n1079 = ~n60 & n91 ;
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  assign n1092 = ( n170 & ~n1072 ) | ( n170 & n1091 ) | ( ~n1072 & n1091 ) ;
  assign n1093 = n41 & ~n1092 ;
  assign n1094 = n60 & n157 ;
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  assign n1110 = n41 | n1107 ;
  assign n1111 = ( ~n42 & n1093 ) | ( ~n42 & n1110 ) | ( n1093 & n1110 ) ;
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  assign n1114 = ~n235 & n438 ;
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  assign n1122 = ( n278 & ~n1112 ) | ( n278 & n1121 ) | ( ~n1112 & n1121 ) ;
  assign n1123 = n1113 & n1122 ;
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  assign n1126 = ~n439 & n1045 ;
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  assign n1135 = n1078 & n1134 ;
  assign n1136 = ~n1124 & n1135 ;
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  assign n1137 = n144 & ~n483 ;
  assign n1138 = ( n1125 & n1136 ) | ( n1125 & n1137 ) | ( n1136 & n1137 ) ;
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  assign n1139 = ( ~n64 & n95 ) | ( ~n64 & n161 ) | ( n95 & n161 ) ;
  assign n1140 = n160 & n194 ;
  assign n1141 = ( n95 & n161 ) | ( n95 & n1140 ) | ( n161 & n1140 ) ;
  assign n1142 = ( n1098 & n1139 ) | ( n1098 & ~n1141 ) | ( n1139 & ~n1141 ) ;
  assign n1143 = n663 & n1081 ;
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  assign n1146 = n129 | n1144 ;
  assign n1147 = ( ~n1142 & n1145 ) | ( ~n1142 & n1146 ) | ( n1145 & n1146 ) ;
  assign n1148 = n34 & ~n1147 ;
  assign n1149 = n66 & n970 ;
  assign n1150 = n34 | n1149 ;
  assign n1151 = ~n1148 & n1150 ;
  buffer buf_n1152( .i (n1151), .o (n1152) );
  assign n1161 = n227 & n705 ;
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  assign n1164 = n366 | n1162 ;
  assign n1165 = ( ~n400 & n1163 ) | ( ~n400 & n1164 ) | ( n1163 & n1164 ) ;
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  assign n1172 = n1152 & n1170 ;
  assign n1173 = n440 & ~n1172 ;
  buffer buf_n1174( .i (n162), .o (n1174) );
  assign n1175 = ( n97 & ~n587 ) | ( n97 & n1174 ) | ( ~n587 & n1174 ) ;
  buffer buf_n1176( .i (n1175), .o (n1176) );
  assign n1177 = ~n199 & n1176 ;
  assign n1178 = ( ~n199 & n589 ) | ( ~n199 & n1176 ) | ( n589 & n1176 ) ;
  assign n1179 = ( n590 & n1177 ) | ( n590 & ~n1178 ) | ( n1177 & ~n1178 ) ;
  assign n1180 = n134 & n1179 ;
  assign n1181 = n440 | n1180 ;
  assign n1182 = ~n1173 & n1181 ;
  assign n1183 = ~n476 & n1182 ;
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  assign n1186 = n475 & n1029 ;
  assign n1187 = ( n442 & n594 ) | ( n442 & ~n1186 ) | ( n594 & ~n1186 ) ;
  assign n1188 = n595 & ~n1187 ;
  assign n1189 = n1184 | n1188 ;
  assign n1190 = ( n107 & n1185 ) | ( n107 & n1189 ) | ( n1185 & n1189 ) ;
  assign n1191 = n278 & n1190 ;
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  assign n1194 = n445 & n754 ;
  assign n1195 = ( n480 & n1159 ) | ( n480 & ~n1194 ) | ( n1159 & ~n1194 ) ;
  assign n1196 = n1160 & ~n1195 ;
  assign n1197 = n1192 | n1196 ;
  assign n1198 = ( n246 & n1193 ) | ( n246 & n1197 ) | ( n1193 & n1197 ) ;
  buffer buf_n1199( .i (n1198), .o (n1199) );
  assign n1200 = ( ~n1058 & n1138 ) | ( ~n1058 & n1199 ) | ( n1138 & n1199 ) ;
  assign n1201 = n520 | n1199 ;
  assign n1202 = ( n1059 & n1200 ) | ( n1059 & n1201 ) | ( n1200 & n1201 ) ;
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  assign n1203 = n133 & ~n1102 ;
  buffer buf_n1204( .i (n36), .o (n1204) );
  assign n1205 = n1203 & n1204 ;
  assign n1206 = n27 & ~n91 ;
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  assign n1215 = n68 & ~n132 ;
  assign n1216 = ( ~n36 & n1214 ) | ( ~n36 & n1215 ) | ( n1214 & n1215 ) ;
  assign n1217 = n1170 & n1216 ;
  assign n1218 = ( n1171 & n1205 ) | ( n1171 & n1217 ) | ( n1205 & n1217 ) ;
  assign n1219 = n93 | n126 ;
  buffer buf_n1220( .i (n1219), .o (n1220) );
  assign n1236 = n93 & ~n126 ;
  buffer buf_n1237( .i (n1236), .o (n1237) );
  assign n1238 = ( ~n95 & n1220 ) | ( ~n95 & n1237 ) | ( n1220 & n1237 ) ;
  buffer buf_n1239( .i (n1238), .o (n1239) );
  assign n1245 = n587 & n1239 ;
  assign n1246 = n436 | n1245 ;
  assign n1247 = n31 | n64 ;
  assign n1248 = n31 & ~n1237 ;
  assign n1249 = n1247 & ~n1248 ;
  assign n1250 = n1166 & n1249 ;
  assign n1251 = n436 & ~n1250 ;
  assign n1252 = n1246 & ~n1251 ;
  assign n1253 = n166 & n1252 ;
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  assign n1256 = n440 | n1254 ;
  assign n1257 = ( n1218 & n1255 ) | ( n1218 & n1256 ) | ( n1255 & n1256 ) ;
  assign n1258 = ~n476 & n1257 ;
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n99), .o (n1261) );
  assign n1262 = n69 | n1261 ;
  assign n1263 = ~n85 & n118 ;
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1283( .i (n68), .o (n1283) );
  assign n1284 = n1277 & n1283 ;
  assign n1285 = ( ~n70 & n1262 ) | ( ~n70 & n1284 ) | ( n1262 & n1284 ) ;
  buffer buf_n1286( .i (n1285), .o (n1286) );
  assign n1290 = n475 & n1286 ;
  assign n1291 = ( n442 & n594 ) | ( n442 & ~n1290 ) | ( n594 & ~n1290 ) ;
  assign n1292 = n595 & ~n1291 ;
  assign n1293 = n1259 | n1292 ;
  assign n1294 = ( n173 & n1260 ) | ( n173 & n1293 ) | ( n1260 & n1293 ) ;
  buffer buf_n1295( .i (n277), .o (n1295) );
  assign n1296 = n1294 & n1295 ;
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  assign n1299 = ( n64 & ~n128 ) | ( n64 & n161 ) | ( ~n128 & n161 ) ;
  buffer buf_n1300( .i (n128), .o (n1300) );
  assign n1301 = ~n1299 & n1300 ;
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  assign n1304 = ~n130 & n1174 ;
  assign n1305 = ( n98 & n1302 ) | ( n98 & n1304 ) | ( n1302 & n1304 ) ;
  assign n1306 = n1303 | n1305 ;
  buffer buf_n1307( .i (n30), .o (n1307) );
  assign n1308 = ~n1220 & n1307 ;
  assign n1309 = n792 & ~n1307 ;
  assign n1310 = ( n32 & ~n1308 ) | ( n32 & n1309 ) | ( ~n1308 & n1309 ) ;
  assign n1311 = n66 & ~n1310 ;
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  assign n1314 = n35 | n1312 ;
  assign n1315 = ( n1306 & n1313 ) | ( n1306 & n1314 ) | ( n1313 & n1314 ) ;
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  assign n1322 = n445 & n1321 ;
  assign n1323 = ( n480 & n755 ) | ( n480 & ~n1322 ) | ( n755 & ~n1322 ) ;
  assign n1324 = n756 & ~n1323 ;
  assign n1325 = n1297 | n1324 ;
  assign n1326 = ( n246 & n1298 ) | ( n246 & n1325 ) | ( n1298 & n1325 ) ;
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  assign n1329 = ~n213 & n1327 ;
  assign n1330 = n159 & ~n465 ;
  assign n1331 = ( n94 & n194 ) | ( n94 & n1330 ) | ( n194 & n1330 ) ;
  assign n1332 = ~n195 & n1331 ;
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  assign n1344 = ~n135 & n237 ;
  assign n1345 = ( n203 & n1280 ) | ( n203 & ~n1344 ) | ( n1280 & ~n1344 ) ;
  buffer buf_n1346( .i (n185), .o (n1346) );
  assign n1347 = n221 & ~n1346 ;
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  assign n1366 = n1278 & n1361 ;
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  assign n1369 = n169 | n1367 ;
  assign n1370 = ( ~n1345 & n1368 ) | ( ~n1345 & n1369 ) | ( n1368 & n1369 ) ;
  assign n1371 = ( n74 & n1341 ) | ( n74 & n1370 ) | ( n1341 & n1370 ) ;
  assign n1372 = n478 & ~n1371 ;
  assign n1373 = ( n479 & n1343 ) | ( n479 & ~n1372 ) | ( n1343 & ~n1372 ) ;
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  assign n1378 = n275 & n595 ;
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  assign n1384 = ( n449 & n1376 ) | ( n449 & ~n1383 ) | ( n1376 & ~n1383 ) ;
  assign n1385 = n1377 & ~n1384 ;
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  assign n1386 = ( n311 & n540 ) | ( n311 & ~n1288 ) | ( n540 & ~n1288 ) ;
  assign n1387 = n1289 & n1386 ;
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  assign n1390 = ( n439 & ~n1045 ) | ( n439 & n1243 ) | ( ~n1045 & n1243 ) ;
  assign n1391 = n1244 & ~n1390 ;
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n475), .o (n1394) );
  assign n1395 = ( ~n170 & n1392 ) | ( ~n170 & n1394 ) | ( n1392 & n1394 ) ;
  assign n1396 = ( n272 & n1115 ) | ( n272 & ~n1316 ) | ( n1115 & ~n1316 ) ;
  assign n1397 = n1317 & n1396 ;
  assign n1398 = ~n1394 & n1397 ;
  assign n1399 = ( n1393 & ~n1395 ) | ( n1393 & n1398 ) | ( ~n1395 & n1398 ) ;
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  assign n1403 = ( n173 & ~n277 ) | ( n173 & n1400 ) | ( ~n277 & n1400 ) ;
  assign n1404 = n1388 & ~n1403 ;
  assign n1405 = ( n1389 & n1402 ) | ( n1389 & ~n1404 ) | ( n1402 & ~n1404 ) ;
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  assign n1408 = ( n211 & n518 ) | ( n211 & ~n1406 ) | ( n518 & ~n1406 ) ;
  buffer buf_n1053( .i (n1052), .o (n1053) );
  assign n1409 = ( n447 & ~n1053 ) | ( n447 & n1374 ) | ( ~n1053 & n1374 ) ;
  assign n1410 = n1375 & ~n1409 ;
  assign n1411 = n518 & n1410 ;
  assign n1412 = ( n1407 & n1408 ) | ( n1407 & n1411 ) | ( n1408 & n1411 ) ;
  assign n1413 = n1385 | n1412 ;
  assign n1414 = ( n1328 & ~n1329 ) | ( n1328 & n1413 ) | ( ~n1329 & n1413 ) ;
  buffer buf_n1415( .i (n166), .o (n1415) );
  assign n1416 = ( n201 & ~n473 ) | ( n201 & n1415 ) | ( ~n473 & n1415 ) ;
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  assign n1419 = ( n135 & n168 ) | ( n135 & n474 ) | ( n168 & n474 ) ;
  assign n1420 = n1417 & ~n1419 ;
  assign n1421 = ( ~n204 & n1418 ) | ( ~n204 & n1420 ) | ( n1418 & n1420 ) ;
  assign n1422 = n89 & ~n155 ;
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  assign n1432 = ( n98 & n198 ) | ( n98 & n1430 ) | ( n198 & n1430 ) ;
  buffer buf_n1433( .i (n1300), .o (n1433) );
  assign n1434 = ( n197 & n1174 ) | ( n197 & n1433 ) | ( n1174 & n1433 ) ;
  assign n1435 = ( n1174 & n1429 ) | ( n1174 & ~n1433 ) | ( n1429 & ~n1433 ) ;
  assign n1436 = n1434 | n1435 ;
  assign n1437 = ( n1431 & ~n1432 ) | ( n1431 & n1436 ) | ( ~n1432 & n1436 ) ;
  assign n1438 = n472 & n1437 ;
  buffer buf_n1439( .i (n1438), .o (n1439) );
  assign n1441 = n71 & n1439 ;
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  assign n1444 = n104 | n1442 ;
  assign n1445 = ( n1421 & n1443 ) | ( n1421 & n1444 ) | ( n1443 & n1444 ) ;
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n444), .o (n1448) );
  assign n1449 = ( ~n1379 & n1446 ) | ( ~n1379 & n1448 ) | ( n1446 & n1448 ) ;
  assign n1450 = n1447 & ~n1449 ;
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  assign n1453 = ~n245 & n1451 ;
  assign n1454 = ( n65 & n96 ) | ( n65 & n196 ) | ( n96 & n196 ) ;
  assign n1455 = n196 & n793 ;
  assign n1456 = ( ~n66 & n1454 ) | ( ~n66 & n1455 ) | ( n1454 & n1455 ) ;
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  assign n1459 = ( ~n85 & n118 ) | ( ~n85 & n185 ) | ( n118 & n185 ) ;
  buffer buf_n1460( .i (n1459), .o (n1460) );
  assign n1481 = n153 & ~n1460 ;
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n1488( .i (n1487), .o (n1488) );
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  assign n1493 = ( ~n21 & n85 ) | ( ~n21 & n185 ) | ( n85 & n185 ) ;
  buffer buf_n1494( .i (n184), .o (n1494) );
  assign n1495 = ( n21 & n118 ) | ( n21 & n1494 ) | ( n118 & n1494 ) ;
  assign n1496 = ~n1493 & n1495 ;
  assign n1497 = ( ~n20 & n117 ) | ( ~n20 & n184 ) | ( n117 & n184 ) ;
  assign n1498 = ~n19 & n149 ;
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1510( .i (n117), .o (n1510) );
  assign n1511 = ( n1497 & n1499 ) | ( n1497 & ~n1510 ) | ( n1499 & ~n1510 ) ;
  buffer buf_n1512( .i (n1511), .o (n1512) );
  assign n1522 = ( n56 & n1496 ) | ( n56 & n1512 ) | ( n1496 & n1512 ) ;
  assign n1523 = ~n623 & n1522 ;
  assign n1524 = ( n58 & n624 ) | ( n58 & n1523 ) | ( n624 & n1523 ) ;
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  assign n1534 = ( ~n1457 & n1492 ) | ( ~n1457 & n1533 ) | ( n1492 & n1533 ) ;
  assign n1535 = n27 | n1525 ;
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1543( .i (n1542), .o (n1543) );
  assign n1544 = ( n1458 & n1534 ) | ( n1458 & n1543 ) | ( n1534 & n1543 ) ;
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  buffer buf_n1549( .i (n1548), .o (n1549) );
  assign n1550 = ( ~n262 & n364 ) | ( ~n262 & n397 ) | ( n364 & n397 ) ;
  buffer buf_n1551( .i (n1550), .o (n1551) );
  assign n1555 = ( n264 & ~n334 ) | ( n264 & n1551 ) | ( ~n334 & n1551 ) ;
  buffer buf_n1556( .i (n1555), .o (n1556) );
  buffer buf_n1557( .i (n1556), .o (n1557) );
  buffer buf_n1558( .i (n1557), .o (n1558) );
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  assign n1561 = ( n266 & n368 ) | ( n266 & ~n1556 ) | ( n368 & ~n1556 ) ;
  assign n1562 = n1554 | n1561 ;
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  assign n1565 = ~n339 & n1563 ;
  assign n1566 = ( ~n1560 & n1564 ) | ( ~n1560 & n1565 ) | ( n1564 & n1565 ) ;
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  assign n1570 = n442 & n1569 ;
  buffer buf_n1571( .i (n1394), .o (n1571) );
  assign n1572 = ( n1548 & ~n1570 ) | ( n1548 & n1571 ) | ( ~n1570 & n1571 ) ;
  assign n1573 = n1549 & ~n1572 ;
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  assign n1576 = ( n243 & n314 ) | ( n243 & ~n1574 ) | ( n314 & ~n1574 ) ;
  buffer buf_n1440( .i (n1439), .o (n1440) );
  assign n1577 = n234 & ~n437 ;
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  assign n1581 = ( n273 & n1440 ) | ( n273 & n1580 ) | ( n1440 & n1580 ) ;
  assign n1582 = ~n274 & n1581 ;
  buffer buf_n1583( .i (n1582), .o (n1583) );
  buffer buf_n1584( .i (n1583), .o (n1584) );
  assign n1585 = ( n75 & n513 ) | ( n75 & ~n1583 ) | ( n513 & ~n1583 ) ;
  buffer buf_n1586( .i (n162), .o (n1586) );
  buffer buf_n1587( .i (n196), .o (n1587) );
  assign n1588 = ( ~n435 & n1586 ) | ( ~n435 & n1587 ) | ( n1586 & n1587 ) ;
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n435), .o (n1591) );
  assign n1592 = ( n131 & n164 ) | ( n131 & n1591 ) | ( n164 & n1591 ) ;
  assign n1593 = n1589 & ~n1592 ;
  buffer buf_n1594( .i (n198), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  assign n1596 = ( n1590 & n1593 ) | ( n1590 & ~n1595 ) | ( n1593 & ~n1595 ) ;
  assign n1597 = ~n271 & n1596 ;
  assign n1598 = n237 & n1597 ;
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  assign n1601 = ( ~n104 & n1394 ) | ( ~n104 & n1599 ) | ( n1394 & n1599 ) ;
  assign n1602 = ( n272 & n1115 ) | ( n272 & ~n1545 ) | ( n1115 & ~n1545 ) ;
  assign n1603 = n1546 & n1602 ;
  buffer buf_n1604( .i (n474), .o (n1604) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  assign n1606 = n1603 & ~n1605 ;
  assign n1607 = ( n1600 & ~n1601 ) | ( n1600 & n1606 ) | ( ~n1601 & n1606 ) ;
  assign n1608 = n513 & n1607 ;
  assign n1609 = ( n1584 & n1585 ) | ( n1584 & n1608 ) | ( n1585 & n1608 ) ;
  assign n1610 = n314 & n1609 ;
  assign n1611 = ( n1575 & n1576 ) | ( n1575 & n1610 ) | ( n1576 & n1610 ) ;
  assign n1612 = n92 & ~n464 ;
  buffer buf_n1613( .i (n1612), .o (n1613) );
  assign n1616 = n94 & ~n1613 ;
  buffer buf_n1617( .i (n1616), .o (n1617) );
  assign n1618 = ~n65 & n1617 ;
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  assign n1619 = ( n1300 & ~n1615 ) | ( n1300 & n1617 ) | ( ~n1615 & n1617 ) ;
  assign n1620 = ( ~n469 & n1618 ) | ( ~n469 & n1619 ) | ( n1618 & n1619 ) ;
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  assign n1627 = n274 & n1626 ;
  buffer buf_n1628( .i (n594), .o (n1628) );
  assign n1629 = ( n443 & ~n1627 ) | ( n443 & n1628 ) | ( ~n1627 & n1628 ) ;
  assign n1630 = n596 & ~n1629 ;
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  assign n1633 = ( ~n243 & n643 ) | ( ~n243 & n1631 ) | ( n643 & n1631 ) ;
  assign n1634 = n231 & ~n266 ;
  assign n1635 = n266 & n434 ;
  assign n1636 = ~n230 & n1307 ;
  assign n1637 = n434 & ~n1636 ;
  assign n1638 = ( n1634 & n1635 ) | ( n1634 & ~n1637 ) | ( n1635 & ~n1637 ) ;
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  assign n1641 = ( n471 & ~n1276 ) | ( n471 & n1639 ) | ( ~n1276 & n1639 ) ;
  assign n1642 = n1640 & ~n1641 ;
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  assign n1646 = n235 & ~n1283 ;
  assign n1647 = n101 & n1646 ;
  assign n1648 = ( ~n272 & n1643 ) | ( ~n272 & n1647 ) | ( n1643 & n1647 ) ;
  assign n1649 = n538 & ~n1648 ;
  assign n1650 = ( n539 & n1645 ) | ( n539 & ~n1649 ) | ( n1645 & ~n1649 ) ;
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  assign n1653 = ( n312 & n513 ) | ( n312 & ~n1651 ) | ( n513 & ~n1651 ) ;
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  assign n1654 = n236 & ~n473 ;
  buffer buf_n1655( .i (n439), .o (n1655) );
  assign n1656 = ( ~n1567 & n1654 ) | ( ~n1567 & n1655 ) | ( n1654 & n1655 ) ;
  assign n1657 = n1568 & n1656 ;
  assign n1658 = ( n104 & n882 ) | ( n104 & n1657 ) | ( n882 & n1657 ) ;
  assign n1659 = ~n105 & n1658 ;
  assign n1660 = n312 & n1659 ;
  assign n1661 = ( n1652 & n1653 ) | ( n1652 & n1660 ) | ( n1653 & n1660 ) ;
  assign n1662 = ~n643 & n1661 ;
  assign n1663 = ( n1632 & ~n1633 ) | ( n1632 & n1662 ) | ( ~n1633 & n1662 ) ;
  assign n1664 = n1611 | n1663 ;
  assign n1665 = ( n1452 & ~n1453 ) | ( n1452 & n1664 ) | ( ~n1453 & n1664 ) ;
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  assign n1669 = n189 & n461 ;
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1673( .i (n190), .o (n1673) );
  assign n1674 = ~n1670 & n1673 ;
  buffer buf_n1675( .i (n1674), .o (n1675) );
  assign n1676 = n93 & n1675 ;
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  assign n1677 = ( n1095 & ~n1672 ) | ( n1095 & n1675 ) | ( ~n1672 & n1675 ) ;
  assign n1678 = ( n466 & n1676 ) | ( n466 & n1677 ) | ( n1676 & n1677 ) ;
  assign n1679 = ~n459 & n1264 ;
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  assign n1683 = ( n58 & ~n843 ) | ( n58 & n1680 ) | ( ~n843 & n1680 ) ;
  assign n1684 = n462 & ~n1683 ;
  assign n1685 = ( n463 & n1682 ) | ( n463 & ~n1684 ) | ( n1682 & ~n1684 ) ;
  assign n1686 = ( n55 & n221 ) | ( n55 & ~n458 ) | ( n221 & ~n458 ) ;
  assign n1687 = ( n152 & n221 ) | ( n152 & n458 ) | ( n221 & n458 ) ;
  assign n1688 = n1686 & n1687 ;
  assign n1689 = n183 & ~n455 ;
  assign n1690 = n51 & ~n217 ;
  assign n1691 = n455 & ~n1690 ;
  assign n1692 = n1689 | n1691 ;
  assign n1693 = n151 & ~n1692 ;
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  assign n1696 = n187 | n1694 ;
  assign n1697 = ( ~n1688 & n1695 ) | ( ~n1688 & n1696 ) | ( n1695 & n1696 ) ;
  assign n1698 = n89 & n1697 ;
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  assign n1701 = n1673 | n1699 ;
  assign n1702 = ( n1685 & n1700 ) | ( n1685 & n1701 ) | ( n1700 & n1701 ) ;
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  assign n1705 = n127 & ~n1703 ;
  assign n1706 = ( n1678 & n1704 ) | ( n1678 & ~n1705 ) | ( n1704 & ~n1705 ) ;
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  assign n1716 = n300 & ~n334 ;
  buffer buf_n1717( .i (n1716), .o (n1717) );
  assign n1718 = ( n302 & n368 ) | ( n302 & n1717 ) | ( n368 & n1717 ) ;
  assign n1719 = ( ~n302 & n368 ) | ( ~n302 & n1717 ) | ( n368 & n1717 ) ;
  assign n1720 = ( n303 & ~n1718 ) | ( n303 & n1719 ) | ( ~n1718 & n1719 ) ;
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  assign n1728 = n1715 & n1727 ;
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  assign n1731 = n157 | n1268 ;
  assign n1732 = ( ~n604 & n1269 ) | ( ~n604 & n1731 ) | ( n1269 & n1731 ) ;
  buffer buf_n1733( .i (n57), .o (n1733) );
  assign n1734 = ( ~n89 & n122 ) | ( ~n89 & n1733 ) | ( n122 & n1733 ) ;
  buffer buf_n1735( .i (n88), .o (n1735) );
  assign n1736 = ( ~n155 & n1733 ) | ( ~n155 & n1735 ) | ( n1733 & n1735 ) ;
  assign n1737 = ~n1734 & n1736 ;
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  assign n1740 = n61 | n1738 ;
  assign n1741 = ( n1732 & n1739 ) | ( n1732 & n1740 ) | ( n1739 & n1740 ) ;
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  assign n1749 = n471 & n1721 ;
  assign n1750 = ( n438 & n1747 ) | ( n438 & ~n1749 ) | ( n1747 & ~n1749 ) ;
  assign n1751 = n1748 & ~n1750 ;
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  assign n1754 = ( n238 & n273 ) | ( n238 & ~n1752 ) | ( n273 & ~n1752 ) ;
  assign n1755 = n86 & n1346 ;
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  assign n1772 = ~n1482 & n1733 ;
  assign n1773 = ( n1483 & n1758 ) | ( n1483 & ~n1772 ) | ( n1758 & ~n1772 ) ;
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  assign n1781 = n323 & ~n388 ;
  assign n1782 = ~n251 & n321 ;
  buffer buf_n1783( .i (n1782), .o (n1783) );
  assign n1804 = ( ~n289 & n323 ) | ( ~n289 & n1783 ) | ( n323 & n1783 ) ;
  assign n1805 = ( n717 & n1781 ) | ( n717 & ~n1804 ) | ( n1781 & ~n1804 ) ;
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  buffer buf_n1813( .i (n1812), .o (n1813) );
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  assign n1818 = ( ~n33 & n1779 ) | ( ~n33 & n1817 ) | ( n1779 & n1817 ) ;
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  assign n1819 = n193 & ~n1207 ;
  assign n1820 = n1009 & ~n1819 ;
  buffer buf_n1821( .i (n63), .o (n1821) );
  assign n1822 = n1820 & n1821 ;
  assign n1823 = ( n65 & n1521 ) | ( n65 & n1822 ) | ( n1521 & n1822 ) ;
  assign n1824 = ~n1817 & n1823 ;
  assign n1825 = ( n1780 & ~n1818 ) | ( n1780 & n1824 ) | ( ~n1818 & n1824 ) ;
  assign n1826 = n424 & ~n1806 ;
  buffer buf_n1827( .i (n1826), .o (n1827) );
  assign n1829 = n188 & n1827 ;
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  assign n1832 = ( ~n26 & n90 ) | ( ~n26 & n1830 ) | ( n90 & n1830 ) ;
  buffer buf_n1828( .i (n1827), .o (n1828) );
  assign n1833 = ( ~n24 & n154 ) | ( ~n24 & n1827 ) | ( n154 & n1827 ) ;
  assign n1834 = n290 & n324 ;
  buffer buf_n1835( .i (n1834), .o (n1835) );
  assign n1855 = n256 & ~n1835 ;
  assign n1856 = ~n425 & n1855 ;
  assign n1857 = ~n154 & n1856 ;
  assign n1858 = ( n1828 & ~n1833 ) | ( n1828 & n1857 ) | ( ~n1833 & n1857 ) ;
  assign n1859 = ~n90 & n1858 ;
  assign n1860 = ( n1831 & ~n1832 ) | ( n1831 & n1859 ) | ( ~n1832 & n1859 ) ;
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  assign n1864 = ( n60 & n1673 ) | ( n60 & ~n1811 ) | ( n1673 & ~n1811 ) ;
  buffer buf_n1865( .i (n156), .o (n1865) );
  assign n1866 = ( n1673 & n1811 ) | ( n1673 & n1865 ) | ( n1811 & n1865 ) ;
  assign n1867 = n1864 & ~n1866 ;
  assign n1868 = ( n29 & n1861 ) | ( n29 & n1867 ) | ( n1861 & n1867 ) ;
  assign n1869 = n432 & ~n1868 ;
  assign n1870 = ( n433 & n1863 ) | ( n433 & ~n1869 ) | ( n1863 & ~n1869 ) ;
  assign n1871 = n1300 & n1870 ;
  buffer buf_n1872( .i (n1871), .o (n1872) );
  buffer buf_n1873( .i (n1872), .o (n1873) );
  assign n1874 = n1591 | n1872 ;
  assign n1875 = ( n1825 & n1873 ) | ( n1825 & n1874 ) | ( n1873 & n1874 ) ;
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  assign n1878 = ( ~n373 & n473 ) | ( ~n373 & n1876 ) | ( n473 & n1876 ) ;
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n1879( .i (n154), .o (n1879) );
  assign n1880 = ( ~n189 & n1735 ) | ( ~n189 & n1879 ) | ( n1735 & n1879 ) ;
  assign n1881 = n123 & ~n1880 ;
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  assign n1884 = ( n1526 & n1774 ) | ( n1526 & ~n1882 ) | ( n1774 & ~n1882 ) ;
  assign n1885 = ( n1536 & n1883 ) | ( n1536 & n1884 ) | ( n1883 & n1884 ) ;
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n1899( .i (n301), .o (n1899) );
  assign n1900 = ( n495 & n1887 ) | ( n495 & n1899 ) | ( n1887 & n1899 ) ;
  assign n1901 = n331 & ~n363 ;
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  assign n1916 = n1887 & n1905 ;
  assign n1917 = ( ~n303 & n1900 ) | ( ~n303 & n1916 ) | ( n1900 & n1916 ) ;
  buffer buf_n1918( .i (n1917), .o (n1918) );
  buffer buf_n1919( .i (n1918), .o (n1919) );
  assign n1920 = ( n269 & n437 ) | ( n269 & ~n1918 ) | ( n437 & ~n1918 ) ;
  assign n1921 = ~n92 & n789 ;
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  assign n1929 = ~n434 & n1845 ;
  assign n1930 = ( n369 & n1925 ) | ( n369 & n1929 ) | ( n1925 & n1929 ) ;
  assign n1931 = ~n370 & n1930 ;
  buffer buf_n1932( .i (n268), .o (n1932) );
  assign n1933 = n1931 & n1932 ;
  assign n1934 = ( n1919 & n1920 ) | ( n1919 & n1933 ) | ( n1920 & n1933 ) ;
  buffer buf_n1935( .i (n472), .o (n1935) );
  assign n1936 = n1934 & ~n1935 ;
  assign n1937 = ( n1877 & ~n1878 ) | ( n1877 & n1936 ) | ( ~n1878 & n1936 ) ;
  assign n1938 = n238 & n1937 ;
  assign n1939 = ( n1753 & n1754 ) | ( n1753 & n1938 ) | ( n1754 & n1938 ) ;
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1941( .i (n1940), .o (n1941) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  assign n1943 = ( n276 & ~n444 ) | ( n276 & n1940 ) | ( ~n444 & n1940 ) ;
  assign n1944 = n1729 & ~n1943 ;
  assign n1945 = ( n1730 & n1942 ) | ( n1730 & ~n1944 ) | ( n1942 & ~n1944 ) ;
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  assign n1952 = n226 & ~n1865 ;
  buffer buf_n1953( .i (n1952), .o (n1953) );
  assign n1960 = n193 | n1953 ;
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1966( .i (n1965), .o (n1966) );
  assign n1967 = ( n437 & ~n1621 ) | ( n437 & n1965 ) | ( ~n1621 & n1965 ) ;
  buffer buf_n1968( .i (n90), .o (n1968) );
  assign n1969 = ( n124 & n226 ) | ( n124 & ~n1968 ) | ( n226 & ~n1968 ) ;
  assign n1970 = ( n226 & n1865 ) | ( n226 & n1968 ) | ( n1865 & n1968 ) ;
  assign n1971 = ~n1969 & n1970 ;
  buffer buf_n1972( .i (n1971), .o (n1972) );
  buffer buf_n1973( .i (n1972), .o (n1973) );
  assign n1974 = ( n123 & n190 ) | ( n123 & ~n225 ) | ( n190 & ~n225 ) ;
  assign n1975 = n1865 & ~n1974 ;
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1986( .i (n1735), .o (n1986) );
  assign n1987 = n225 & ~n1986 ;
  assign n1988 = n124 & n1987 ;
  buffer buf_n1989( .i (n1988), .o (n1989) );
  assign n1999 = ( n465 & n1976 ) | ( n465 & n1989 ) | ( n1976 & n1989 ) ;
  assign n2000 = ~n1972 & n1999 ;
  assign n2001 = ( n467 & n1973 ) | ( n467 & n2000 ) | ( n1973 & n2000 ) ;
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n1821), .o (n2004) );
  buffer buf_n2005( .i (n2004), .o (n2005) );
  assign n2006 = n2002 & ~n2005 ;
  assign n2007 = n461 | n1735 ;
  assign n2008 = n57 & n121 ;
  assign n2009 = n461 & ~n2008 ;
  assign n2010 = n2007 & ~n2009 ;
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n2012( .i (n2011), .o (n2012) );
  assign n2013 = ~n227 & n2011 ;
  assign n2014 = ( ~n159 & n2012 ) | ( ~n159 & n2013 ) | ( n2012 & n2013 ) ;
  buffer buf_n2015( .i (n2014), .o (n2015) );
  buffer buf_n2016( .i (n2015), .o (n2016) );
  assign n2017 = ( ~n92 & n227 ) | ( ~n92 & n464 ) | ( n227 & n464 ) ;
  buffer buf_n2018( .i (n1968), .o (n2018) );
  assign n2019 = ( ~n125 & n464 ) | ( ~n125 & n2018 ) | ( n464 & n2018 ) ;
  assign n2020 = ~n2017 & n2019 ;
  buffer buf_n2021( .i (n225), .o (n2021) );
  assign n2022 = n463 & ~n2021 ;
  assign n2023 = ( n61 & n158 ) | ( n61 & n2022 ) | ( n158 & n2022 ) ;
  buffer buf_n2024( .i (n158), .o (n2024) );
  assign n2025 = n2023 & ~n2024 ;
  assign n2026 = ( n194 & n2020 ) | ( n194 & n2025 ) | ( n2020 & n2025 ) ;
  assign n2027 = ~n2015 & n2026 ;
  buffer buf_n2028( .i (n195), .o (n2028) );
  assign n2029 = ( n2016 & n2027 ) | ( n2016 & n2028 ) | ( n2027 & n2028 ) ;
  assign n2030 = n1333 | n2029 ;
  assign n2031 = ( n2003 & ~n2006 ) | ( n2003 & n2030 ) | ( ~n2006 & n2030 ) ;
  buffer buf_n2032( .i (n1591), .o (n2032) );
  assign n2033 = n2031 & ~n2032 ;
  assign n2034 = ( n1966 & ~n1967 ) | ( n1966 & n2033 ) | ( ~n1967 & n2033 ) ;
  buffer buf_n2035( .i (n2034), .o (n2035) );
  buffer buf_n340( .i (n339), .o (n340) );
  assign n2037 = n328 & n360 ;
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  assign n2052 = n340 & ~n2048 ;
  buffer buf_n2053( .i (n2052), .o (n2053) );
  assign n2054 = n2035 & n2053 ;
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2055( .i (n160), .o (n2055) );
  assign n2056 = n1272 & ~n2055 ;
  buffer buf_n2057( .i (n433), .o (n2057) );
  assign n2058 = n2056 & ~n2057 ;
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  assign n2061 = n433 & n1886 ;
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  assign n2071 = n467 & n1742 ;
  assign n2072 = ~n2057 & n2071 ;
  buffer buf_n2073( .i (n2072), .o (n2073) );
  assign n2076 = ( ~n2059 & n2063 ) | ( ~n2059 & n2073 ) | ( n2063 & n2073 ) ;
  assign n2077 = n470 & ~n2073 ;
  assign n2078 = ( n2060 & n2076 ) | ( n2060 & ~n2077 ) | ( n2076 & ~n2077 ) ;
  assign n2079 = ~n435 & n1707 ;
  buffer buf_n2080( .i (n2079), .o (n2080) );
  buffer buf_n2081( .i (n2080), .o (n2081) );
  buffer buf_n2086( .i (n233), .o (n2086) );
  assign n2087 = n2080 | n2086 ;
  assign n2088 = ( n2078 & n2081 ) | ( n2078 & n2087 ) | ( n2081 & n2087 ) ;
  buffer buf_n2089( .i (n2088), .o (n2089) );
  assign n2090 = ( ~n2050 & n2053 ) | ( ~n2050 & n2089 ) | ( n2053 & n2089 ) ;
  assign n2091 = ( n375 & n2054 ) | ( n375 & n2090 ) | ( n2054 & n2090 ) ;
  assign n2092 = n274 & ~n2091 ;
  buffer buf_n2036( .i (n2035), .o (n2036) );
  assign n2093 = n375 & n2036 ;
  buffer buf_n2094( .i (n273), .o (n2094) );
  assign n2095 = n2093 | n2094 ;
  assign n2096 = ~n2092 & n2095 ;
  assign n2097 = n312 & n2096 ;
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n2099( .i (n2098), .o (n2099) );
  buffer buf_n1888( .i (n1887), .o (n1888) );
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  assign n2100 = n238 | n375 ;
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n2101( .i (n237), .o (n2101) );
  buffer buf_n2102( .i (n374), .o (n2102) );
  assign n2103 = ( n703 & n2101 ) | ( n703 & ~n2102 ) | ( n2101 & ~n2102 ) ;
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1907( .i (n1906), .o (n1907) );
  buffer buf_n1908( .i (n1907), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  assign n2104 = n304 | n403 ;
  assign n2105 = ( n305 & n371 ) | ( n305 & ~n2104 ) | ( n371 & ~n2104 ) ;
  buffer buf_n2106( .i (n2105), .o (n2106) );
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n341( .i (n340), .o (n341) );
  assign n2108 = ( ~n341 & n373 ) | ( ~n341 & n2106 ) | ( n373 & n2106 ) ;
  assign n2109 = ( n1911 & ~n2107 ) | ( n1911 & n2108 ) | ( ~n2107 & n2108 ) ;
  assign n2110 = n2101 & n2109 ;
  assign n2111 = ( n2100 & ~n2103 ) | ( n2100 & n2110 ) | ( ~n2103 & n2110 ) ;
  assign n2112 = n443 & n2111 ;
  assign n2113 = ( n478 & n1897 ) | ( n478 & ~n2112 ) | ( n1897 & ~n2112 ) ;
  assign n2114 = n1898 & ~n2113 ;
  assign n2115 = n2098 | n2114 ;
  assign n2116 = ( n279 & n2099 ) | ( n279 & n2115 ) | ( n2099 & n2115 ) ;
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  buffer buf_n2119( .i (n2118), .o (n2119) );
  buffer buf_n2120( .i (n2119), .o (n2120) );
  buffer buf_n2121( .i (n2120), .o (n2121) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n2064( .i (n2063), .o (n2064) );
  buffer buf_n2065( .i (n2064), .o (n2065) );
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  assign n2122 = ~n1604 & n2068 ;
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  assign n2129 = ( n382 & n560 ) | ( n382 & n2128 ) | ( n560 & n2128 ) ;
  assign n2130 = ~n383 & n2129 ;
  buffer buf_n2131( .i (n2130), .o (n2131) );
  buffer buf_n2132( .i (n2131), .o (n2132) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n2133( .i (n271), .o (n2133) );
  assign n2134 = ( n374 & n2089 ) | ( n374 & n2133 ) | ( n2089 & n2133 ) ;
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  buffer buf_n2137( .i (n2136), .o (n2137) );
  buffer buf_n2138( .i (n2137), .o (n2138) );
  assign n2139 = ~n376 & n2135 ;
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n275), .o (n2142) );
  buffer buf_n2143( .i (n311), .o (n2143) );
  assign n2144 = ( n2140 & ~n2142 ) | ( n2140 & n2143 ) | ( ~n2142 & n2143 ) ;
  assign n2145 = ( n2138 & n2141 ) | ( n2138 & n2144 ) | ( n2141 & n2144 ) ;
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n363), .o (n2148) );
  assign n2149 = n397 & n2148 ;
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  buffer buf_n2152( .i (n2151), .o (n2152) );
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n2155( .i (n2154), .o (n2155) );
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  assign n2158 = ( ~n373 & n2066 ) | ( ~n373 & n2157 ) | ( n2066 & n2157 ) ;
  buffer buf_n2159( .i (n2158), .o (n2159) );
  buffer buf_n2160( .i (n2159), .o (n2160) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  assign n2161 = n270 & n1928 ;
  buffer buf_n2162( .i (n372), .o (n2162) );
  buffer buf_n2163( .i (n438), .o (n2163) );
  assign n2164 = ( n2161 & n2162 ) | ( n2161 & n2163 ) | ( n2162 & n2163 ) ;
  assign n2165 = ~n1655 & n2164 ;
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n2075( .i (n2074), .o (n2075) );
  assign n2166 = n372 & n2075 ;
  assign n2167 = n271 & n2166 ;
  buffer buf_n2168( .i (n2167), .o (n2168) );
  assign n2169 = ( ~n2159 & n2165 ) | ( ~n2159 & n2168 ) | ( n2165 & n2168 ) ;
  assign n2170 = n1604 & ~n2168 ;
  assign n2171 = ( n2160 & n2169 ) | ( n2160 & ~n2170 ) | ( n2169 & ~n2170 ) ;
  buffer buf_n2172( .i (n2171), .o (n2172) );
  buffer buf_n2173( .i (n2172), .o (n2173) );
  assign n2174 = ( ~n241 & n2143 ) | ( ~n241 & n2172 ) | ( n2143 & n2172 ) ;
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  assign n2175 = n376 & n2085 ;
  assign n2176 = n275 & n2175 ;
  assign n2177 = ~n2143 & n2176 ;
  assign n2178 = ( n2173 & ~n2174 ) | ( n2173 & n2177 ) | ( ~n2174 & n2177 ) ;
  assign n2179 = n377 & n2123 ;
  assign n2180 = ( n241 & n2142 ) | ( n241 & n2179 ) | ( n2142 & n2179 ) ;
  assign n2181 = ~n242 & n2180 ;
  assign n2182 = ( n348 & n2178 ) | ( n348 & n2181 ) | ( n2178 & n2181 ) ;
  assign n2183 = ~n2146 & n2182 ;
  assign n2184 = ( n350 & n2147 ) | ( n350 & n2183 ) | ( n2147 & n2183 ) ;
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  buffer buf_n2187( .i (n2186), .o (n2187) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n282( .i (n281), .o (n282) );
  assign n2188 = ( n247 & ~n282 ) | ( n247 & n2185 ) | ( ~n282 & n2185 ) ;
  assign n2189 = n2131 & ~n2188 ;
  assign n2190 = ( n2132 & n2187 ) | ( n2132 & ~n2189 ) | ( n2187 & ~n2189 ) ;
  assign n2191 = ( n232 & n337 ) | ( n232 & n2062 ) | ( n337 & n2062 ) ;
  assign n2192 = n334 & n1922 ;
  buffer buf_n2193( .i (n432), .o (n2193) );
  assign n2194 = ( n367 & n2192 ) | ( n367 & n2193 ) | ( n2192 & n2193 ) ;
  assign n2195 = ~n2057 & n2194 ;
  assign n2196 = n232 & n2195 ;
  assign n2197 = ( ~n338 & n2191 ) | ( ~n338 & n2196 ) | ( n2191 & n2196 ) ;
  buffer buf_n2198( .i (n2197), .o (n2198) );
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n2200( .i (n2199), .o (n2200) );
  buffer buf_n2201( .i (n96), .o (n2201) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  assign n2203 = ( n610 & ~n1591 ) | ( n610 & n2202 ) | ( ~n1591 & n2202 ) ;
  buffer buf_n2204( .i (n2021), .o (n2204) );
  assign n2205 = n125 & n2204 ;
  assign n2206 = n2024 & n2205 ;
  buffer buf_n2207( .i (n2206), .o (n2207) );
  assign n2215 = n195 & ~n2207 ;
  assign n2216 = ( n1011 & ~n2028 ) | ( n1011 & n2215 ) | ( ~n2028 & n2215 ) ;
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2219( .i (n2057), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  assign n2221 = ( n2202 & ~n2217 ) | ( n2202 & n2220 ) | ( ~n2217 & n2220 ) ;
  assign n2222 = n2203 & ~n2221 ;
  assign n2223 = ( n340 & n2198 ) | ( n340 & n2222 ) | ( n2198 & n2222 ) ;
  assign n2224 = n2162 & ~n2223 ;
  assign n2225 = ( n374 & n2200 ) | ( n374 & ~n2224 ) | ( n2200 & ~n2224 ) ;
  assign n2226 = ~n309 & n2225 ;
  buffer buf_n2227( .i (n2226), .o (n2227) );
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  assign n2229 = n99 & ~n2218 ;
  buffer buf_n2230( .i (n128), .o (n2230) );
  assign n2231 = n1962 & n2230 ;
  buffer buf_n2232( .i (n2231), .o (n2232) );
  assign n2239 = ~n2202 & n2232 ;
  buffer buf_n2240( .i (n2239), .o (n2240) );
  assign n2246 = ( n1261 & ~n2229 ) | ( n1261 & n2240 ) | ( ~n2229 & n2240 ) ;
  assign n2247 = ( n341 & n2162 ) | ( n341 & ~n2246 ) | ( n2162 & ~n2246 ) ;
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  assign n2250 = n343 & ~n2248 ;
  assign n2251 = ( n376 & ~n2249 ) | ( n376 & n2250 ) | ( ~n2249 & n2250 ) ;
  assign n2252 = n2227 | n2251 ;
  assign n2253 = ( ~n444 & n2228 ) | ( ~n444 & n2252 ) | ( n2228 & n2252 ) ;
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  assign n2256 = ~n1295 & n2254 ;
  assign n2257 = ( n270 & ~n340 ) | ( n270 & n372 ) | ( ~n340 & n372 ) ;
  assign n2258 = n341 & ~n2257 ;
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2162), .o (n2261) );
  assign n2262 = ~n342 & n2261 ;
  assign n2263 = ( n309 & n2259 ) | ( n309 & n2262 ) | ( n2259 & n2262 ) ;
  assign n2264 = n2260 | n2263 ;
  buffer buf_n2265( .i (n441), .o (n2265) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  assign n2267 = n2264 & n2266 ;
  buffer buf_n2268( .i (n240), .o (n2268) );
  assign n2269 = ( ~n1897 & n2267 ) | ( ~n1897 & n2268 ) | ( n2267 & n2268 ) ;
  assign n2270 = n1898 & n2269 ;
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n1915( .i (n1914), .o (n1915) );
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  assign n2271 = ( ~n101 & n134 ) | ( ~n101 & n1415 ) | ( n134 & n1415 ) ;
  assign n2272 = n653 & ~n2271 ;
  buffer buf_n2273( .i (n202), .o (n2273) );
  assign n2274 = ( n654 & n2272 ) | ( n654 & ~n2273 ) | ( n2272 & ~n2273 ) ;
  assign n2275 = ~n2244 & n2274 ;
  assign n2276 = ( n834 & n2245 ) | ( n834 & n2275 ) | ( n2245 & n2275 ) ;
  assign n2277 = ( ~n1915 & n2142 ) | ( ~n1915 & n2276 ) | ( n2142 & n2276 ) ;
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  assign n2278 = ( n239 & n2069 ) | ( n239 & ~n2094 ) | ( n2069 & ~n2094 ) ;
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  assign n2279 = n1127 & n1771 ;
  assign n2280 = ~n239 & n2279 ;
  assign n2281 = ( n2070 & ~n2278 ) | ( n2070 & n2280 ) | ( ~n2278 & n2280 ) ;
  assign n2282 = ~n1915 & n2281 ;
  buffer buf_n2283( .i (n2142), .o (n2283) );
  assign n2284 = ( n2277 & n2282 ) | ( n2277 & ~n2283 ) | ( n2282 & ~n2283 ) ;
  assign n2285 = n2270 | n2284 ;
  assign n2286 = ( n2255 & ~n2256 ) | ( n2255 & n2285 ) | ( ~n2256 & n2285 ) ;
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  assign n2289 = ( ~n416 & n483 ) | ( ~n416 & n2287 ) | ( n483 & n2287 ) ;
  buffer buf_n2290( .i (n135), .o (n2290) );
  assign n2291 = ( ~n72 & n2101 ) | ( ~n72 & n2290 ) | ( n2101 & n2290 ) ;
  buffer buf_n2292( .i (n59), .o (n2292) );
  buffer buf_n2293( .i (n156), .o (n2293) );
  assign n2294 = ( n2021 & n2292 ) | ( n2021 & n2293 ) | ( n2292 & n2293 ) ;
  buffer buf_n2295( .i (n2294), .o (n2295) );
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n2297( .i (n2296), .o (n2297) );
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  assign n2307 = ~n2291 & n2306 ;
  buffer buf_n2308( .i (n2307), .o (n2308) );
  buffer buf_n2309( .i (n2308), .o (n2309) );
  buffer buf_n2310( .i (n224), .o (n2310) );
  assign n2311 = n190 & ~n2310 ;
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n2321( .i (n2320), .o (n2321) );
  buffer buf_n2322( .i (n2321), .o (n2322) );
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2325( .i (n2324), .o (n2325) );
  assign n2326 = ( ~n170 & n204 ) | ( ~n170 & n239 ) | ( n204 & n239 ) ;
  assign n2327 = n72 & n2101 ;
  buffer buf_n2328( .i (n2327), .o (n2328) );
  assign n2329 = ( n2325 & n2326 ) | ( n2325 & ~n2328 ) | ( n2326 & ~n2328 ) ;
  assign n2330 = n201 & ~n855 ;
  buffer buf_n2331( .i (n2330), .o (n2331) );
  buffer buf_n2332( .i (n2331), .o (n2332) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  buffer buf_n1983( .i (n1982), .o (n1983) );
  buffer buf_n1984( .i (n1983), .o (n1984) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n1990( .i (n1989), .o (n1990) );
  buffer buf_n1991( .i (n1990), .o (n1991) );
  buffer buf_n1992( .i (n1991), .o (n1992) );
  buffer buf_n1993( .i (n1992), .o (n1993) );
  buffer buf_n1994( .i (n1993), .o (n1994) );
  buffer buf_n1995( .i (n1994), .o (n1995) );
  buffer buf_n1996( .i (n1995), .o (n1996) );
  buffer buf_n1997( .i (n1996), .o (n1997) );
  buffer buf_n1998( .i (n1997), .o (n1998) );
  assign n2333 = ( n71 & n1985 ) | ( n71 & n1998 ) | ( n1985 & n1998 ) ;
  assign n2334 = ~n2331 & n2333 ;
  assign n2335 = ( n73 & n2332 ) | ( n73 & n2334 ) | ( n2332 & n2334 ) ;
  buffer buf_n2336( .i (n2335), .o (n2336) );
  assign n2337 = ( ~n2308 & n2329 ) | ( ~n2308 & n2336 ) | ( n2329 & n2336 ) ;
  assign n2338 = n106 | n2336 ;
  assign n2339 = ( n2309 & n2337 ) | ( n2309 & n2338 ) | ( n2337 & n2338 ) ;
  buffer buf_n2340( .i (n2339), .o (n2340) );
  buffer buf_n2341( .i (n2340), .o (n2341) );
  buffer buf_n2342( .i (n2094), .o (n2342) );
  buffer buf_n2343( .i (n2342), .o (n2343) );
  assign n2344 = ( n346 & n378 ) | ( n346 & n2343 ) | ( n378 & n2343 ) ;
  buffer buf_n2345( .i (n310), .o (n2345) );
  assign n2346 = ( n377 & ~n2342 ) | ( n377 & n2345 ) | ( ~n2342 & n2345 ) ;
  assign n2347 = n346 & n2346 ;
  assign n2348 = ( n1051 & n2344 ) | ( n1051 & ~n2347 ) | ( n2344 & ~n2347 ) ;
  buffer buf_n2349( .i (n479), .o (n2349) );
  assign n2350 = n2348 & n2349 ;
  assign n2351 = ( n447 & n2340 ) | ( n447 & ~n2350 ) | ( n2340 & ~n2350 ) ;
  assign n2352 = n2341 & ~n2351 ;
  assign n2353 = n416 & n2352 ;
  assign n2354 = ( n2288 & ~n2289 ) | ( n2288 & n2353 ) | ( ~n2289 & n2353 ) ;
  buffer buf_n2355( .i (n2354), .o (n2355) );
  buffer buf_n2356( .i (n2355), .o (n2356) );
  buffer buf_n111( .i (n110), .o (n111) );
  assign n2357 = ( n261 & n297 ) | ( n261 & n363 ) | ( n297 & n363 ) ;
  assign n2358 = ( ~n332 & n2148 ) | ( ~n332 & n2357 ) | ( n2148 & n2357 ) ;
  buffer buf_n2359( .i (n2358), .o (n2359) );
  buffer buf_n2362( .i (n365), .o (n2362) );
  assign n2363 = ~n2359 & n2362 ;
  buffer buf_n2364( .i (n2363), .o (n2364) );
  buffer buf_n2365( .i (n2364), .o (n2365) );
  buffer buf_n2360( .i (n2359), .o (n2360) );
  buffer buf_n2361( .i (n2360), .o (n2361) );
  assign n2366 = n2361 | n2364 ;
  assign n2367 = ( ~n369 & n2365 ) | ( ~n369 & n2366 ) | ( n2365 & n2366 ) ;
  buffer buf_n2368( .i (n2367), .o (n2368) );
  buffer buf_n2369( .i (n2368), .o (n2369) );
  assign n2374 = ( ~n1067 & n2032 ) | ( ~n1067 & n2368 ) | ( n2032 & n2368 ) ;
  assign n2375 = n2369 & ~n2374 ;
  buffer buf_n2376( .i (n2375), .o (n2376) );
  buffer buf_n2377( .i (n2376), .o (n2377) );
  assign n2378 = ( n261 & ~n297 ) | ( n261 & n331 ) | ( ~n297 & n331 ) ;
  buffer buf_n2379( .i (n2378), .o (n2379) );
  buffer buf_n2380( .i (n2379), .o (n2380) );
  assign n2381 = ( n299 & n365 ) | ( n299 & ~n2379 ) | ( n365 & ~n2379 ) ;
  assign n2382 = n2380 & ~n2381 ;
  assign n2383 = n1039 | n2382 ;
  buffer buf_n2384( .i (n2383), .o (n2384) );
  buffer buf_n2385( .i (n2384), .o (n2385) );
  buffer buf_n2386( .i (n2385), .o (n2386) );
  buffer buf_n2387( .i (n2386), .o (n2387) );
  buffer buf_n2388( .i (n2387), .o (n2388) );
  assign n2392 = n35 & n2032 ;
  assign n2393 = ( n1261 & ~n2387 ) | ( n1261 & n2392 ) | ( ~n2387 & n2392 ) ;
  assign n2394 = n2388 & n2393 ;
  assign n2395 = ( n33 & n2005 ) | ( n33 & n2384 ) | ( n2005 & n2384 ) ;
  assign n2396 = ( n33 & n1587 ) | ( n33 & ~n2384 ) | ( n1587 & ~n2384 ) ;
  assign n2397 = n2395 & ~n2396 ;
  assign n2398 = n2032 & n2397 ;
  assign n2399 = n1261 & n2398 ;
  buffer buf_n2400( .i (n2399), .o (n2400) );
  assign n2401 = ( ~n2376 & n2394 ) | ( ~n2376 & n2400 ) | ( n2394 & n2400 ) ;
  buffer buf_n2402( .i (n133), .o (n2402) );
  buffer buf_n2403( .i (n2402), .o (n2403) );
  assign n2404 = ~n2400 & n2403 ;
  assign n2405 = ( n2377 & n2401 ) | ( n2377 & ~n2404 ) | ( n2401 & ~n2404 ) ;
  buffer buf_n2406( .i (n169), .o (n2406) );
  assign n2407 = n2405 & n2406 ;
  buffer buf_n2408( .i (n2407), .o (n2408) );
  buffer buf_n2409( .i (n2408), .o (n2409) );
  assign n2410 = n70 | n798 ;
  assign n2411 = n201 & n1204 ;
  assign n2412 = ( n799 & ~n2410 ) | ( n799 & n2411 ) | ( ~n2410 & n2411 ) ;
  buffer buf_n2413( .i (n2412), .o (n2413) );
  buffer buf_n2414( .i (n2413), .o (n2414) );
  assign n2415 = ( n36 & ~n1283 ) | ( n36 & n1595 ) | ( ~n1283 & n1595 ) ;
  buffer buf_n2416( .i (n2415), .o (n2416) );
  assign n2417 = ( n202 & n2403 ) | ( n202 & ~n2416 ) | ( n2403 & ~n2416 ) ;
  assign n2418 = ( ~n38 & n2403 ) | ( ~n38 & n2416 ) | ( n2403 & n2416 ) ;
  assign n2419 = n2417 & ~n2418 ;
  assign n2420 = ~n2413 & n2419 ;
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2391( .i (n2390), .o (n2391) );
  assign n2421 = n2265 & n2391 ;
  assign n2422 = ( n2414 & n2420 ) | ( n2414 & n2421 ) | ( n2420 & n2421 ) ;
  assign n2423 = n2408 | n2422 ;
  assign n2424 = ( n107 & n2409 ) | ( n107 & n2423 ) | ( n2409 & n2423 ) ;
  assign n2425 = n413 & n2424 ;
  buffer buf_n2426( .i (n2425), .o (n2426) );
  buffer buf_n2427( .i (n2426), .o (n2427) );
  assign n2428 = ( n345 & n410 ) | ( n345 & n2342 ) | ( n410 & n2342 ) ;
  buffer buf_n2429( .i (n308), .o (n2429) );
  assign n2430 = n2102 | n2429 ;
  buffer buf_n2431( .i (n2430), .o (n2431) );
  assign n2439 = n345 & ~n2431 ;
  assign n2440 = ( ~n411 & n2428 ) | ( ~n411 & n2439 ) | ( n2428 & n2439 ) ;
  buffer buf_n2441( .i (n2440), .o (n2441) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  assign n2443 = n741 & ~n2441 ;
  buffer buf_n2444( .i (n1586), .o (n2444) );
  assign n2445 = ~n610 & n2444 ;
  assign n2446 = n1587 & ~n2005 ;
  assign n2447 = ( n610 & ~n2444 ) | ( n610 & n2446 ) | ( ~n2444 & n2446 ) ;
  assign n2448 = n2445 | n2447 ;
  assign n2449 = ( n28 & ~n125 ) | ( n28 & n192 ) | ( ~n125 & n192 ) ;
  buffer buf_n2450( .i (n2449), .o (n2450) );
  buffer buf_n2451( .i (n2450), .o (n2451) );
  assign n2452 = n1307 & n2451 ;
  buffer buf_n2453( .i (n2024), .o (n2453) );
  assign n2454 = ( n30 & ~n2450 ) | ( n30 & n2453 ) | ( ~n2450 & n2453 ) ;
  assign n2455 = n2451 | n2454 ;
  assign n2456 = ~n2452 & n2455 ;
  assign n2457 = n2005 & n2456 ;
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  assign n2460 = n35 | n2458 ;
  assign n2461 = ( n2448 & n2459 ) | ( n2448 & n2460 ) | ( n2459 & n2460 ) ;
  buffer buf_n2462( .i (n2461), .o (n2462) );
  assign n2470 = n1655 & n2462 ;
  buffer buf_n2471( .i (n2470), .o (n2471) );
  buffer buf_n2472( .i (n2471), .o (n2472) );
  buffer buf_n2473( .i (n2472), .o (n2473) );
  buffer buf_n2474( .i (n2473), .o (n2474) );
  buffer buf_n2475( .i (n2474), .o (n2475) );
  buffer buf_n2476( .i (n2475), .o (n2476) );
  assign n2477 = ( n2442 & n2443 ) | ( n2442 & n2476 ) | ( n2443 & n2476 ) ;
  assign n2478 = n2426 | n2477 ;
  assign n2479 = ( n111 & n2427 ) | ( n111 & n2478 ) | ( n2427 & n2478 ) ;
  buffer buf_n2480( .i (n2479), .o (n2480) );
  buffer buf_n2481( .i (n2480), .o (n2481) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  assign n2482 = ( ~n248 & n485 ) | ( ~n248 & n2480 ) | ( n485 & n2480 ) ;
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  assign n2483 = n919 | n1230 ;
  buffer buf_n2484( .i (n2483), .o (n2484) );
  buffer buf_n2485( .i (n2484), .o (n2485) );
  assign n2486 = n410 | n2431 ;
  buffer buf_n2487( .i (n2266), .o (n2487) );
  assign n2488 = n2486 | n2487 ;
  assign n2489 = ( n242 & ~n2484 ) | ( n242 & n2488 ) | ( ~n2484 & n2488 ) ;
  buffer buf_n2490( .i (n103), .o (n2490) );
  assign n2491 = ( ~n511 & n2471 ) | ( ~n511 & n2490 ) | ( n2471 & n2490 ) ;
  assign n2492 = n512 & n2491 ;
  assign n2493 = n306 & ~n1595 ;
  assign n2494 = ~n1226 & n2493 ;
  assign n2495 = n2050 & n2494 ;
  buffer buf_n2496( .i (n1655), .o (n2496) );
  assign n2497 = ( n408 & n2495 ) | ( n408 & n2496 ) | ( n2495 & n2496 ) ;
  assign n2498 = ~n2265 & n2497 ;
  assign n2499 = n2342 & n2498 ;
  assign n2500 = ( n2343 & n2492 ) | ( n2343 & n2499 ) | ( n2492 & n2499 ) ;
  assign n2501 = ~n242 & n2500 ;
  assign n2502 = ( n2485 & n2489 ) | ( n2485 & ~n2501 ) | ( n2489 & ~n2501 ) ;
  buffer buf_n2503( .i (n2502), .o (n2503) );
  buffer buf_n2504( .i (n2503), .o (n2504) );
  buffer buf_n2505( .i (n2504), .o (n2505) );
  buffer buf_n2463( .i (n2462), .o (n2463) );
  buffer buf_n2464( .i (n2463), .o (n2464) );
  buffer buf_n2465( .i (n2464), .o (n2465) );
  buffer buf_n2466( .i (n2465), .o (n2466) );
  buffer buf_n2467( .i (n2466), .o (n2467) );
  buffer buf_n2468( .i (n2467), .o (n2468) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  assign n2506 = ~n409 & n2265 ;
  buffer buf_n2507( .i (n2506), .o (n2507) );
  buffer buf_n2508( .i (n2507), .o (n2508) );
  buffer buf_n2509( .i (n2508), .o (n2509) );
  assign n2510 = ( n380 & ~n2468 ) | ( n380 & n2509 ) | ( ~n2468 & n2509 ) ;
  assign n2511 = n2469 & n2510 ;
  buffer buf_n2512( .i (n109), .o (n2512) );
  assign n2513 = ( ~n2503 & n2511 ) | ( ~n2503 & n2512 ) | ( n2511 & n2512 ) ;
  assign n2514 = n281 & ~n2513 ;
  assign n2515 = ( ~n282 & n2505 ) | ( ~n282 & n2514 ) | ( n2505 & n2514 ) ;
  assign n2516 = n485 | n2515 ;
  assign n2517 = ( n2481 & ~n2482 ) | ( n2481 & ~n2516 ) | ( ~n2482 & ~n2516 ) ;
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n2518( .i (n165), .o (n2518) );
  assign n2519 = n270 & n2518 ;
  buffer buf_n2520( .i (n2519), .o (n2520) );
  buffer buf_n2521( .i (n2520), .o (n2521) );
  buffer buf_n2522( .i (n2521), .o (n2522) );
  buffer buf_n2523( .i (n2522), .o (n2523) );
  buffer buf_n2524( .i (n2523), .o (n2524) );
  buffer buf_n2525( .i (n2524), .o (n2525) );
  assign n2526 = ( n207 & n1232 ) | ( n207 & n2525 ) | ( n1232 & n2525 ) ;
  assign n2527 = ~n1233 & n2526 ;
  buffer buf_n2528( .i (n2527), .o (n2528) );
  buffer buf_n2529( .i (n2528), .o (n2529) );
  buffer buf_n315( .i (n314), .o (n315) );
  assign n2530 = ~n378 & n411 ;
  assign n2531 = ~n1448 & n2530 ;
  assign n2532 = ~n348 & n2531 ;
  assign n2533 = n315 & n2532 ;
  assign n2534 = ( n482 & n2528 ) | ( n482 & ~n2533 ) | ( n2528 & ~n2533 ) ;
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  assign n2535 = ( n126 & n1061 ) | ( n126 & ~n1080 ) | ( n1061 & ~n1080 ) ;
  assign n2536 = ~n121 & n188 ;
  buffer buf_n2537( .i (n2536), .o (n2537) );
  assign n2546 = ( n59 & n1986 ) | ( n59 & n2537 ) | ( n1986 & n2537 ) ;
  assign n2547 = ~n1968 & n2546 ;
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  assign n2550 = n2024 | n2548 ;
  assign n2551 = ( ~n2535 & n2549 ) | ( ~n2535 & n2550 ) | ( n2549 & n2550 ) ;
  buffer buf_n2552( .i (n2551), .o (n2552) );
  buffer buf_n2564( .i (n2193), .o (n2564) );
  assign n2565 = n2552 & n2564 ;
  buffer buf_n2566( .i (n2565), .o (n2566) );
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n2568( .i (n2567), .o (n2568) );
  buffer buf_n2569( .i (n2568), .o (n2569) );
  buffer buf_n2570( .i (n2569), .o (n2570) );
  buffer buf_n2571( .i (n2570), .o (n2571) );
  buffer buf_n2572( .i (n2571), .o (n2572) );
  buffer buf_n2573( .i (n2572), .o (n2573) );
  buffer buf_n2574( .i (n2573), .o (n2574) );
  buffer buf_n2575( .i (n2574), .o (n2575) );
  buffer buf_n2576( .i (n2575), .o (n2576) );
  assign n2577 = ( n44 & ~n765 ) | ( n44 & n2576 ) | ( ~n765 & n2576 ) ;
  assign n2578 = n766 & n2577 ;
  assign n2579 = ~n482 & n2578 ;
  assign n2580 = ( n2529 & ~n2534 ) | ( n2529 & n2579 ) | ( ~n2534 & n2579 ) ;
  buffer buf_n2581( .i (n2580), .o (n2581) );
  buffer buf_n2582( .i (n2581), .o (n2582) );
  buffer buf_n2583( .i (n2293), .o (n2583) );
  buffer buf_n2584( .i (n2583), .o (n2584) );
  assign n2585 = n62 | n2584 ;
  assign n2586 = ~n1061 & n2584 ;
  assign n2587 = n2585 & ~n2586 ;
  buffer buf_n2588( .i (n2587), .o (n2588) );
  buffer buf_n2589( .i (n2588), .o (n2589) );
  buffer buf_n2590( .i (n2589), .o (n2590) );
  buffer buf_n2591( .i (n2590), .o (n2591) );
  buffer buf_n2592( .i (n2591), .o (n2592) );
  buffer buf_n2593( .i (n2592), .o (n2593) );
  buffer buf_n2594( .i (n2593), .o (n2594) );
  buffer buf_n2595( .i (n2594), .o (n2595) );
  buffer buf_n2596( .i (n2595), .o (n2596) );
  buffer buf_n2597( .i (n2596), .o (n2597) );
  buffer buf_n2598( .i (n2597), .o (n2598) );
  buffer buf_n2599( .i (n2598), .o (n2599) );
  assign n2600 = n1448 & n2599 ;
  assign n2601 = ( n765 & n2349 ) | ( n765 & ~n2600 ) | ( n2349 & ~n2600 ) ;
  assign n2602 = n766 & ~n2601 ;
  buffer buf_n2603( .i (n2602), .o (n2603) );
  buffer buf_n2604( .i (n2603), .o (n2604) );
  buffer buf_n47( .i (n46), .o (n47) );
  assign n2605 = ( n47 & n144 ) | ( n47 & ~n2603 ) | ( n144 & ~n2603 ) ;
  buffer buf_n2606( .i (n1932), .o (n2606) );
  buffer buf_n2607( .i (n589), .o (n2607) );
  assign n2608 = n2606 & ~n2607 ;
  assign n2609 = n305 & n506 ;
  assign n2610 = n2606 | n2609 ;
  assign n2611 = ~n2608 & n2610 ;
  buffer buf_n2612( .i (n2611), .o (n2612) );
  assign n2613 = n169 | n2612 ;
  assign n2614 = ~n295 & n329 ;
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  buffer buf_n2617( .i (n2616), .o (n2617) );
  buffer buf_n2618( .i (n2617), .o (n2618) );
  buffer buf_n2619( .i (n2618), .o (n2619) );
  buffer buf_n2620( .i (n2619), .o (n2620) );
  buffer buf_n2621( .i (n2620), .o (n2621) );
  buffer buf_n2622( .i (n2621), .o (n2622) );
  buffer buf_n2623( .i (n2622), .o (n2623) );
  buffer buf_n2624( .i (n2623), .o (n2624) );
  buffer buf_n2625( .i (n2624), .o (n2625) );
  assign n2633 = n2157 & n2625 ;
  assign n2634 = ~n916 & n2633 ;
  buffer buf_n2635( .i (n168), .o (n2635) );
  assign n2636 = ~n2634 & n2635 ;
  assign n2637 = n2613 & ~n2636 ;
  buffer buf_n2638( .i (n2637), .o (n2638) );
  buffer buf_n2639( .i (n2638), .o (n2639) );
  buffer buf_n2640( .i (n362), .o (n2640) );
  assign n2641 = n396 | n2640 ;
  buffer buf_n2642( .i (n2641), .o (n2642) );
  buffer buf_n2643( .i (n2642), .o (n2643) );
  buffer buf_n2644( .i (n2643), .o (n2644) );
  buffer buf_n2645( .i (n2644), .o (n2645) );
  buffer buf_n2646( .i (n2645), .o (n2646) );
  buffer buf_n2647( .i (n2646), .o (n2647) );
  buffer buf_n2648( .i (n2647), .o (n2648) );
  buffer buf_n2649( .i (n2648), .o (n2649) );
  buffer buf_n2650( .i (n2649), .o (n2650) );
  buffer buf_n2651( .i (n2650), .o (n2651) );
  buffer buf_n2652( .i (n2651), .o (n2652) );
  buffer buf_n2653( .i (n2652), .o (n2653) );
  buffer buf_n2654( .i (n2653), .o (n2654) );
  buffer buf_n2370( .i (n2369), .o (n2370) );
  assign n2658 = n403 & ~n2444 ;
  buffer buf_n2659( .i (n2658), .o (n2659) );
  assign n2663 = ( n1595 & n2369 ) | ( n1595 & ~n2659 ) | ( n2369 & ~n2659 ) ;
  assign n2664 = n2370 & ~n2663 ;
  buffer buf_n2665( .i (n2664), .o (n2665) );
  buffer buf_n2666( .i (n2665), .o (n2666) );
  buffer buf_n2667( .i (n2666), .o (n2667) );
  buffer buf_n2626( .i (n2625), .o (n2626) );
  buffer buf_n2627( .i (n2626), .o (n2627) );
  assign n2668 = ~n263 & n2584 ;
  buffer buf_n2669( .i (n2668), .o (n2669) );
  buffer buf_n2670( .i (n2669), .o (n2670) );
  buffer buf_n2671( .i (n2670), .o (n2671) );
  buffer buf_n2672( .i (n2671), .o (n2672) );
  buffer buf_n2673( .i (n2672), .o (n2673) );
  buffer buf_n2674( .i (n2673), .o (n2674) );
  buffer buf_n2675( .i (n2674), .o (n2675) );
  buffer buf_n2676( .i (n1594), .o (n2676) );
  buffer buf_n2677( .i (n2676), .o (n2677) );
  assign n2678 = n2675 & n2677 ;
  buffer buf_n2679( .i (n2678), .o (n2679) );
  assign n2682 = ( n2627 & n2665 ) | ( n2627 & n2679 ) | ( n2665 & n2679 ) ;
  assign n2683 = n2653 | n2682 ;
  assign n2684 = ( ~n2654 & n2667 ) | ( ~n2654 & n2683 ) | ( n2667 & n2683 ) ;
  assign n2685 = n73 & n1605 ;
  buffer buf_n2686( .i (n2685), .o (n2686) );
  buffer buf_n2687( .i (n1571), .o (n2687) );
  assign n2688 = ( n2684 & ~n2686 ) | ( n2684 & n2687 ) | ( ~n2686 & n2687 ) ;
  assign n2689 = ( n2638 & ~n2686 ) | ( n2638 & n2687 ) | ( ~n2686 & n2687 ) ;
  assign n2690 = ( n2639 & n2688 ) | ( n2639 & ~n2689 ) | ( n2688 & ~n2689 ) ;
  buffer buf_n2691( .i (n2690), .o (n2691) );
  buffer buf_n2692( .i (n2691), .o (n2692) );
  assign n2693 = ( ~n109 & n447 ) | ( ~n109 & n2691 ) | ( n447 & n2691 ) ;
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  assign n2694 = n377 & n2629 ;
  assign n2695 = ( n411 & n2687 ) | ( n411 & n2694 ) | ( n2687 & n2694 ) ;
  assign n2696 = ~n479 & n2695 ;
  assign n2697 = n103 | n638 ;
  assign n2698 = n1604 & n2612 ;
  assign n2699 = ( n639 & ~n2697 ) | ( n639 & n2698 ) | ( ~n2697 & n2698 ) ;
  assign n2700 = n74 & n2699 ;
  buffer buf_n2701( .i (n2700), .o (n2701) );
  buffer buf_n2702( .i (n2701), .o (n2702) );
  buffer buf_n920( .i (n919), .o (n920) );
  assign n2703 = ~n105 & n171 ;
  assign n2704 = ~n920 & n2703 ;
  assign n2705 = n2701 | n2704 ;
  assign n2706 = ( n2696 & n2702 ) | ( n2696 & n2705 ) | ( n2702 & n2705 ) ;
  buffer buf_n2707( .i (n446), .o (n2707) );
  assign n2708 = n2706 & ~n2707 ;
  assign n2709 = ( n2692 & ~n2693 ) | ( n2692 & n2708 ) | ( ~n2693 & n2708 ) ;
  assign n2710 = n144 & n2709 ;
  assign n2711 = ( n2604 & n2605 ) | ( n2604 & n2710 ) | ( n2605 & n2710 ) ;
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  assign n2712 = ( n34 & ~n505 ) | ( n34 & n2566 ) | ( ~n505 & n2566 ) ;
  assign n2713 = n506 & n2712 ;
  buffer buf_n2714( .i (n2713), .o (n2714) );
  buffer buf_n2715( .i (n2714), .o (n2715) );
  buffer buf_n2716( .i (n2715), .o (n2716) );
  buffer buf_n1846( .i (n1845), .o (n1846) );
  buffer buf_n1847( .i (n1846), .o (n1847) );
  assign n2717 = n370 & n1847 ;
  buffer buf_n2718( .i (n2220), .o (n2718) );
  assign n2719 = ( n404 & n2717 ) | ( n404 & n2718 ) | ( n2717 & n2718 ) ;
  buffer buf_n2720( .i (n2718), .o (n2720) );
  assign n2721 = n2719 & ~n2720 ;
  assign n2722 = ( ~n1226 & n2714 ) | ( ~n1226 & n2721 ) | ( n2714 & n2721 ) ;
  assign n2723 = n1017 | n2722 ;
  assign n2724 = ( ~n1018 & n2716 ) | ( ~n1018 & n2723 ) | ( n2716 & n2723 ) ;
  buffer buf_n2725( .i (n2724), .o (n2725) );
  buffer buf_n2726( .i (n2725), .o (n2726) );
  buffer buf_n2727( .i (n236), .o (n2727) );
  buffer buf_n2728( .i (n2727), .o (n2728) );
  buffer buf_n2729( .i (n2728), .o (n2729) );
  buffer buf_n2730( .i (n2729), .o (n2730) );
  buffer buf_n2731( .i (n2094), .o (n2731) );
  assign n2732 = ( n2725 & n2730 ) | ( n2725 & ~n2731 ) | ( n2730 & ~n2731 ) ;
  assign n2733 = n265 | n301 ;
  buffer buf_n2734( .i (n2733), .o (n2734) );
  buffer buf_n2735( .i (n2734), .o (n2735) );
  buffer buf_n2736( .i (n2735), .o (n2736) );
  buffer buf_n2737( .i (n2736), .o (n2737) );
  assign n2742 = n405 | n2737 ;
  buffer buf_n2743( .i (n371), .o (n2743) );
  buffer buf_n2744( .i (n2743), .o (n2744) );
  assign n2745 = ( n2163 & n2742 ) | ( n2163 & ~n2744 ) | ( n2742 & ~n2744 ) ;
  assign n2746 = n2261 | n2745 ;
  assign n2747 = n1018 | n2746 ;
  assign n2748 = n1229 | n2747 ;
  assign n2749 = n2730 | n2748 ;
  assign n2750 = ( ~n2726 & n2732 ) | ( ~n2726 & n2749 ) | ( n2732 & n2749 ) ;
  buffer buf_n2751( .i (n2750), .o (n2751) );
  buffer buf_n2752( .i (n2751), .o (n2752) );
  buffer buf_n2753( .i (n2752), .o (n2753) );
  buffer buf_n2553( .i (n2552), .o (n2553) );
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2555( .i (n2554), .o (n2555) );
  buffer buf_n2556( .i (n2555), .o (n2556) );
  buffer buf_n2557( .i (n2556), .o (n2557) );
  buffer buf_n2558( .i (n2557), .o (n2558) );
  buffer buf_n2559( .i (n2558), .o (n2559) );
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  buffer buf_n2563( .i (n2562), .o (n2563) );
  assign n2754 = ( n378 & n2507 ) | ( n378 & ~n2562 ) | ( n2507 & ~n2562 ) ;
  assign n2755 = n2563 & n2754 ;
  assign n2756 = ( n44 & ~n2751 ) | ( n44 & n2755 ) | ( ~n2751 & n2755 ) ;
  assign n2757 = n279 & ~n2756 ;
  assign n2758 = ( ~n280 & n2753 ) | ( ~n280 & n2757 ) | ( n2753 & n2757 ) ;
  assign n2759 = n32 & ~n468 ;
  assign n2760 = ( n2219 & ~n2589 ) | ( n2219 & n2759 ) | ( ~n2589 & n2759 ) ;
  assign n2761 = n2590 & n2760 ;
  buffer buf_n2762( .i (n2761), .o (n2762) );
  buffer buf_n2763( .i (n2762), .o (n2763) );
  buffer buf_n2764( .i (n153), .o (n2764) );
  assign n2765 = ~n223 & n2764 ;
  buffer buf_n2766( .i (n2765), .o (n2766) );
  assign n2780 = n59 & ~n2766 ;
  assign n2781 = n990 & ~n2780 ;
  assign n2782 = n2018 & n2781 ;
  buffer buf_n2783( .i (n2782), .o (n2783) );
  buffer buf_n2784( .i (n2783), .o (n2784) );
  assign n2785 = ( n192 & n2312 ) | ( n192 & ~n2583 ) | ( n2312 & ~n2583 ) ;
  buffer buf_n2786( .i (n2785), .o (n2786) );
  assign n2790 = n2783 | n2786 ;
  assign n2791 = ( n1821 & n2784 ) | ( n1821 & n2790 ) | ( n2784 & n2790 ) ;
  buffer buf_n2792( .i (n2791), .o (n2792) );
  assign n2794 = n469 & n2792 ;
  assign n2795 = ~n2220 & n2794 ;
  buffer buf_n2796( .i (n2795), .o (n2796) );
  buffer buf_n2793( .i (n2792), .o (n2793) );
  assign n2800 = n468 & ~n1845 ;
  assign n2801 = ( n2219 & n2792 ) | ( n2219 & ~n2800 ) | ( n2792 & ~n2800 ) ;
  assign n2802 = n2793 & ~n2801 ;
  buffer buf_n2803( .i (n2802), .o (n2803) );
  assign n2804 = ( ~n2762 & n2796 ) | ( ~n2762 & n2803 ) | ( n2796 & n2803 ) ;
  assign n2805 = n405 & ~n2803 ;
  assign n2806 = ( n2763 & n2804 ) | ( n2763 & ~n2805 ) | ( n2804 & ~n2805 ) ;
  assign n2807 = n2261 & ~n2806 ;
  buffer buf_n2797( .i (n2796), .o (n2797) );
  buffer buf_n2808( .i (n339), .o (n2808) );
  buffer buf_n2809( .i (n2808), .o (n2809) );
  assign n2810 = n2797 & n2809 ;
  assign n2811 = n2261 | n2810 ;
  assign n2812 = ~n2807 & n2811 ;
  buffer buf_n2813( .i (n2133), .o (n2813) );
  buffer buf_n2814( .i (n2813), .o (n2814) );
  assign n2815 = n2812 & n2814 ;
  buffer buf_n2816( .i (n2815), .o (n2816) );
  buffer buf_n2817( .i (n2816), .o (n2817) );
  assign n2818 = ( n890 & n2220 ) | ( n890 & ~n2590 ) | ( n2220 & ~n2590 ) ;
  assign n2819 = n2591 & n2818 ;
  assign n2820 = ~n235 & n2819 ;
  assign n2821 = n1204 & n2820 ;
  buffer buf_n2822( .i (n2821), .o (n2822) );
  buffer buf_n2823( .i (n2822), .o (n2823) );
  buffer buf_n2824( .i (n2823), .o (n2824) );
  buffer buf_n2798( .i (n2797), .o (n2798) );
  buffer buf_n2799( .i (n2798), .o (n2799) );
  assign n2825 = ( n2799 & ~n2813 ) | ( n2799 & n2822 ) | ( ~n2813 & n2822 ) ;
  assign n2826 = n310 & ~n2825 ;
  assign n2827 = ( n2345 & n2824 ) | ( n2345 & ~n2826 ) | ( n2824 & ~n2826 ) ;
  assign n2828 = n2816 | n2827 ;
  assign n2829 = ( n514 & n2817 ) | ( n514 & n2828 ) | ( n2817 & n2828 ) ;
  assign n2830 = n141 & n2829 ;
  buffer buf_n2831( .i (n2830), .o (n2831) );
  buffer buf_n2832( .i (n2831), .o (n2832) );
  assign n2833 = n482 & ~n2831 ;
  assign n2834 = ( n2758 & ~n2832 ) | ( n2758 & n2833 ) | ( ~n2832 & n2833 ) ;
  buffer buf_n2835( .i (n2834), .o (n2835) );
  assign n2836 = ( n2581 & ~n2711 ) | ( n2581 & n2835 ) | ( ~n2711 & n2835 ) ;
  assign n2837 = ~n248 & n2835 ;
  assign n2838 = ( n2582 & ~n2836 ) | ( n2582 & ~n2837 ) | ( ~n2836 & ~n2837 ) ;
  buffer buf_n2839( .i (n481), .o (n2839) );
  assign n2840 = n415 | n2839 ;
  assign n2841 = n449 | n2840 ;
  buffer buf_n2842( .i (n2841), .o (n2842) );
  assign n2843 = n300 | n575 ;
  buffer buf_n2844( .i (n2843), .o (n2844) );
  buffer buf_n2845( .i (n2844), .o (n2845) );
  buffer buf_n2846( .i (n2845), .o (n2846) );
  buffer buf_n2847( .i (n2846), .o (n2847) );
  buffer buf_n2848( .i (n2847), .o (n2848) );
  buffer buf_n2849( .i (n2848), .o (n2849) );
  buffer buf_n2850( .i (n2849), .o (n2850) );
  buffer buf_n2851( .i (n2850), .o (n2851) );
  buffer buf_n2852( .i (n2851), .o (n2852) );
  buffer buf_n2853( .i (n2852), .o (n2853) );
  buffer buf_n2854( .i (n2853), .o (n2854) );
  buffer buf_n2855( .i (n2854), .o (n2855) );
  buffer buf_n2856( .i (n2855), .o (n2856) );
  buffer buf_n2857( .i (n2856), .o (n2857) );
  buffer buf_n2858( .i (n2857), .o (n2858) );
  buffer buf_n2859( .i (n2858), .o (n2859) );
  buffer buf_n2860( .i (n2859), .o (n2860) );
  buffer buf_n2861( .i (n2860), .o (n2861) );
  assign n2862 = n2842 | n2861 ;
  assign n2863 = ~n328 & n523 ;
  assign n2864 = n1349 & n2863 ;
  buffer buf_n2865( .i (n2864), .o (n2865) );
  buffer buf_n2866( .i (n2865), .o (n2866) );
  buffer buf_n2867( .i (n2866), .o (n2867) );
  assign n2868 = ( n224 & n329 ) | ( n224 & ~n427 ) | ( n329 & ~n427 ) ;
  buffer buf_n2869( .i (n460), .o (n2869) );
  assign n2870 = ( n224 & n329 ) | ( n224 & ~n2869 ) | ( n329 & ~n2869 ) ;
  assign n2871 = ~n2868 & n2870 ;
  assign n2872 = ( ~n27 & n2865 ) | ( ~n27 & n2871 ) | ( n2865 & n2871 ) ;
  buffer buf_n2873( .i (n188), .o (n2873) );
  buffer buf_n2874( .i (n2873), .o (n2874) );
  buffer buf_n2875( .i (n2874), .o (n2875) );
  buffer buf_n2876( .i (n2875), .o (n2876) );
  assign n2877 = ~n2872 & n2876 ;
  assign n2878 = ( n193 & n2867 ) | ( n193 & ~n2877 ) | ( n2867 & ~n2877 ) ;
  buffer buf_n2879( .i (n2878), .o (n2879) );
  buffer buf_n2880( .i (n2879), .o (n2880) );
  assign n2881 = n261 & ~n2640 ;
  buffer buf_n2882( .i (n2881), .o (n2882) );
  buffer buf_n2883( .i (n2882), .o (n2883) );
  buffer buf_n2884( .i (n2883), .o (n2884) );
  buffer buf_n2886( .i (n299), .o (n2886) );
  buffer buf_n2887( .i (n2886), .o (n2887) );
  assign n2888 = ( ~n2879 & n2884 ) | ( ~n2879 & n2887 ) | ( n2884 & n2887 ) ;
  assign n2889 = n2880 & n2888 ;
  buffer buf_n2890( .i (n2889), .o (n2890) );
  buffer buf_n2891( .i (n2890), .o (n2891) );
  buffer buf_n2892( .i (n2891), .o (n2892) );
  assign n2893 = n1357 & ~n2734 ;
  assign n2894 = ( n533 & n2890 ) | ( n533 & n2893 ) | ( n2890 & n2893 ) ;
  assign n2895 = n2047 & ~n2894 ;
  assign n2896 = ( n2048 & n2892 ) | ( n2048 & ~n2895 ) | ( n2892 & ~n2895 ) ;
  assign n2897 = n70 & n2896 ;
  buffer buf_n2898( .i (n2897), .o (n2898) );
  buffer buf_n2899( .i (n2898), .o (n2899) );
  buffer buf_n2371( .i (n2370), .o (n2371) );
  assign n2900 = ( ~n1578 & n1935 ) | ( ~n1578 & n2370 ) | ( n1935 & n2370 ) ;
  assign n2901 = n2371 & ~n2900 ;
  assign n2902 = n2898 | n2901 ;
  assign n2903 = ( ~n204 & n2899 ) | ( ~n204 & n2902 ) | ( n2899 & n2902 ) ;
  assign n2904 = n171 | n2903 ;
  buffer buf_n2905( .i (n331), .o (n2905) );
  assign n2906 = n262 & ~n2905 ;
  buffer buf_n2907( .i (n2906), .o (n2907) );
  buffer buf_n2908( .i (n260), .o (n2908) );
  buffer buf_n2909( .i (n330), .o (n2909) );
  assign n2910 = n2908 | n2909 ;
  buffer buf_n2911( .i (n2910), .o (n2911) );
  buffer buf_n2912( .i (n2911), .o (n2912) );
  assign n2913 = ( ~n264 & n2907 ) | ( ~n264 & n2912 ) | ( n2907 & n2912 ) ;
  buffer buf_n2914( .i (n2913), .o (n2914) );
  buffer buf_n2915( .i (n2914), .o (n2915) );
  buffer buf_n2916( .i (n2915), .o (n2916) );
  buffer buf_n2917( .i (n2916), .o (n2917) );
  buffer buf_n2918( .i (n2917), .o (n2918) );
  assign n2922 = ~n370 & n470 ;
  assign n2923 = ( n2718 & n2917 ) | ( n2718 & ~n2922 ) | ( n2917 & ~n2922 ) ;
  assign n2924 = n2918 & ~n2923 ;
  assign n2925 = n307 & n2924 ;
  buffer buf_n2926( .i (n2677), .o (n2926) );
  assign n2927 = ( n2727 & n2925 ) | ( n2727 & n2926 ) | ( n2925 & n2926 ) ;
  assign n2928 = ~n2273 & n2927 ;
  assign n2929 = ~n73 & n2928 ;
  buffer buf_n2930( .i (n2406), .o (n2930) );
  assign n2931 = ~n2929 & n2930 ;
  assign n2932 = n2904 & ~n2931 ;
  assign n2933 = n107 & ~n2932 ;
  buffer buf_n2919( .i (n2918), .o (n2919) );
  buffer buf_n2920( .i (n2919), .o (n2920) );
  assign n2934 = n472 | n2743 ;
  assign n2935 = ( n2163 & n2919 ) | ( n2163 & n2934 ) | ( n2919 & n2934 ) ;
  assign n2936 = n2920 & ~n2935 ;
  assign n2937 = n2429 & n2936 ;
  buffer buf_n2938( .i (n2273), .o (n2938) );
  assign n2939 = ( n2729 & n2937 ) | ( n2729 & n2938 ) | ( n2937 & n2938 ) ;
  assign n2940 = ~n205 & n2939 ;
  assign n2941 = n172 & n2940 ;
  buffer buf_n2942( .i (n106), .o (n2942) );
  assign n2943 = n2941 | n2942 ;
  assign n2944 = ~n2933 & n2943 ;
  assign n2945 = n142 & ~n2944 ;
  assign n2946 = n257 & n293 ;
  buffer buf_n2947( .i (n2946), .o (n2947) );
  buffer buf_n2948( .i (n2947), .o (n2948) );
  buffer buf_n2949( .i (n2948), .o (n2949) );
  buffer buf_n2950( .i (n2949), .o (n2950) );
  buffer buf_n2951( .i (n2950), .o (n2951) );
  buffer buf_n2952( .i (n2951), .o (n2952) );
  buffer buf_n2953( .i (n2952), .o (n2953) );
  buffer buf_n2954( .i (n2953), .o (n2954) );
  buffer buf_n2955( .i (n2954), .o (n2955) );
  buffer buf_n2956( .i (n2955), .o (n2956) );
  buffer buf_n2957( .i (n2956), .o (n2957) );
  assign n2964 = ~n2086 & n2957 ;
  buffer buf_n2965( .i (n2964), .o (n2965) );
  buffer buf_n2966( .i (n2965), .o (n2966) );
  buffer buf_n2967( .i (n2966), .o (n2967) );
  buffer buf_n2968( .i (n2967), .o (n2968) );
  buffer buf_n2969( .i (n474), .o (n2969) );
  assign n2970 = ( n1018 & n2967 ) | ( n1018 & n2969 ) | ( n2967 & n2969 ) ;
  buffer buf_n2738( .i (n2737), .o (n2738) );
  buffer buf_n2739( .i (n2738), .o (n2739) );
  assign n2971 = n230 & n2055 ;
  buffer buf_n2972( .i (n2971), .o (n2972) );
  buffer buf_n2973( .i (n2972), .o (n2973) );
  buffer buf_n2974( .i (n2973), .o (n2974) );
  buffer buf_n2975( .i (n2974), .o (n2975) );
  buffer buf_n2976( .i (n2975), .o (n2976) );
  assign n2980 = ( n2677 & n2738 ) | ( n2677 & n2976 ) | ( n2738 & n2976 ) ;
  assign n2981 = ~n2739 & n2980 ;
  assign n2982 = ~n2969 & n2981 ;
  assign n2983 = ( n2968 & ~n2970 ) | ( n2968 & n2982 ) | ( ~n2970 & n2982 ) ;
  assign n2984 = n345 & n2983 ;
  buffer buf_n2985( .i (n2102), .o (n2985) );
  buffer buf_n2986( .i (n2985), .o (n2986) );
  buffer buf_n2987( .i (n2986), .o (n2987) );
  assign n2988 = ( n2487 & n2984 ) | ( n2487 & n2987 ) | ( n2984 & n2987 ) ;
  assign n2989 = ~n1448 & n2988 ;
  assign n2990 = ~n108 & n2989 ;
  assign n2991 = n142 | n2990 ;
  assign n2992 = ~n2945 & n2991 ;
  assign n2993 = n416 & n2992 ;
  buffer buf_n2994( .i (n2993), .o (n2994) );
  buffer buf_n2995( .i (n2994), .o (n2995) );
  assign n2996 = n1229 | n2729 ;
  buffer buf_n2997( .i (n2996), .o (n2997) );
  buffer buf_n2998( .i (n2997), .o (n2998) );
  buffer buf_n2999( .i (n2998), .o (n2999) );
  buffer buf_n3000( .i (n2999), .o (n3000) );
  buffer buf_n3001( .i (n3000), .o (n3001) );
  buffer buf_n3002( .i (n3001), .o (n3002) );
  assign n3003 = ( ~n211 & n281 ) | ( ~n211 & n3002 ) | ( n281 & n3002 ) ;
  assign n3004 = n212 | n3003 ;
  assign n3005 = ~n2994 & n3004 ;
  assign n3006 = ( ~n2862 & n2995 ) | ( ~n2862 & ~n3005 ) | ( n2995 & ~n3005 ) ;
  buffer buf_n2432( .i (n2431), .o (n2432) );
  buffer buf_n2433( .i (n2432), .o (n2433) );
  buffer buf_n2434( .i (n2433), .o (n2434) );
  buffer buf_n2435( .i (n2434), .o (n2435) );
  buffer buf_n2436( .i (n2435), .o (n2436) );
  buffer buf_n2437( .i (n2436), .o (n2437) );
  buffer buf_n2438( .i (n2437), .o (n2438) );
  assign n3007 = n282 | n2438 ;
  assign n3008 = n2842 | n3007 ;
  buffer buf_n2630( .i (n2629), .o (n2630) );
  buffer buf_n2680( .i (n2679), .o (n2680) );
  buffer buf_n2681( .i (n2680), .o (n2681) );
  buffer buf_n3009( .i (n2744), .o (n3009) );
  buffer buf_n3010( .i (n2163), .o (n3010) );
  assign n3011 = n3009 & ~n3010 ;
  assign n3012 = ~n2969 & n3011 ;
  buffer buf_n3013( .i (n3012), .o (n3013) );
  assign n3015 = n2681 & n3013 ;
  assign n3016 = ( n1231 & n2630 ) | ( n1231 & n3015 ) | ( n2630 & n3015 ) ;
  assign n3017 = ~n1232 & n3016 ;
  buffer buf_n3018( .i (n3017), .o (n3018) );
  buffer buf_n3019( .i (n3018), .o (n3019) );
  assign n3020 = ( n29 & n333 ) | ( n29 & ~n365 ) | ( n333 & ~n365 ) ;
  assign n3021 = ( ~n2362 & n2453 ) | ( ~n2362 & n3020 ) | ( n2453 & n3020 ) ;
  buffer buf_n3022( .i (n3021), .o (n3022) );
  buffer buf_n3025( .i (n2362), .o (n3025) );
  buffer buf_n3026( .i (n3025), .o (n3026) );
  assign n3027 = n3022 & n3026 ;
  buffer buf_n3028( .i (n3027), .o (n3028) );
  buffer buf_n3029( .i (n3028), .o (n3029) );
  buffer buf_n3023( .i (n3022), .o (n3023) );
  buffer buf_n3024( .i (n3023), .o (n3024) );
  assign n3030 = n3024 & ~n3028 ;
  buffer buf_n3031( .i (n369), .o (n3031) );
  buffer buf_n3032( .i (n3031), .o (n3032) );
  assign n3033 = ( ~n3029 & n3030 ) | ( ~n3029 & n3032 ) | ( n3030 & n3032 ) ;
  buffer buf_n3034( .i (n3033), .o (n3034) );
  buffer buf_n3035( .i (n3034), .o (n3035) );
  buffer buf_n3036( .i (n471), .o (n3036) );
  assign n3037 = n306 & ~n3036 ;
  buffer buf_n3038( .i (n2720), .o (n3038) );
  assign n3039 = ( n3034 & n3037 ) | ( n3034 & n3038 ) | ( n3037 & n3038 ) ;
  assign n3040 = ~n3035 & n3039 ;
  buffer buf_n3041( .i (n3040), .o (n3041) );
  buffer buf_n3042( .i (n3041), .o (n3042) );
  buffer buf_n3043( .i (n102), .o (n3043) );
  assign n3044 = n2813 & n3043 ;
  assign n3045 = ( n2938 & ~n3041 ) | ( n2938 & n3044 ) | ( ~n3041 & n3044 ) ;
  assign n3046 = n3042 & n3045 ;
  buffer buf_n3047( .i (n3046), .o (n3047) );
  buffer buf_n3048( .i (n3047), .o (n3048) );
  buffer buf_n3049( .i (n74), .o (n3049) );
  buffer buf_n3050( .i (n3049), .o (n3050) );
  assign n3051 = ( n140 & ~n3047 ) | ( n140 & n3050 ) | ( ~n3047 & n3050 ) ;
  buffer buf_n2372( .i (n2371), .o (n2372) );
  buffer buf_n2373( .i (n2372), .o (n2373) );
  assign n3052 = ( ~n638 & n2372 ) | ( ~n638 & n2969 ) | ( n2372 & n2969 ) ;
  assign n3053 = n2373 & ~n3052 ;
  assign n3054 = ( n105 & ~n2266 ) | ( n105 & n3053 ) | ( ~n2266 & n3053 ) ;
  assign n3055 = n469 & n2621 ;
  assign n3056 = n3031 & n3055 ;
  buffer buf_n3057( .i (n152), .o (n3057) );
  assign n3058 = ~n56 & n3057 ;
  buffer buf_n3059( .i (n3058), .o (n3059) );
  buffer buf_n3060( .i (n3059), .o (n3060) );
  buffer buf_n3061( .i (n3060), .o (n3061) );
  buffer buf_n3062( .i (n3061), .o (n3062) );
  buffer buf_n3063( .i (n3062), .o (n3063) );
  buffer buf_n3064( .i (n3063), .o (n3064) );
  buffer buf_n3065( .i (n3064), .o (n3065) );
  buffer buf_n3066( .i (n3065), .o (n3066) );
  buffer buf_n3067( .i (n3066), .o (n3067) );
  buffer buf_n3068( .i (n3067), .o (n3068) );
  buffer buf_n3069( .i (n3068), .o (n3069) );
  assign n3072 = n3056 & n3069 ;
  assign n3073 = ~n914 & n3072 ;
  buffer buf_n3074( .i (n3073), .o (n3074) );
  buffer buf_n3075( .i (n3074), .o (n3075) );
  buffer buf_n3076( .i (n3075), .o (n3076) );
  assign n3077 = ~n330 & n462 ;
  assign n3078 = ~n2640 & n3077 ;
  buffer buf_n3079( .i (n3078), .o (n3079) );
  buffer buf_n3080( .i (n3079), .o (n3080) );
  buffer buf_n3081( .i (n3080), .o (n3081) );
  buffer buf_n3082( .i (n3081), .o (n3082) );
  buffer buf_n3083( .i (n3082), .o (n3083) );
  buffer buf_n3084( .i (n3083), .o (n3084) );
  buffer buf_n3085( .i (n2004), .o (n3085) );
  assign n3086 = n632 & ~n3085 ;
  assign n3087 = n3084 & n3086 ;
  buffer buf_n3088( .i (n3087), .o (n3088) );
  assign n3089 = ( n1283 & n3036 ) | ( n1283 & ~n3088 ) | ( n3036 & ~n3088 ) ;
  buffer buf_n3090( .i (n2148), .o (n3090) );
  assign n3091 = ( n333 & n2584 ) | ( n333 & ~n3090 ) | ( n2584 & ~n3090 ) ;
  buffer buf_n3092( .i (n2876), .o (n3092) );
  buffer buf_n3093( .i (n3092), .o (n3093) );
  assign n3094 = ( ~n2362 & n3091 ) | ( ~n2362 & n3093 ) | ( n3091 & n3093 ) ;
  buffer buf_n3095( .i (n3094), .o (n3095) );
  assign n3098 = n3026 & n3095 ;
  buffer buf_n3099( .i (n3098), .o (n3099) );
  buffer buf_n3100( .i (n3099), .o (n3100) );
  buffer buf_n3096( .i (n3095), .o (n3096) );
  buffer buf_n3097( .i (n3096), .o (n3097) );
  assign n3101 = n3097 & ~n3099 ;
  assign n3102 = ( n3032 & ~n3100 ) | ( n3032 & n3101 ) | ( ~n3100 & n3101 ) ;
  assign n3103 = ~n3088 & n3102 ;
  buffer buf_n3104( .i (n68), .o (n3104) );
  buffer buf_n3105( .i (n3104), .o (n3105) );
  assign n3106 = ( n3089 & n3103 ) | ( n3089 & ~n3105 ) | ( n3103 & ~n3105 ) ;
  assign n3107 = ( n2133 & n3074 ) | ( n2133 & ~n3106 ) | ( n3074 & ~n3106 ) ;
  assign n3108 = n2429 & ~n3107 ;
  assign n3109 = ( n310 & n3076 ) | ( n310 & ~n3108 ) | ( n3076 & ~n3108 ) ;
  buffer buf_n3110( .i (n2490), .o (n3110) );
  assign n3111 = ( n2266 & ~n3109 ) | ( n2266 & n3110 ) | ( ~n3109 & n3110 ) ;
  assign n3112 = n3054 & ~n3111 ;
  assign n3113 = n140 & n3112 ;
  assign n3114 = ( n3048 & n3051 ) | ( n3048 & n3113 ) | ( n3051 & n3113 ) ;
  buffer buf_n2767( .i (n2766), .o (n2767) );
  buffer buf_n2768( .i (n2767), .o (n2768) );
  buffer buf_n2769( .i (n2768), .o (n2769) );
  buffer buf_n2770( .i (n2769), .o (n2770) );
  buffer buf_n2771( .i (n2770), .o (n2771) );
  buffer buf_n2772( .i (n2771), .o (n2772) );
  buffer buf_n2773( .i (n2772), .o (n2773) );
  buffer buf_n2774( .i (n2773), .o (n2774) );
  buffer buf_n2775( .i (n2774), .o (n2775) );
  buffer buf_n2776( .i (n2775), .o (n2776) );
  buffer buf_n2777( .i (n2776), .o (n2777) );
  buffer buf_n2778( .i (n2777), .o (n2778) );
  buffer buf_n2779( .i (n2778), .o (n2779) );
  assign n3115 = ( ~n1228 & n2273 ) | ( ~n1228 & n2779 ) | ( n2273 & n2779 ) ;
  assign n3116 = ~n2938 & n3115 ;
  buffer buf_n3117( .i (n3116), .o (n3117) );
  buffer buf_n3118( .i (n3117), .o (n3118) );
  buffer buf_n3014( .i (n3013), .o (n3014) );
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  assign n3119 = n1854 & n2731 ;
  assign n3120 = ( n3014 & ~n3117 ) | ( n3014 & n3119 ) | ( ~n3117 & n3119 ) ;
  assign n3121 = n3118 & n3120 ;
  buffer buf_n3122( .i (n3121), .o (n3122) );
  assign n3123 = ( ~n3018 & n3114 ) | ( ~n3018 & n3122 ) | ( n3114 & n3122 ) ;
  assign n3124 = n244 | n3122 ;
  assign n3125 = ( n3019 & n3123 ) | ( n3019 & n3124 ) | ( n3123 & n3124 ) ;
  assign n3126 = n416 & n3125 ;
  buffer buf_n3127( .i (n3126), .o (n3127) );
  buffer buf_n3128( .i (n3127), .o (n3128) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  assign n3129 = n210 | n1235 ;
  assign n3130 = ( ~n177 & n246 ) | ( ~n177 & n3129 ) | ( n246 & n3129 ) ;
  assign n3131 = n178 | n3130 ;
  assign n3132 = ~n3127 & n3131 ;
  assign n3133 = ( ~n3008 & n3128 ) | ( ~n3008 & ~n3132 ) | ( n3128 & ~n3132 ) ;
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  assign n3134 = n303 & n2045 ;
  buffer buf_n3135( .i (n3134), .o (n3135) );
  buffer buf_n3136( .i (n3135), .o (n3136) );
  buffer buf_n3137( .i (n3136), .o (n3137) );
  buffer buf_n3138( .i (n3137), .o (n3138) );
  buffer buf_n3139( .i (n3138), .o (n3139) );
  buffer buf_n3140( .i (n3139), .o (n3140) );
  buffer buf_n3141( .i (n3140), .o (n3141) );
  buffer buf_n3142( .i (n3141), .o (n3142) );
  buffer buf_n3143( .i (n2926), .o (n3143) );
  assign n3144 = n2813 & ~n3143 ;
  assign n3145 = ~n2729 & n3144 ;
  buffer buf_n3146( .i (n2496), .o (n3146) );
  buffer buf_n3147( .i (n3146), .o (n3147) );
  assign n3148 = ( n3141 & ~n3145 ) | ( n3141 & n3147 ) | ( ~n3145 & n3147 ) ;
  buffer buf_n2977( .i (n2976), .o (n2977) );
  buffer buf_n2978( .i (n2977), .o (n2978) );
  assign n3149 = ( ~n2372 & n2978 ) | ( ~n2372 & n3143 ) | ( n2978 & n3143 ) ;
  assign n3150 = n2373 & n3149 ;
  assign n3151 = ~n3147 & n3150 ;
  assign n3152 = ( n3142 & ~n3148 ) | ( n3142 & n3151 ) | ( ~n3148 & n3151 ) ;
  buffer buf_n3153( .i (n2687), .o (n3153) );
  assign n3154 = ( n2942 & n3152 ) | ( n2942 & ~n3153 ) | ( n3152 & ~n3153 ) ;
  assign n3155 = n101 & ~n1016 ;
  assign n3156 = ( n38 & n71 ) | ( n38 & n3155 ) | ( n71 & n3155 ) ;
  assign n3157 = ~n39 & n3156 ;
  buffer buf_n3158( .i (n3157), .o (n3158) );
  buffer buf_n3159( .i (n3158), .o (n3159) );
  assign n3160 = ~n343 & n2496 ;
  assign n3161 = n2985 & n3160 ;
  buffer buf_n2740( .i (n2739), .o (n2740) );
  buffer buf_n2741( .i (n2740), .o (n2741) );
  buffer buf_n3162( .i (n2728), .o (n3162) );
  assign n3163 = ~n2741 & n3162 ;
  assign n3164 = ( ~n3158 & n3161 ) | ( ~n3158 & n3163 ) | ( n3161 & n3163 ) ;
  assign n3165 = n3159 & n3164 ;
  assign n3166 = ~n3153 & n3165 ;
  assign n3167 = ( ~n108 & n3154 ) | ( ~n108 & n3166 ) | ( n3154 & n3166 ) ;
  assign n3168 = ~n142 & n3167 ;
  buffer buf_n3169( .i (n468), .o (n3169) );
  assign n3170 = n3085 & ~n3169 ;
  buffer buf_n3171( .i (n3026), .o (n3171) );
  assign n3172 = n2219 | n3171 ;
  assign n3173 = ( n67 & ~n3170 ) | ( n67 & n3172 ) | ( ~n3170 & n3172 ) ;
  assign n3174 = n305 | n3173 ;
  buffer buf_n3175( .i (n2086), .o (n3175) );
  assign n3176 = ( n2808 & n3174 ) | ( n2808 & ~n3175 ) | ( n3174 & ~n3175 ) ;
  buffer buf_n3177( .i (n3175), .o (n3177) );
  assign n3178 = n3176 | n3177 ;
  buffer buf_n3179( .i (n3178), .o (n3179) );
  buffer buf_n3180( .i (n3179), .o (n3180) );
  assign n3181 = n187 & n327 ;
  buffer buf_n3182( .i (n3181), .o (n3182) );
  assign n3187 = ( n361 & n2869 ) | ( n361 & n3182 ) | ( n2869 & n3182 ) ;
  buffer buf_n3188( .i (n2869), .o (n3188) );
  assign n3189 = n3187 & ~n3188 ;
  buffer buf_n3190( .i (n3189), .o (n3190) );
  buffer buf_n3191( .i (n3190), .o (n3191) );
  buffer buf_n3192( .i (n3191), .o (n3192) );
  assign n3193 = ( n61 & n2876 ) | ( n61 & ~n3190 ) | ( n2876 & ~n3190 ) ;
  assign n3194 = n3079 & n3193 ;
  assign n3195 = ( n3080 & n3192 ) | ( n3080 & ~n3194 ) | ( n3192 & ~n3194 ) ;
  buffer buf_n3196( .i (n3195), .o (n3196) );
  buffer buf_n3197( .i (n3196), .o (n3197) );
  assign n3198 = ( ~n162 & n2564 ) | ( ~n162 & n3196 ) | ( n2564 & n3196 ) ;
  assign n3199 = n1008 | n3090 ;
  buffer buf_n3200( .i (n333), .o (n3200) );
  assign n3201 = ( n466 & n3199 ) | ( n466 & ~n3200 ) | ( n3199 & ~n3200 ) ;
  assign n3202 = n335 | n3201 ;
  assign n3203 = n2564 | n3202 ;
  assign n3204 = ( ~n3197 & n3198 ) | ( ~n3197 & n3203 ) | ( n3198 & n3203 ) ;
  buffer buf_n3205( .i (n3204), .o (n3205) );
  buffer buf_n3206( .i (n3205), .o (n3206) );
  buffer buf_n3207( .i (n304), .o (n3207) );
  assign n3208 = ( n2086 & n3205 ) | ( n2086 & n3207 ) | ( n3205 & n3207 ) ;
  assign n3209 = n222 & n327 ;
  buffer buf_n3210( .i (n3209), .o (n3210) );
  assign n3225 = n361 & n3210 ;
  assign n3226 = ( n156 & ~n525 ) | ( n156 & n3225 ) | ( ~n525 & n3225 ) ;
  assign n3227 = n526 & n3226 ;
  buffer buf_n3228( .i (n3227), .o (n3228) );
  buffer buf_n3229( .i (n3228), .o (n3229) );
  buffer buf_n3230( .i (n3229), .o (n3230) );
  assign n3231 = n2038 & n2310 ;
  assign n3232 = n23 & ~n3057 ;
  buffer buf_n3233( .i (n3232), .o (n3233) );
  assign n3236 = n25 & ~n3233 ;
  buffer buf_n3237( .i (n3236), .o (n3237) );
  assign n3238 = n3231 & n3237 ;
  buffer buf_n3234( .i (n3233), .o (n3234) );
  buffer buf_n3235( .i (n3234), .o (n3235) );
  assign n3239 = ( n222 & n327 ) | ( n222 & n359 ) | ( n327 & n359 ) ;
  buffer buf_n3240( .i (n3239), .o (n3240) );
  buffer buf_n3241( .i (n3240), .o (n3241) );
  buffer buf_n3242( .i (n223), .o (n3242) );
  assign n3243 = ~n3240 & n3242 ;
  assign n3244 = ( n330 & ~n3241 ) | ( n330 & n3243 ) | ( ~n3241 & n3243 ) ;
  assign n3245 = ( ~n3235 & n3237 ) | ( ~n3235 & n3244 ) | ( n3237 & n3244 ) ;
  assign n3246 = ( ~n2583 & n3238 ) | ( ~n2583 & n3245 ) | ( n3238 & n3245 ) ;
  assign n3247 = ( ~n465 & n3228 ) | ( ~n465 & n3246 ) | ( n3228 & n3246 ) ;
  assign n3248 = n432 & ~n3247 ;
  assign n3249 = ( n2193 & n3230 ) | ( n2193 & ~n3248 ) | ( n3230 & ~n3248 ) ;
  buffer buf_n3250( .i (n3249), .o (n3250) );
  buffer buf_n3251( .i (n3250), .o (n3251) );
  assign n3252 = ( n1587 & n3085 ) | ( n1587 & ~n3250 ) | ( n3085 & ~n3250 ) ;
  assign n3253 = n529 & n1354 ;
  assign n3254 = ( ~n576 & n2055 ) | ( ~n576 & n3253 ) | ( n2055 & n3253 ) ;
  buffer buf_n3255( .i (n2055), .o (n3255) );
  assign n3256 = n3254 & ~n3255 ;
  assign n3257 = n3085 & n3256 ;
  assign n3258 = ( n3251 & n3252 ) | ( n3251 & n3257 ) | ( n3252 & n3257 ) ;
  assign n3259 = n3207 & n3258 ;
  assign n3260 = ( ~n3206 & n3208 ) | ( ~n3206 & n3259 ) | ( n3208 & n3259 ) ;
  buffer buf_n3261( .i (n3260), .o (n3261) );
  buffer buf_n3262( .i (n3261), .o (n3262) );
  buffer buf_n3263( .i (n3262), .o (n3263) );
  assign n3264 = ( n168 & n2926 ) | ( n168 & ~n3261 ) | ( n2926 & ~n3261 ) ;
  assign n3265 = ~n3179 & n3264 ;
  assign n3266 = ( n3180 & ~n3263 ) | ( n3180 & n3265 ) | ( ~n3263 & n3265 ) ;
  buffer buf_n3267( .i (n3266), .o (n3267) );
  buffer buf_n3268( .i (n3267), .o (n3268) );
  assign n3269 = ( n106 & n2343 ) | ( n106 & n3267 ) | ( n2343 & n3267 ) ;
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  assign n3270 = ( n304 & n1100 ) | ( n304 & n3031 ) | ( n1100 & n3031 ) ;
  buffer buf_n3271( .i (n2004), .o (n3271) );
  buffer buf_n3272( .i (n1899), .o (n3272) );
  assign n3273 = ( ~n1099 & n3271 ) | ( ~n1099 & n3272 ) | ( n3271 & n3272 ) ;
  assign n3274 = ( n2444 & n3031 ) | ( n2444 & n3273 ) | ( n3031 & n3273 ) ;
  assign n3275 = ~n3270 & n3274 ;
  assign n3276 = n3036 & ~n3275 ;
  assign n3277 = n298 | n2583 ;
  buffer buf_n3278( .i (n3277), .o (n3278) );
  buffer buf_n3279( .i (n3278), .o (n3279) );
  buffer buf_n3280( .i (n3279), .o (n3280) );
  buffer buf_n3281( .i (n3280), .o (n3281) );
  buffer buf_n3282( .i (n3281), .o (n3282) );
  buffer buf_n3283( .i (n3282), .o (n3283) );
  assign n3284 = n3032 & ~n3283 ;
  assign n3285 = n3036 | n3284 ;
  assign n3286 = ~n3276 & n3285 ;
  buffer buf_n3287( .i (n3286), .o (n3287) );
  buffer buf_n3288( .i (n3287), .o (n3288) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  assign n3289 = ( ~n1803 & n2496 ) | ( ~n1803 & n3287 ) | ( n2496 & n3287 ) ;
  assign n3290 = n3288 & ~n3289 ;
  assign n3291 = n1365 & n3290 ;
  buffer buf_n3292( .i (n3110), .o (n3292) );
  assign n3293 = n3291 & n3292 ;
  assign n3294 = ( ~n3268 & n3269 ) | ( ~n3268 & n3293 ) | ( n3269 & n3293 ) ;
  buffer buf_n3295( .i (n326), .o (n3295) );
  buffer buf_n3296( .i (n3295), .o (n3296) );
  assign n3297 = n258 & n3296 ;
  buffer buf_n3298( .i (n3297), .o (n3298) );
  buffer buf_n3299( .i (n3298), .o (n3299) );
  buffer buf_n3300( .i (n3299), .o (n3300) );
  buffer buf_n3301( .i (n3300), .o (n3301) );
  buffer buf_n3302( .i (n3301), .o (n3302) );
  buffer buf_n3303( .i (n3302), .o (n3303) );
  buffer buf_n3304( .i (n3303), .o (n3304) );
  buffer buf_n3305( .i (n3304), .o (n3305) );
  buffer buf_n3306( .i (n3305), .o (n3306) );
  buffer buf_n3307( .i (n3306), .o (n3307) );
  buffer buf_n3308( .i (n3307), .o (n3308) );
  assign n3309 = ( n306 & n2743 ) | ( n306 & ~n3308 ) | ( n2743 & ~n3308 ) ;
  assign n3310 = ( ~n1932 & n3207 ) | ( ~n1932 & n3307 ) | ( n3207 & n3307 ) ;
  assign n3311 = ( n2743 & ~n2808 ) | ( n2743 & n3310 ) | ( ~n2808 & n3310 ) ;
  assign n3312 = n3309 & ~n3311 ;
  buffer buf_n3313( .i (n3312), .o (n3313) );
  buffer buf_n3314( .i (n3313), .o (n3314) );
  buffer buf_n3315( .i (n1935), .o (n3315) );
  buffer buf_n3316( .i (n3315), .o (n3316) );
  assign n3317 = ( ~n1580 & n3313 ) | ( ~n1580 & n3316 ) | ( n3313 & n3316 ) ;
  assign n3318 = n3314 & ~n3317 ;
  assign n3319 = ~n205 & n3318 ;
  assign n3320 = ( n172 & n3292 ) | ( n172 & n3319 ) | ( n3292 & n3319 ) ;
  assign n3321 = ~n2942 & n3320 ;
  assign n3322 = n3294 | n3321 ;
  buffer buf_n3323( .i (n141), .o (n3323) );
  assign n3324 = n3322 & n3323 ;
  assign n3325 = n3168 | n3324 ;
  buffer buf_n3326( .i (n415), .o (n3326) );
  assign n3327 = n3325 & n3326 ;
  buffer buf_n3328( .i (n3327), .o (n3328) );
  buffer buf_n3329( .i (n3328), .o (n3329) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n3211( .i (n3210), .o (n3211) );
  buffer buf_n3212( .i (n3211), .o (n3212) );
  buffer buf_n3213( .i (n3212), .o (n3213) );
  buffer buf_n3214( .i (n3213), .o (n3214) );
  buffer buf_n3215( .i (n3214), .o (n3215) );
  buffer buf_n3216( .i (n3215), .o (n3216) );
  buffer buf_n3217( .i (n3216), .o (n3217) );
  buffer buf_n3218( .i (n3217), .o (n3218) );
  buffer buf_n3219( .i (n3218), .o (n3219) );
  buffer buf_n3220( .i (n3219), .o (n3220) );
  buffer buf_n3221( .i (n3220), .o (n3221) );
  buffer buf_n3222( .i (n3221), .o (n3222) );
  buffer buf_n3223( .i (n3222), .o (n3223) );
  buffer buf_n3224( .i (n3223), .o (n3224) );
  buffer buf_n3330( .i (n3105), .o (n3330) );
  assign n3331 = n3315 | n3330 ;
  assign n3332 = ( n72 & n3224 ) | ( n72 & ~n3331 ) | ( n3224 & ~n3331 ) ;
  buffer buf_n3333( .i (n3332), .o (n3333) );
  buffer buf_n3334( .i (n3333), .o (n3334) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  assign n3335 = ( n617 & n2930 ) | ( n617 & ~n3333 ) | ( n2930 & ~n3333 ) ;
  assign n3336 = n3334 & n3335 ;
  buffer buf_n3337( .i (n3336), .o (n3337) );
  buffer buf_n3338( .i (n3337), .o (n3338) );
  assign n3339 = ( ~n108 & n446 ) | ( ~n108 & n3337 ) | ( n446 & n3337 ) ;
  buffer buf_n3340( .i (n1571), .o (n3340) );
  assign n3341 = ( ~n206 & n2997 ) | ( ~n206 & n3340 ) | ( n2997 & n3340 ) ;
  assign n3342 = n207 | n3341 ;
  buffer buf_n3343( .i (n2487), .o (n3343) );
  buffer buf_n3344( .i (n3343), .o (n3344) );
  assign n3345 = n3342 | n3344 ;
  assign n3346 = ( ~n3338 & n3339 ) | ( ~n3338 & n3345 ) | ( n3339 & n3345 ) ;
  assign n3347 = n382 | n3346 ;
  assign n3348 = ( ~n317 & n3326 ) | ( ~n317 & n3347 ) | ( n3326 & n3347 ) ;
  assign n3349 = n318 | n3348 ;
  assign n3350 = ~n3328 & n3349 ;
  assign n3351 = ( ~n284 & n3329 ) | ( ~n284 & ~n3350 ) | ( n3329 & ~n3350 ) ;
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  assign n3352 = ~n137 & n1477 ;
  buffer buf_n3353( .i (n3352), .o (n3353) );
  buffer buf_n3354( .i (n3353), .o (n3354) );
  assign n3355 = ( n172 & ~n206 ) | ( n172 & n3353 ) | ( ~n206 & n3353 ) ;
  assign n3356 = ( n1480 & n3354 ) | ( n1480 & n3355 ) | ( n3354 & n3355 ) ;
  buffer buf_n3357( .i (n3356), .o (n3357) );
  buffer buf_n3358( .i (n3357), .o (n3358) );
  buffer buf_n2958( .i (n2957), .o (n2958) );
  buffer buf_n2959( .i (n2958), .o (n2959) );
  buffer buf_n2960( .i (n2959), .o (n2960) );
  buffer buf_n2961( .i (n2960), .o (n2961) );
  buffer buf_n2962( .i (n2961), .o (n2962) );
  buffer buf_n2963( .i (n2962), .o (n2963) );
  assign n3359 = n2150 & n3200 ;
  buffer buf_n3360( .i (n3359), .o (n3360) );
  buffer buf_n3361( .i (n3360), .o (n3361) );
  buffer buf_n3362( .i (n3361), .o (n3362) );
  buffer buf_n3363( .i (n3362), .o (n3363) );
  buffer buf_n3364( .i (n3363), .o (n3364) );
  buffer buf_n3365( .i (n3364), .o (n3365) );
  buffer buf_n3366( .i (n3365), .o (n3366) );
  buffer buf_n3367( .i (n3366), .o (n3367) );
  buffer buf_n3368( .i (n3367), .o (n3368) );
  buffer buf_n3369( .i (n3368), .o (n3369) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  assign n3370 = n585 | n3368 ;
  assign n3371 = ( n2963 & n3369 ) | ( n2963 & ~n3370 ) | ( n3369 & ~n3370 ) ;
  buffer buf_n3372( .i (n3371), .o (n3372) );
  buffer buf_n3373( .i (n3372), .o (n3373) );
  buffer buf_n3374( .i (n2268), .o (n3374) );
  assign n3375 = n3372 & ~n3374 ;
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  assign n3376 = n205 | n1282 ;
  buffer buf_n3377( .i (n2930), .o (n3377) );
  assign n3378 = n3376 | n3377 ;
  buffer buf_n496( .i (n495), .o (n496) );
  assign n3379 = n496 & ~n2734 ;
  buffer buf_n3380( .i (n3379), .o (n3380) );
  buffer buf_n3381( .i (n3380), .o (n3381) );
  buffer buf_n3382( .i (n3381), .o (n3382) );
  buffer buf_n3383( .i (n3382), .o (n3383) );
  buffer buf_n3384( .i (n3383), .o (n3384) );
  buffer buf_n3385( .i (n3384), .o (n3385) );
  buffer buf_n3386( .i (n3385), .o (n3386) );
  buffer buf_n3387( .i (n3386), .o (n3387) );
  assign n3388 = n262 | n2204 ;
  buffer buf_n3389( .i (n3388), .o (n3389) );
  buffer buf_n3390( .i (n3389), .o (n3390) );
  buffer buf_n3391( .i (n3390), .o (n3391) );
  buffer buf_n3392( .i (n3391), .o (n3392) );
  buffer buf_n3393( .i (n3392), .o (n3393) );
  buffer buf_n3394( .i (n3393), .o (n3394) );
  buffer buf_n3395( .i (n3394), .o (n3395) );
  buffer buf_n3396( .i (n3395), .o (n3396) );
  buffer buf_n3397( .i (n3396), .o (n3397) );
  buffer buf_n3398( .i (n3397), .o (n3398) );
  buffer buf_n3399( .i (n3398), .o (n3399) );
  assign n3400 = ( ~n1913 & n3162 ) | ( ~n1913 & n3399 ) | ( n3162 & n3399 ) ;
  assign n3401 = n41 & n3400 ;
  assign n3402 = ~n3387 & n3401 ;
  assign n3403 = n3378 & n3402 ;
  assign n3404 = ( ~n3373 & n3375 ) | ( ~n3373 & n3403 ) | ( n3375 & n3403 ) ;
  assign n3405 = n2650 & n3177 ;
  assign n3406 = ( n2651 & n2926 ) | ( n2651 & n3405 ) | ( n2926 & n3405 ) ;
  buffer buf_n3407( .i (n2133), .o (n3407) );
  assign n3408 = n3406 & ~n3407 ;
  assign n3409 = ~n399 & n3093 ;
  buffer buf_n3410( .i (n3093), .o (n3410) );
  assign n3411 = ( n335 & n3409 ) | ( n335 & ~n3410 ) | ( n3409 & ~n3410 ) ;
  buffer buf_n3412( .i (n3411), .o (n3412) );
  buffer buf_n3413( .i (n3412), .o (n3413) );
  assign n3414 = ( n337 & n3171 ) | ( n337 & n3412 ) | ( n3171 & n3412 ) ;
  assign n3415 = ( n579 & n3413 ) | ( n579 & ~n3414 ) | ( n3413 & ~n3414 ) ;
  buffer buf_n3416( .i (n3415), .o (n3416) );
  buffer buf_n3417( .i (n3416), .o (n3417) );
  buffer buf_n3418( .i (n132), .o (n3418) );
  assign n3419 = ~n3416 & n3418 ;
  assign n3420 = n579 | n1766 ;
  assign n3421 = ( n1767 & ~n3363 ) | ( n1767 & n3420 ) | ( ~n3363 & n3420 ) ;
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n3422( .i (n30), .o (n3422) );
  assign n3423 = ( ~n576 & n1509 ) | ( ~n576 & n3422 ) | ( n1509 & n3422 ) ;
  buffer buf_n3424( .i (n3423), .o (n3424) );
  buffer buf_n3425( .i (n3424), .o (n3425) );
  buffer buf_n3426( .i (n3425), .o (n3426) );
  buffer buf_n3427( .i (n3422), .o (n3427) );
  buffer buf_n3428( .i (n3427), .o (n3428) );
  assign n3429 = ( n3361 & n3424 ) | ( n3361 & ~n3428 ) | ( n3424 & ~n3428 ) ;
  buffer buf_n3430( .i (n2028), .o (n3430) );
  buffer buf_n3431( .i (n3430), .o (n3431) );
  assign n3432 = ~n3429 & n3431 ;
  assign n3433 = ( n1594 & n3426 ) | ( n1594 & ~n3432 ) | ( n3426 & ~n3432 ) ;
  assign n3434 = n3421 & ~n3433 ;
  assign n3435 = ( n3417 & n3419 ) | ( n3417 & n3434 ) | ( n3419 & n3434 ) ;
  assign n3436 = n2727 & ~n3435 ;
  assign n3437 = n3407 & ~n3436 ;
  assign n3438 = n3408 | n3437 ;
  buffer buf_n3439( .i (n3438), .o (n3439) );
  buffer buf_n3440( .i (n3439), .o (n3440) );
  assign n3441 = n2143 | n3439 ;
  buffer buf_n3442( .i (n231), .o (n3442) );
  assign n3443 = ( n3171 & n3430 ) | ( n3171 & ~n3442 ) | ( n3430 & ~n3442 ) ;
  assign n3444 = n131 & n3443 ;
  buffer buf_n3445( .i (n131), .o (n3445) );
  assign n3446 = ( n1594 & n3444 ) | ( n1594 & ~n3445 ) | ( n3444 & ~n3445 ) ;
  buffer buf_n3447( .i (n3446), .o (n3447) );
  buffer buf_n3448( .i (n3447), .o (n3448) );
  assign n3449 = n1204 & ~n3447 ;
  assign n3450 = n268 & n3431 ;
  buffer buf_n3451( .i (n233), .o (n3451) );
  assign n3452 = n3450 & n3451 ;
  assign n3453 = n2155 & n3207 ;
  assign n3454 = n3452 & n3453 ;
  assign n3455 = n785 & ~n3454 ;
  assign n3456 = ( n3448 & n3449 ) | ( n3448 & n3455 ) | ( n3449 & n3455 ) ;
  buffer buf_n3457( .i (n3456), .o (n3457) );
  buffer buf_n3458( .i (n3457), .o (n3458) );
  assign n3459 = ( n344 & ~n2406 ) | ( n344 & n3457 ) | ( ~n2406 & n3457 ) ;
  assign n3460 = n229 | n1903 ;
  buffer buf_n3461( .i (n3460), .o (n3461) );
  buffer buf_n3462( .i (n3461), .o (n3462) );
  buffer buf_n3464( .i (n2018), .o (n3464) );
  buffer buf_n3465( .i (n298), .o (n3465) );
  assign n3466 = n3464 & ~n3465 ;
  buffer buf_n3467( .i (n263), .o (n3467) );
  assign n3468 = ( n2150 & n3466 ) | ( n2150 & n3467 ) | ( n3466 & n3467 ) ;
  assign n3469 = ~n265 & n3468 ;
  assign n3470 = n3461 & ~n3469 ;
  assign n3471 = ( n3428 & n3462 ) | ( n3428 & ~n3470 ) | ( n3462 & ~n3470 ) ;
  buffer buf_n3472( .i (n3471), .o (n3472) );
  buffer buf_n3473( .i (n3472), .o (n3473) );
  buffer buf_n3474( .i (n3428), .o (n3474) );
  buffer buf_n3475( .i (n3474), .o (n3475) );
  assign n3476 = ( n3445 & n3472 ) | ( n3445 & n3475 ) | ( n3472 & n3475 ) ;
  assign n3477 = ( n878 & n3473 ) | ( n878 & ~n3476 ) | ( n3473 & ~n3476 ) ;
  buffer buf_n3478( .i (n3477), .o (n3478) );
  buffer buf_n3479( .i (n3478), .o (n3479) );
  buffer buf_n3480( .i (n2677), .o (n3480) );
  assign n3481 = ~n3478 & n3480 ;
  buffer buf_n3482( .i (n1733), .o (n3482) );
  assign n3483 = n26 & n3482 ;
  buffer buf_n3484( .i (n1986), .o (n3484) );
  buffer buf_n3485( .i (n123), .o (n3485) );
  assign n3486 = ( n3483 & n3484 ) | ( n3483 & n3485 ) | ( n3484 & n3485 ) ;
  buffer buf_n3487( .i (n3485), .o (n3487) );
  assign n3488 = n3486 & ~n3487 ;
  buffer buf_n3489( .i (n3488), .o (n3489) );
  buffer buf_n3490( .i (n3489), .o (n3490) );
  buffer buf_n3491( .i (n3490), .o (n3491) );
  buffer buf_n3492( .i (n3491), .o (n3492) );
  buffer buf_n3493( .i (n3492), .o (n3493) );
  assign n3494 = ( n2954 & n3427 ) | ( n2954 & ~n3491 ) | ( n3427 & ~n3491 ) ;
  assign n3495 = n1433 & n3494 ;
  buffer buf_n3496( .i (n1433), .o (n3496) );
  assign n3497 = ( n3493 & ~n3495 ) | ( n3493 & n3496 ) | ( ~n3495 & n3496 ) ;
  buffer buf_n3498( .i (n3497), .o (n3498) );
  buffer buf_n3499( .i (n3498), .o (n3499) );
  buffer buf_n3500( .i (n3032), .o (n3500) );
  assign n3501 = n3498 & ~n3500 ;
  buffer buf_n3502( .i (n2676), .o (n3502) );
  assign n3503 = ( n3499 & n3501 ) | ( n3499 & n3502 ) | ( n3501 & n3502 ) ;
  buffer buf_n3504( .i (n3431), .o (n3504) );
  buffer buf_n3505( .i (n3171), .o (n3505) );
  buffer buf_n3506( .i (n3505), .o (n3506) );
  assign n3507 = ( n3445 & ~n3504 ) | ( n3445 & n3506 ) | ( ~n3504 & n3506 ) ;
  assign n3508 = ( n1277 & n2676 ) | ( n1277 & n3507 ) | ( n2676 & n3507 ) ;
  buffer buf_n3463( .i (n3462), .o (n3463) );
  assign n3509 = n127 | n3489 ;
  assign n3510 = ( ~n3422 & n3490 ) | ( ~n3422 & n3509 ) | ( n3490 & n3509 ) ;
  buffer buf_n3511( .i (n3510), .o (n3511) );
  buffer buf_n3512( .i (n3511), .o (n3512) );
  assign n3513 = ~n402 & n3511 ;
  assign n3514 = ( ~n3463 & n3512 ) | ( ~n3463 & n3513 ) | ( n3512 & n3513 ) ;
  buffer buf_n3515( .i (n3514), .o (n3515) );
  buffer buf_n3516( .i (n3515), .o (n3516) );
  buffer buf_n3517( .i (n3475), .o (n3517) );
  assign n3518 = ~n3515 & n3517 ;
  assign n3519 = ( n3508 & n3516 ) | ( n3508 & ~n3518 ) | ( n3516 & ~n3518 ) ;
  assign n3520 = n3503 | n3519 ;
  assign n3521 = ( n3479 & n3481 ) | ( n3479 & ~n3520 ) | ( n3481 & ~n3520 ) ;
  assign n3522 = n2406 | n3521 ;
  assign n3523 = ( n3458 & ~n3459 ) | ( n3458 & n3522 ) | ( ~n3459 & n3522 ) ;
  assign n3524 = n56 & n87 ;
  buffer buf_n3525( .i (n3524), .o (n3525) );
  buffer buf_n3526( .i (n3525), .o (n3526) );
  buffer buf_n3527( .i (n3526), .o (n3527) );
  buffer buf_n3528( .i (n3527), .o (n3528) );
  buffer buf_n3529( .i (n3528), .o (n3529) );
  buffer buf_n3530( .i (n3529), .o (n3530) );
  buffer buf_n3540( .i (n29), .o (n3540) );
  assign n3541 = n3530 & n3540 ;
  buffer buf_n3542( .i (n3541), .o (n3542) );
  assign n3544 = n969 & n3542 ;
  assign n3545 = ( n337 & n3430 ) | ( n337 & n3544 ) | ( n3430 & n3544 ) ;
  assign n3546 = ~n338 & n3545 ;
  buffer buf_n3547( .i (n3546), .o (n3547) );
  buffer buf_n3548( .i (n3547), .o (n3548) );
  buffer buf_n3549( .i (n3548), .o (n3549) );
  assign n3550 = ( ~n405 & n2808 ) | ( ~n405 & n3547 ) | ( n2808 & n3547 ) ;
  assign n3551 = n2738 | n3550 ;
  assign n3552 = ( ~n2739 & n3549 ) | ( ~n2739 & n3551 ) | ( n3549 & n3551 ) ;
  buffer buf_n3553( .i (n3552), .o (n3553) );
  buffer buf_n3554( .i (n3553), .o (n3554) );
  assign n3555 = ~n2985 & n3553 ;
  assign n3556 = ( n2616 & n2905 ) | ( n2616 & ~n3487 ) | ( n2905 & ~n3487 ) ;
  buffer buf_n3557( .i (n2908), .o (n3557) );
  buffer buf_n3558( .i (n3557), .o (n3558) );
  assign n3559 = ~n3556 & n3558 ;
  assign n3560 = n777 & ~n3558 ;
  buffer buf_n3561( .i (n3090), .o (n3561) );
  assign n3562 = ( n3559 & ~n3560 ) | ( n3559 & n3561 ) | ( ~n3560 & n3561 ) ;
  buffer buf_n3563( .i (n3562), .o (n3563) );
  buffer buf_n3564( .i (n265), .o (n3564) );
  assign n3565 = ( n3026 & n3563 ) | ( n3026 & ~n3564 ) | ( n3563 & ~n3564 ) ;
  buffer buf_n3566( .i (n399), .o (n3566) );
  assign n3567 = ( n494 & n3410 ) | ( n494 & n3566 ) | ( n3410 & n3566 ) ;
  assign n3568 = n3563 & n3567 ;
  assign n3569 = ( n267 & n3565 ) | ( n267 & n3568 ) | ( n3565 & n3568 ) ;
  buffer buf_n3570( .i (n3569), .o (n3570) );
  assign n3571 = ( n1908 & n1932 ) | ( n1908 & n3570 ) | ( n1932 & n3570 ) ;
  buffer buf_n3572( .i (n2202), .o (n3572) );
  assign n3573 = n3570 & n3572 ;
  assign n3574 = ( ~n1909 & n3571 ) | ( ~n1909 & n3573 ) | ( n3571 & n3573 ) ;
  buffer buf_n3575( .i (n3574), .o (n3575) );
  buffer buf_n3576( .i (n3575), .o (n3576) );
  assign n3577 = n911 & ~n1906 ;
  buffer buf_n3578( .i (n3577), .o (n3578) );
  buffer buf_n3579( .i (n3578), .o (n3579) );
  assign n3580 = n165 & ~n3578 ;
  assign n3581 = ( n3517 & ~n3579 ) | ( n3517 & n3580 ) | ( ~n3579 & n3580 ) ;
  buffer buf_n3543( .i (n3542), .o (n3543) );
  assign n3582 = ( n608 & n3255 ) | ( n608 & ~n3542 ) | ( n3255 & ~n3542 ) ;
  assign n3583 = n3543 & n3582 ;
  buffer buf_n3584( .i (n3583), .o (n3584) );
  buffer buf_n3585( .i (n3584), .o (n3585) );
  buffer buf_n3589( .i (n267), .o (n3589) );
  buffer buf_n3590( .i (n3589), .o (n3590) );
  assign n3591 = n1908 | n3590 ;
  assign n3592 = ( n1909 & ~n3585 ) | ( n1909 & n3591 ) | ( ~n3585 & n3591 ) ;
  assign n3593 = ( n3177 & ~n3581 ) | ( n3177 & n3592 ) | ( ~n3581 & n3592 ) ;
  assign n3594 = n3575 & ~n3593 ;
  assign n3595 = ( n2728 & n3576 ) | ( n2728 & ~n3594 ) | ( n3576 & ~n3594 ) ;
  buffer buf_n3586( .i (n3585), .o (n3586) );
  buffer buf_n3587( .i (n3586), .o (n3587) );
  buffer buf_n3588( .i (n3587), .o (n3588) );
  assign n3596 = ~n294 & n487 ;
  assign n3597 = ~n903 & n3596 ;
  buffer buf_n3598( .i (n3597), .o (n3598) );
  buffer buf_n3599( .i (n3598), .o (n3599) );
  buffer buf_n3600( .i (n3599), .o (n3600) );
  assign n3601 = ( n601 & n1879 ) | ( n601 & n2947 ) | ( n1879 & n2947 ) ;
  assign n3602 = ~n2948 & n3601 ;
  assign n3603 = ( n2292 & n3598 ) | ( n2292 & n3602 ) | ( n3598 & n3602 ) ;
  assign n3604 = n2018 & ~n3603 ;
  assign n3605 = ( n3464 & n3600 ) | ( n3464 & ~n3604 ) | ( n3600 & ~n3604 ) ;
  assign n3606 = n3540 & n3605 ;
  buffer buf_n3607( .i (n3606), .o (n3607) );
  buffer buf_n3608( .i (n3607), .o (n3608) );
  assign n3609 = ( n1423 & ~n2875 ) | ( n1423 & n3485 ) | ( ~n2875 & n3485 ) ;
  assign n3610 = ~n3487 & n3609 ;
  buffer buf_n3611( .i (n3610), .o (n3611) );
  buffer buf_n3612( .i (n3611), .o (n3612) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  assign n3613 = ( n688 & ~n3200 ) | ( n688 & n3611 ) | ( ~n3200 & n3611 ) ;
  assign n3614 = ~n3612 & n3613 ;
  assign n3615 = n3607 | n3614 ;
  buffer buf_n3616( .i (n3564), .o (n3616) );
  assign n3617 = ( n3608 & n3615 ) | ( n3608 & ~n3616 ) | ( n3615 & ~n3616 ) ;
  buffer buf_n3618( .i (n3617), .o (n3618) );
  assign n3619 = ( n3380 & ~n3584 ) | ( n3380 & n3618 ) | ( ~n3584 & n3618 ) ;
  assign n3620 = n3506 & ~n3618 ;
  assign n3621 = ( n3585 & n3619 ) | ( n3585 & ~n3620 ) | ( n3619 & ~n3620 ) ;
  buffer buf_n3622( .i (n3621), .o (n3622) );
  assign n3623 = ( n583 & n3587 ) | ( n583 & ~n3622 ) | ( n3587 & ~n3622 ) ;
  assign n3624 = n407 & ~n3622 ;
  assign n3625 = ( ~n3588 & n3623 ) | ( ~n3588 & n3624 ) | ( n3623 & n3624 ) ;
  assign n3626 = n3595 & n3625 ;
  assign n3627 = ( ~n3554 & n3555 ) | ( ~n3554 & n3626 ) | ( n3555 & n3626 ) ;
  assign n3628 = n3523 & n3627 ;
  assign n3629 = ( n3440 & ~n3441 ) | ( n3440 & n3628 ) | ( ~n3441 & n3628 ) ;
  buffer buf_n3630( .i (n3629), .o (n3630) );
  assign n3631 = ( n3357 & n3404 ) | ( n3357 & n3630 ) | ( n3404 & n3630 ) ;
  buffer buf_n78( .i (n77), .o (n78) );
  assign n3632 = n78 & n3630 ;
  assign n3633 = ( ~n3358 & n3631 ) | ( ~n3358 & n3632 ) | ( n3631 & n3632 ) ;
  assign n3634 = n449 & ~n3633 ;
  assign n3635 = ~n297 & n2021 ;
  buffer buf_n3636( .i (n3635), .o (n3636) );
  buffer buf_n3637( .i (n3636), .o (n3637) );
  buffer buf_n3638( .i (n3637), .o (n3638) );
  buffer buf_n3639( .i (n3638), .o (n3639) );
  buffer buf_n3640( .i (n3639), .o (n3640) );
  buffer buf_n3641( .i (n3640), .o (n3641) );
  buffer buf_n3642( .i (n3641), .o (n3642) );
  buffer buf_n3643( .i (n3642), .o (n3643) );
  buffer buf_n3644( .i (n3643), .o (n3644) );
  buffer buf_n3645( .i (n3644), .o (n3645) );
  assign n3646 = ( n1415 & n1769 ) | ( n1415 & ~n3644 ) | ( n1769 & ~n3644 ) ;
  assign n3647 = n3645 & n3646 ;
  buffer buf_n3648( .i (n3647), .o (n3648) );
  buffer buf_n3649( .i (n3648), .o (n3649) );
  buffer buf_n3650( .i (n3649), .o (n3650) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  assign n3651 = ( n572 & ~n3162 ) | ( n572 & n3648 ) | ( ~n3162 & n3648 ) ;
  assign n3652 = n2731 & ~n3651 ;
  assign n3653 = ( n2343 & n3650 ) | ( n2343 & ~n3652 ) | ( n3650 & ~n3652 ) ;
  buffer buf_n3654( .i (n3653), .o (n3654) );
  buffer buf_n3655( .i (n3654), .o (n3655) );
  assign n3656 = ( n141 & n380 ) | ( n141 & ~n3654 ) | ( n380 & ~n3654 ) ;
  assign n3657 = n3451 | n3504 ;
  buffer buf_n3658( .i (n3657), .o (n3658) );
  buffer buf_n3659( .i (n3658), .o (n3659) );
  buffer buf_n3660( .i (n3659), .o (n3660) );
  buffer buf_n3661( .i (n3660), .o (n3661) );
  buffer buf_n3662( .i (n3661), .o (n3662) );
  assign n3663 = n2741 & n2938 ;
  buffer buf_n3664( .i (n3143), .o (n3664) );
  buffer buf_n3665( .i (n3664), .o (n3665) );
  assign n3666 = ( n3662 & n3663 ) | ( n3662 & ~n3665 ) | ( n3663 & ~n3665 ) ;
  assign n3667 = ( n339 & n3451 ) | ( n339 & n3590 ) | ( n3451 & n3590 ) ;
  buffer buf_n3668( .i (n3667), .o (n3668) );
  buffer buf_n3669( .i (n3668), .o (n3669) );
  buffer buf_n3670( .i (n404), .o (n3670) );
  assign n3671 = ( ~n2606 & n3175 ) | ( ~n2606 & n3670 ) | ( n3175 & n3670 ) ;
  assign n3672 = n3668 | n3671 ;
  assign n3673 = ( ~n342 & n3669 ) | ( ~n342 & n3672 ) | ( n3669 & n3672 ) ;
  assign n3674 = ( n2102 & ~n3043 ) | ( n2102 & n3673 ) | ( ~n3043 & n3673 ) ;
  assign n3675 = n3217 & n3255 ;
  assign n3676 = n2201 & n3675 ;
  buffer buf_n3677( .i (n3676), .o (n3677) );
  buffer buf_n3678( .i (n3677), .o (n3678) );
  buffer buf_n3679( .i (n338), .o (n3679) );
  assign n3680 = ~n3677 & n3679 ;
  assign n3681 = ( n2606 & n3678 ) | ( n2606 & ~n3680 ) | ( n3678 & ~n3680 ) ;
  assign n3682 = n307 & n3681 ;
  assign n3683 = n3480 & n3682 ;
  buffer buf_n3684( .i (n3009), .o (n3684) );
  assign n3685 = n3683 & ~n3684 ;
  assign n3686 = ( n2490 & n3674 ) | ( n2490 & ~n3685 ) | ( n3674 & ~n3685 ) ;
  buffer buf_n3687( .i (n3686), .o (n3687) );
  assign n3688 = ( n3292 & n3666 ) | ( n3292 & n3687 ) | ( n3666 & n3687 ) ;
  assign n3689 = ( ~n396 & n2908 ) | ( ~n396 & n2909 ) | ( n2908 & n2909 ) ;
  buffer buf_n3690( .i (n3689), .o (n3690) );
  buffer buf_n3691( .i (n3690), .o (n3691) );
  buffer buf_n3692( .i (n3691), .o (n3692) );
  buffer buf_n3693( .i (n3692), .o (n3693) );
  buffer buf_n3694( .i (n3693), .o (n3694) );
  buffer buf_n3695( .i (n3694), .o (n3695) );
  buffer buf_n3696( .i (n3695), .o (n3696) );
  buffer buf_n3697( .i (n3696), .o (n3697) );
  buffer buf_n3698( .i (n3697), .o (n3698) );
  buffer buf_n3699( .i (n3590), .o (n3699) );
  buffer buf_n3700( .i (n3699), .o (n3700) );
  assign n3701 = ( n307 & n3698 ) | ( n307 & ~n3700 ) | ( n3698 & ~n3700 ) ;
  buffer buf_n3702( .i (n3272), .o (n3702) );
  buffer buf_n3703( .i (n3702), .o (n3703) );
  buffer buf_n3704( .i (n3703), .o (n3704) );
  buffer buf_n3705( .i (n3704), .o (n3705) );
  assign n3706 = ( n406 & n3698 ) | ( n406 & ~n3705 ) | ( n3698 & ~n3705 ) ;
  assign n3707 = n3701 & n3706 ;
  buffer buf_n3708( .i (n3707), .o (n3708) );
  buffer buf_n3709( .i (n3708), .o (n3709) );
  buffer buf_n2979( .i (n2978), .o (n2979) );
  assign n3710 = ( n2979 & n3664 ) | ( n2979 & n3708 ) | ( n3664 & n3708 ) ;
  assign n3711 = ~n3709 & n3710 ;
  assign n3712 = ( n3292 & ~n3687 ) | ( n3292 & n3711 ) | ( ~n3687 & n3711 ) ;
  assign n3713 = n3688 & ~n3712 ;
  buffer buf_n3714( .i (n140), .o (n3714) );
  assign n3715 = ~n3713 & n3714 ;
  assign n3716 = ( n3655 & n3656 ) | ( n3655 & n3715 ) | ( n3656 & n3715 ) ;
  assign n3717 = n2728 & n3367 ;
  assign n3718 = n2962 & n3717 ;
  buffer buf_n3719( .i (n3718), .o (n3719) );
  buffer buf_n3720( .i (n3719), .o (n3720) );
  buffer buf_n3721( .i (n3720), .o (n3721) );
  buffer buf_n3722( .i (n2429), .o (n3722) );
  assign n3723 = n2653 & ~n3722 ;
  assign n3724 = n2049 & n3700 ;
  buffer buf_n3725( .i (n3724), .o (n3725) );
  buffer buf_n3726( .i (n3725), .o (n3726) );
  assign n3727 = n3722 & ~n3726 ;
  assign n3728 = n3723 | n3727 ;
  buffer buf_n3729( .i (n3110), .o (n3729) );
  assign n3730 = ( n3719 & n3728 ) | ( n3719 & ~n3729 ) | ( n3728 & ~n3729 ) ;
  assign n3731 = n3374 | n3730 ;
  assign n3732 = ( ~n243 & n3721 ) | ( ~n243 & n3731 ) | ( n3721 & n3731 ) ;
  assign n3733 = ~n404 & n3445 ;
  assign n3734 = ( ~n2676 & n3418 ) | ( ~n2676 & n3733 ) | ( n3418 & n3733 ) ;
  assign n3735 = n581 & n3699 ;
  buffer buf_n3736( .i (n3442), .o (n3736) );
  assign n3737 = ~n3505 & n3736 ;
  assign n3738 = ( n3451 & ~n3504 ) | ( n3451 & n3737 ) | ( ~n3504 & n3737 ) ;
  assign n3739 = n3699 | n3738 ;
  assign n3740 = ( n3734 & n3735 ) | ( n3734 & n3739 ) | ( n3735 & n3739 ) ;
  buffer buf_n3741( .i (n3740), .o (n3741) );
  buffer buf_n3742( .i (n3741), .o (n3742) );
  buffer buf_n3743( .i (n308), .o (n3743) );
  assign n3744 = ~n3741 & n3743 ;
  assign n3745 = n296 & ~n362 ;
  buffer buf_n3746( .i (n3745), .o (n3746) );
  buffer buf_n3747( .i (n3746), .o (n3747) );
  assign n3748 = ( n2616 & ~n3300 ) | ( n2616 & n3746 ) | ( ~n3300 & n3746 ) ;
  assign n3749 = ( n3090 & n3747 ) | ( n3090 & n3748 ) | ( n3747 & n3748 ) ;
  buffer buf_n3750( .i (n3749), .o (n3750) );
  buffer buf_n3751( .i (n3750), .o (n3751) );
  assign n3752 = n230 | n3750 ;
  buffer buf_n3753( .i (n2905), .o (n3753) );
  assign n3754 = ( n3465 & ~n3558 ) | ( n3465 & n3753 ) | ( ~n3558 & n3753 ) ;
  assign n3755 = ( n3200 & n3389 ) | ( n3200 & ~n3754 ) | ( n3389 & ~n3754 ) ;
  assign n3756 = ( n326 & ~n358 ) | ( n326 & n391 ) | ( ~n358 & n391 ) ;
  assign n3757 = n293 & n3756 ;
  assign n3758 = ( ~n294 & n393 ) | ( ~n294 & n3757 ) | ( n393 & n3757 ) ;
  buffer buf_n3759( .i (n3758), .o (n3759) );
  assign n3760 = ( n296 & ~n362 ) | ( n296 & n3759 ) | ( ~n362 & n3759 ) ;
  assign n3761 = n2310 & n3759 ;
  buffer buf_n3762( .i (n295), .o (n3762) );
  buffer buf_n3763( .i (n3762), .o (n3763) );
  assign n3764 = ( n3760 & n3761 ) | ( n3760 & ~n3763 ) | ( n3761 & ~n3763 ) ;
  buffer buf_n3765( .i (n3764), .o (n3765) );
  buffer buf_n3766( .i (n3765), .o (n3766) );
  assign n3767 = ~n3753 & n3765 ;
  assign n3768 = ( n3637 & n3766 ) | ( n3637 & n3767 ) | ( n3766 & n3767 ) ;
  assign n3769 = n3755 & n3768 ;
  assign n3770 = ( n3751 & ~n3752 ) | ( n3751 & n3769 ) | ( ~n3752 & n3769 ) ;
  buffer buf_n3771( .i (n3770), .o (n3771) );
  buffer buf_n3772( .i (n336), .o (n3772) );
  buffer buf_n3773( .i (n3772), .o (n3773) );
  assign n3774 = ( ~n3702 & n3771 ) | ( ~n3702 & n3773 ) | ( n3771 & n3773 ) ;
  assign n3775 = n3496 & n3771 ;
  assign n3776 = ( n3703 & n3774 ) | ( n3703 & n3775 ) | ( n3774 & n3775 ) ;
  buffer buf_n3777( .i (n3776), .o (n3777) );
  buffer buf_n3778( .i (n3777), .o (n3778) );
  assign n3779 = ( n1415 & n3502 ) | ( n1415 & ~n3777 ) | ( n3502 & ~n3777 ) ;
  assign n3780 = ( ~n1847 & n2647 ) | ( ~n1847 & n3505 ) | ( n2647 & n3505 ) ;
  assign n3781 = ( n401 & n1899 ) | ( n401 & ~n3564 ) | ( n1899 & ~n3564 ) ;
  buffer buf_n3782( .i (n2453), .o (n3782) );
  buffer buf_n3783( .i (n575), .o (n3783) );
  assign n3784 = ( n2669 & n3782 ) | ( n2669 & ~n3783 ) | ( n3782 & ~n3783 ) ;
  assign n3785 = ~n1899 & n3784 ;
  assign n3786 = ( n3616 & n3781 ) | ( n3616 & ~n3785 ) | ( n3781 & ~n3785 ) ;
  buffer buf_n3787( .i (n3786), .o (n3787) );
  assign n3788 = ( n3590 & n3780 ) | ( n3590 & n3787 ) | ( n3780 & n3787 ) ;
  assign n3789 = n402 & ~n1846 ;
  assign n3790 = ( n579 & ~n2154 ) | ( n579 & n3789 ) | ( ~n2154 & n3789 ) ;
  buffer buf_n3791( .i (n3589), .o (n3791) );
  assign n3792 = ( n3787 & n3790 ) | ( n3787 & ~n3791 ) | ( n3790 & ~n3791 ) ;
  assign n3793 = n3788 & n3792 ;
  assign n3794 = n3502 | n3793 ;
  assign n3795 = ( n3778 & n3779 ) | ( n3778 & n3794 ) | ( n3779 & n3794 ) ;
  assign n3796 = ( ~n335 & n3638 ) | ( ~n335 & n3782 ) | ( n3638 & n3782 ) ;
  assign n3797 = n187 & n293 ;
  buffer buf_n3798( .i (n3797), .o (n3798) );
  buffer buf_n3799( .i (n3798), .o (n3799) );
  buffer buf_n3800( .i (n3799), .o (n3800) );
  buffer buf_n3801( .i (n3800), .o (n3801) );
  buffer buf_n3802( .i (n3801), .o (n3802) );
  buffer buf_n3803( .i (n3802), .o (n3803) );
  assign n3804 = n398 & ~n3802 ;
  assign n3805 = ( n229 & ~n3803 ) | ( n229 & n3804 ) | ( ~n3803 & n3804 ) ;
  buffer buf_n3806( .i (n3753), .o (n3806) );
  buffer buf_n3807( .i (n3806), .o (n3807) );
  assign n3808 = n3805 | n3807 ;
  assign n3809 = ( n3639 & ~n3796 ) | ( n3639 & n3808 ) | ( ~n3796 & n3808 ) ;
  assign n3810 = n3616 & n3809 ;
  assign n3811 = n231 | n495 ;
  assign n3812 = ~n3616 & n3811 ;
  assign n3813 = n3810 | n3812 ;
  assign n3814 = n3506 | n3813 ;
  buffer buf_n3815( .i (n3814), .o (n3815) );
  buffer buf_n3816( .i (n3815), .o (n3816) );
  assign n3817 = ~n2965 & n3815 ;
  assign n3818 = ( ~n3366 & n3816 ) | ( ~n3366 & n3817 ) | ( n3816 & n3817 ) ;
  assign n3819 = n3795 & n3818 ;
  assign n3820 = ( n3742 & n3744 ) | ( n3742 & n3819 ) | ( n3744 & n3819 ) ;
  buffer buf_n3821( .i (n229), .o (n3821) );
  buffer buf_n3822( .i (n3821), .o (n3822) );
  assign n3823 = ( ~n401 & n3255 ) | ( ~n401 & n3822 ) | ( n3255 & n3822 ) ;
  buffer buf_n3824( .i (n3566), .o (n3824) );
  assign n3825 = ( n2028 & n3822 ) | ( n2028 & n3824 ) | ( n3822 & n3824 ) ;
  assign n3826 = ~n3823 & n3825 ;
  buffer buf_n3827( .i (n3826), .o (n3827) );
  buffer buf_n3828( .i (n3827), .o (n3828) );
  assign n3829 = n3505 & n3589 ;
  assign n3830 = ( n3679 & ~n3827 ) | ( n3679 & n3829 ) | ( ~n3827 & n3829 ) ;
  assign n3831 = n3828 & n3830 ;
  buffer buf_n3832( .i (n3831), .o (n3832) );
  buffer buf_n3833( .i (n3832), .o (n3833) );
  assign n3834 = ~n3303 & n3807 ;
  buffer buf_n3835( .i (n3834), .o (n3835) );
  assign n3836 = n3442 & n3835 ;
  assign n3837 = ( n3305 & n3430 ) | ( n3305 & ~n3835 ) | ( n3430 & ~n3835 ) ;
  assign n3838 = ( n3589 & n3836 ) | ( n3589 & ~n3837 ) | ( n3836 & ~n3837 ) ;
  buffer buf_n3839( .i (n3838), .o (n3839) );
  buffer buf_n3840( .i (n3839), .o (n3840) );
  assign n3841 = ( n3418 & n3500 ) | ( n3418 & n3839 ) | ( n3500 & n3839 ) ;
  assign n3842 = ( n1961 & ~n3566 ) | ( n1961 & n3807 ) | ( ~n3566 & n3807 ) ;
  assign n3843 = ( n696 & n3304 ) | ( n696 & ~n3842 ) | ( n3304 & ~n3842 ) ;
  buffer buf_n3844( .i (n3843), .o (n3844) );
  buffer buf_n3845( .i (n3844), .o (n3845) );
  assign n3846 = n3736 & n3844 ;
  assign n3847 = ( ~n2917 & n3845 ) | ( ~n2917 & n3846 ) | ( n3845 & n3846 ) ;
  assign n3848 = n3500 | n3847 ;
  assign n3849 = ( ~n3840 & n3841 ) | ( ~n3840 & n3848 ) | ( n3841 & n3848 ) ;
  buffer buf_n3850( .i (n2293), .o (n3850) );
  buffer buf_n3851( .i (n3850), .o (n3851) );
  assign n3852 = ( n2642 & ~n3753 ) | ( n2642 & n3851 ) | ( ~n3753 & n3851 ) ;
  assign n3853 = ( n3278 & n3806 ) | ( n3278 & n3852 ) | ( n3806 & n3852 ) ;
  buffer buf_n3854( .i (n3853), .o (n3854) );
  buffer buf_n3855( .i (n2887), .o (n3855) );
  assign n3856 = ( ~n503 & n3854 ) | ( ~n503 & n3855 ) | ( n3854 & n3855 ) ;
  assign n3857 = n3822 & n3854 ;
  assign n3858 = ( n504 & n3856 ) | ( n504 & n3857 ) | ( n3856 & n3857 ) ;
  buffer buf_n3859( .i (n228), .o (n3859) );
  assign n3860 = ( ~n2886 & n3561 ) | ( ~n2886 & n3859 ) | ( n3561 & n3859 ) ;
  buffer buf_n3183( .i (n3182), .o (n3183) );
  buffer buf_n3184( .i (n3183), .o (n3184) );
  buffer buf_n3185( .i (n3184), .o (n3185) );
  buffer buf_n3186( .i (n3185), .o (n3186) );
  assign n3861 = ( n2148 & n2905 ) | ( n2148 & ~n3487 ) | ( n2905 & ~n3487 ) ;
  buffer buf_n3862( .i (n3485), .o (n3862) );
  buffer buf_n3863( .i (n3862), .o (n3863) );
  assign n3864 = ( n3186 & n3861 ) | ( n3186 & n3863 ) | ( n3861 & n3863 ) ;
  assign n3865 = ( n2886 & n3859 ) | ( n2886 & n3864 ) | ( n3859 & n3864 ) ;
  assign n3866 = n3860 & ~n3865 ;
  buffer buf_n3867( .i (n3866), .o (n3867) );
  buffer buf_n3868( .i (n3867), .o (n3868) );
  buffer buf_n3869( .i (n3410), .o (n3869) );
  buffer buf_n3870( .i (n3869), .o (n3870) );
  assign n3871 = n3867 | n3870 ;
  assign n3872 = ( ~n3858 & n3868 ) | ( ~n3858 & n3871 ) | ( n3868 & n3871 ) ;
  assign n3873 = n3791 | n3872 ;
  buffer buf_n2787( .i (n2786), .o (n2787) );
  buffer buf_n2788( .i (n2787), .o (n2788) );
  buffer buf_n2789( .i (n2788), .o (n2789) );
  buffer buf_n3874( .i (n3025), .o (n3874) );
  assign n3875 = n3639 & ~n3874 ;
  buffer buf_n3876( .i (n3874), .o (n3876) );
  assign n3877 = ( n2789 & n3875 ) | ( n2789 & ~n3876 ) | ( n3875 & ~n3876 ) ;
  assign n3878 = ~n3773 & n3877 ;
  assign n3879 = n3791 & ~n3878 ;
  assign n3880 = n3873 & ~n3879 ;
  buffer buf_n3881( .i (n3880), .o (n3881) );
  assign n3882 = ( n3832 & n3849 ) | ( n3832 & ~n3881 ) | ( n3849 & ~n3881 ) ;
  assign n3883 = n308 | n3881 ;
  assign n3884 = ( n3833 & ~n3882 ) | ( n3833 & n3883 ) | ( ~n3882 & n3883 ) ;
  buffer buf_n3885( .i (n3884), .o (n3885) );
  assign n3886 = ( n3110 & ~n3820 ) | ( n3110 & n3885 ) | ( ~n3820 & n3885 ) ;
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  buffer buf_n2235( .i (n2234), .o (n2235) );
  buffer buf_n2236( .i (n2235), .o (n2236) );
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  assign n3887 = n3700 & ~n3705 ;
  buffer buf_n3888( .i (n3705), .o (n3888) );
  assign n3889 = ( ~n552 & n3887 ) | ( ~n552 & n3888 ) | ( n3887 & n3888 ) ;
  assign n3890 = n2237 | n3889 ;
  assign n3891 = ( n406 & ~n2738 ) | ( n406 & n3177 ) | ( ~n2738 & n3177 ) ;
  assign n3892 = n3135 & n3791 ;
  buffer buf_n3893( .i (n3504), .o (n3893) );
  assign n3894 = n3892 & n3893 ;
  assign n3895 = n406 & n3894 ;
  assign n3896 = ( ~n2727 & n3891 ) | ( ~n2727 & n3895 ) | ( n3891 & n3895 ) ;
  buffer buf_n3897( .i (n3863), .o (n3897) );
  buffer buf_n3898( .i (n3897), .o (n3898) );
  assign n3899 = n2043 | n3898 ;
  assign n3900 = ( ~n631 & n2044 ) | ( ~n631 & n3899 ) | ( n2044 & n3899 ) ;
  buffer buf_n3901( .i (n3900), .o (n3901) );
  buffer buf_n3902( .i (n3901), .o (n3902) );
  assign n3903 = ( n778 & n2453 ) | ( n778 & n3897 ) | ( n2453 & n3897 ) ;
  buffer buf_n3904( .i (n3903), .o (n3904) );
  buffer buf_n3905( .i (n3782), .o (n3905) );
  assign n3906 = ( n2152 & n3904 ) | ( n2152 & ~n3905 ) | ( n3904 & ~n3905 ) ;
  assign n3907 = n3564 & n3904 ;
  assign n3908 = ( n1586 & n3906 ) | ( n1586 & n3907 ) | ( n3906 & n3907 ) ;
  assign n3909 = n2640 | n3299 ;
  assign n3910 = ( n298 & n3300 ) | ( n298 & n3909 ) | ( n3300 & n3909 ) ;
  assign n3911 = ~n397 & n3850 ;
  assign n3912 = ( ~n790 & n3910 ) | ( ~n790 & n3911 ) | ( n3910 & n3911 ) ;
  buffer buf_n3913( .i (n3912), .o (n3913) );
  buffer buf_n3914( .i (n3913), .o (n3914) );
  assign n3915 = n3410 & n3913 ;
  assign n3916 = ( n2643 & ~n2907 ) | ( n2643 & n3467 ) | ( ~n2907 & n3467 ) ;
  assign n3917 = n398 | n3863 ;
  assign n3918 = ( ~n1843 & n3897 ) | ( ~n1843 & n3917 ) | ( n3897 & n3917 ) ;
  assign n3919 = n3916 & n3918 ;
  assign n3920 = ( ~n3914 & n3915 ) | ( ~n3914 & n3919 ) | ( n3915 & n3919 ) ;
  buffer buf_n3921( .i (n3920), .o (n3921) );
  assign n3922 = ( ~n3901 & n3908 ) | ( ~n3901 & n3921 ) | ( n3908 & n3921 ) ;
  assign n3923 = n3702 & n3921 ;
  assign n3924 = ( n3902 & n3922 ) | ( n3902 & n3923 ) | ( n3922 & n3923 ) ;
  buffer buf_n3925( .i (n3924), .o (n3925) );
  buffer buf_n3926( .i (n3925), .o (n3926) );
  buffer buf_n3927( .i (n3175), .o (n3927) );
  assign n3928 = n3925 | n3927 ;
  assign n3929 = n2882 & ~n3851 ;
  buffer buf_n3930( .i (n3929), .o (n3930) );
  buffer buf_n3931( .i (n3930), .o (n3931) );
  buffer buf_n3932( .i (n3931), .o (n3932) );
  buffer buf_n2885( .i (n2884), .o (n2885) );
  buffer buf_n3933( .i (n3093), .o (n3933) );
  assign n3934 = ( n3782 & n3930 ) | ( n3782 & ~n3933 ) | ( n3930 & ~n3933 ) ;
  assign n3935 = ( n2230 & n2885 ) | ( n2230 & ~n3934 ) | ( n2885 & ~n3934 ) ;
  assign n3936 = ~n3932 & n3935 ;
  buffer buf_n3937( .i (n3936), .o (n3937) );
  buffer buf_n3938( .i (n3937), .o (n3938) );
  assign n3939 = ( ~n3679 & n3703 ) | ( ~n3679 & n3937 ) | ( n3703 & n3937 ) ;
  buffer buf_n2538( .i (n2537), .o (n2538) );
  buffer buf_n2539( .i (n2538), .o (n2539) );
  buffer buf_n2540( .i (n2539), .o (n2540) );
  buffer buf_n2541( .i (n2540), .o (n2541) );
  buffer buf_n2542( .i (n2541), .o (n2542) );
  buffer buf_n2543( .i (n2542), .o (n2543) );
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n3940( .i (n3467), .o (n3940) );
  buffer buf_n3941( .i (n3940), .o (n3941) );
  buffer buf_n3942( .i (n3941), .o (n3942) );
  buffer buf_n3943( .i (n3942), .o (n3943) );
  assign n3944 = ( n2545 & n3306 ) | ( n2545 & ~n3943 ) | ( n3306 & ~n3943 ) ;
  assign n3945 = n3703 & n3944 ;
  assign n3946 = ( ~n3938 & n3939 ) | ( ~n3938 & n3945 ) | ( n3939 & n3945 ) ;
  assign n3947 = ~n2844 & n3941 ;
  buffer buf_n3948( .i (n3947), .o (n3948) );
  buffer buf_n3949( .i (n3948), .o (n3949) );
  buffer buf_n3950( .i (n3949), .o (n3950) );
  assign n3951 = ( n1846 & n2972 ) | ( n1846 & n3442 ) | ( n2972 & n3442 ) ;
  assign n3952 = ( n3496 & ~n3948 ) | ( n3496 & n3951 ) | ( ~n3948 & n3951 ) ;
  buffer buf_n3953( .i (n3431), .o (n3953) );
  assign n3954 = n3952 & n3953 ;
  assign n3955 = ( n3893 & n3950 ) | ( n3893 & ~n3954 ) | ( n3950 & ~n3954 ) ;
  assign n3956 = n3946 | n3955 ;
  assign n3957 = ( ~n3926 & n3928 ) | ( ~n3926 & n3956 ) | ( n3928 & n3956 ) ;
  assign n3958 = n3896 | n3957 ;
  assign n3959 = ( ~n2238 & n3890 ) | ( ~n2238 & n3958 ) | ( n3890 & n3958 ) ;
  buffer buf_n3960( .i (n2490), .o (n3960) );
  assign n3961 = ( n3885 & n3959 ) | ( n3885 & ~n3960 ) | ( n3959 & ~n3960 ) ;
  assign n3962 = n3886 | n3961 ;
  buffer buf_n3963( .i (n3962), .o (n3963) );
  buffer buf_n3964( .i (n3963), .o (n3964) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  assign n3965 = n620 & ~n3963 ;
  assign n3966 = ( n3732 & n3964 ) | ( n3732 & ~n3965 ) | ( n3964 & ~n3965 ) ;
  assign n3967 = n3716 | n3966 ;
  buffer buf_n3968( .i (n448), .o (n3968) );
  assign n3969 = n3967 & ~n3968 ;
  assign n3970 = n3634 | n3969 ;
  assign n3971 = n485 | n3970 ;
  buffer buf_n450( .i (n449), .o (n450) );
  assign n3972 = ~n1106 & n2814 ;
  buffer buf_n3531( .i (n3530), .o (n3531) );
  buffer buf_n3532( .i (n3531), .o (n3532) );
  buffer buf_n3533( .i (n3532), .o (n3533) );
  buffer buf_n3534( .i (n3533), .o (n3534) );
  buffer buf_n3535( .i (n3534), .o (n3535) );
  buffer buf_n3536( .i (n3535), .o (n3536) );
  buffer buf_n3537( .i (n3536), .o (n3537) );
  buffer buf_n3538( .i (n3537), .o (n3538) );
  buffer buf_n3539( .i (n3538), .o (n3539) );
  buffer buf_n2208( .i (n2207), .o (n2208) );
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n2211( .i (n2210), .o (n2211) );
  buffer buf_n2212( .i (n2211), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  buffer buf_n2214( .i (n2213), .o (n2214) );
  assign n3973 = ( n2214 & n2651 ) | ( n2214 & ~n3538 ) | ( n2651 & ~n3538 ) ;
  assign n3974 = n2650 & ~n3700 ;
  buffer buf_n3975( .i (n3974), .o (n3975) );
  assign n3977 = ( n3539 & n3973 ) | ( n3539 & n3975 ) | ( n3973 & n3975 ) ;
  buffer buf_n3978( .i (n3927), .o (n3978) );
  assign n3979 = n2520 & n3978 ;
  assign n3980 = n84 & n117 ;
  buffer buf_n3981( .i (n3980), .o (n3981) );
  buffer buf_n3982( .i (n3981), .o (n3982) );
  buffer buf_n3983( .i (n3982), .o (n3983) );
  buffer buf_n3984( .i (n3983), .o (n3984) );
  buffer buf_n3985( .i (n3984), .o (n3985) );
  buffer buf_n3986( .i (n3985), .o (n3986) );
  buffer buf_n3987( .i (n3986), .o (n3987) );
  buffer buf_n3988( .i (n3987), .o (n3988) );
  buffer buf_n3989( .i (n3988), .o (n3989) );
  buffer buf_n3990( .i (n3989), .o (n3990) );
  buffer buf_n3991( .i (n3990), .o (n3991) );
  buffer buf_n3992( .i (n3991), .o (n3992) );
  buffer buf_n3993( .i (n3992), .o (n3993) );
  buffer buf_n3994( .i (n3993), .o (n3994) );
  buffer buf_n3995( .i (n3994), .o (n3995) );
  buffer buf_n3996( .i (n3995), .o (n3996) );
  buffer buf_n3997( .i (n3996), .o (n3997) );
  assign n3998 = n3330 & n3997 ;
  assign n3999 = n3979 & n3998 ;
  assign n4000 = n3977 | n3999 ;
  assign n4001 = ( n1107 & n3972 ) | ( n1107 & ~n4000 ) | ( n3972 & ~n4000 ) ;
  buffer buf_n4002( .i (n4001), .o (n4002) );
  buffer buf_n4003( .i (n4002), .o (n4003) );
  assign n4004 = ( n207 & ~n313 ) | ( n207 & n4002 ) | ( ~n313 & n4002 ) ;
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2660), .o (n2661) );
  buffer buf_n2662( .i (n2661), .o (n2662) );
  assign n4005 = ( n407 & n3009 ) | ( n407 & n3330 ) | ( n3009 & n3330 ) ;
  buffer buf_n4006( .i (n3330), .o (n4006) );
  assign n4007 = ( n2662 & n4005 ) | ( n2662 & ~n4006 ) | ( n4005 & ~n4006 ) ;
  assign n4008 = ( n402 & ~n3271 ) | ( n402 & n3876 ) | ( ~n3271 & n3876 ) ;
  buffer buf_n4009( .i (n3822), .o (n4009) );
  buffer buf_n4010( .i (n3824), .o (n4010) );
  assign n4011 = ~n4009 & n4010 ;
  assign n4012 = ( n67 & n4008 ) | ( n67 & n4011 ) | ( n4008 & n4011 ) ;
  buffer buf_n4013( .i (n4012), .o (n4013) );
  buffer buf_n4014( .i (n4013), .o (n4014) );
  assign n4015 = n2518 & ~n4013 ;
  assign n4016 = n3221 & n3995 ;
  assign n4017 = ( n4014 & n4015 ) | ( n4014 & n4016 ) | ( n4015 & n4016 ) ;
  buffer buf_n4018( .i (n4017), .o (n4018) );
  buffer buf_n4019( .i (n4018), .o (n4019) );
  assign n4020 = n3143 & n4018 ;
  assign n4021 = ( n4007 & n4019 ) | ( n4007 & n4020 ) | ( n4019 & n4020 ) ;
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n3070( .i (n3069), .o (n3070) );
  buffer buf_n3071( .i (n3070), .o (n3071) );
  buffer buf_n1954( .i (n1953), .o (n1954) );
  buffer buf_n1955( .i (n1954), .o (n1955) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  assign n4022 = ( n1959 & n3069 ) | ( n1959 & n3535 ) | ( n3069 & n3535 ) ;
  assign n4023 = n3418 & ~n4022 ;
  assign n4024 = ( n2402 & n3071 ) | ( n2402 & ~n4023 ) | ( n3071 & ~n4023 ) ;
  assign n4025 = ~n3480 & n4024 ;
  assign n4026 = ( ~n2051 & n3725 ) | ( ~n2051 & n4025 ) | ( n3725 & n4025 ) ;
  buffer buf_n4027( .i (n4026), .o (n4027) );
  assign n4028 = ( n2731 & n4021 ) | ( n2731 & ~n4027 ) | ( n4021 & ~n4027 ) ;
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  assign n4029 = n1005 & ~n3684 ;
  assign n4030 = ~n344 & n4029 ;
  buffer buf_n4031( .i (n2814), .o (n4031) );
  assign n4032 = ( n4027 & n4030 ) | ( n4027 & n4031 ) | ( n4030 & n4031 ) ;
  assign n4033 = n4028 & ~n4032 ;
  assign n4034 = n313 | n4033 ;
  assign n4035 = ( n4003 & ~n4004 ) | ( n4003 & n4034 ) | ( ~n4004 & n4034 ) ;
  buffer buf_n4036( .i (n4035), .o (n4036) );
  buffer buf_n4037( .i (n4036), .o (n4037) );
  buffer buf_n2631( .i (n2630), .o (n2631) );
  buffer buf_n2632( .i (n2631), .o (n2632) );
  buffer buf_n2655( .i (n2654), .o (n2655) );
  buffer buf_n2656( .i (n2655), .o (n2656) );
  buffer buf_n2657( .i (n2656), .o (n2657) );
  assign n4038 = ( ~n1295 & n2632 ) | ( ~n1295 & n2657 ) | ( n2632 & n2657 ) ;
  assign n4039 = n3060 | n3526 ;
  assign n4040 = ( n788 & n3061 ) | ( n788 & n4039 ) | ( n3061 & n4039 ) ;
  buffer buf_n4041( .i (n4040), .o (n4041) );
  buffer buf_n4042( .i (n4041), .o (n4042) );
  buffer buf_n4043( .i (n4042), .o (n4043) );
  buffer buf_n4044( .i (n4043), .o (n4044) );
  buffer buf_n4045( .i (n4044), .o (n4045) );
  buffer buf_n4046( .i (n4045), .o (n4046) );
  buffer buf_n4047( .i (n4046), .o (n4047) );
  buffer buf_n4048( .i (n4047), .o (n4048) );
  buffer buf_n4049( .i (n4048), .o (n4049) );
  buffer buf_n4050( .i (n4049), .o (n4050) );
  buffer buf_n4051( .i (n4050), .o (n4051) );
  buffer buf_n4052( .i (n4051), .o (n4052) );
  buffer buf_n4053( .i (n4052), .o (n4053) );
  buffer buf_n4054( .i (n4053), .o (n4054) );
  assign n4055 = n2987 & n4054 ;
  buffer buf_n4056( .i (n206), .o (n4056) );
  assign n4057 = n4055 & ~n4056 ;
  assign n4058 = ~n2632 & n4057 ;
  assign n4059 = ( n279 & n4038 ) | ( n279 & ~n4058 ) | ( n4038 & ~n4058 ) ;
  buffer buf_n3976( .i (n3975), .o (n3976) );
  assign n4060 = n3366 & n3888 ;
  assign n4061 = n3407 & ~n4060 ;
  assign n4062 = n3976 | n4061 ;
  buffer buf_n4063( .i (n4062), .o (n4063) );
  buffer buf_n4064( .i (n4063), .o (n4064) );
  buffer buf_n4065( .i (n4064), .o (n4065) );
  assign n4066 = n2328 & n3665 ;
  assign n4067 = ( n979 & n4063 ) | ( n979 & n4066 ) | ( n4063 & n4066 ) ;
  assign n4068 = n2942 & ~n4067 ;
  buffer buf_n4069( .i (n3729), .o (n4069) );
  buffer buf_n4070( .i (n4069), .o (n4070) );
  assign n4071 = ( n4065 & ~n4068 ) | ( n4065 & n4070 ) | ( ~n4068 & n4070 ) ;
  buffer buf_n4072( .i (n3699), .o (n4072) );
  buffer buf_n4073( .i (n4072), .o (n4073) );
  assign n4074 = ( ~n3480 & n3978 ) | ( ~n3480 & n4073 ) | ( n3978 & n4073 ) ;
  buffer buf_n4075( .i (n3502), .o (n4075) );
  assign n4076 = ( ~n1911 & n4073 ) | ( ~n1911 & n4075 ) | ( n4073 & n4075 ) ;
  assign n4077 = n4074 | n4076 ;
  buffer buf_n4078( .i (n4077), .o (n4078) );
  buffer buf_n4079( .i (n4078), .o (n4079) );
  buffer buf_n4080( .i (n4079), .o (n4080) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  assign n4081 = n501 & ~n3009 ;
  assign n4082 = ~n3743 & n4081 ;
  buffer buf_n4083( .i (n2290), .o (n4083) );
  assign n4084 = n4082 & n4083 ;
  assign n4085 = ( n3665 & n4078 ) | ( n3665 & n4084 ) | ( n4078 & n4084 ) ;
  assign n4086 = ~n2268 & n4085 ;
  assign n4087 = ( n3374 & n4080 ) | ( n3374 & n4086 ) | ( n4080 & n4086 ) ;
  buffer buf_n4088( .i (n3893), .o (n4088) );
  assign n4089 = ( n858 & ~n3927 ) | ( n858 & n4088 ) | ( ~n3927 & n4088 ) ;
  assign n4090 = ( n856 & n859 ) | ( n856 & n4089 ) | ( n859 & n4089 ) ;
  buffer buf_n4091( .i (n4090), .o (n4091) );
  buffer buf_n4092( .i (n4091), .o (n4092) );
  buffer buf_n2921( .i (n2920), .o (n2921) );
  buffer buf_n4093( .i (n2744), .o (n4093) );
  assign n4094 = n2920 & n4093 ;
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  assign n4095 = ( n805 & ~n2402 ) | ( n805 & n3658 ) | ( ~n2402 & n3658 ) ;
  buffer buf_n4096( .i (n3105), .o (n4096) );
  assign n4097 = n4095 & n4096 ;
  assign n4098 = ( ~n2921 & n4094 ) | ( ~n2921 & n4097 ) | ( n4094 & n4097 ) ;
  assign n4099 = ( n67 & n1958 ) | ( n67 & n2916 ) | ( n1958 & n2916 ) ;
  assign n4100 = n2916 & ~n3496 ;
  buffer buf_n4101( .i (n3271), .o (n4101) );
  buffer buf_n4102( .i (n4101), .o (n4102) );
  assign n4103 = ( n4099 & n4100 ) | ( n4099 & ~n4102 ) | ( n4100 & ~n4102 ) ;
  buffer buf_n4104( .i (n4103), .o (n4104) );
  buffer buf_n4105( .i (n4104), .o (n4105) );
  assign n4106 = ( n632 & n3272 ) | ( n632 & n3772 ) | ( n3272 & n3772 ) ;
  assign n4107 = n3772 & ~n4009 ;
  assign n4108 = ( ~n633 & n4106 ) | ( ~n633 & n4107 ) | ( n4106 & n4107 ) ;
  assign n4109 = ( n3242 & n3798 ) | ( n3242 & ~n3984 ) | ( n3798 & ~n3984 ) ;
  assign n4110 = n3985 & n4109 ;
  buffer buf_n4111( .i (n4110), .o (n4111) );
  buffer buf_n4112( .i (n4111), .o (n4112) );
  buffer buf_n4113( .i (n4112), .o (n4113) );
  assign n4114 = ( n2876 & n3557 ) | ( n2876 & ~n4111 ) | ( n3557 & ~n4111 ) ;
  buffer buf_n4115( .i (n2909), .o (n4115) );
  buffer buf_n4116( .i (n4115), .o (n4116) );
  assign n4117 = n4114 & n4116 ;
  assign n4118 = ( n3806 & n4113 ) | ( n3806 & ~n4117 ) | ( n4113 & ~n4117 ) ;
  buffer buf_n4119( .i (n4118), .o (n4119) );
  buffer buf_n4120( .i (n4119), .o (n4120) );
  assign n4121 = ( n2004 & n3905 ) | ( n2004 & ~n4119 ) | ( n3905 & ~n4119 ) ;
  assign n4122 = ~n909 & n1844 ;
  buffer buf_n4123( .i (n1821), .o (n4123) );
  assign n4124 = n4122 & n4123 ;
  assign n4125 = ( n4120 & n4121 ) | ( n4120 & n4124 ) | ( n4121 & n4124 ) ;
  buffer buf_n4126( .i (n4125), .o (n4126) );
  buffer buf_n4127( .i (n3943), .o (n4127) );
  assign n4128 = ( n4108 & n4126 ) | ( n4108 & ~n4127 ) | ( n4126 & ~n4127 ) ;
  assign n4129 = ( n1957 & n3271 ) | ( n1957 & ~n3772 ) | ( n3271 & ~n3772 ) ;
  assign n4130 = n3279 & n3821 ;
  assign n4131 = ( n62 & n3465 ) | ( n62 & ~n3851 ) | ( n3465 & ~n3851 ) ;
  assign n4132 = n398 | n3851 ;
  assign n4133 = ( n63 & ~n4131 ) | ( n63 & n4132 ) | ( ~n4131 & n4132 ) ;
  buffer buf_n4134( .i (n3092), .o (n4134) );
  assign n4135 = n399 & ~n4134 ;
  assign n4136 = n4133 & n4135 ;
  assign n4137 = ( ~n3280 & n4130 ) | ( ~n3280 & n4136 ) | ( n4130 & n4136 ) ;
  buffer buf_n4138( .i (n336), .o (n4138) );
  assign n4139 = n4137 | n4138 ;
  assign n4140 = ( n1958 & ~n4129 ) | ( n1958 & n4139 ) | ( ~n4129 & n4139 ) ;
  assign n4141 = ( n4126 & n4127 ) | ( n4126 & ~n4140 ) | ( n4127 & ~n4140 ) ;
  assign n4142 = n4128 | n4141 ;
  assign n4143 = n62 & ~n2295 ;
  buffer buf_n4144( .i (n3850), .o (n4144) );
  buffer buf_n4145( .i (n4144), .o (n4145) );
  assign n4146 = ( ~n2296 & n4143 ) | ( ~n2296 & n4145 ) | ( n4143 & n4145 ) ;
  assign n4147 = ( ~n2911 & n3690 ) | ( ~n2911 & n4041 ) | ( n3690 & n4041 ) ;
  assign n4148 = n1836 & n3982 ;
  assign n4149 = ( n57 & n2764 ) | ( n57 & n4148 ) | ( n2764 & n4148 ) ;
  assign n4150 = ~n1879 & n4149 ;
  buffer buf_n4151( .i (n4150), .o (n4151) );
  buffer buf_n4152( .i (n4151), .o (n4152) );
  buffer buf_n4153( .i (n4152), .o (n4153) );
  buffer buf_n4154( .i (n122), .o (n4154) );
  buffer buf_n4155( .i (n4154), .o (n4155) );
  assign n4156 = ( n2292 & ~n4151 ) | ( n2292 & n4155 ) | ( ~n4151 & n4155 ) ;
  assign n4157 = n3850 & n4156 ;
  assign n4158 = ( n4144 & n4153 ) | ( n4144 & ~n4157 ) | ( n4153 & ~n4157 ) ;
  assign n4159 = n4147 | n4158 ;
  assign n4160 = n4146 | n4159 ;
  assign n4161 = ~n3869 & n4160 ;
  buffer buf_n4162( .i (n4161), .o (n4162) );
  buffer buf_n4163( .i (n4162), .o (n4163) );
  assign n4164 = ( n396 & ~n2908 ) | ( n396 & n2909 ) | ( ~n2908 & n2909 ) ;
  assign n4165 = ( n2616 & n3557 ) | ( n2616 & n4164 ) | ( n3557 & n4164 ) ;
  assign n4166 = n228 & ~n4165 ;
  assign n4167 = n4134 & n4166 ;
  buffer buf_n4168( .i (n4167), .o (n4168) );
  buffer buf_n4169( .i (n4168), .o (n4169) );
  buffer buf_n4170( .i (n94), .o (n4170) );
  buffer buf_n4171( .i (n4145), .o (n4171) );
  assign n4172 = n4170 & n4171 ;
  assign n4173 = ( n2230 & ~n4168 ) | ( n2230 & n4172 ) | ( ~n4168 & n4172 ) ;
  assign n4174 = n4169 & n4173 ;
  assign n4175 = n4162 | n4174 ;
  assign n4176 = ( n4102 & n4163 ) | ( n4102 & n4175 ) | ( n4163 & n4175 ) ;
  buffer buf_n4177( .i (n4176), .o (n4177) );
  assign n4178 = ( ~n4104 & n4142 ) | ( ~n4104 & n4177 ) | ( n4142 & n4177 ) ;
  assign n4179 = n2744 & ~n4177 ;
  assign n4180 = ( n4105 & n4178 ) | ( n4105 & ~n4179 ) | ( n4178 & ~n4179 ) ;
  buffer buf_n4181( .i (n4180), .o (n4181) );
  assign n4182 = ( n4091 & n4098 ) | ( n4091 & ~n4181 ) | ( n4098 & ~n4181 ) ;
  buffer buf_n4183( .i (n3043), .o (n4183) );
  assign n4184 = ~n4181 & n4183 ;
  assign n4185 = ( ~n4092 & n4182 ) | ( ~n4092 & n4184 ) | ( n4182 & n4184 ) ;
  buffer buf_n4186( .i (n4185), .o (n4186) );
  buffer buf_n4187( .i (n4186), .o (n4187) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  assign n4188 = n1109 & n4186 ;
  assign n4189 = ( n4087 & n4187 ) | ( n4087 & n4188 ) | ( n4187 & n4188 ) ;
  assign n4190 = n4071 & n4189 ;
  assign n4191 = ( ~n4036 & n4059 ) | ( ~n4036 & n4190 ) | ( n4059 & n4190 ) ;
  assign n4192 = n4037 & n4191 ;
  assign n4193 = n450 | n4192 ;
  assign n4194 = n485 & n4193 ;
  assign n4195 = n3971 & ~n4194 ;
  assign y0 = n967 ;
  assign y1 = n1202 ;
  assign y2 = n1414 ;
  assign y3 = n1668 ;
  assign y4 = n1951 ;
  assign y5 = n2121 ;
  assign y6 = n2190 ;
  assign y7 = n2356 ;
  assign y8 = n2517 ;
  assign y9 = n2838 ;
  assign y10 = n3006 ;
  assign y11 = n3133 ;
  assign y12 = n3351 ;
  assign y13 = n4195 ;
endmodule
