module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 ;
  buffer buf_n7( .i (x0), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (x1), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n77( .i (x4), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n42( .i (x2), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n59( .i (x3), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  assign n113 = ( n32 & n49 ) | ( n32 & n66 ) | ( n49 & n66 ) ;
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  assign n121 = n92 & ~n120 ;
  assign n122 = ( n41 & n93 ) | ( n41 & ~n121 ) | ( n93 & ~n121 ) ;
  assign n123 = n24 & n122 ;
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  assign n124 = n35 & ~n52 ;
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  assign n130 = n71 & ~n89 ;
  assign n131 = ( n55 & ~n72 ) | ( n55 & n130 ) | ( ~n72 & n130 ) ;
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  assign n134 = ( ~n40 & n57 ) | ( ~n40 & n132 ) | ( n57 & n132 ) ;
  assign n135 = ( n129 & ~n133 ) | ( n129 & n134 ) | ( ~n133 & n134 ) ;
  assign n136 = n24 & ~n135 ;
  assign n137 = ( n20 & n72 ) | ( n20 & n90 ) | ( n72 & n90 ) ;
  buffer buf_n94( .i (x5), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  assign n138 = ( n9 & n61 ) | ( n9 & ~n96 ) | ( n61 & ~n96 ) ;
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  assign n150 = n137 & ~n149 ;
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  assign n153 = n51 & ~n86 ;
  assign n154 = n69 & n153 ;
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  assign n157 = n31 | n65 ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n159 = ( n15 & ~n50 ) | ( n15 & n158 ) | ( ~n50 & n158 ) ;
  assign n160 = ( n15 & n67 ) | ( n15 & ~n158 ) | ( n67 & ~n158 ) ;
  assign n161 = ( n34 & ~n159 ) | ( n34 & n160 ) | ( ~n159 & n160 ) ;
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  assign n165 = ( n18 & ~n36 ) | ( n18 & n162 ) | ( ~n36 & n162 ) ;
  assign n166 = n155 & ~n165 ;
  assign n167 = ( n156 & n164 ) | ( n156 & ~n166 ) | ( n164 & ~n166 ) ;
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  assign n171 = ( n40 & ~n57 ) | ( n40 & n168 ) | ( ~n57 & n168 ) ;
  assign n172 = n151 & ~n171 ;
  assign n173 = ( n152 & n170 ) | ( n152 & ~n172 ) | ( n170 & ~n172 ) ;
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  assign n174 = ( n34 & ~n68 ) | ( n34 & n103 ) | ( ~n68 & n103 ) ;
  buffer buf_n175( .i (n174), .o (n175) );
  assign n176 = ( n53 & ~n105 ) | ( n53 & n175 ) | ( ~n105 & n175 ) ;
  assign n177 = ( n36 & n53 ) | ( n36 & ~n175 ) | ( n53 & ~n175 ) ;
  assign n178 = n176 & ~n177 ;
  assign n179 = n20 & ~n178 ;
  assign n180 = ~n51 & n68 ;
  buffer buf_n181( .i (n180), .o (n181) );
  assign n188 = ~n105 & n181 ;
  assign n189 = n37 & n188 ;
  assign n190 = n20 | n189 ;
  assign n191 = ~n179 & n190 ;
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  assign n194 = ~n93 & n192 ;
  assign n195 = ( n15 & ~n50 ) | ( n15 & n67 ) | ( ~n50 & n67 ) ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n201 = ( ~n17 & n35 ) | ( ~n17 & n196 ) | ( n35 & n196 ) ;
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  assign n206 = ( ~n54 & n71 ) | ( ~n54 & n202 ) | ( n71 & n202 ) ;
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  assign n209 = ~n200 & n207 ;
  assign n210 = ( ~n205 & n208 ) | ( ~n205 & n209 ) | ( n208 & n209 ) ;
  assign n211 = ( n33 & ~n50 ) | ( n33 & n67 ) | ( ~n50 & n67 ) ;
  buffer buf_n212( .i (n211), .o (n212) );
  assign n215 = n34 & n86 ;
  assign n216 = ( n69 & ~n212 ) | ( n69 & n215 ) | ( ~n212 & n215 ) ;
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n219 = ( ~n89 & n214 ) | ( ~n89 & n217 ) | ( n214 & n217 ) ;
  assign n220 = ( ~n72 & n218 ) | ( ~n72 & n219 ) | ( n218 & n219 ) ;
  assign n221 = n21 & ~n220 ;
  buffer buf_n182( .i (n181), .o (n182) );
  assign n222 = ~n89 & n182 ;
  assign n223 = n38 & n222 ;
  assign n224 = n21 | n223 ;
  assign n225 = ~n221 & n224 ;
  assign n226 = n210 | n225 ;
  assign n227 = ( n193 & ~n194 ) | ( n193 & n226 ) | ( ~n194 & n226 ) ;
  buffer buf_n228( .i (n49), .o (n228) );
  assign n229 = ( n33 & ~n102 ) | ( n33 & n228 ) | ( ~n102 & n228 ) ;
  assign n230 = n114 | n229 ;
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  assign n233 = n105 & n231 ;
  assign n234 = ( ~n117 & n232 ) | ( ~n117 & n233 ) | ( n232 & n233 ) ;
  assign n235 = n90 & ~n234 ;
  assign n236 = ~n69 & n104 ;
  buffer buf_n237( .i (n104), .o (n237) );
  assign n238 = ( n36 & n236 ) | ( n36 & n237 ) | ( n236 & n237 ) ;
  assign n239 = n54 & n238 ;
  assign n240 = n90 | n239 ;
  assign n241 = ~n235 & n240 ;
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  assign n244 = ~n23 & n242 ;
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n245( .i (n88), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  assign n247 = ~n107 & n246 ;
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n73( .i (n72), .o (n73) );
  assign n252 = ~n19 & n37 ;
  assign n253 = ~n55 & n252 ;
  assign n254 = n73 & n253 ;
  assign n255 = n248 & n254 ;
  buffer buf_n256( .i (n33), .o (n256) );
  assign n257 = ( n16 & n51 ) | ( n16 & ~n256 ) | ( n51 & ~n256 ) ;
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  assign n260 = n54 | n259 ;
  assign n261 = ( n18 & ~n70 ) | ( n18 & n258 ) | ( ~n70 & n258 ) ;
  buffer buf_n262( .i (n53), .o (n262) );
  assign n263 = n261 & n262 ;
  assign n264 = n260 & ~n263 ;
  assign n265 = n91 & ~n264 ;
  buffer buf_n266( .i (n35), .o (n266) );
  buffer buf_n267( .i (n52), .o (n267) );
  assign n268 = n266 | n267 ;
  assign n269 = ( ~n37 & n125 ) | ( ~n37 & n268 ) | ( n125 & n268 ) ;
  buffer buf_n270( .i (n71), .o (n270) );
  assign n271 = n269 & n270 ;
  assign n272 = n91 | n271 ;
  assign n273 = ~n265 & n272 ;
  assign n274 = n255 | n273 ;
  assign n275 = ( n243 & ~n244 ) | ( n243 & n274 ) | ( ~n244 & n274 ) ;
  assign n276 = n70 | n267 ;
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n279( .i (n19), .o (n279) );
  assign n280 = ( ~n55 & n277 ) | ( ~n55 & n279 ) | ( n277 & n279 ) ;
  assign n281 = ( ~n38 & n277 ) | ( ~n38 & n279 ) | ( n277 & n279 ) ;
  assign n282 = ( n127 & ~n280 ) | ( n127 & n281 ) | ( ~n280 & n281 ) ;
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  assign n285 = ~n93 & n283 ;
  buffer buf_n286( .i (n70), .o (n286) );
  assign n287 = n262 & ~n286 ;
  buffer buf_n288( .i (n287), .o (n288) );
  assign n289 = ( n21 & ~n91 ) | ( n21 & n288 ) | ( ~n91 & n288 ) ;
  assign n290 = ~n22 & n289 ;
  assign n291 = ( n13 & ~n65 ) | ( n13 & n100 ) | ( ~n65 & n100 ) ;
  assign n292 = ( ~n32 & n101 ) | ( ~n32 & n291 ) | ( n101 & n291 ) ;
  buffer buf_n293( .i (n292), .o (n293) );
  assign n296 = n103 & ~n293 ;
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  assign n299 = n295 | n297 ;
  assign n300 = ( ~n106 & n298 ) | ( ~n106 & n299 ) | ( n298 & n299 ) ;
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  assign n303 = ~n56 & n301 ;
  assign n304 = n237 & ~n267 ;
  buffer buf_n305( .i (n266), .o (n305) );
  assign n306 = ( n19 & n304 ) | ( n19 & n305 ) | ( n304 & n305 ) ;
  assign n307 = ~n38 & n306 ;
  assign n308 = ( n46 & n98 ) | ( n46 & n139 ) | ( n98 & n139 ) ;
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  assign n313 = ( n13 & n65 ) | ( n13 & n309 ) | ( n65 & n309 ) ;
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  assign n316 = n143 & ~n314 ;
  assign n317 = ( n312 & ~n315 ) | ( n312 & n316 ) | ( ~n315 & n316 ) ;
  assign n318 = n87 & ~n317 ;
  assign n319 = n49 | n101 ;
  buffer buf_n320( .i (n64), .o (n320) );
  assign n321 = n100 | n320 ;
  buffer buf_n322( .i (n48), .o (n322) );
  assign n323 = ~n321 & n322 ;
  assign n324 = ( ~n228 & n319 ) | ( ~n228 & n323 ) | ( n319 & n323 ) ;
  assign n325 = n16 & n324 ;
  assign n326 = n87 | n325 ;
  assign n327 = ~n318 & n326 ;
  assign n328 = n305 & ~n327 ;
  buffer buf_n329( .i (n228), .o (n329) );
  assign n330 = ( n86 & n103 ) | ( n86 & n329 ) | ( n103 & n329 ) ;
  buffer buf_n331( .i (n85), .o (n331) );
  buffer buf_n332( .i (n102), .o (n332) );
  assign n333 = ( ~n68 & n331 ) | ( ~n68 & n332 ) | ( n331 & n332 ) ;
  assign n334 = n330 & ~n333 ;
  assign n335 = n18 & n334 ;
  assign n336 = n305 | n335 ;
  assign n337 = ~n328 & n336 ;
  assign n338 = n307 | n337 ;
  assign n339 = ( n302 & ~n303 ) | ( n302 & n338 ) | ( ~n303 & n338 ) ;
  assign n340 = n290 | n339 ;
  assign n341 = ( n284 & ~n285 ) | ( n284 & n340 ) | ( ~n285 & n340 ) ;
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  assign n342 = ( n245 & n262 ) | ( n245 & n286 ) | ( n262 & n286 ) ;
  buffer buf_n343( .i (n342), .o (n343) );
  assign n344 = n39 & ~n343 ;
  assign n345 = ~n39 & n343 ;
  assign n346 = n344 | n345 ;
  assign n347 = n110 & ~n346 ;
  buffer buf_n278( .i (n277), .o (n278) );
  assign n348 = ( ~n56 & n278 ) | ( ~n56 & n288 ) | ( n278 & n288 ) ;
  assign n349 = n92 & n348 ;
  assign n350 = n110 | n349 ;
  assign n351 = ~n347 & n350 ;
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  assign n352 = ( n58 & n75 ) | ( n58 & n110 ) | ( n75 & n110 ) ;
  assign n353 = n74 & n92 ;
  buffer buf_n354( .i (n109), .o (n354) );
  assign n355 = ( n75 & n353 ) | ( n75 & n354 ) | ( n353 & n354 ) ;
  assign n356 = ( n187 & n352 ) | ( n187 & ~n355 ) | ( n352 & ~n355 ) ;
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n357( .i (n246), .o (n357) );
  assign n358 = ( n73 & n108 ) | ( n73 & n357 ) | ( n108 & n357 ) ;
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  assign n361 = ~n93 & n359 ;
  assign n362 = ( ~n76 & n360 ) | ( ~n76 & n361 ) | ( n360 & n361 ) ;
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  assign y0 = n123 ;
  assign y1 = n136 ;
  assign y2 = n173 ;
  assign y3 = n227 ;
  assign y4 = n275 ;
  assign y5 = n341 ;
  assign y6 = n351 ;
  assign y7 = n356 ;
  assign y8 = n362 ;
  assign y9 = n251 ;
  assign y10 = 1'b0 ;
  assign y11 = n112 ;
endmodule
