module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n8 , n10 , n11 , n12 , n13 , n14 , n15 , n17 , n18 , n19 , n20 , n21 , n22 , n24 , n25 , n26 , n27 , n28 , n29 , n31 , n32 , n33 , n34 , n35 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 ;
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n10( .i (x1), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  assign n46 = n5 & n13 ;
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n31( .i (x4), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  assign n48 = n3 & n32 ;
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n17( .i (x2), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n24( .i (x3), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  assign n51 = n19 & n26 ;
  buffer buf_n52( .i (n51), .o (n52) );
  assign n54 = n50 & n52 ;
  assign n55 = n47 | n54 ;
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  assign n58 = n24 & n31 ;
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  assign n61 = ~n10 & n17 ;
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  assign n64 = n60 & n63 ;
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  assign n68 = n15 & ~n22 ;
  assign n69 = n8 & ~n68 ;
  assign n70 = ~n67 & n69 ;
  buffer buf_n37( .i (x5), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  assign n71 = n11 & n38 ;
  buffer buf_n72( .i (n71), .o (n72) );
  assign n75 = n60 & n72 ;
  assign n76 = ~n59 & n62 ;
  assign n77 = n11 & n25 ;
  assign n78 = n4 & n77 ;
  assign n79 = ( n5 & n76 ) | ( n5 & n78 ) | ( n76 & n78 ) ;
  assign n80 = n75 | n79 ;
  buffer buf_n81( .i (n80), .o (n81) );
  assign n82 = ~n18 & n38 ;
  buffer buf_n83( .i (n82), .o (n83) );
  assign n84 = n49 & n83 ;
  buffer buf_n85( .i (n84), .o (n85) );
  assign n86 = ( n5 & n13 ) | ( n5 & n20 ) | ( n13 & n20 ) ;
  assign n87 = ~n6 & n86 ;
  assign n88 = ( n15 & n85 ) | ( n15 & n87 ) | ( n85 & n87 ) ;
  assign n89 = n81 | n88 ;
  buffer buf_n90( .i (n89), .o (n90) );
  assign n91 = n25 & ~n32 ;
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  assign n95 = n47 & n94 ;
  assign n96 = n31 & n37 ;
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  assign n99 = n11 | n25 ;
  buffer buf_n100( .i (n99), .o (n100) );
  assign n101 = n98 | n100 ;
  buffer buf_n102( .i (n101), .o (n102) );
  assign n103 = ~n65 & n102 ;
  assign n104 = ~n95 & n103 ;
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  assign n105 = n21 & ~n50 ;
  assign n106 = ( ~n29 & n85 ) | ( ~n29 & n105 ) | ( n85 & n105 ) ;
  assign n107 = n60 & n83 ;
  buffer buf_n108( .i (n107), .o (n108) );
  assign n109 = n6 | n14 ;
  assign n110 = ( n7 & ~n108 ) | ( n7 & n109 ) | ( ~n108 & n109 ) ;
  assign n111 = ~n106 & n110 ;
  assign n112 = n104 & n111 ;
  assign n113 = n32 & ~n38 ;
  buffer buf_n114( .i (n113), .o (n114) );
  assign n120 = ~n100 & n114 ;
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n33( .i (n32), .o (n33) );
  assign n121 = n19 & ~n33 ;
  assign n122 = n40 & n121 ;
  assign n123 = n120 | n122 ;
  assign n124 = n7 & n123 ;
  assign n125 = n4 & n97 ;
  assign n126 = ~n33 & n62 ;
  assign n127 = n125 | n126 ;
  assign n128 = n28 & n127 ;
  assign n129 = ~n20 & n92 ;
  assign n130 = n20 & n98 ;
  assign n131 = ( n14 & n129 ) | ( n14 & n130 ) | ( n129 & n130 ) ;
  assign n132 = n128 | n131 ;
  assign n133 = n124 | n132 ;
  buffer buf_n134( .i (n4), .o (n134) );
  buffer buf_n135( .i (n19), .o (n135) );
  assign n136 = n134 & n135 ;
  buffer buf_n137( .i (n10), .o (n137) );
  buffer buf_n138( .i (n24), .o (n138) );
  buffer buf_n139( .i (n31), .o (n139) );
  assign n140 = ( n137 & n138 ) | ( n137 & ~n139 ) | ( n138 & ~n139 ) ;
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n143( .i (n18), .o (n143) );
  assign n144 = n39 & n143 ;
  assign n145 = ( n72 & ~n141 ) | ( n72 & n144 ) | ( ~n141 & n144 ) ;
  assign n146 = ( n6 & n136 ) | ( n6 & n145 ) | ( n136 & n145 ) ;
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  assign n147 = ( n12 & n26 ) | ( n12 & n143 ) | ( n26 & n143 ) ;
  assign n148 = ~n83 & n147 ;
  buffer buf_n149( .i (n134), .o (n149) );
  assign n150 = ( n35 & n148 ) | ( n35 & n149 ) | ( n148 & n149 ) ;
  assign n151 = ~n146 & n150 ;
  assign n152 = ~n81 & n151 ;
  assign n153 = n133 | n152 ;
  buffer buf_n142( .i (n141), .o (n142) );
  assign n154 = ( n14 & n21 ) | ( n14 & ~n142 ) | ( n21 & ~n142 ) ;
  buffer buf_n155( .i (n154), .o (n155) );
  assign n156 = n8 & ~n155 ;
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  assign n157 = ( n8 & n43 ) | ( n8 & ~n155 ) | ( n43 & ~n155 ) ;
  assign n158 = n26 | n33 ;
  buffer buf_n159( .i (n158), .o (n159) );
  assign n160 = n21 & ~n159 ;
  buffer buf_n161( .i (n13), .o (n161) );
  buffer buf_n162( .i (n135), .o (n162) );
  assign n163 = n161 & n162 ;
  assign n164 = ( n35 & n161 ) | ( n35 & n162 ) | ( n161 & n162 ) ;
  assign n165 = ( n160 & ~n163 ) | ( n160 & n164 ) | ( ~n163 & n164 ) ;
  assign n166 = n43 | n165 ;
  assign n167 = ( n156 & ~n157 ) | ( n156 & n166 ) | ( ~n157 & n166 ) ;
  assign n168 = ( n18 & n138 ) | ( n18 & n139 ) | ( n138 & n139 ) ;
  buffer buf_n169( .i (n168), .o (n169) );
  assign n172 = n72 & ~n169 ;
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  assign n175 = n41 & n52 ;
  assign n176 = ( ~n53 & n171 ) | ( ~n53 & n175 ) | ( n171 & n175 ) ;
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  assign n177 = n74 & ~n173 ;
  assign n178 = ( n174 & n176 ) | ( n174 & ~n177 ) | ( n176 & ~n177 ) ;
  buffer buf_n179( .i (n178), .o (n179) );
  assign n180 = n22 | n29 ;
  assign n181 = ( n22 & n29 ) | ( n22 & ~n42 ) | ( n29 & ~n42 ) ;
  assign n182 = ~n42 & n94 ;
  assign n183 = ( n180 & ~n181 ) | ( n180 & n182 ) | ( ~n181 & n182 ) ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n185 = n40 & ~n60 ;
  assign n186 = n159 & n185 ;
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  assign y0 = n57 ;
  assign y1 = n70 ;
  assign y2 = n90 ;
  assign y3 = n112 ;
  assign y4 = n153 ;
  assign y5 = n167 ;
  assign y6 = n179 ;
  assign y7 = n184 ;
  assign y8 = n189 ;
  assign y9 = n119 ;
  assign y10 = 1'b0 ;
  assign y11 = n45 ;
endmodule
