module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( b_4_ , a_1_ , a_2_ , b_1_ , b_7_ , a_6_ , a_4_ , b_2_ , a_7_ , a_5_ , b_5_ , b_3_ , b_6_ , b_0_ , a_3_ , a_0_ , s_1_ , s_8_ , s_3_ , s_5_ , s_9_ , s_2_ , s_11_ , s_15_ , s_4_ , s_10_ , s_14_ , s_7_ , s_13_ , s_12_ , s_6_ , s_0_ );
  input b_4_ , a_1_ , a_2_ , b_1_ , b_7_ , a_6_ , a_4_ , b_2_ , a_7_ , a_5_ , b_5_ , b_3_ , b_6_ , b_0_ , a_3_ , a_0_ ;
  output s_1_ , s_8_ , s_3_ , s_5_ , s_9_ , s_2_ , s_11_ , s_15_ , s_4_ , s_10_ , s_14_ , s_7_ , s_13_ , s_12_ , s_6_ , s_0_ ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 ;
  assign n17 = a_1_ & b_0_ ;
  buffer buf_n18( .i (n17), .o (n18) );
  assign n19 = b_1_ & a_0_ ;
  buffer buf_n20( .i (n19), .o (n20) );
  assign n21 = n18 & n20 ;
  buffer buf_n22( .i (n21), .o (n22) );
  assign n23 = n18 | n20 ;
  buffer buf_n24( .i (n23), .o (n24) );
  assign n25 = ~n22 & n24 ;
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  assign n84 = a_1_ & b_6_ ;
  buffer buf_n85( .i (n84), .o (n85) );
  assign n86 = b_4_ & a_2_ ;
  buffer buf_n87( .i (n86), .o (n87) );
  assign n88 = b_3_ & a_3_ ;
  buffer buf_n89( .i (n88), .o (n89) );
  assign n90 = n87 & n89 ;
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  assign n96 = a_1_ & b_5_ ;
  buffer buf_n97( .i (n96), .o (n97) );
  assign n98 = n87 | n89 ;
  buffer buf_n99( .i (n98), .o (n99) );
  assign n100 = ~n91 & n99 ;
  buffer buf_n101( .i (n100), .o (n101) );
  assign n102 = n97 & n101 ;
  buffer buf_n103( .i (n102), .o (n103) );
  assign n104 = n95 | n103 ;
  buffer buf_n105( .i (n104), .o (n105) );
  assign n106 = n85 & n105 ;
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  assign n112 = b_7_ & a_0_ ;
  buffer buf_n113( .i (n112), .o (n113) );
  assign n114 = n85 | n105 ;
  buffer buf_n115( .i (n114), .o (n115) );
  assign n116 = ~n107 & n115 ;
  buffer buf_n117( .i (n116), .o (n117) );
  assign n118 = n113 & n117 ;
  buffer buf_n119( .i (n118), .o (n119) );
  assign n120 = n111 | n119 ;
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  assign n130 = a_1_ & b_7_ ;
  buffer buf_n131( .i (n130), .o (n131) );
  assign n132 = a_2_ & b_6_ ;
  buffer buf_n133( .i (n132), .o (n133) );
  assign n134 = b_4_ & a_3_ ;
  buffer buf_n135( .i (n134), .o (n135) );
  assign n136 = a_4_ & b_3_ ;
  buffer buf_n137( .i (n136), .o (n137) );
  assign n138 = n135 & n137 ;
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  assign n144 = n135 | n137 ;
  buffer buf_n145( .i (n144), .o (n145) );
  assign n146 = ~n139 & n145 ;
  buffer buf_n147( .i (n146), .o (n147) );
  assign n148 = a_2_ & b_5_ ;
  buffer buf_n149( .i (n148), .o (n149) );
  assign n150 = n147 & n149 ;
  buffer buf_n151( .i (n150), .o (n151) );
  assign n152 = n143 | n151 ;
  buffer buf_n153( .i (n152), .o (n153) );
  assign n154 = n133 & n153 ;
  buffer buf_n155( .i (n154), .o (n155) );
  assign n160 = n133 | n153 ;
  buffer buf_n161( .i (n160), .o (n161) );
  assign n162 = ~n155 & n161 ;
  buffer buf_n163( .i (n162), .o (n163) );
  assign n164 = n131 & n163 ;
  buffer buf_n165( .i (n164), .o (n165) );
  assign n166 = n131 | n163 ;
  buffer buf_n167( .i (n166), .o (n167) );
  assign n168 = ~n165 & n167 ;
  buffer buf_n169( .i (n168), .o (n169) );
  assign n170 = b_5_ & a_3_ ;
  buffer buf_n171( .i (n170), .o (n171) );
  assign n172 = b_4_ & a_4_ ;
  buffer buf_n173( .i (n172), .o (n173) );
  assign n174 = a_5_ & b_3_ ;
  buffer buf_n175( .i (n174), .o (n175) );
  assign n176 = n173 & n175 ;
  buffer buf_n177( .i (n176), .o (n177) );
  assign n182 = n173 | n175 ;
  buffer buf_n183( .i (n182), .o (n183) );
  assign n184 = ~n177 & n183 ;
  buffer buf_n185( .i (n184), .o (n185) );
  assign n186 = n171 & n185 ;
  buffer buf_n187( .i (n186), .o (n187) );
  assign n188 = n171 | n185 ;
  buffer buf_n189( .i (n188), .o (n189) );
  assign n190 = ~n187 & n189 ;
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  assign n197 = b_1_ & a_6_ ;
  buffer buf_n198( .i (n197), .o (n198) );
  assign n203 = a_7_ & b_0_ ;
  buffer buf_n204( .i (n203), .o (n204) );
  assign n205 = n198 & n204 ;
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  assign n211 = b_2_ & a_5_ ;
  buffer buf_n212( .i (n211), .o (n212) );
  assign n213 = n198 | n204 ;
  buffer buf_n214( .i (n213), .o (n214) );
  assign n215 = ~n206 & n214 ;
  buffer buf_n216( .i (n215), .o (n216) );
  assign n217 = n212 & n216 ;
  buffer buf_n218( .i (n217), .o (n218) );
  assign n219 = n210 | n218 ;
  buffer buf_n220( .i (n219), .o (n220) );
  assign n221 = b_1_ & a_7_ ;
  assign n222 = a_6_ & b_2_ ;
  assign n223 = n221 | n222 ;
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  assign n224 = b_2_ & a_7_ ;
  buffer buf_n225( .i (n224), .o (n225) );
  assign n226 = n202 & n225 ;
  buffer buf_n227( .i (n226), .o (n227) );
  assign n231 = n223 & ~n227 ;
  buffer buf_n232( .i (n231), .o (n232) );
  assign n233 = n220 & n232 ;
  buffer buf_n234( .i (n233), .o (n234) );
  assign n239 = n220 | n232 ;
  buffer buf_n240( .i (n239), .o (n240) );
  assign n241 = ~n234 & n240 ;
  buffer buf_n242( .i (n241), .o (n242) );
  assign n243 = n196 & n242 ;
  buffer buf_n244( .i (n243), .o (n244) );
  assign n245 = n196 | n242 ;
  buffer buf_n246( .i (n245), .o (n246) );
  assign n247 = ~n244 & n246 ;
  buffer buf_n248( .i (n247), .o (n248) );
  assign n249 = n212 | n216 ;
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = ~n218 & n250 ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n253 = a_5_ & b_0_ ;
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  assign n256 = n198 & n255 ;
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  assign n262 = a_4_ & b_2_ ;
  buffer buf_n263( .i (n262), .o (n263) );
  assign n264 = b_1_ & a_5_ ;
  assign n265 = a_6_ & b_0_ ;
  assign n266 = n264 | n265 ;
  assign n267 = ~n257 & n266 ;
  buffer buf_n268( .i (n267), .o (n268) );
  assign n269 = n263 & n268 ;
  buffer buf_n270( .i (n269), .o (n270) );
  assign n271 = n261 | n270 ;
  buffer buf_n272( .i (n271), .o (n272) );
  assign n273 = n252 & n272 ;
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  assign n279 = n147 | n149 ;
  buffer buf_n280( .i (n279), .o (n280) );
  assign n281 = ~n151 & n280 ;
  buffer buf_n282( .i (n281), .o (n282) );
  assign n283 = n252 | n272 ;
  buffer buf_n284( .i (n283), .o (n284) );
  assign n285 = ~n274 & n284 ;
  buffer buf_n286( .i (n285), .o (n286) );
  assign n287 = n282 & n286 ;
  buffer buf_n288( .i (n287), .o (n288) );
  assign n289 = n278 | n288 ;
  buffer buf_n290( .i (n289), .o (n290) );
  assign n291 = n248 & n290 ;
  buffer buf_n292( .i (n291), .o (n292) );
  assign n297 = n248 | n290 ;
  buffer buf_n298( .i (n297), .o (n298) );
  assign n299 = ~n292 & n298 ;
  buffer buf_n300( .i (n299), .o (n300) );
  assign n301 = n169 & n300 ;
  buffer buf_n302( .i (n301), .o (n302) );
  assign n303 = n169 | n300 ;
  buffer buf_n304( .i (n303), .o (n304) );
  assign n305 = ~n302 & n304 ;
  buffer buf_n306( .i (n305), .o (n306) );
  assign n307 = n282 | n286 ;
  buffer buf_n308( .i (n307), .o (n308) );
  assign n309 = ~n288 & n308 ;
  buffer buf_n310( .i (n309), .o (n310) );
  assign n311 = n263 | n268 ;
  buffer buf_n312( .i (n311), .o (n312) );
  assign n313 = ~n270 & n312 ;
  buffer buf_n314( .i (n313), .o (n314) );
  assign n315 = b_1_ & a_4_ ;
  buffer buf_n316( .i (n315), .o (n316) );
  assign n317 = n254 & n316 ;
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  assign n323 = b_2_ & a_3_ ;
  buffer buf_n324( .i (n323), .o (n324) );
  assign n325 = n254 | n316 ;
  buffer buf_n326( .i (n325), .o (n326) );
  assign n327 = ~n318 & n326 ;
  buffer buf_n328( .i (n327), .o (n328) );
  assign n329 = n324 & n328 ;
  buffer buf_n330( .i (n329), .o (n330) );
  assign n331 = n322 | n330 ;
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  assign n334 = n314 & n333 ;
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  assign n340 = n97 | n101 ;
  buffer buf_n341( .i (n340), .o (n341) );
  assign n342 = ~n103 & n341 ;
  buffer buf_n343( .i (n342), .o (n343) );
  assign n344 = n314 | n333 ;
  buffer buf_n345( .i (n344), .o (n345) );
  assign n346 = ~n335 & n345 ;
  buffer buf_n347( .i (n346), .o (n347) );
  assign n348 = n343 & n347 ;
  buffer buf_n349( .i (n348), .o (n349) );
  assign n350 = n339 | n349 ;
  buffer buf_n351( .i (n350), .o (n351) );
  assign n352 = n310 & n351 ;
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  assign n358 = n113 | n117 ;
  buffer buf_n359( .i (n358), .o (n359) );
  assign n360 = ~n119 & n359 ;
  buffer buf_n361( .i (n360), .o (n361) );
  assign n362 = n310 | n351 ;
  buffer buf_n363( .i (n362), .o (n363) );
  assign n364 = ~n353 & n363 ;
  buffer buf_n365( .i (n364), .o (n365) );
  assign n366 = n361 & n365 ;
  buffer buf_n367( .i (n366), .o (n367) );
  assign n368 = n357 | n367 ;
  buffer buf_n369( .i (n368), .o (n369) );
  assign n370 = n306 & n369 ;
  buffer buf_n371( .i (n370), .o (n371) );
  assign n376 = n306 | n369 ;
  buffer buf_n377( .i (n376), .o (n377) );
  assign n378 = ~n371 & n377 ;
  buffer buf_n379( .i (n378), .o (n379) );
  assign n380 = n129 & n379 ;
  buffer buf_n381( .i (n380), .o (n381) );
  assign n382 = n129 | n379 ;
  buffer buf_n383( .i (n382), .o (n383) );
  assign n384 = ~n381 & n383 ;
  buffer buf_n385( .i (n384), .o (n385) );
  assign n386 = n361 | n365 ;
  buffer buf_n387( .i (n386), .o (n387) );
  assign n388 = ~n367 & n387 ;
  buffer buf_n389( .i (n388), .o (n389) );
  assign n390 = n343 | n347 ;
  buffer buf_n391( .i (n390), .o (n391) );
  assign n392 = ~n349 & n391 ;
  buffer buf_n393( .i (n392), .o (n393) );
  assign n394 = n324 | n328 ;
  buffer buf_n395( .i (n394), .o (n395) );
  assign n396 = ~n330 & n395 ;
  buffer buf_n397( .i (n396), .o (n397) );
  assign n398 = a_4_ & b_0_ ;
  buffer buf_n399( .i (n398), .o (n399) );
  assign n400 = b_1_ & a_3_ ;
  buffer buf_n401( .i (n400), .o (n401) );
  assign n402 = n399 & n401 ;
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  assign n408 = a_2_ & b_2_ ;
  buffer buf_n409( .i (n408), .o (n409) );
  assign n410 = n399 | n401 ;
  buffer buf_n411( .i (n410), .o (n411) );
  assign n412 = ~n403 & n411 ;
  buffer buf_n413( .i (n412), .o (n413) );
  assign n414 = n409 & n413 ;
  buffer buf_n415( .i (n414), .o (n415) );
  assign n416 = n407 | n415 ;
  buffer buf_n417( .i (n416), .o (n417) );
  assign n418 = n397 & n417 ;
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  assign n424 = b_5_ & a_0_ ;
  buffer buf_n425( .i (n424), .o (n425) );
  assign n426 = b_4_ & a_1_ ;
  buffer buf_n427( .i (n426), .o (n427) );
  assign n428 = a_2_ & b_3_ ;
  buffer buf_n429( .i (n428), .o (n429) );
  assign n430 = n427 | n429 ;
  buffer buf_n431( .i (n430), .o (n431) );
  assign n432 = n427 & n429 ;
  buffer buf_n433( .i (n432), .o (n433) );
  assign n438 = n431 & ~n433 ;
  buffer buf_n439( .i (n438), .o (n439) );
  assign n440 = n425 & n439 ;
  buffer buf_n441( .i (n440), .o (n441) );
  assign n442 = n425 | n439 ;
  buffer buf_n443( .i (n442), .o (n443) );
  assign n444 = ~n441 & n443 ;
  buffer buf_n445( .i (n444), .o (n445) );
  assign n446 = n397 | n417 ;
  buffer buf_n447( .i (n446), .o (n447) );
  assign n448 = ~n419 & n447 ;
  buffer buf_n449( .i (n448), .o (n449) );
  assign n450 = n445 & n449 ;
  buffer buf_n451( .i (n450), .o (n451) );
  assign n452 = n423 | n451 ;
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  assign n455 = n393 & n454 ;
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  assign n461 = b_6_ & a_0_ ;
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  assign n463 = n437 | n441 ;
  buffer buf_n464( .i (n463), .o (n464) );
  assign n465 = n462 & n464 ;
  buffer buf_n466( .i (n465), .o (n466) );
  assign n482 = n462 | n464 ;
  buffer buf_n483( .i (n482), .o (n483) );
  assign n484 = ~n466 & n483 ;
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  assign n491 = n393 | n454 ;
  buffer buf_n492( .i (n491), .o (n492) );
  assign n493 = ~n456 & n492 ;
  buffer buf_n494( .i (n493), .o (n494) );
  assign n495 = n490 & n494 ;
  buffer buf_n496( .i (n495), .o (n496) );
  assign n497 = n460 | n496 ;
  buffer buf_n498( .i (n497), .o (n498) );
  assign n499 = n389 & n498 ;
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  assign n505 = n389 | n498 ;
  buffer buf_n506( .i (n505), .o (n506) );
  assign n507 = ~n500 & n506 ;
  buffer buf_n508( .i (n507), .o (n508) );
  assign n509 = n481 & n508 ;
  buffer buf_n510( .i (n509), .o (n510) );
  assign n511 = n504 | n510 ;
  buffer buf_n512( .i (n511), .o (n512) );
  assign n513 = n385 | n512 ;
  buffer buf_n514( .i (n513), .o (n514) );
  assign n515 = n385 & n512 ;
  buffer buf_n516( .i (n515), .o (n516) );
  assign n525 = n514 & ~n516 ;
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  assign n531 = n481 | n508 ;
  buffer buf_n532( .i (n531), .o (n532) );
  assign n533 = ~n510 & n532 ;
  buffer buf_n534( .i (n533), .o (n534) );
  assign n535 = n490 | n494 ;
  buffer buf_n536( .i (n535), .o (n536) );
  assign n537 = ~n496 & n536 ;
  buffer buf_n538( .i (n537), .o (n538) );
  assign n539 = n445 | n449 ;
  buffer buf_n540( .i (n539), .o (n540) );
  assign n541 = ~n451 & n540 ;
  buffer buf_n542( .i (n541), .o (n542) );
  assign n543 = n409 | n413 ;
  buffer buf_n544( .i (n543), .o (n544) );
  assign n545 = ~n415 & n544 ;
  buffer buf_n546( .i (n545), .o (n546) );
  assign n547 = a_2_ & b_1_ ;
  buffer buf_n548( .i (n547), .o (n548) );
  assign n549 = b_0_ & a_3_ ;
  buffer buf_n550( .i (n549), .o (n550) );
  assign n551 = n548 & n550 ;
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  assign n557 = a_1_ & b_2_ ;
  buffer buf_n558( .i (n557), .o (n558) );
  assign n559 = n548 | n550 ;
  buffer buf_n560( .i (n559), .o (n560) );
  assign n561 = ~n552 & n560 ;
  buffer buf_n562( .i (n561), .o (n562) );
  assign n563 = n558 & n562 ;
  buffer buf_n564( .i (n563), .o (n564) );
  assign n565 = n556 | n564 ;
  buffer buf_n566( .i (n565), .o (n566) );
  assign n567 = n546 & n566 ;
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  assign n573 = a_1_ & b_3_ ;
  assign n574 = b_4_ & a_0_ ;
  assign n575 = n573 | n574 ;
  assign n576 = b_3_ & a_0_ ;
  buffer buf_n577( .i (n576), .o (n577) );
  assign n586 = n427 & n577 ;
  buffer buf_n587( .i (n586), .o (n587) );
  assign n602 = n575 & ~n587 ;
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  assign n608 = n546 | n566 ;
  buffer buf_n609( .i (n608), .o (n609) );
  assign n610 = ~n568 & n609 ;
  buffer buf_n611( .i (n610), .o (n611) );
  assign n612 = n607 & n611 ;
  buffer buf_n613( .i (n612), .o (n613) );
  assign n614 = n572 | n613 ;
  buffer buf_n615( .i (n614), .o (n615) );
  assign n616 = n542 & n615 ;
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  assign n622 = n542 | n615 ;
  buffer buf_n623( .i (n622), .o (n623) );
  assign n624 = ~n617 & n623 ;
  buffer buf_n625( .i (n624), .o (n625) );
  assign n626 = n601 & n625 ;
  buffer buf_n627( .i (n626), .o (n627) );
  assign n628 = n621 | n627 ;
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  assign n631 = n538 & n630 ;
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  assign n639 = n534 & n638 ;
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  assign n645 = n534 | n638 ;
  buffer buf_n646( .i (n645), .o (n646) );
  assign n647 = ~n640 & n646 ;
  buffer buf_n648( .i (n647), .o (n648) );
  assign n649 = n538 | n630 ;
  buffer buf_n650( .i (n649), .o (n650) );
  assign n651 = ~n632 & n650 ;
  buffer buf_n652( .i (n651), .o (n652) );
  assign n653 = n601 | n625 ;
  buffer buf_n654( .i (n653), .o (n654) );
  assign n655 = ~n627 & n654 ;
  buffer buf_n656( .i (n655), .o (n656) );
  assign n657 = n607 | n611 ;
  buffer buf_n658( .i (n657), .o (n658) );
  assign n659 = ~n613 & n658 ;
  buffer buf_n660( .i (n659), .o (n660) );
  assign n661 = a_1_ & b_1_ ;
  buffer buf_n662( .i (n661), .o (n662) );
  assign n663 = a_2_ & b_0_ ;
  buffer buf_n664( .i (n663), .o (n664) );
  assign n665 = n662 & n664 ;
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  assign n671 = b_2_ & a_0_ ;
  buffer buf_n672( .i (n671), .o (n672) );
  assign n673 = n662 | n664 ;
  buffer buf_n674( .i (n673), .o (n674) );
  assign n675 = ~n666 & n674 ;
  buffer buf_n676( .i (n675), .o (n676) );
  assign n677 = n672 & n676 ;
  buffer buf_n678( .i (n677), .o (n678) );
  assign n679 = n670 | n678 ;
  buffer buf_n680( .i (n679), .o (n680) );
  assign n681 = n558 | n562 ;
  buffer buf_n682( .i (n681), .o (n682) );
  assign n683 = ~n564 & n682 ;
  buffer buf_n684( .i (n683), .o (n684) );
  assign n685 = n680 & n684 ;
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  assign n691 = n680 | n684 ;
  buffer buf_n692( .i (n691), .o (n692) );
  assign n693 = ~n686 & n692 ;
  buffer buf_n694( .i (n693), .o (n694) );
  assign n695 = n585 & n694 ;
  buffer buf_n696( .i (n695), .o (n696) );
  assign n697 = n690 | n696 ;
  buffer buf_n698( .i (n697), .o (n698) );
  assign n699 = n660 & n698 ;
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  assign n707 = n656 & n706 ;
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  assign n712 = n652 & n711 ;
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  assign n718 = n652 | n711 ;
  buffer buf_n719( .i (n718), .o (n719) );
  assign n720 = ~n713 & n719 ;
  buffer buf_n721( .i (n720), .o (n721) );
  assign n722 = n656 | n706 ;
  buffer buf_n723( .i (n722), .o (n723) );
  assign n724 = ~n708 & n723 ;
  buffer buf_n725( .i (n724), .o (n725) );
  assign n726 = n660 | n698 ;
  buffer buf_n727( .i (n726), .o (n727) );
  assign n728 = ~n700 & n727 ;
  buffer buf_n729( .i (n728), .o (n729) );
  assign n730 = n672 | n676 ;
  buffer buf_n731( .i (n730), .o (n731) );
  assign n732 = ~n678 & n731 ;
  buffer buf_n733( .i (n732), .o (n733) );
  assign n734 = n22 & n733 ;
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  assign n742 = n585 | n694 ;
  buffer buf_n743( .i (n742), .o (n743) );
  assign n744 = ~n696 & n743 ;
  buffer buf_n745( .i (n744), .o (n745) );
  assign n746 = n741 & n745 ;
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  assign n750 = n729 & n749 ;
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  assign n758 = n725 & n757 ;
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  assign n763 = n721 & n762 ;
  buffer buf_n764( .i (n763), .o (n764) );
  assign n765 = n717 | n764 ;
  buffer buf_n766( .i (n765), .o (n766) );
  assign n767 = n648 & n766 ;
  buffer buf_n768( .i (n767), .o (n768) );
  assign n769 = n644 | n768 ;
  buffer buf_n770( .i (n769), .o (n770) );
  assign n771 = n530 & n770 ;
  buffer buf_n772( .i (n771), .o (n772) );
  assign n773 = n530 | n770 ;
  buffer buf_n774( .i (n773), .o (n774) );
  assign n775 = ~n772 & n774 ;
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  assign n799 = n741 | n745 ;
  buffer buf_n800( .i (n799), .o (n800) );
  assign n801 = ~n747 & n800 ;
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  assign n850 = n725 | n757 ;
  buffer buf_n851( .i (n850), .o (n851) );
  assign n852 = ~n759 & n851 ;
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  assign n889 = n524 | n772 ;
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  assign n891 = n375 | n381 ;
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  assign n893 = n159 | n165 ;
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  assign n903 = a_2_ & b_7_ ;
  buffer buf_n904( .i (n903), .o (n904) );
  assign n905 = b_6_ & a_3_ ;
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  assign n907 = n181 | n187 ;
  buffer buf_n908( .i (n907), .o (n908) );
  assign n909 = n906 & n908 ;
  buffer buf_n910( .i (n909), .o (n910) );
  assign n915 = n906 | n908 ;
  buffer buf_n916( .i (n915), .o (n916) );
  assign n917 = ~n910 & n916 ;
  buffer buf_n918( .i (n917), .o (n918) );
  assign n919 = n904 & n918 ;
  buffer buf_n920( .i (n919), .o (n920) );
  assign n921 = n904 | n918 ;
  buffer buf_n922( .i (n921), .o (n922) );
  assign n923 = ~n920 & n922 ;
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  assign n930 = a_4_ & b_5_ ;
  buffer buf_n931( .i (n930), .o (n931) );
  assign n932 = b_4_ & a_5_ ;
  assign n933 = a_6_ & b_3_ ;
  buffer buf_n934( .i (n933), .o (n934) );
  assign n935 = n932 | n934 ;
  buffer buf_n936( .i (n935), .o (n936) );
  assign n937 = b_4_ & a_6_ ;
  buffer buf_n938( .i (n937), .o (n938) );
  assign n939 = n175 & n938 ;
  buffer buf_n940( .i (n939), .o (n940) );
  assign n945 = n936 & ~n940 ;
  buffer buf_n946( .i (n945), .o (n946) );
  assign n947 = n931 & n946 ;
  buffer buf_n948( .i (n947), .o (n948) );
  assign n949 = n931 | n946 ;
  buffer buf_n950( .i (n949), .o (n950) );
  assign n951 = ~n948 & n950 ;
  buffer buf_n952( .i (n951), .o (n952) );
  assign n953 = ~n202 & n225 ;
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  assign n956 = n952 & n955 ;
  buffer buf_n957( .i (n956), .o (n957) );
  assign n958 = n952 | n955 ;
  buffer buf_n959( .i (n958), .o (n959) );
  assign n960 = ~n957 & n959 ;
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  assign n967 = n238 | n244 ;
  buffer buf_n968( .i (n967), .o (n968) );
  assign n969 = n966 & n968 ;
  buffer buf_n970( .i (n969), .o (n970) );
  assign n975 = n966 | n968 ;
  buffer buf_n976( .i (n975), .o (n976) );
  assign n977 = ~n970 & n976 ;
  buffer buf_n978( .i (n977), .o (n978) );
  assign n979 = n929 & n978 ;
  buffer buf_n980( .i (n979), .o (n980) );
  assign n981 = n929 | n978 ;
  buffer buf_n982( .i (n981), .o (n982) );
  assign n983 = ~n980 & n982 ;
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  assign n985 = n296 | n302 ;
  buffer buf_n986( .i (n985), .o (n986) );
  assign n987 = n984 & n986 ;
  buffer buf_n988( .i (n987), .o (n988) );
  assign n993 = n984 | n986 ;
  buffer buf_n994( .i (n993), .o (n994) );
  assign n995 = ~n988 & n994 ;
  buffer buf_n996( .i (n995), .o (n996) );
  assign n997 = n902 & n996 ;
  buffer buf_n998( .i (n997), .o (n998) );
  assign n999 = n902 | n996 ;
  buffer buf_n1000( .i (n999), .o (n1000) );
  assign n1001 = ~n998 & n1000 ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  assign n1003 = n892 & n1002 ;
  buffer buf_n1004( .i (n1003), .o (n1004) );
  assign n1015 = n892 | n1002 ;
  buffer buf_n1016( .i (n1015), .o (n1016) );
  assign n1028 = ~n1004 & n1016 ;
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  assign n1038 = n890 | n1037 ;
  assign n1039 = n890 & n1037 ;
  assign n1040 = n1038 & ~n1039 ;
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1061 = n22 | n733 ;
  buffer buf_n1062( .i (n1061), .o (n1062) );
  assign n1063 = ~n735 & n1062 ;
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  assign n1120 = n944 | n948 ;
  buffer buf_n1121( .i (n1120), .o (n1121) );
  assign n1122 = a_4_ & b_6_ ;
  buffer buf_n1123( .i (n1122), .o (n1123) );
  assign n1124 = n1121 & n1123 ;
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  assign n1130 = b_7_ & a_3_ ;
  buffer buf_n1131( .i (n1130), .o (n1131) );
  assign n1132 = n1121 | n1123 ;
  buffer buf_n1133( .i (n1132), .o (n1133) );
  assign n1134 = ~n1125 & n1133 ;
  buffer buf_n1135( .i (n1134), .o (n1135) );
  assign n1136 = n1131 & n1135 ;
  buffer buf_n1137( .i (n1136), .o (n1137) );
  assign n1138 = n1129 | n1137 ;
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  assign n1148 = a_7_ & b_5_ ;
  buffer buf_n1149( .i (n1148), .o (n1149) );
  assign n1160 = n938 & n1149 ;
  buffer buf_n1161( .i (n1160), .o (n1161) );
  assign n1162 = b_4_ & a_7_ ;
  buffer buf_n1163( .i (n1162), .o (n1163) );
  assign n1164 = a_6_ & b_5_ ;
  assign n1165 = n1163 | n1164 ;
  buffer buf_n1166( .i (n1165), .o (n1166) );
  assign n1167 = ~n1161 & n1166 ;
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  assign n1181 = b_7_ & a_4_ ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  assign n1183 = n934 & n1163 ;
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  assign n1189 = a_5_ & b_5_ ;
  buffer buf_n1190( .i (n1189), .o (n1190) );
  assign n1191 = a_7_ & b_3_ ;
  assign n1192 = n938 | n1191 ;
  buffer buf_n1193( .i (n1192), .o (n1193) );
  assign n1194 = ~n1184 & n1193 ;
  buffer buf_n1195( .i (n1194), .o (n1195) );
  assign n1196 = n1190 & n1195 ;
  buffer buf_n1197( .i (n1196), .o (n1197) );
  assign n1198 = n1188 | n1197 ;
  buffer buf_n1199( .i (n1198), .o (n1199) );
  assign n1200 = a_5_ & b_6_ ;
  buffer buf_n1201( .i (n1200), .o (n1201) );
  assign n1202 = n1199 & n1201 ;
  buffer buf_n1203( .i (n1202), .o (n1203) );
  assign n1208 = n1199 | n1201 ;
  buffer buf_n1209( .i (n1208), .o (n1209) );
  assign n1210 = ~n1203 & n1209 ;
  buffer buf_n1211( .i (n1210), .o (n1211) );
  assign n1212 = n1182 & n1211 ;
  buffer buf_n1213( .i (n1212), .o (n1213) );
  assign n1214 = n1182 | n1211 ;
  buffer buf_n1215( .i (n1214), .o (n1215) );
  assign n1216 = ~n1213 & n1215 ;
  buffer buf_n1217( .i (n1216), .o (n1217) );
  assign n1218 = n1180 & n1217 ;
  buffer buf_n1219( .i (n1218), .o (n1219) );
  assign n1220 = n1180 | n1217 ;
  buffer buf_n1221( .i (n1220), .o (n1221) );
  assign n1222 = ~n1219 & n1221 ;
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  assign n1224 = n230 | n957 ;
  buffer buf_n1225( .i (n1224), .o (n1225) );
  assign n1226 = n1190 | n1195 ;
  buffer buf_n1227( .i (n1226), .o (n1227) );
  assign n1228 = ~n1197 & n1227 ;
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  assign n1234 = n1225 & n1233 ;
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  assign n1240 = n1225 | n1233 ;
  buffer buf_n1241( .i (n1240), .o (n1241) );
  assign n1242 = ~n1235 & n1241 ;
  buffer buf_n1243( .i (n1242), .o (n1243) );
  assign n1244 = n1131 | n1135 ;
  buffer buf_n1245( .i (n1244), .o (n1245) );
  assign n1246 = ~n1137 & n1245 ;
  buffer buf_n1247( .i (n1246), .o (n1247) );
  assign n1248 = n1243 & n1247 ;
  buffer buf_n1249( .i (n1248), .o (n1249) );
  assign n1250 = n1239 | n1249 ;
  buffer buf_n1251( .i (n1250), .o (n1251) );
  assign n1252 = n1223 & n1251 ;
  buffer buf_n1253( .i (n1252), .o (n1253) );
  assign n1258 = n1223 | n1251 ;
  buffer buf_n1259( .i (n1258), .o (n1259) );
  assign n1260 = ~n1253 & n1259 ;
  buffer buf_n1261( .i (n1260), .o (n1261) );
  assign n1262 = n1147 & n1261 ;
  buffer buf_n1263( .i (n1262), .o (n1263) );
  assign n1264 = n1147 | n1261 ;
  buffer buf_n1265( .i (n1264), .o (n1265) );
  assign n1266 = ~n1263 & n1265 ;
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  assign n1273 = n974 | n980 ;
  buffer buf_n1274( .i (n1273), .o (n1274) );
  assign n1275 = n1243 | n1247 ;
  buffer buf_n1276( .i (n1275), .o (n1276) );
  assign n1277 = ~n1249 & n1276 ;
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  assign n1284 = n1274 & n1283 ;
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  assign n1290 = n914 | n920 ;
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  assign n1305 = n1274 | n1283 ;
  buffer buf_n1306( .i (n1305), .o (n1306) );
  assign n1307 = ~n1285 & n1306 ;
  buffer buf_n1308( .i (n1307), .o (n1308) );
  assign n1309 = n1304 & n1308 ;
  buffer buf_n1310( .i (n1309), .o (n1310) );
  assign n1311 = n1289 | n1310 ;
  buffer buf_n1312( .i (n1311), .o (n1312) );
  assign n1313 = n1272 & n1312 ;
  buffer buf_n1314( .i (n1313), .o (n1314) );
  assign n1334 = n1272 | n1312 ;
  buffer buf_n1335( .i (n1334), .o (n1335) );
  assign n1336 = ~n1314 & n1335 ;
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  assign n1353 = n992 | n998 ;
  buffer buf_n1354( .i (n1353), .o (n1354) );
  assign n1355 = n1304 | n1308 ;
  buffer buf_n1356( .i (n1355), .o (n1356) );
  assign n1357 = ~n1310 & n1356 ;
  buffer buf_n1358( .i (n1357), .o (n1358) );
  assign n1359 = n1354 & n1358 ;
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  assign n1376 = n890 | n1014 ;
  assign n1377 = n1027 & n1376 ;
  buffer buf_n1378( .i (n1377), .o (n1378) );
  assign n1379 = n1354 | n1358 ;
  buffer buf_n1380( .i (n1379), .o (n1380) );
  assign n1381 = ~n1360 & n1380 ;
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  assign n1394 = n1378 & n1393 ;
  buffer buf_n1395( .i (n1394), .o (n1395) );
  assign n1396 = n1375 | n1395 ;
  buffer buf_n1397( .i (n1396), .o (n1397) );
  assign n1398 = n1352 | n1397 ;
  buffer buf_n1399( .i (n1398), .o (n1399) );
  assign n1400 = n1352 & n1397 ;
  buffer buf_n1401( .i (n1400), .o (n1401) );
  assign n1402 = n1399 & ~n1401 ;
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  assign n1415 = a_6_ & b_6_ ;
  buffer buf_n1416( .i (n1415), .o (n1416) );
  assign n1417 = b_7_ & a_7_ ;
  buffer buf_n1418( .i (n1417), .o (n1418) );
  assign n1419 = n1416 & n1418 ;
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  assign n1439 = ~n1416 & n1418 ;
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  buffer buf_n1455( .i (n1454), .o (n1455) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  assign n1457 = a_7_ & b_6_ ;
  assign n1458 = b_7_ & a_6_ ;
  assign n1459 = n1457 | n1458 ;
  assign n1460 = ~n1420 & n1459 ;
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  assign n1468 = b_7_ & a_5_ ;
  buffer buf_n1469( .i (n1468), .o (n1469) );
  assign n1470 = b_6_ & n1161 ;
  buffer buf_n1471( .i (n1470), .o (n1471) );
  assign n1476 = n1161 | n1416 ;
  buffer buf_n1477( .i (n1476), .o (n1477) );
  assign n1478 = ~n1471 & n1477 ;
  buffer buf_n1479( .i (n1478), .o (n1479) );
  assign n1480 = n1469 & n1479 ;
  buffer buf_n1481( .i (n1480), .o (n1481) );
  assign n1482 = n1469 | n1479 ;
  buffer buf_n1483( .i (n1482), .o (n1483) );
  assign n1484 = ~n1481 & n1483 ;
  buffer buf_n1485( .i (n1484), .o (n1485) );
  assign n1486 = n1159 & n1485 ;
  buffer buf_n1487( .i (n1486), .o (n1487) );
  assign n1488 = n1467 & n1487 ;
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  assign n1494 = n1475 | n1481 ;
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  assign n1502 = n1467 | n1487 ;
  buffer buf_n1503( .i (n1502), .o (n1503) );
  assign n1504 = ~n1489 & n1503 ;
  buffer buf_n1505( .i (n1504), .o (n1505) );
  assign n1506 = n1501 & n1505 ;
  buffer buf_n1507( .i (n1506), .o (n1507) );
  assign n1508 = n1493 | n1507 ;
  buffer buf_n1509( .i (n1508), .o (n1509) );
  assign n1510 = n1456 & n1509 ;
  buffer buf_n1511( .i (n1510), .o (n1511) );
  assign n1512 = n1438 | n1511 ;
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n1522( .i (n1521), .o (n1522) );
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  buffer buf_n1534( .i (n1533), .o (n1534) );
  buffer buf_n1535( .i (n1534), .o (n1535) );
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  assign n1556 = n1456 | n1509 ;
  buffer buf_n1557( .i (n1556), .o (n1557) );
  assign n1558 = ~n1511 & n1557 ;
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  assign n1600 = n1501 | n1505 ;
  buffer buf_n1601( .i (n1600), .o (n1601) );
  assign n1602 = ~n1507 & n1601 ;
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  assign n1610 = n1159 | n1485 ;
  buffer buf_n1611( .i (n1610), .o (n1611) );
  assign n1612 = ~n1487 & n1611 ;
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  assign n1618 = n1219 & n1617 ;
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  assign n1624 = n1207 | n1213 ;
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  assign n1632 = n1219 | n1617 ;
  buffer buf_n1633( .i (n1632), .o (n1633) );
  assign n1634 = ~n1619 & n1633 ;
  buffer buf_n1635( .i (n1634), .o (n1635) );
  assign n1636 = n1631 & n1635 ;
  buffer buf_n1637( .i (n1636), .o (n1637) );
  assign n1638 = n1623 | n1637 ;
  buffer buf_n1639( .i (n1638), .o (n1639) );
  assign n1640 = n1609 & n1639 ;
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  buffer buf_n1658( .i (n1657), .o (n1658) );
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  assign n1676 = n1609 | n1639 ;
  buffer buf_n1677( .i (n1676), .o (n1677) );
  assign n1678 = ~n1641 & n1677 ;
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  assign n1710 = n1631 | n1635 ;
  buffer buf_n1711( .i (n1710), .o (n1711) );
  assign n1712 = ~n1637 & n1711 ;
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  assign n1716 = n1257 | n1263 ;
  buffer buf_n1717( .i (n1716), .o (n1717) );
  assign n1718 = n1715 & n1717 ;
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  assign n1748 = n1715 | n1717 ;
  buffer buf_n1749( .i (n1748), .o (n1749) );
  assign n1750 = ~n1719 & n1749 ;
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  assign n1776 = n1333 | n1401 ;
  buffer buf_n1777( .i (n1776), .o (n1777) );
  assign n1778 = n1775 & n1777 ;
  buffer buf_n1779( .i (n1778), .o (n1779) );
  assign n1780 = n1747 | n1779 ;
  buffer buf_n1781( .i (n1780), .o (n1781) );
  assign n1782 = n1709 & n1781 ;
  buffer buf_n1783( .i (n1782), .o (n1783) );
  assign n1784 = n1675 | n1783 ;
  buffer buf_n1785( .i (n1784), .o (n1785) );
  assign n1786 = n1599 & n1785 ;
  buffer buf_n1787( .i (n1786), .o (n1787) );
  assign n1788 = n1555 | n1787 ;
  assign n1789 = n729 | n749 ;
  buffer buf_n1790( .i (n1789), .o (n1790) );
  assign n1791 = ~n751 & n1790 ;
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  buffer buf_n1813( .i (n1812), .o (n1813) );
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  buffer buf_n1821( .i (n1820), .o (n1821) );
  buffer buf_n1822( .i (n1821), .o (n1822) );
  buffer buf_n1823( .i (n1822), .o (n1823) );
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1825( .i (n1824), .o (n1825) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  assign n1836 = n1378 | n1393 ;
  buffer buf_n1837( .i (n1836), .o (n1837) );
  assign n1838 = ~n1395 & n1837 ;
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  buffer buf_n1846( .i (n1845), .o (n1846) );
  buffer buf_n1847( .i (n1846), .o (n1847) );
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  assign n1855 = n1599 | n1785 ;
  buffer buf_n1856( .i (n1855), .o (n1856) );
  assign n1857 = ~n1787 & n1856 ;
  assign n1858 = n648 | n766 ;
  buffer buf_n1859( .i (n1858), .o (n1859) );
  assign n1860 = ~n768 & n1859 ;
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  buffer buf_n1872( .i (n1871), .o (n1872) );
  buffer buf_n1873( .i (n1872), .o (n1873) );
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  buffer buf_n1879( .i (n1878), .o (n1879) );
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  assign n1888 = n1709 | n1781 ;
  buffer buf_n1889( .i (n1888), .o (n1889) );
  assign n1890 = ~n1783 & n1889 ;
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  assign n1895 = n1775 | n1777 ;
  buffer buf_n1896( .i (n1895), .o (n1896) );
  assign n1897 = ~n1779 & n1896 ;
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  assign n1906 = n721 | n762 ;
  buffer buf_n1907( .i (n1906), .o (n1907) );
  assign n1908 = ~n764 & n1907 ;
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n1915( .i (n1914), .o (n1915) );
  buffer buf_n1916( .i (n1915), .o (n1916) );
  buffer buf_n1917( .i (n1916), .o (n1917) );
  buffer buf_n1918( .i (n1917), .o (n1918) );
  buffer buf_n1919( .i (n1918), .o (n1919) );
  buffer buf_n1920( .i (n1919), .o (n1920) );
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  buffer buf_n1930( .i (n1929), .o (n1930) );
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n1934( .i (n1933), .o (n1934) );
  buffer buf_n1935( .i (n1934), .o (n1935) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  assign n1940 = b_0_ & a_0_ ;
  assign s_1_ = n83 ;
  assign s_8_ = n798 ;
  assign s_3_ = n849 ;
  assign s_5_ = n888 ;
  assign s_9_ = n1060 ;
  assign s_2_ = n1119 ;
  assign s_11_ = n1414 ;
  assign s_15_ = n1788 ;
  assign s_4_ = n1835 ;
  assign s_10_ = n1854 ;
  assign s_14_ = n1857 ;
  assign s_7_ = n1887 ;
  assign s_13_ = n1894 ;
  assign s_12_ = n1905 ;
  assign s_6_ = n1939 ;
  assign s_0_ = n1940 ;
endmodule
