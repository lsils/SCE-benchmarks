module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 ;
  buffer buf_n103( .i (x4), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n57( .i (x2), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n34( .i (x1), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n126( .i (x5), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n173( .i (x7), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n196 = n139 & ~n186 ;
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  assign n200 = n50 & n198 ;
  assign n201 = ( n74 & n120 ) | ( n74 & n200 ) | ( n120 & n200 ) ;
  assign n202 = ~n121 & n201 ;
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  assign n205 = ( n43 & n66 ) | ( n43 & n135 ) | ( n66 & n135 ) ;
  buffer buf_n206( .i (n205), .o (n206) );
  assign n211 = ( ~n68 & n114 ) | ( ~n68 & n206 ) | ( n114 & n206 ) ;
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  assign n216 = ( n47 & n139 ) | ( n47 & n212 ) | ( n139 & n212 ) ;
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  assign n219 = ~n210 & n217 ;
  assign n220 = ( ~n215 & n218 ) | ( ~n215 & n219 ) | ( n218 & n219 ) ;
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n150( .i (x6), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  assign n223 = ( n168 & ~n191 ) | ( n168 & n221 ) | ( ~n191 & n221 ) ;
  assign n224 = ~n45 & n68 ;
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n140( .i (n139), .o (n140) );
  assign n231 = ~n140 & n164 ;
  buffer buf_n232( .i (n231), .o (n232) );
  assign n235 = n119 & n232 ;
  assign n236 = n229 & n235 ;
  assign n237 = n191 & n236 ;
  assign n238 = ( n222 & ~n223 ) | ( n222 & n237 ) | ( ~n223 & n237 ) ;
  buffer buf_n9( .i (x0), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  assign n239 = ~n23 & n71 ;
  assign n240 = n49 & n239 ;
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  assign n243 = n164 & ~n187 ;
  buffer buf_n244( .i (n243), .o (n244) );
  assign n250 = n142 & n244 ;
  assign n251 = ( n120 & ~n241 ) | ( n120 & n250 ) | ( ~n241 & n250 ) ;
  assign n252 = n242 & n251 ;
  buffer buf_n253( .i (n252), .o (n253) );
  assign n254 = ( ~n203 & n238 ) | ( ~n203 & n253 ) | ( n238 & n253 ) ;
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  assign n255 = n29 | n253 ;
  assign n256 = ( n204 & n254 ) | ( n204 & n255 ) | ( n254 & n255 ) ;
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n79( .i (x3), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  assign n259 = ~n102 & n257 ;
  assign n260 = n21 & n69 ;
  buffer buf_n261( .i (n260), .o (n261) );
  assign n266 = n48 & n261 ;
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  assign n274 = n137 & n184 ;
  buffer buf_n275( .i (n274), .o (n275) );
  assign n280 = ( n116 & n163 ) | ( n116 & n275 ) | ( n163 & n275 ) ;
  assign n281 = ~n117 & n280 ;
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  assign n289 = n273 & n288 ;
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  assign n290 = ( n52 & ~n75 ) | ( n52 & n144 ) | ( ~n75 & n144 ) ;
  assign n291 = ( n42 & n134 ) | ( n42 & ~n158 ) | ( n134 & ~n158 ) ;
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  assign n302 = ~n290 & n301 ;
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  assign n305 = ( n30 & n124 ) | ( n30 & ~n303 ) | ( n124 & ~n303 ) ;
  assign n306 = ( n52 & n144 ) | ( n52 & n168 ) | ( n144 & n168 ) ;
  assign n307 = n28 & ~n306 ;
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  assign n308 = n167 & n279 ;
  assign n309 = n52 & n308 ;
  assign n310 = n28 | n309 ;
  assign n311 = ~n307 & n310 ;
  assign n312 = n124 & n311 ;
  assign n313 = ( n304 & n305 ) | ( n304 & n312 ) | ( n305 & n312 ) ;
  assign n314 = n289 | n313 ;
  assign n315 = ( n258 & ~n259 ) | ( n258 & n314 ) | ( ~n259 & n314 ) ;
  buffer buf_n316( .i (n315), .o (n316) );
  assign n317 = ( ~n93 & n117 ) | ( ~n93 & n140 ) | ( n117 & n140 ) ;
  buffer buf_n318( .i (n317), .o (n318) );
  assign n319 = ( n73 & ~n142 ) | ( n73 & n318 ) | ( ~n142 & n318 ) ;
  assign n320 = ( n73 & n119 ) | ( n73 & ~n318 ) | ( n119 & ~n318 ) ;
  assign n321 = n319 & ~n320 ;
  assign n322 = n27 & ~n321 ;
  assign n323 = ~n113 & n136 ;
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  assign n329 = n95 & n328 ;
  assign n330 = n74 & n329 ;
  assign n331 = n27 | n330 ;
  assign n332 = ~n322 & n331 ;
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  assign n335 = ( ~n55 & n171 ) | ( ~n55 & n333 ) | ( n171 & n333 ) ;
  buffer buf_n76( .i (n75), .o (n76) );
  assign n336 = ~n27 & n97 ;
  assign n337 = ~n76 & n336 ;
  assign n338 = n135 & n159 ;
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  assign n348 = ~n122 & n347 ;
  assign n349 = n337 & n348 ;
  assign n350 = n55 & n349 ;
  assign n351 = ( n334 & ~n335 ) | ( n334 & n350 ) | ( ~n335 & n350 ) ;
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  assign n354 = ~n121 & n269 ;
  assign n355 = ( n98 & n347 ) | ( n98 & n354 ) | ( n347 & n354 ) ;
  assign n356 = ~n99 & n355 ;
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  assign n359 = ( ~n18 & n43 ) | ( ~n18 & n135 ) | ( n43 & n135 ) ;
  buffer buf_n360( .i (n359), .o (n360) );
  assign n365 = ( n20 & ~n161 ) | ( n20 & n360 ) | ( ~n161 & n360 ) ;
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  assign n370 = ( n47 & n139 ) | ( n47 & n366 ) | ( n139 & n366 ) ;
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  assign n373 = ~n364 & n371 ;
  assign n374 = ( ~n369 & n372 ) | ( ~n369 & n373 ) | ( n372 & n373 ) ;
  assign n375 = n74 | n374 ;
  assign n376 = n23 & ~n48 ;
  buffer buf_n377( .i (n376), .o (n377) );
  assign n381 = n232 & n377 ;
  buffer buf_n382( .i (n73), .o (n382) );
  assign n383 = ~n381 & n382 ;
  assign n384 = n375 & ~n383 ;
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  assign n387 = ( n99 & n123 ) | ( n99 & ~n385 ) | ( n123 & ~n385 ) ;
  assign n388 = ~n92 & n341 ;
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  assign n394 = ~n16 & n41 ;
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  assign n406 = n393 & n405 ;
  assign n407 = n123 & n406 ;
  assign n408 = ( n386 & n387 ) | ( n386 & n407 ) | ( n387 & n407 ) ;
  assign n409 = ( n89 & n160 ) | ( n89 & n292 ) | ( n160 & n292 ) ;
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  assign n414 = ( n46 & n138 ) | ( n46 & n410 ) | ( n138 & n410 ) ;
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  assign n417 = ~n296 & n415 ;
  assign n418 = ( ~n413 & n416 ) | ( ~n413 & n417 ) | ( n416 & n417 ) ;
  buffer buf_n419( .i (n72), .o (n419) );
  assign n420 = ~n418 & n419 ;
  assign n421 = n49 & n389 ;
  assign n422 = n419 | n421 ;
  assign n423 = ~n420 & n422 ;
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n26), .o (n426) );
  assign n427 = n191 & ~n426 ;
  assign n428 = ( n122 & n424 ) | ( n122 & ~n427 ) | ( n424 & ~n427 ) ;
  assign n429 = n425 & ~n428 ;
  buffer buf_n430( .i (n429), .o (n430) );
  assign n431 = ( ~n357 & n408 ) | ( ~n357 & n430 ) | ( n408 & n430 ) ;
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  assign n432 = n195 & ~n430 ;
  assign n433 = ( n358 & n431 ) | ( n358 & ~n432 ) | ( n431 & ~n432 ) ;
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n145( .i (n144), .o (n145) );
  assign n434 = ( ~n120 & n143 ) | ( ~n120 & n382 ) | ( n143 & n382 ) ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n436 = ( n145 & n169 ) | ( n145 & ~n435 ) | ( n169 & ~n435 ) ;
  assign n437 = ( ~n76 & n169 ) | ( ~n76 & n435 ) | ( n169 & n435 ) ;
  assign n438 = n436 & ~n437 ;
  assign n439 = n29 & ~n99 ;
  assign n440 = ( n55 & n438 ) | ( n55 & n439 ) | ( n438 & n439 ) ;
  assign n441 = ~n56 & n440 ;
  assign n442 = ( n119 & n142 ) | ( n119 & ~n419 ) | ( n142 & ~n419 ) ;
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n51), .o (n444) );
  assign n445 = ( ~n144 & n443 ) | ( ~n144 & n444 ) | ( n443 & n444 ) ;
  assign n446 = ( n121 & ~n443 ) | ( n121 & n444 ) | ( ~n443 & n444 ) ;
  assign n447 = n445 & ~n446 ;
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  assign n450 = ~n30 & n448 ;
  assign n451 = n28 & ~n122 ;
  assign n452 = n51 & n143 ;
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n426), .o (n455) );
  buffer buf_n456( .i (n118), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  assign n460 = ( n453 & ~n455 ) | ( n453 & n459 ) | ( ~n455 & n459 ) ;
  assign n461 = ( n451 & ~n454 ) | ( n451 & n460 ) | ( ~n454 & n460 ) ;
  assign n462 = ( n115 & ~n138 ) | ( n115 & n162 ) | ( ~n138 & n162 ) ;
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  assign n467 = n117 & ~n463 ;
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  assign n470 = ( n166 & n419 ) | ( n166 & n468 ) | ( n419 & n468 ) ;
  assign n471 = ( ~n466 & n469 ) | ( ~n466 & n470 ) | ( n469 & n470 ) ;
  assign n472 = n444 & n471 ;
  assign n473 = n455 | n472 ;
  buffer buf_n230( .i (n229), .o (n230) );
  assign n474 = n114 & ~n137 ;
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  assign n480 = ~n167 & n479 ;
  assign n481 = n230 & n480 ;
  assign n482 = n455 & ~n481 ;
  assign n483 = n473 & ~n482 ;
  assign n484 = n461 | n483 ;
  assign n485 = ( n449 & ~n450 ) | ( n449 & n484 ) | ( ~n450 & n484 ) ;
  assign n486 = n441 | n485 ;
  assign n487 = ( ~n352 & n433 ) | ( ~n352 & n486 ) | ( n433 & n486 ) ;
  assign n488 = n353 | n487 ;
  assign n489 = ( n65 & ~n111 ) | ( n65 & n181 ) | ( ~n111 & n181 ) ;
  assign n490 = ( ~n88 & n182 ) | ( ~n88 & n489 ) | ( n182 & n489 ) ;
  buffer buf_n491( .i (n490), .o (n491) );
  assign n494 = n184 & ~n491 ;
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  assign n497 = n493 | n495 ;
  assign n498 = ( ~n187 & n496 ) | ( ~n187 & n497 ) | ( n496 & n497 ) ;
  assign n499 = ( ~n24 & n141 ) | ( ~n24 & n498 ) | ( n141 & n498 ) ;
  assign n500 = n70 & n116 ;
  assign n501 = n92 | n186 ;
  assign n502 = ( n71 & ~n500 ) | ( n71 & n501 ) | ( ~n500 & n501 ) ;
  assign n503 = ( n24 & n141 ) | ( n24 & ~n502 ) | ( n141 & ~n502 ) ;
  assign n504 = n499 & n503 ;
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  assign n508 = ( n71 & ~n140 ) | ( n71 & n187 ) | ( ~n140 & n187 ) ;
  buffer buf_n509( .i (n508), .o (n509) );
  assign n512 = ( ~n189 & n456 ) | ( ~n189 & n509 ) | ( n456 & n509 ) ;
  buffer buf_n513( .i (n72), .o (n513) );
  assign n514 = ( n456 & ~n509 ) | ( n456 & n513 ) | ( ~n509 & n513 ) ;
  assign n515 = n512 & ~n514 ;
  assign n516 = ( ~n426 & n505 ) | ( ~n426 & n515 ) | ( n505 & n515 ) ;
  assign n517 = n98 & ~n516 ;
  buffer buf_n518( .i (n98), .o (n518) );
  assign n519 = ( n507 & ~n517 ) | ( n507 & n518 ) | ( ~n517 & n518 ) ;
  buffer buf_n520( .i (n54), .o (n520) );
  assign n521 = ( ~n171 & n519 ) | ( ~n171 & n520 ) | ( n519 & n520 ) ;
  assign n522 = n69 & ~n91 ;
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n528( .i (n116), .o (n528) );
  assign n529 = n523 & ~n528 ;
  assign n530 = ( n24 & n197 ) | ( n24 & n529 ) | ( n197 & n529 ) ;
  assign n531 = ~n25 & n530 ;
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n70), .o (n535) );
  buffer buf_n536( .i (n186), .o (n536) );
  assign n537 = ( n528 & n535 ) | ( n528 & ~n536 ) | ( n535 & ~n536 ) ;
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n141), .o (n539) );
  assign n540 = ( ~n513 & n538 ) | ( ~n513 & n539 ) | ( n538 & n539 ) ;
  assign n541 = ( n189 & n538 ) | ( n189 & ~n539 ) | ( n538 & ~n539 ) ;
  assign n542 = n540 & n541 ;
  assign n543 = ( n426 & n532 ) | ( n426 & n542 ) | ( n532 & n542 ) ;
  buffer buf_n544( .i (n97), .o (n544) );
  assign n545 = ~n543 & n544 ;
  assign n546 = ( n518 & n534 ) | ( n518 & ~n545 ) | ( n534 & ~n545 ) ;
  assign n547 = ( n171 & n520 ) | ( n171 & n546 ) | ( n520 & n546 ) ;
  assign n548 = n521 & n547 ;
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  assign n551 = n380 & n544 ;
  assign n552 = n77 & n551 ;
  assign n553 = n249 & n552 ;
  assign n554 = ( n125 & n148 ) | ( n125 & n553 ) | ( n148 & n553 ) ;
  assign n555 = ~n149 & n554 ;
  assign n556 = ( n47 & n70 ) | ( n47 & ~n163 ) | ( n70 & ~n163 ) ;
  buffer buf_n557( .i (n556), .o (n557) );
  assign n558 = ( n72 & n118 ) | ( n72 & ~n557 ) | ( n118 & ~n557 ) ;
  assign n559 = ( ~n49 & n118 ) | ( ~n49 & n557 ) | ( n118 & n557 ) ;
  assign n560 = n558 & ~n559 ;
  assign n561 = n26 | n560 ;
  assign n562 = ~n68 & n114 ;
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  assign n566 = ~n165 & n565 ;
  assign n567 = ~n50 & n566 ;
  assign n568 = n26 & ~n567 ;
  assign n569 = n561 & ~n568 ;
  assign n570 = ( n145 & n192 ) | ( n145 & n569 ) | ( n192 & n569 ) ;
  buffer buf_n571( .i (n570), .o (n571) );
  assign n572 = ( n100 & ~n147 ) | ( n100 & n571 ) | ( ~n147 & n571 ) ;
  assign n573 = ( n100 & n194 ) | ( n100 & ~n571 ) | ( n194 & ~n571 ) ;
  assign n574 = n572 & ~n573 ;
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n575( .i (n138), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  assign n577 = ( n48 & n528 ) | ( n48 & ~n576 ) | ( n528 & ~n576 ) ;
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  assign n581 = ( n50 & n456 ) | ( n50 & ~n578 ) | ( n456 & ~n578 ) ;
  assign n582 = ( n167 & n457 ) | ( n167 & n581 ) | ( n457 & n581 ) ;
  assign n583 = ( n346 & n580 ) | ( n346 & ~n582 ) | ( n580 & ~n582 ) ;
  assign n584 = n455 & n583 ;
  buffer buf_n585( .i (n46), .o (n585) );
  buffer buf_n586( .i (n115), .o (n586) );
  assign n587 = ( n163 & n585 ) | ( n163 & ~n586 ) | ( n585 & ~n586 ) ;
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n113), .o (n592) );
  assign n593 = ( n137 & n161 ) | ( n137 & ~n592 ) | ( n161 & ~n592 ) ;
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  assign n597 = n588 & n596 ;
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  assign n600 = n143 & ~n598 ;
  assign n601 = ( n591 & ~n599 ) | ( n591 & n600 ) | ( ~n599 & n600 ) ;
  buffer buf_n602( .i (n25), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  assign n605 = n601 | n604 ;
  assign n606 = ( ~n29 & n584 ) | ( ~n29 & n605 ) | ( n584 & n605 ) ;
  buffer buf_n607( .i (n136), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  assign n609 = ( n46 & n91 ) | ( n46 & n608 ) | ( n91 & n608 ) ;
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  assign n612 = ( n16 & n110 ) | ( n16 & n157 ) | ( n110 & n157 ) ;
  assign n613 = ( ~n65 & n158 ) | ( ~n65 & n612 ) | ( n158 & n612 ) ;
  buffer buf_n614( .i (n613), .o (n614) );
  assign n617 = n160 & ~n614 ;
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  assign n620 = n616 | n618 ;
  buffer buf_n621( .i (n162), .o (n621) );
  assign n622 = ( n619 & n620 ) | ( n619 & ~n621 ) | ( n620 & ~n621 ) ;
  assign n623 = n92 | n585 ;
  assign n624 = ( n576 & n622 ) | ( n576 & n623 ) | ( n622 & n623 ) ;
  assign n625 = ~n611 & n624 ;
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  assign n629 = ( n86 & n133 ) | ( n86 & n157 ) | ( n133 & n157 ) ;
  buffer buf_n630( .i (n629), .o (n630) );
  assign n639 = ( ~n112 & n159 ) | ( ~n112 & n630 ) | ( n159 & n630 ) ;
  buffer buf_n640( .i (n639), .o (n640) );
  assign n643 = n161 & ~n640 ;
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  assign n646 = n642 | n644 ;
  assign n647 = ( ~n164 & n645 ) | ( ~n164 & n646 ) | ( n645 & n646 ) ;
  buffer buf_n648( .i (n585), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  assign n650 = n647 | n649 ;
  assign n651 = ~n162 & n324 ;
  buffer buf_n652( .i (n651), .o (n652) );
  assign n654 = ~n93 & n652 ;
  assign n655 = n649 & ~n654 ;
  assign n656 = n650 & ~n655 ;
  assign n657 = ( n602 & n626 ) | ( n602 & n656 ) | ( n626 & n656 ) ;
  assign n658 = n75 & ~n657 ;
  assign n659 = ( n76 & n628 ) | ( n76 & ~n658 ) | ( n628 & ~n658 ) ;
  buffer buf_n660( .i (n659), .o (n660) );
  assign n661 = ( n78 & n606 ) | ( n78 & n660 ) | ( n606 & n660 ) ;
  buffer buf_n662( .i (n539), .o (n662) );
  assign n663 = ~n51 & n662 ;
  buffer buf_n664( .i (n649), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  assign n666 = ( ~n457 & n662 ) | ( ~n457 & n665 ) | ( n662 & n665 ) ;
  assign n667 = ( n345 & ~n457 ) | ( n345 & n662 ) | ( ~n457 & n662 ) ;
  assign n668 = ( n663 & n666 ) | ( n663 & ~n667 ) | ( n666 & ~n667 ) ;
  buffer buf_n669( .i (n45), .o (n669) );
  buffer buf_n670( .i (n160), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  assign n672 = n669 & ~n671 ;
  assign n673 = ~n41 & n110 ;
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  assign n679 = n115 & ~n671 ;
  assign n680 = ( n672 & n678 ) | ( n672 & ~n679 ) | ( n678 & ~n679 ) ;
  assign n681 = ( n23 & n576 ) | ( n23 & ~n680 ) | ( n576 & ~n680 ) ;
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  assign n684 = n25 & ~n682 ;
  assign n685 = ( n662 & ~n683 ) | ( n662 & n684 ) | ( ~n683 & n684 ) ;
  buffer buf_n686( .i (n685), .o (n686) );
  assign n687 = ( ~n604 & n668 ) | ( ~n604 & n686 ) | ( n668 & n686 ) ;
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  assign n688 = ~n528 & n648 ;
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n539), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  assign n694 = ( n234 & n691 ) | ( n234 & n693 ) | ( n691 & n693 ) ;
  assign n695 = ( n604 & n686 ) | ( n604 & n694 ) | ( n686 & n694 ) ;
  assign n696 = n687 | n695 ;
  assign n697 = ( ~n78 & n660 ) | ( ~n78 & n696 ) | ( n660 & n696 ) ;
  assign n698 = n661 | n697 ;
  assign n699 = n574 | n698 ;
  assign n700 = ( ~n549 & n555 ) | ( ~n549 & n699 ) | ( n555 & n699 ) ;
  assign n701 = n550 | n700 ;
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n172( .i (n171), .o (n172) );
  assign n702 = ( n69 & n91 ) | ( n69 & n185 ) | ( n91 & n185 ) ;
  buffer buf_n703( .i (n90), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  assign n705 = ( ~n575 & n702 ) | ( ~n575 & n704 ) | ( n702 & n704 ) ;
  buffer buf_n706( .i (n705), .o (n706) );
  assign n709 = n94 & ~n706 ;
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  assign n712 = n708 | n710 ;
  assign n713 = ( ~n97 & n711 ) | ( ~n97 & n712 ) | ( n711 & n712 ) ;
  assign n714 = ( ~n53 & n459 ) | ( ~n53 & n713 ) | ( n459 & n713 ) ;
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  assign n715 = ( n96 & n382 ) | ( n96 & ~n692 ) | ( n382 & ~n692 ) ;
  assign n716 = n511 & ~n715 ;
  assign n717 = ( n53 & n459 ) | ( n53 & n716 ) | ( n459 & n716 ) ;
  assign n718 = n714 & n717 ;
  assign n719 = n77 | n193 ;
  buffer buf_n720( .i (n586), .o (n720) );
  assign n721 = ( n93 & n610 ) | ( n93 & ~n720 ) | ( n610 & ~n720 ) ;
  buffer buf_n722( .i (n721), .o (n722) );
  assign n725 = n95 & ~n722 ;
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  assign n728 = n724 | n726 ;
  assign n729 = ( ~n544 & n727 ) | ( ~n544 & n728 ) | ( n727 & n728 ) ;
  assign n730 = ( n77 & n193 ) | ( n77 & ~n729 ) | ( n193 & ~n729 ) ;
  assign n731 = ( n718 & n719 ) | ( n718 & ~n730 ) | ( n719 & ~n730 ) ;
  assign n732 = n172 & ~n731 ;
  buffer buf_n733( .i (n185), .o (n733) );
  assign n734 = ( n575 & n704 ) | ( n575 & ~n733 ) | ( n704 & ~n733 ) ;
  assign n735 = ( n576 & ~n648 ) | ( n576 & n734 ) | ( ~n648 & n734 ) ;
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  assign n739 = ( ~n95 & n664 ) | ( ~n95 & n736 ) | ( n664 & n736 ) ;
  assign n740 = n190 | n739 ;
  assign n741 = ( ~n693 & n738 ) | ( ~n693 & n740 ) | ( n738 & n740 ) ;
  buffer buf_n742( .i (n75), .o (n742) );
  assign n743 = n741 & ~n742 ;
  buffer buf_n199( .i (n198), .o (n199) );
  assign n744 = n96 & n199 ;
  assign n745 = n444 & n744 ;
  assign n746 = n742 & ~n745 ;
  assign n747 = n743 | n746 ;
  assign n748 = n124 & ~n747 ;
  assign n749 = n172 | n748 ;
  assign n750 = ~n732 & n749 ;
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n751( .i (n22), .o (n751) );
  buffer buf_n752( .i (n575), .o (n752) );
  assign n753 = ( ~n635 & n751 ) | ( ~n635 & n752 ) | ( n751 & n752 ) ;
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n757( .i (n752), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  assign n759 = ( n166 & n754 ) | ( n166 & ~n758 ) | ( n754 & ~n758 ) ;
  assign n760 = n638 | n759 ;
  assign n761 = ( ~n603 & n756 ) | ( ~n603 & n760 ) | ( n756 & n760 ) ;
  assign n762 = n742 & n761 ;
  buffer buf_n763( .i (n94), .o (n763) );
  assign n764 = ~n166 & n763 ;
  assign n765 = n692 & n764 ;
  assign n766 = n603 & n765 ;
  assign n767 = n742 | n766 ;
  assign n768 = ~n762 & n767 ;
  assign n769 = ( n43 & n66 ) | ( n43 & n159 ) | ( n66 & n159 ) ;
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n67), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  assign n775 = n608 & ~n774 ;
  assign n776 = n670 & n770 ;
  assign n777 = ( n608 & n669 ) | ( n608 & n776 ) | ( n669 & n776 ) ;
  assign n778 = ( n772 & n775 ) | ( n772 & ~n777 ) | ( n775 & ~n777 ) ;
  assign n779 = n720 | n778 ;
  assign n780 = n225 & n341 ;
  assign n781 = n720 & ~n780 ;
  assign n782 = n779 & ~n781 ;
  assign n783 = n763 & n782 ;
  buffer buf_n784( .i (n158), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  assign n786 = n67 | n785 ;
  buffer buf_n787( .i (n786), .o (n787) );
  assign n788 = ( n608 & ~n774 ) | ( n608 & n787 ) | ( ~n774 & n787 ) ;
  buffer buf_n789( .i (n592), .o (n789) );
  buffer buf_n790( .i (n607), .o (n790) );
  assign n791 = ( n787 & ~n789 ) | ( n787 & n790 ) | ( ~n789 & n790 ) ;
  assign n792 = ( n563 & ~n788 ) | ( n563 & n791 ) | ( ~n788 & n791 ) ;
  assign n793 = n648 & n792 ;
  assign n794 = ( n671 & n774 ) | ( n671 & n789 ) | ( n774 & n789 ) ;
  assign n795 = ( n592 & n607 ) | ( n592 & n670 ) | ( n607 & n670 ) ;
  assign n796 = n774 | n795 ;
  assign n797 = ~n794 & n796 ;
  buffer buf_n798( .i (n585), .o (n798) );
  assign n799 = n797 | n798 ;
  assign n800 = ( ~n649 & n793 ) | ( ~n649 & n799 ) | ( n793 & n799 ) ;
  assign n801 = n763 | n800 ;
  assign n802 = ( ~n96 & n783 ) | ( ~n96 & n801 ) | ( n783 & n801 ) ;
  assign n803 = n603 & n802 ;
  assign n804 = ( n86 & ~n110 ) | ( n86 & n157 ) | ( ~n110 & n157 ) ;
  assign n805 = ( n87 & ~n134 ) | ( n87 & n804 ) | ( ~n134 & n804 ) ;
  buffer buf_n806( .i (n805), .o (n806) );
  assign n809 = n89 & ~n806 ;
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  assign n812 = n808 | n810 ;
  assign n813 = ( ~n704 & n811 ) | ( ~n704 & n812 ) | ( n811 & n812 ) ;
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n798), .o (n816) );
  buffer buf_n817( .i (n535), .o (n817) );
  assign n818 = ( ~n814 & n816 ) | ( ~n814 & n817 ) | ( n816 & n817 ) ;
  assign n819 = n340 & n789 ;
  buffer buf_n820( .i (n669), .o (n820) );
  assign n821 = ( n704 & n819 ) | ( n704 & n820 ) | ( n819 & n820 ) ;
  assign n822 = ~n798 & n821 ;
  assign n823 = n817 & n822 ;
  assign n824 = ( n815 & n818 ) | ( n815 & n823 ) | ( n818 & n823 ) ;
  assign n825 = n586 | n594 ;
  buffer buf_n826( .i (n621), .o (n826) );
  assign n827 = ( n595 & n825 ) | ( n595 & ~n826 ) | ( n825 & ~n826 ) ;
  assign n828 = n45 & n773 ;
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n832( .i (n773), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  assign n834 = ~n829 & n833 ;
  buffer buf_n835( .i (n834), .o (n835) );
  assign n836 = ~n827 & n835 ;
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  assign n837 = ( n653 & ~n831 ) | ( n653 & n835 ) | ( ~n831 & n835 ) ;
  assign n838 = ( n664 & n836 ) | ( n664 & n837 ) | ( n836 & n837 ) ;
  assign n839 = n824 | n838 ;
  buffer buf_n840( .i (n602), .o (n840) );
  assign n841 = n839 & ~n840 ;
  assign n842 = n803 | n841 ;
  buffer buf_n843( .i (n842), .o (n843) );
  assign n844 = ( n520 & n768 ) | ( n520 & n843 ) | ( n768 & n843 ) ;
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n845( .i (n165), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  assign n847 = ( ~n382 & n526 ) | ( ~n382 & n846 ) | ( n526 & n846 ) ;
  assign n848 = ( n526 & n602 ) | ( n526 & n846 ) | ( n602 & n846 ) ;
  assign n849 = ( n265 & n847 ) | ( n265 & ~n848 ) | ( n847 & ~n848 ) ;
  assign n850 = n145 | n849 ;
  assign n851 = ~n763 & n845 ;
  buffer buf_n852( .i (n513), .o (n852) );
  assign n853 = ( n846 & n851 ) | ( n846 & ~n852 ) | ( n851 & ~n852 ) ;
  assign n854 = ~n840 & n853 ;
  buffer buf_n855( .i (n693), .o (n855) );
  assign n856 = ~n854 & n855 ;
  assign n857 = n850 & ~n856 ;
  assign n858 = ( ~n520 & n843 ) | ( ~n520 & n857 ) | ( n843 & n857 ) ;
  assign n859 = n844 | n858 ;
  buffer buf_n860( .i (n859), .o (n860) );
  assign n861 = ( n33 & n750 ) | ( n33 & n860 ) | ( n750 & n860 ) ;
  buffer buf_n862( .i (n703), .o (n862) );
  assign n863 = ( n733 & ~n833 ) | ( n733 & n862 ) | ( ~n833 & n862 ) ;
  assign n864 = ( n535 & n752 ) | ( n535 & ~n863 ) | ( n752 & ~n863 ) ;
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  assign n868 = ( n189 & ~n758 ) | ( n189 & n865 ) | ( ~n758 & n865 ) ;
  buffer buf_n869( .i (n94), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  assign n871 = n868 & n870 ;
  buffer buf_n872( .i (n852), .o (n872) );
  assign n873 = ( n867 & n871 ) | ( n867 & ~n872 ) | ( n871 & ~n872 ) ;
  assign n874 = ( n165 & n197 ) | ( n165 & n524 ) | ( n197 & n524 ) ;
  assign n875 = ~n845 & n874 ;
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  assign n878 = n168 | n876 ;
  assign n879 = ( n873 & n877 ) | ( n873 & n878 ) | ( n877 & n878 ) ;
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n54), .o (n882) );
  buffer buf_n883( .i (n123), .o (n883) );
  assign n884 = ( n880 & ~n882 ) | ( n880 & n883 ) | ( ~n882 & n883 ) ;
  buffer buf_n527( .i (n526), .o (n527) );
  assign n885 = n527 & ~n693 ;
  assign n886 = ( n53 & n247 ) | ( n53 & n885 ) | ( n247 & n885 ) ;
  assign n887 = ~n54 & n886 ;
  assign n888 = ~n883 & n887 ;
  assign n889 = ( n881 & ~n884 ) | ( n881 & n888 ) | ( ~n884 & n888 ) ;
  assign n890 = n172 | n195 ;
  assign n891 = n513 & n869 ;
  buffer buf_n892( .i (n720), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  assign n895 = ( ~n665 & n891 ) | ( ~n665 & n894 ) | ( n891 & n894 ) ;
  buffer buf_n896( .i (n895), .o (n896) );
  assign n897 = n459 | n896 ;
  buffer buf_n898( .i (n458), .o (n898) );
  assign n899 = n896 & n898 ;
  assign n900 = n897 & ~n899 ;
  assign n901 = n664 & ~n758 ;
  assign n902 = ( n852 & n894 ) | ( n852 & n901 ) | ( n894 & n901 ) ;
  assign n903 = ~n872 & n902 ;
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  assign n906 = n146 | n904 ;
  assign n907 = ( n900 & n905 ) | ( n900 & n906 ) | ( n905 & n906 ) ;
  assign n908 = ( n172 & n195 ) | ( n172 & ~n907 ) | ( n195 & ~n907 ) ;
  assign n909 = ( n889 & n890 ) | ( n889 & ~n908 ) | ( n890 & ~n908 ) ;
  assign n910 = ( ~n33 & n860 ) | ( ~n33 & n909 ) | ( n860 & n909 ) ;
  assign n911 = n861 | n910 ;
  assign n912 = ( n44 & ~n113 ) | ( n44 & n183 ) | ( ~n113 & n183 ) ;
  buffer buf_n913( .i (n912), .o (n913) );
  assign n917 = ( n789 & n832 ) | ( n789 & n913 ) | ( n832 & n913 ) ;
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n921( .i (n586), .o (n921) );
  assign n922 = ( n536 & ~n918 ) | ( n536 & n921 ) | ( ~n918 & n921 ) ;
  assign n923 = n916 & n922 ;
  buffer buf_n924( .i (n817), .o (n924) );
  assign n925 = ( ~n920 & n923 ) | ( ~n920 & n924 ) | ( n923 & n924 ) ;
  assign n926 = n870 & ~n925 ;
  assign n927 = n188 & n892 ;
  assign n928 = n228 & n927 ;
  assign n929 = n870 | n928 ;
  assign n930 = ~n926 & n929 ;
  assign n931 = ( n604 & n855 ) | ( n604 & ~n930 ) | ( n855 & ~n930 ) ;
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  assign n934 = n30 & ~n932 ;
  assign n935 = ( n148 & ~n933 ) | ( n148 & n934 ) | ( ~n933 & n934 ) ;
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  assign n938 = ( ~n61 & n130 ) | ( ~n61 & n177 ) | ( n130 & n177 ) ;
  buffer buf_n939( .i (n938), .o (n939) );
  assign n951 = ( n40 & n179 ) | ( n40 & ~n939 ) | ( n179 & ~n939 ) ;
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  assign n956 = ( n65 & ~n134 ) | ( n65 & n952 ) | ( ~n134 & n952 ) ;
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  assign n959 = n943 & n957 ;
  assign n960 = ( ~n955 & n958 ) | ( ~n955 & n959 ) | ( n958 & n959 ) ;
  buffer buf_n961( .i (n592), .o (n961) );
  assign n962 = n960 & ~n961 ;
  assign n963 = ~n22 & n962 ;
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  assign n966 = n475 & ~n733 ;
  buffer buf_n967( .i (n966), .o (n967) );
  assign n971 = n964 | n967 ;
  assign n972 = ( n267 & n965 ) | ( n267 & n971 ) | ( n965 & n971 ) ;
  assign n973 = ( n846 & n870 ) | ( n846 & ~n972 ) | ( n870 & ~n972 ) ;
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  assign n976 = n544 & ~n974 ;
  assign n977 = ( n170 & ~n975 ) | ( n170 & n976 ) | ( ~n975 & n976 ) ;
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  assign n980 = n41 & ~n64 ;
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n990( .i (n64), .o (n990) );
  assign n991 = n17 & ~n990 ;
  assign n992 = ( n395 & ~n981 ) | ( n395 & n991 ) | ( ~n981 & n991 ) ;
  assign n993 = ( n136 & n183 ) | ( n136 & n992 ) | ( n183 & n992 ) ;
  buffer buf_n994( .i (n993), .o (n994) );
  assign n995 = ( ~n185 & n671 ) | ( ~n185 & n994 ) | ( n671 & n994 ) ;
  buffer buf_n996( .i (n670), .o (n996) );
  assign n997 = ( n790 & ~n994 ) | ( n790 & n996 ) | ( ~n994 & n996 ) ;
  assign n998 = n995 & ~n997 ;
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n785), .o (n1002) );
  assign n1003 = ( n184 & n773 ) | ( n184 & ~n1002 ) | ( n773 & ~n1002 ) ;
  buffer buf_n1004( .i (n1003), .o (n1004) );
  assign n1005 = ( ~n733 & n820 ) | ( ~n733 & n1004 ) | ( n820 & n1004 ) ;
  assign n1006 = ( n820 & n833 ) | ( n820 & ~n1004 ) | ( n833 & ~n1004 ) ;
  assign n1007 = n1005 & ~n1006 ;
  buffer buf_n1008( .i (n751), .o (n1008) );
  assign n1009 = ( n999 & n1007 ) | ( n999 & n1008 ) | ( n1007 & n1008 ) ;
  assign n1010 = n758 & ~n1009 ;
  assign n1011 = ( n692 & n1001 ) | ( n692 & ~n1010 ) | ( n1001 & ~n1010 ) ;
  assign n1012 = n458 | n1011 ;
  assign n1013 = ~n44 & n183 ;
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n790), .o (n1016) );
  assign n1017 = ( n621 & n1015 ) | ( n621 & ~n1016 ) | ( n1015 & ~n1016 ) ;
  buffer buf_n1018( .i (n182), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  assign n1021 = ( n996 & ~n1014 ) | ( n996 & n1020 ) | ( ~n1014 & n1020 ) ;
  assign n1022 = ( n820 & n1016 ) | ( n820 & ~n1021 ) | ( n1016 & ~n1021 ) ;
  assign n1023 = n1017 | n1022 ;
  assign n1024 = n817 & n1023 ;
  buffer buf_n1025( .i (n133), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  assign n1028 = ( n785 & n1018 ) | ( n785 & n1027 ) | ( n1018 & n1027 ) ;
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  assign n1031 = n790 & ~n1029 ;
  buffer buf_n1032( .i (n1020), .o (n1032) );
  assign n1033 = ( ~n1030 & n1031 ) | ( ~n1030 & n1032 ) | ( n1031 & n1032 ) ;
  assign n1034 = n798 & n1033 ;
  buffer buf_n1035( .i (n535), .o (n1035) );
  assign n1036 = n1034 | n1035 ;
  assign n1037 = ~n1024 & n1036 ;
  buffer buf_n1038( .i (n1008), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  assign n1040 = n1037 & n1039 ;
  assign n1041 = n458 & ~n1040 ;
  assign n1042 = n1012 & ~n1041 ;
  assign n1043 = n518 | n1042 ;
  assign n1044 = ( n182 & ~n674 ) | ( n182 & n1026 ) | ( ~n674 & n1026 ) ;
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1049( .i (n112), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  assign n1051 = n1045 & n1050 ;
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  assign n1055 = ( n678 & ~n1016 ) | ( n678 & n1052 ) | ( ~n1016 & n1052 ) ;
  buffer buf_n1056( .i (n669), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  assign n1058 = ( n1048 & n1055 ) | ( n1048 & ~n1057 ) | ( n1055 & ~n1057 ) ;
  assign n1059 = ( ~n188 & n1054 ) | ( ~n188 & n1058 ) | ( n1054 & n1058 ) ;
  assign n1060 = n924 | n1059 ;
  assign n1061 = ( n607 & n1019 ) | ( n607 & n1050 ) | ( n1019 & n1050 ) ;
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n961), .o (n1064) );
  assign n1065 = ~n1062 & n1064 ;
  assign n1066 = ( n752 & ~n1063 ) | ( n752 & n1065 ) | ( ~n1063 & n1065 ) ;
  assign n1067 = ~n816 & n1066 ;
  assign n1068 = n924 & ~n1067 ;
  assign n1069 = n1060 & ~n1068 ;
  assign n1070 = n1018 | n1027 ;
  assign n1071 = n1002 | n1070 ;
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  assign n1074 = n1056 & n1064 ;
  buffer buf_n1075( .i (n833), .o (n1075) );
  assign n1076 = ( ~n1073 & n1074 ) | ( ~n1073 & n1075 ) | ( n1074 & n1075 ) ;
  assign n1077 = ~n1035 & n1076 ;
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n845), .o (n1080) );
  assign n1081 = n1078 | n1080 ;
  assign n1082 = ( n1069 & n1079 ) | ( n1069 & n1081 ) | ( n1079 & n1081 ) ;
  buffer buf_n1083( .i (n840), .o (n1083) );
  assign n1084 = n1082 & n1083 ;
  assign n1085 = n518 & ~n1084 ;
  assign n1086 = n1043 & ~n1085 ;
  buffer buf_n1087( .i (n832), .o (n1087) );
  assign n1088 = ( n862 & n1016 ) | ( n862 & ~n1087 ) | ( n1016 & ~n1087 ) ;
  assign n1089 = ( n621 & ~n862 ) | ( n621 & n1087 ) | ( ~n862 & n1087 ) ;
  assign n1090 = n1088 & n1089 ;
  assign n1091 = n816 & ~n1090 ;
  buffer buf_n1092( .i (n1027), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  assign n1094 = n703 & ~n1093 ;
  buffer buf_n1095( .i (n996), .o (n1095) );
  assign n1096 = n1094 & ~n1095 ;
  assign n1097 = ~n1075 & n1096 ;
  assign n1098 = n816 | n1097 ;
  assign n1099 = ~n1091 & n1098 ;
  assign n1100 = ( n190 & ~n1039 ) | ( n190 & n1099 ) | ( ~n1039 & n1099 ) ;
  buffer buf_n1101( .i (n1100), .o (n1101) );
  assign n1102 = ( ~n192 & n898 ) | ( ~n192 & n1101 ) | ( n898 & n1101 ) ;
  assign n1103 = ( ~n898 & n1083 ) | ( ~n898 & n1101 ) | ( n1083 & n1101 ) ;
  assign n1104 = n1102 & n1103 ;
  assign n1105 = n1064 & ~n1072 ;
  buffer buf_n1106( .i (n862), .o (n1106) );
  assign n1107 = ( n751 & n1105 ) | ( n751 & n1106 ) | ( n1105 & n1106 ) ;
  assign n1108 = ~n1008 & n1107 ;
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  assign n1112 = ( n18 & ~n88 ) | ( n18 & n784 ) | ( ~n88 & n784 ) ;
  buffer buf_n1113( .i (n1112), .o (n1113) );
  assign n1118 = ( n20 & n1092 ) | ( n20 & ~n1113 ) | ( n1092 & ~n1113 ) ;
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n703), .o (n1123) );
  assign n1124 = ( ~n1095 & n1119 ) | ( ~n1095 & n1123 ) | ( n1119 & n1123 ) ;
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  assign n1127 = n1117 & n1125 ;
  assign n1128 = ( ~n1122 & n1126 ) | ( ~n1122 & n1127 ) | ( n1126 & n1127 ) ;
  assign n1129 = ( ~n894 & n1109 ) | ( ~n894 & n1128 ) | ( n1109 & n1128 ) ;
  buffer buf_n1130( .i (n190), .o (n1130) );
  assign n1131 = ~n1129 & n1130 ;
  assign n1132 = ( n192 & n1111 ) | ( n192 & ~n1131 ) | ( n1111 & ~n1131 ) ;
  buffer buf_n1133( .i (n1106), .o (n1133) );
  assign n1134 = n1008 & n1133 ;
  assign n1135 = ( n282 & n924 ) | ( n282 & n1134 ) | ( n924 & n1134 ) ;
  assign n1136 = ~n852 & n1135 ;
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n872), .o (n1139) );
  assign n1140 = n1137 | n1139 ;
  assign n1141 = ( n1132 & n1138 ) | ( n1132 & n1140 ) | ( n1138 & n1140 ) ;
  assign n1142 = n1104 | n1141 ;
  assign n1143 = ( ~n978 & n1086 ) | ( ~n978 & n1142 ) | ( n1086 & n1142 ) ;
  assign n1144 = n979 | n1143 ;
  buffer buf_n1145( .i (n188), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  assign n1147 = n690 & ~n1146 ;
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n1148( .i (n1057), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1035), .o (n1150) );
  assign n1151 = ( n689 & ~n1149 ) | ( n689 & n1150 ) | ( ~n1149 & n1150 ) ;
  assign n1152 = ( n989 & n1146 ) | ( n989 & n1151 ) | ( n1146 & n1151 ) ;
  assign n1153 = ( n1130 & n1147 ) | ( n1130 & ~n1152 ) | ( n1147 & ~n1152 ) ;
  buffer buf_n1154( .i (n869), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  assign n1157 = ( n855 & n1153 ) | ( n855 & n1156 ) | ( n1153 & n1156 ) ;
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1083), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  assign n1161 = ( ~n147 & n1158 ) | ( ~n147 & n1160 ) | ( n1158 & n1160 ) ;
  assign n1162 = ( n100 & ~n1158 ) | ( n100 & n1160 ) | ( ~n1158 & n1160 ) ;
  assign n1163 = n1161 & ~n1162 ;
  buffer buf_n1164( .i (n536), .o (n1164) );
  assign n1165 = ( ~n1035 & n1148 ) | ( ~n1035 & n1164 ) | ( n1148 & n1164 ) ;
  assign n1166 = ~n536 & n1075 ;
  assign n1167 = ( n757 & n1148 ) | ( n757 & ~n1166 ) | ( n1148 & ~n1166 ) ;
  assign n1168 = ~n1165 & n1167 ;
  assign n1169 = n1039 & n1168 ;
  buffer buf_n1170( .i (n1075), .o (n1170) );
  assign n1171 = n1164 & n1170 ;
  buffer buf_n1172( .i (n1093), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  assign n1174 = n1057 | n1173 ;
  assign n1175 = n1164 & n1174 ;
  assign n1176 = ( n988 & n1171 ) | ( n988 & ~n1175 ) | ( n1171 & ~n1175 ) ;
  assign n1177 = n1039 | n1176 ;
  assign n1178 = ( ~n840 & n1169 ) | ( ~n840 & n1177 ) | ( n1169 & n1177 ) ;
  assign n1179 = n898 & ~n1178 ;
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n1180( .i (n1032), .o (n1180) );
  assign n1181 = ~n947 & n1180 ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  assign n1184 = ( n1149 & n1150 ) | ( n1149 & ~n1182 ) | ( n1150 & ~n1182 ) ;
  assign n1185 = ( n950 & ~n1183 ) | ( n950 & n1184 ) | ( ~n1183 & n1184 ) ;
  buffer buf_n1186( .i (n1038), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  assign n1188 = ~n1185 & n1187 ;
  buffer buf_n1189( .i (n894), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  assign n1191 = n1188 | n1190 ;
  assign n1192 = ~n1179 & n1191 ;
  assign n1193 = ( n19 & n89 ) | ( n19 & n1027 ) | ( n89 & n1027 ) ;
  assign n1194 = ( ~n1050 & n1092 ) | ( ~n1050 & n1193 ) | ( n1092 & n1193 ) ;
  buffer buf_n1195( .i (n1194), .o (n1195) );
  assign n1198 = n1172 & ~n1195 ;
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  assign n1201 = n1197 | n1199 ;
  buffer buf_n1202( .i (n757), .o (n1202) );
  assign n1203 = ( n1200 & n1201 ) | ( n1200 & ~n1202 ) | ( n1201 & ~n1202 ) ;
  assign n1204 = ~n1146 & n1203 ;
  buffer buf_n1205( .i (n665), .o (n1205) );
  assign n1206 = ~n1204 & n1205 ;
  assign n1207 = n921 & n1173 ;
  assign n1208 = ( n1133 & n1164 ) | ( n1133 & ~n1207 ) | ( n1164 & ~n1207 ) ;
  assign n1209 = n318 & n1208 ;
  assign n1210 = ~n1186 & n1209 ;
  assign n1211 = n1205 | n1210 ;
  assign n1212 = ~n1206 & n1211 ;
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1156), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  assign n1216 = ( n1192 & n1213 ) | ( n1192 & n1215 ) | ( n1213 & n1215 ) ;
  buffer buf_n1217( .i (n44), .o (n1217) );
  assign n1218 = ( n944 & ~n1092 ) | ( n944 & n1217 ) | ( ~n1092 & n1217 ) ;
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  assign n1223 = ( n1032 & ~n1087 ) | ( n1032 & n1219 ) | ( ~n1087 & n1219 ) ;
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  assign n1226 = ~n948 & n1224 ;
  assign n1227 = ( ~n1222 & n1225 ) | ( ~n1222 & n1226 ) | ( n1225 & n1226 ) ;
  buffer buf_n1228( .i (n893), .o (n1228) );
  assign n1229 = ~n1227 & n1228 ;
  buffer buf_n1230( .i (n1087), .o (n1230) );
  assign n1231 = n1057 | n1230 ;
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1235( .i (n1180), .o (n1235) );
  assign n1236 = ~n757 & n1235 ;
  assign n1237 = ~n1232 & n1236 ;
  assign n1238 = n1228 | n1237 ;
  assign n1239 = ~n1229 & n1238 ;
  assign n1240 = n1083 | n1239 ;
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  assign n1241 = n970 & ~n1234 ;
  buffer buf_n1242( .i (n1187), .o (n1242) );
  assign n1243 = ~n1241 & n1242 ;
  assign n1244 = n1240 & ~n1243 ;
  assign n1245 = ( n1213 & ~n1215 ) | ( n1213 & n1244 ) | ( ~n1215 & n1244 ) ;
  assign n1246 = n1216 | n1245 ;
  assign n1247 = n1163 | n1246 ;
  assign n1248 = ( ~n936 & n1144 ) | ( ~n936 & n1247 ) | ( n1144 & n1247 ) ;
  assign n1249 = n937 | n1248 ;
  assign y0 = n316 ;
  assign y1 = n488 ;
  assign y2 = n701 ;
  assign y3 = n911 ;
  assign y4 = n1249 ;
endmodule
