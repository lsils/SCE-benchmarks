module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n2 , n4 , n5 , n6 , n7 , n8 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n18 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n33 , n34 , n35 , n36 , n37 , n38 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n49 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n66 , n67 , n68 , n69 , n70 , n71 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n82 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n99 , n100 , n101 , n102 , n103 , n104 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n115 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n132 , n133 , n134 , n135 , n136 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n146 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n162 , n163 , n164 , n165 , n166 , n168 , n169 , n170 , n171 , n172 , n173 , n175 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n189 , n190 , n191 , n192 , n194 , n195 , n196 , n197 , n198 , n199 , n201 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n216 , n217 , n218 , n219 , n220 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n230 , n231 , n232 , n233 , n234 , n235 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n251 , n252 , n253 , n255 , n256 , n257 , n258 , n259 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 ;
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n4( .i (x1), .o (n4) );
  assign n264 = ~n2 & n4 ;
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n82( .i (x11), .o (n82) );
  buffer buf_n99( .i (x13), .o (n99) );
  assign n272 = ~n82 & n99 ;
  buffer buf_n273( .i (n272), .o (n273) );
  assign n280 = n265 | n273 ;
  buffer buf_n18( .i (x3), .o (n18) );
  buffer buf_n33( .i (x5), .o (n33) );
  assign n281 = ~n18 & n33 ;
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n146( .i (x19), .o (n146) );
  buffer buf_n162( .i (x21), .o (n162) );
  assign n290 = ~n146 & n162 ;
  buffer buf_n291( .i (n290), .o (n291) );
  assign n300 = n282 | n291 ;
  assign n301 = n280 | n300 ;
  buffer buf_n49( .i (x7), .o (n49) );
  buffer buf_n66( .i (x9), .o (n66) );
  assign n302 = ~n49 & n66 ;
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n201( .i (x27), .o (n201) );
  buffer buf_n216( .i (x29), .o (n216) );
  assign n311 = ~n201 & n216 ;
  buffer buf_n312( .i (n311), .o (n312) );
  assign n320 = n303 | n312 ;
  buffer buf_n115( .i (x15), .o (n115) );
  buffer buf_n132( .i (x17), .o (n132) );
  assign n321 = ~n115 & n132 ;
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n175( .i (x23), .o (n175) );
  buffer buf_n189( .i (x25), .o (n189) );
  assign n330 = ~n175 & n189 ;
  buffer buf_n331( .i (n330), .o (n331) );
  assign n336 = n322 | n331 ;
  assign n337 = n320 | n336 ;
  assign n338 = n301 | n337 ;
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n230( .i (x31), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n251( .i (x33), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  assign n345 = ~n231 & n252 ;
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  assign n350 = n339 | n349 ;
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n168( .i (x22), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n292( .i (n291), .o (n292) );
  assign n370 = ( n165 & n292 ) | ( n165 & ~n346 ) | ( n292 & ~n346 ) ;
  buffer buf_n371( .i (n370), .o (n371) );
  assign n377 = ~n173 & n371 ;
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n166( .i (n165), .o (n166) );
  assign n379 = n166 & ~n172 ;
  assign n380 = n294 & n379 ;
  buffer buf_n381( .i (n380), .o (n381) );
  assign n382 = ( ~n340 & n378 ) | ( ~n340 & n381 ) | ( n378 & n381 ) ;
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n106( .i (x14), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  assign n394 = n100 & ~n107 ;
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n10( .i (x2), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  assign n396 = n5 & ~n11 ;
  buffer buf_n397( .i (n396), .o (n397) );
  assign n398 = n395 | n397 ;
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n40( .i (x6), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  assign n399 = n34 & ~n41 ;
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  assign n402 = n398 | n401 ;
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n73( .i (x10), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  assign n403 = n67 & ~n74 ;
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n138( .i (x18), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  assign n405 = n133 & ~n139 ;
  buffer buf_n406( .i (n405), .o (n406) );
  assign n407 = n404 | n406 ;
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n222( .i (x30), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  assign n408 = n217 & ~n223 ;
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n255( .i (x34), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  assign n410 = n253 & ~n257 ;
  assign n411 = n409 | n410 ;
  assign n412 = n407 | n411 ;
  assign n413 = n402 | n412 ;
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  assign n416 = ~n351 & n415 ;
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n258( .i (n257), .o (n258) );
  assign n418 = ~n258 & n346 ;
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n323( .i (n322), .o (n323) );
  assign n420 = n323 & n406 ;
  buffer buf_n421( .i (n420), .o (n421) );
  assign n425 = n419 | n421 ;
  buffer buf_n313( .i (n312), .o (n313) );
  assign n426 = n313 & n409 ;
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  assign n431 = n425 | n428 ;
  buffer buf_n274( .i (n273), .o (n274) );
  assign n432 = n274 & n395 ;
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n304( .i (n303), .o (n304) );
  assign n437 = n304 & n404 ;
  buffer buf_n438( .i (n437), .o (n438) );
  assign n443 = n433 | n438 ;
  buffer buf_n283( .i (n282), .o (n283) );
  assign n444 = n283 & n400 ;
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n266( .i (n265), .o (n266) );
  assign n450 = n266 & n397 ;
  buffer buf_n451( .i (n450), .o (n451) );
  assign n454 = n445 | n451 ;
  assign n455 = n443 | n454 ;
  assign n456 = n431 | n455 ;
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n194( .i (x26), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n332( .i (n331), .o (n332) );
  assign n458 = ( n192 & n332 ) | ( n192 & ~n346 ) | ( n332 & ~n346 ) ;
  buffer buf_n459( .i (n458), .o (n459) );
  assign n461 = ~n199 & n459 ;
  buffer buf_n333( .i (n332), .o (n333) );
  assign n462 = n192 & ~n197 ;
  assign n463 = n333 & n462 ;
  buffer buf_n464( .i (n463), .o (n464) );
  assign n465 = ( ~n339 & n461 ) | ( ~n339 & n464 ) | ( n461 & n464 ) ;
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  assign n469 = n457 | n467 ;
  assign n470 = n417 | n469 ;
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  assign n479 = n393 | n478 ;
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n460( .i (n459), .o (n460) );
  assign n486 = ( n335 & ~n339 ) | ( n335 & n460 ) | ( ~n339 & n460 ) ;
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  assign n489 = ( ~n457 & n467 ) | ( ~n457 & n488 ) | ( n467 & n488 ) ;
  assign n490 = ( ~n417 & n468 ) | ( ~n417 & n489 ) | ( n468 & n489 ) ;
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n203( .i (x28), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n497 = n384 & ~n468 ;
  assign n498 = n214 | n497 ;
  assign n499 = n491 & ~n498 ;
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n177( .i (x24), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  assign n503 = ~n187 & n299 ;
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  assign n504 = ~n187 & n376 ;
  assign n505 = ( ~n344 & n503 ) | ( ~n344 & n504 ) | ( n503 & n504 ) ;
  assign n506 = ~n184 & n381 ;
  assign n507 = ~n184 & n378 ;
  assign n508 = ( ~n341 & n506 ) | ( ~n341 & n507 ) | ( n506 & n507 ) ;
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  assign n512 = ( ~n471 & n505 ) | ( ~n471 & n511 ) | ( n505 & n511 ) ;
  buffer buf_n513( .i (n512), .o (n513) );
  assign n515 = n500 | n513 ;
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n117( .i (x16), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  assign n520 = ( n104 & n276 ) | ( n104 & ~n348 ) | ( n276 & ~n348 ) ;
  buffer buf_n521( .i (n520), .o (n521) );
  assign n523 = ~n113 & n521 ;
  assign n524 = ( ~n341 & n436 ) | ( ~n341 & n523 ) | ( n436 & n523 ) ;
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  assign n529 = ~n130 & n528 ;
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n522( .i (n521), .o (n522) );
  assign n530 = ( n279 & ~n341 ) | ( n279 & n522 ) | ( ~n341 & n522 ) ;
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  assign n533 = ( ~n385 & n526 ) | ( ~n385 & n532 ) | ( n526 & n532 ) ;
  buffer buf_n534( .i (n533), .o (n534) );
  assign n535 = ~n130 & n534 ;
  assign n536 = ( ~n473 & n529 ) | ( ~n473 & n535 ) | ( n529 & n535 ) ;
  buffer buf_n537( .i (n536), .o (n537) );
  assign n539 = n516 | n537 ;
  buffer buf_n84( .i (x12), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  assign n540 = ( n71 & n306 ) | ( n71 & ~n348 ) | ( n306 & ~n348 ) ;
  buffer buf_n541( .i (n540), .o (n541) );
  assign n544 = ~n80 & n541 ;
  buffer buf_n545( .i (n544), .o (n545) );
  assign n546 = ( ~n342 & n442 ) | ( ~n342 & n545 ) | ( n442 & n545 ) ;
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  assign n550 = ~n97 & n549 ;
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  assign n551 = ( n310 & ~n342 ) | ( n310 & n543 ) | ( ~n342 & n543 ) ;
  buffer buf_n552( .i (n551), .o (n552) );
  assign n553 = ( ~n385 & n547 ) | ( ~n385 & n552 ) | ( n547 & n552 ) ;
  buffer buf_n554( .i (n553), .o (n554) );
  assign n555 = ~n97 & n554 ;
  assign n556 = ( ~n473 & n550 ) | ( ~n473 & n555 ) | ( n550 & n555 ) ;
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n51( .i (x8), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  assign n561 = ( n38 & n285 ) | ( n38 & ~n348 ) | ( n285 & ~n348 ) ;
  buffer buf_n562( .i (n561), .o (n562) );
  assign n565 = ~n47 & n562 ;
  buffer buf_n566( .i (n565), .o (n566) );
  assign n567 = ( ~n342 & n449 ) | ( ~n342 & n566 ) | ( n449 & n566 ) ;
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  assign n571 = ~n64 & n570 ;
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n572( .i (n340), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  assign n574 = ( n289 & n564 ) | ( n289 & ~n573 ) | ( n564 & ~n573 ) ;
  buffer buf_n575( .i (n574), .o (n575) );
  assign n576 = ( ~n385 & n568 ) | ( ~n385 & n575 ) | ( n568 & n575 ) ;
  buffer buf_n577( .i (n576), .o (n577) );
  assign n578 = ~n64 & n577 ;
  assign n579 = ( ~n473 & n571 ) | ( ~n473 & n578 ) | ( n571 & n578 ) ;
  buffer buf_n580( .i (n579), .o (n580) );
  assign n584 = n557 | n580 ;
  assign n585 = n539 | n584 ;
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n20( .i (x4), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n267( .i (n266), .o (n267) );
  assign n588 = ( n8 & n267 ) | ( n8 & ~n347 ) | ( n267 & ~n347 ) ;
  buffer buf_n589( .i (n588), .o (n589) );
  assign n592 = ~n16 & n589 ;
  assign n593 = ( ~n340 & n453 ) | ( ~n340 & n592 ) | ( n453 & n592 ) ;
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  assign n601 = ~n31 & n596 ;
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  assign n602 = ( n271 & ~n572 ) | ( n271 & n591 ) | ( ~n572 & n591 ) ;
  assign n603 = ( ~n383 & n594 ) | ( ~n383 & n602 ) | ( n594 & n602 ) ;
  buffer buf_n604( .i (n603), .o (n604) );
  assign n609 = ~n31 & n604 ;
  assign n610 = ( ~n471 & n601 ) | ( ~n471 & n609 ) | ( n601 & n609 ) ;
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n261( .i (x35), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  assign n617 = n253 & ~n263 ;
  buffer buf_n618( .i (n617), .o (n618) );
  assign n625 = ~n259 & n618 ;
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  assign n630 = n233 | n258 ;
  assign n631 = n618 & ~n630 ;
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  assign n636 = ( ~n573 & n629 ) | ( ~n573 & n635 ) | ( n629 & n635 ) ;
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  assign n640 = ~n235 & n619 ;
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  assign n645 = ( ~n343 & n624 ) | ( ~n343 & n644 ) | ( n624 & n644 ) ;
  buffer buf_n646( .i (n645), .o (n646) );
  assign n647 = ( ~n386 & n638 ) | ( ~n386 & n646 ) | ( n638 & n646 ) ;
  assign n648 = ( ~n472 & n639 ) | ( ~n472 & n647 ) | ( n639 & n647 ) ;
  assign n649 = n611 | n648 ;
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n148( .i (x20), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n324( .i (n323), .o (n324) );
  assign n653 = ( n136 & n324 ) | ( n136 & ~n347 ) | ( n324 & ~n347 ) ;
  buffer buf_n654( .i (n653), .o (n654) );
  assign n658 = ~n144 & n654 ;
  buffer buf_n659( .i (n658), .o (n659) );
  assign n660 = ( n424 & ~n572 ) | ( n424 & n659 ) | ( ~n572 & n659 ) ;
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  assign n665 = ~n160 & n663 ;
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  assign n666 = ( n329 & ~n573 ) | ( n329 & n657 ) | ( ~n573 & n657 ) ;
  assign n667 = ( ~n384 & n661 ) | ( ~n384 & n666 ) | ( n661 & n666 ) ;
  buffer buf_n668( .i (n667), .o (n668) );
  assign n670 = ~n160 & n668 ;
  assign n671 = ( ~n472 & n665 ) | ( ~n472 & n670 ) | ( n665 & n670 ) ;
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n237( .i (x32), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n314( .i (n313), .o (n314) );
  assign n675 = ( n220 & n314 ) | ( n220 & ~n347 ) | ( n314 & ~n347 ) ;
  buffer buf_n676( .i (n675), .o (n676) );
  assign n680 = ~n228 & n676 ;
  buffer buf_n681( .i (n680), .o (n681) );
  assign n682 = ( n430 & ~n572 ) | ( n430 & n681 ) | ( ~n572 & n681 ) ;
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  assign n689 = ~n249 & n685 ;
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  assign n690 = ( n319 & ~n573 ) | ( n319 & n679 ) | ( ~n573 & n679 ) ;
  assign n691 = ( ~n384 & n683 ) | ( ~n384 & n690 ) | ( n683 & n690 ) ;
  buffer buf_n692( .i (n691), .o (n692) );
  assign n696 = ~n249 & n692 ;
  assign n697 = ( ~n472 & n689 ) | ( ~n472 & n696 ) | ( n689 & n696 ) ;
  buffer buf_n698( .i (n697), .o (n698) );
  assign n703 = n672 | n698 ;
  assign n704 = n650 | n703 ;
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  assign n709 = n587 | n707 ;
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n715( .i (n471), .o (n715) );
  assign n716 = ( n549 & n554 ) | ( n549 & ~n715 ) | ( n554 & ~n715 ) ;
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  assign n719 = ~n537 & n718 ;
  assign n720 = ~n517 & n719 ;
  assign n721 = ~n705 & n720 ;
  assign n722 = n560 | n721 ;
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  assign n724 = ( n570 & n577 ) | ( n570 & ~n715 ) | ( n577 & ~n715 ) ;
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  assign n729 = ( n582 & ~n705 ) | ( n582 & n728 ) | ( ~n705 & n728 ) ;
  assign n730 = ( n583 & ~n586 ) | ( n583 & n729 ) | ( ~n586 & n729 ) ;
  buffer buf_n731( .i (n730), .o (n731) );
  assign n733 = n723 | n731 ;
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  assign n735 = n538 | n674 ;
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  assign n740 = n519 & ~n736 ;
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n669( .i (n668), .o (n669) );
  assign n743 = ( n664 & n669 ) | ( n664 & ~n715 ) | ( n669 & ~n715 ) ;
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  assign n748 = ( n528 & n534 ) | ( n528 & ~n715 ) | ( n534 & ~n715 ) ;
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  assign n753 = n747 | n752 ;
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  assign n756 = ~n741 & n755 ;
  buffer buf_n708( .i (n707), .o (n708) );
  assign n757 = n708 & ~n738 ;
  assign n758 = ( n739 & n756 ) | ( n739 & ~n757 ) | ( n756 & ~n757 ) ;
  assign n759 = n734 | n758 ;
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  assign n762 = ( ~n474 & n600 ) | ( ~n474 & n608 ) | ( n600 & n608 ) ;
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  assign n765 = ( n615 & ~n705 ) | ( n615 & n764 ) | ( ~n705 & n764 ) ;
  assign n766 = ( ~n586 & n616 ) | ( ~n586 & n765 ) | ( n616 & n765 ) ;
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  assign n772 = ( n299 & ~n343 ) | ( n299 & n376 ) | ( ~n343 & n376 ) ;
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  assign n777 = ( n389 & ~n474 ) | ( n389 & n776 ) | ( ~n474 & n776 ) ;
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  assign n779 = n218 | n253 ;
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  assign n791 = n493 | n790 ;
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  assign n794 = n778 | n793 ;
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  assign n798 = ~n767 & n797 ;
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  assign n802 = ( n760 & ~n771 ) | ( n760 & n801 ) | ( ~n771 & n801 ) ;
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  assign n803 = n496 | n778 ;
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  assign n806 = ~n754 & n805 ;
  assign n807 = ~n708 & n806 ;
  assign n808 = n742 | n807 ;
  assign n809 = n734 | n808 ;
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n514( .i (n513), .o (n514) );
  assign n812 = n514 & ~n672 ;
  buffer buf_n813( .i (n812), .o (n813) );
  assign n814 = n538 | n813 ;
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  assign n818 = ~n746 & n778 ;
  assign n819 = ~n652 & n818 ;
  assign n820 = n702 | n819 ;
  assign n821 = n651 | n674 ;
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  assign n823 = ( ~n474 & n688 ) | ( ~n474 & n695 ) | ( n688 & n695 ) ;
  buffer buf_n824( .i (n823), .o (n824) );
  assign n825 = ~n496 & n824 ;
  assign n826 = n752 | n825 ;
  assign n827 = ~n822 & n826 ;
  assign n828 = n820 | n827 ;
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  assign n829 = n502 & ~n537 ;
  assign n830 = ~n813 & n829 ;
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  assign n834 = ( n817 & n828 ) | ( n817 & ~n833 ) | ( n828 & ~n833 ) ;
  assign n835 = n723 & ~n731 ;
  assign n836 = ( n732 & n834 ) | ( n732 & ~n835 ) | ( n834 & ~n835 ) ;
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  assign y0 = n369 ;
  assign y1 = n485 ;
  assign y2 = n714 ;
  assign y3 = n802 ;
  assign y4 = n761 ;
  assign y5 = n811 ;
  assign y6 = n839 ;
endmodule
