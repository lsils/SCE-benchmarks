module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G158 , G159 , G16 , G160 , G161 , G162 , G163 , G164 , G165 , G166 , G167 , G168 , G169 , G17 , G170 , G171 , G172 , G173 , G174 , G175 , G176 , G177 , G178 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 , G5193 , G5194 , G5195 , G5196 , G5197 , G5198 , G5199 , G5200 , G5201 , G5202 , G5203 , G5204 , G5205 , G5206 , G5207 , G5208 , G5209 , G5210 , G5211 , G5212 , G5213 , G5214 , G5215 , G5216 , G5217 , G5218 , G5219 , G5220 , G5221 , G5222 , G5223 , G5224 , G5225 , G5226 , G5227 , G5228 , G5229 , G5230 , G5231 , G5232 , G5233 , G5234 , G5235 , G5236 , G5237 , G5238 , G5239 , G5240 , G5241 , G5242 , G5243 , G5244 , G5245 , G5246 , G5247 , G5248 , G5249 , G5250 , G5251 , G5252 , G5253 , G5254 , G5255 , G5256 , G5257 , G5258 , G5259 , G5260 , G5261 , G5262 , G5263 , G5264 , G5265 , G5266 , G5267 , G5268 , G5269 , G5270 , G5271 , G5272 , G5273 , G5274 , G5275 , G5276 , G5277 , G5278 , G5279 , G5280 , G5281 , G5282 , G5283 , G5284 , G5285 , G5286 , G5287 , G5288 , G5289 , G5290 , G5291 , G5292 , G5293 , G5294 , G5295 , G5296 , G5297 , G5298 , G5299 , G5300 , G5301 , G5302 , G5303 , G5304 , G5305 , G5306 , G5307 , G5308 , G5309 , G5310 , G5311 , G5312 , G5313 , G5314 , G5315 );
  input G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G158 , G159 , G16 , G160 , G161 , G162 , G163 , G164 , G165 , G166 , G167 , G168 , G169 , G17 , G170 , G171 , G172 , G173 , G174 , G175 , G176 , G177 , G178 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 ;
  output G5193 , G5194 , G5195 , G5196 , G5197 , G5198 , G5199 , G5200 , G5201 , G5202 , G5203 , G5204 , G5205 , G5206 , G5207 , G5208 , G5209 , G5210 , G5211 , G5212 , G5213 , G5214 , G5215 , G5216 , G5217 , G5218 , G5219 , G5220 , G5221 , G5222 , G5223 , G5224 , G5225 , G5226 , G5227 , G5228 , G5229 , G5230 , G5231 , G5232 , G5233 , G5234 , G5235 , G5236 , G5237 , G5238 , G5239 , G5240 , G5241 , G5242 , G5243 , G5244 , G5245 , G5246 , G5247 , G5248 , G5249 , G5250 , G5251 , G5252 , G5253 , G5254 , G5255 , G5256 , G5257 , G5258 , G5259 , G5260 , G5261 , G5262 , G5263 , G5264 , G5265 , G5266 , G5267 , G5268 , G5269 , G5270 , G5271 , G5272 , G5273 , G5274 , G5275 , G5276 , G5277 , G5278 , G5279 , G5280 , G5281 , G5282 , G5283 , G5284 , G5285 , G5286 , G5287 , G5288 , G5289 , G5290 , G5291 , G5292 , G5293 , G5294 , G5295 , G5296 , G5297 , G5298 , G5299 , G5300 , G5301 , G5302 , G5303 , G5304 , G5305 , G5306 , G5307 , G5308 , G5309 , G5310 , G5311 , G5312 , G5313 , G5314 , G5315 ;
  wire n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 ;
  buffer buf_n1024( .i (G66), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  inverter inv_n1026( .i (n1025), .o (n1026) );
  buffer buf_n288( .i (G113), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  inverter inv_n312( .i (n311), .o (n312) );
  buffer buf_n941( .i (G165), .o (n941) );
  inverter inv_n942( .i (n941), .o (n942) );
  inverter inv_n889( .i (G151), .o (n889) );
  buffer buf_n496( .i (G127), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  inverter inv_n529( .i (n528), .o (n529) );
  buffer buf_n607( .i (G131), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  inverter inv_n640( .i (n639), .o (n640) );
  buffer buf_n892( .i (G153), .o (n892) );
  buffer buf_n908( .i (G156), .o (n908) );
  assign n1183 = n892 & n908 ;
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n890( .i (G152), .o (n890) );
  inverter inv_n891( .i (n890), .o (n891) );
  buffer buf_n444( .i (G125), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  inverter inv_n474( .i (n473), .o (n474) );
  buffer buf_n553( .i (G129), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  inverter inv_n588( .i (n587), .o (n588) );
  assign n1190 = G67 & n1025 ;
  buffer buf_n1175( .i (G99), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n1181( .i (n1180), .o (n1181) );
  inverter inv_n1182( .i (n1181), .o (n1182) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  inverter inv_n899( .i (n898), .o (n899) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  inverter inv_n915( .i (n914), .o (n915) );
  buffer buf_n900( .i (G155), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  inverter inv_n907( .i (n906), .o (n907) );
  buffer buf_n179( .i (G1), .o (n179) );
  assign n1191 = G134 & n179 ;
  assign n1192 = G63 & ~n941 ;
  buffer buf_n280( .i (G11), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  assign n1193 = G164 | ~n285 ;
  assign n1194 = G136 & G154 ;
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  inverter inv_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1020( .i (G64), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1235( .i (n1024), .o (n1235) );
  buffer buf_n4222( .i (n1235), .o (n4222) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n4223( .i (n890), .o (n4223) );
  buffer buf_n313( .i (G114), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  assign n1202 = G12 & n280 ;
  buffer buf_n1203( .i (n1202), .o (n1203) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  assign n1208 = ~G65 | ~n1206 ;
  inverter inv_n1207( .i (n1206), .o (n1207) );
  inverter inv_n4224( .i (n179), .o (n4224) );
  inverter inv_n4225( .i (n336), .o (n4225) );
  buffer buf_n938( .i (G163), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  assign n1209 = G34 & n940 ;
  assign n1210 = G33 & ~n940 ;
  assign n1211 = n1209 | n1210 ;
  assign n1212 = ~n1206 | ~n1211 ;
  assign n1213 = G13 & n939 ;
  assign n1214 = G35 & ~n939 ;
  assign n1215 = n1213 | n1214 ;
  assign n1216 = n1205 & n1215 ;
  inverter inv_n1217( .i (n1216), .o (n1217) );
  assign n1218 = ~G32 | ~n1206 ;
  assign n1219 = G9 & ~n940 ;
  assign n1220 = G8 & n939 ;
  assign n1221 = n1204 & ~n1220 ;
  assign n1222 = ~n1219 & n1221 ;
  assign n1223 = n1025 & ~n1222 ;
  assign n1224 = G30 & ~n940 ;
  buffer buf_n1225( .i (n938), .o (n1225) );
  assign n1226 = G10 & n1225 ;
  assign n1227 = n1204 & ~n1226 ;
  assign n1228 = ~n1224 & n1227 ;
  assign n1229 = n1025 & ~n1228 ;
  buffer buf_n1230( .i (n1225), .o (n1230) );
  assign n1231 = G7 & ~n1230 ;
  assign n1232 = G28 & n1225 ;
  assign n1233 = n1204 & ~n1232 ;
  assign n1234 = ~n1231 & n1233 ;
  assign n1236 = ~n1234 & n1235 ;
  assign n1237 = G29 & ~n1230 ;
  assign n1238 = G31 & n1225 ;
  buffer buf_n1239( .i (n1203), .o (n1239) );
  assign n1240 = ~n1238 & n1239 ;
  assign n1241 = ~n1237 & n1240 ;
  assign n1242 = n1235 & ~n1241 ;
  buffer buf_n818( .i (G145), .o (n818) );
  buffer buf_n181( .i (G100), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n349( .i (G117), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  assign n1243 = n182 | n350 ;
  buffer buf_n185( .i (G101), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n1244 = ~n186 & n350 ;
  assign n1245 = n1243 & ~n1244 ;
  assign n1246 = n818 & ~n1245 ;
  buffer buf_n189( .i (G102), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  assign n1247 = n190 & n350 ;
  buffer buf_n1171( .i (G98), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1248( .i (n349), .o (n1248) );
  assign n1249 = n1172 & ~n1248 ;
  assign n1250 = n1247 | n1249 ;
  assign n1251 = ~n818 & n1250 ;
  assign n1252 = n1246 | n1251 ;
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n821( .i (G146), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n363( .i (G119), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  assign n1263 = n182 | n366 ;
  assign n1264 = ~n186 & n366 ;
  assign n1265 = n1263 & ~n1264 ;
  assign n1266 = n823 & ~n1265 ;
  assign n1267 = n190 & n366 ;
  buffer buf_n1268( .i (n365), .o (n1268) );
  assign n1269 = n1172 & ~n1268 ;
  assign n1270 = n1267 | n1269 ;
  assign n1271 = ~n823 & n1270 ;
  assign n1272 = n1266 | n1271 ;
  buffer buf_n1273( .i (n1272), .o (n1273) );
  assign n1283 = n1253 & n1273 ;
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n870( .i (G150), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n530( .i (G128), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n952( .i (G169), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  assign n1294 = n549 | n953 ;
  buffer buf_n949( .i (G168), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  assign n1295 = n549 & ~n950 ;
  assign n1296 = n1294 & ~n1295 ;
  assign n1297 = n888 & ~n1296 ;
  buffer buf_n946( .i (G167), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  assign n1298 = n549 & n947 ;
  buffer buf_n943( .i (G166), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n1299( .i (n548), .o (n1299) );
  assign n1300 = n944 & ~n1299 ;
  assign n1301 = n1298 | n1300 ;
  assign n1302 = ~n888 & n1301 ;
  assign n1303 = n1297 | n1302 ;
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  assign n1305 = n289 | n1174 ;
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  assign n1306 = ~n192 & n289 ;
  assign n1307 = n1305 & ~n1306 ;
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n338( .i (G115), .o (n338) );
  assign n1324 = n184 | n338 ;
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  assign n1325 = ~n188 & n338 ;
  assign n1326 = n1324 & ~n1325 ;
  buffer buf_n1327( .i (n1326), .o (n1327) );
  assign n1338 = n1308 & ~n1327 ;
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n589( .i (G130), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  assign n1346 = n182 | n597 ;
  assign n1347 = ~n186 & n597 ;
  assign n1348 = n1346 & ~n1347 ;
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n839( .i (G148), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  assign n1362 = ~n851 & n944 ;
  assign n1363 = n851 & ~n953 ;
  assign n1364 = n1362 | n1363 ;
  buffer buf_n1365( .i (n1364), .o (n1365) );
  assign n1366 = ~n1358 & n1365 ;
  assign n1367 = n1345 & n1366 ;
  assign n1368 = n1304 & n1367 ;
  buffer buf_n824( .i (G147), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n379( .i (G121), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  assign n1369 = n394 | n953 ;
  assign n1370 = n394 & ~n950 ;
  assign n1371 = n1369 & ~n1370 ;
  assign n1372 = n838 & ~n1371 ;
  assign n1373 = n394 & n947 ;
  buffer buf_n1374( .i (n393), .o (n1374) );
  assign n1375 = n944 & ~n1374 ;
  assign n1376 = n1373 | n1375 ;
  assign n1377 = ~n838 & n1376 ;
  assign n1378 = n1372 | n1377 ;
  buffer buf_n1379( .i (n1378), .o (n1379) );
  buffer buf_n852( .i (G149), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n475( .i (G126), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n1380( .i (n952), .o (n1380) );
  assign n1381 = n492 | n1380 ;
  assign n1382 = n492 & ~n950 ;
  assign n1383 = n1381 & ~n1382 ;
  assign n1384 = n868 & ~n1383 ;
  assign n1385 = n492 & n947 ;
  buffer buf_n1386( .i (n491), .o (n1386) );
  buffer buf_n1387( .i (n943), .o (n1387) );
  assign n1388 = ~n1386 & n1387 ;
  assign n1389 = n1385 | n1388 ;
  assign n1390 = ~n868 & n1389 ;
  assign n1391 = n1384 | n1390 ;
  buffer buf_n1392( .i (n1391), .o (n1392) );
  assign n1393 = n1379 & n1392 ;
  assign n1394 = n1368 & n1393 ;
  assign n1395 = n1293 & n1394 ;
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n722( .i (G140), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n1125( .i (G94), .o (n1125) );
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  assign n1404 = n1147 | n1380 ;
  buffer buf_n1405( .i (n949), .o (n1405) );
  assign n1406 = n1147 & ~n1405 ;
  assign n1407 = n1404 & ~n1406 ;
  assign n1408 = n743 & ~n1407 ;
  buffer buf_n1409( .i (n946), .o (n1409) );
  assign n1410 = n1147 & n1409 ;
  buffer buf_n1411( .i (n1146), .o (n1411) );
  assign n1412 = n1387 & ~n1411 ;
  assign n1413 = n1410 | n1412 ;
  assign n1414 = ~n743 & n1413 ;
  assign n1415 = n1408 | n1414 ;
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n775( .i (G143), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n1072( .i (G90), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  assign n1420 = n1092 | n1380 ;
  assign n1421 = n1092 & ~n1405 ;
  assign n1422 = n1420 & ~n1421 ;
  assign n1423 = n794 & ~n1422 ;
  assign n1424 = n1092 & n1409 ;
  buffer buf_n1425( .i (n1091), .o (n1425) );
  assign n1426 = n1387 & ~n1425 ;
  assign n1427 = n1424 | n1426 ;
  assign n1428 = ~n794 & n1427 ;
  assign n1429 = n1423 | n1428 ;
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n795( .i (G144), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n1097( .i (G92), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  assign n1433 = n1120 | n1380 ;
  assign n1434 = n1120 & ~n1405 ;
  assign n1435 = n1433 & ~n1434 ;
  assign n1436 = n817 & ~n1435 ;
  assign n1437 = n1120 & n1409 ;
  buffer buf_n1438( .i (n1119), .o (n1438) );
  assign n1439 = n1387 & ~n1438 ;
  assign n1440 = n1437 | n1439 ;
  assign n1441 = ~n817 & n1440 ;
  assign n1442 = n1436 | n1441 ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  assign n1446 = n1432 & n1445 ;
  assign n1447 = n1419 & n1446 ;
  buffer buf_n644( .i (G135), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n259( .i (G109), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n954( .i (n953), .o (n954) );
  assign n1448 = n279 | n954 ;
  buffer buf_n951( .i (n950), .o (n951) );
  assign n1449 = n279 & ~n951 ;
  assign n1450 = n1448 & ~n1449 ;
  assign n1451 = n663 & ~n1450 ;
  buffer buf_n948( .i (n947), .o (n948) );
  assign n1452 = n279 & n948 ;
  buffer buf_n945( .i (n944), .o (n945) );
  assign n1453 = ~n279 & n945 ;
  assign n1454 = n1452 | n1453 ;
  assign n1455 = ~n663 & n1454 ;
  assign n1456 = n1451 | n1455 ;
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n744( .i (G141), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n1152( .i (G96), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  assign n1459 = n954 | n1170 ;
  assign n1460 = ~n951 & n1170 ;
  assign n1461 = n1459 & ~n1460 ;
  assign n1462 = n761 & ~n1461 ;
  assign n1463 = n948 & n1170 ;
  assign n1464 = n945 & ~n1170 ;
  assign n1465 = n1463 | n1464 ;
  assign n1466 = ~n761 & n1465 ;
  assign n1467 = n1462 | n1466 ;
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  assign n1470 = n1458 & n1469 ;
  buffer buf_n701( .i (G139), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n235( .i (G107), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  assign n1471 = n255 | n954 ;
  assign n1472 = n255 & ~n951 ;
  assign n1473 = n1471 & ~n1472 ;
  assign n1474 = n720 & ~n1473 ;
  assign n1475 = n255 & n948 ;
  buffer buf_n1476( .i (n254), .o (n1476) );
  assign n1477 = n945 & ~n1476 ;
  assign n1478 = n1475 | n1477 ;
  assign n1479 = ~n720 & n1478 ;
  assign n1480 = n1474 | n1479 ;
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n762( .i (G142), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n1047( .i (G88), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1482 = n188 | n1060 ;
  assign n1483 = ~n184 & n1060 ;
  assign n1484 = n1482 & ~n1483 ;
  assign n1485 = n774 & ~n1484 ;
  assign n1486 = n1060 & n1174 ;
  buffer buf_n1487( .i (n1059), .o (n1487) );
  assign n1488 = n192 & ~n1487 ;
  assign n1489 = n1486 | n1488 ;
  assign n1490 = ~n774 & n1489 ;
  assign n1491 = n1485 | n1490 ;
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  assign n1502 = n1481 & n1500 ;
  buffer buf_n664( .i (G137), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n193( .i (G103), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  assign n1503 = n211 | n954 ;
  assign n1504 = n211 & ~n951 ;
  assign n1505 = n1503 & ~n1504 ;
  assign n1506 = n681 & ~n1505 ;
  assign n1507 = n211 & n948 ;
  assign n1508 = ~n211 & n945 ;
  assign n1509 = n1507 | n1508 ;
  assign n1510 = ~n681 & n1509 ;
  assign n1511 = n1506 | n1510 ;
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n682( .i (G138), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n212( .i (G105), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n1513( .i (n952), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  assign n1515 = n231 | n1514 ;
  buffer buf_n1516( .i (n1405), .o (n1516) );
  assign n1517 = n231 & ~n1516 ;
  assign n1518 = n1515 & ~n1517 ;
  assign n1519 = n700 & ~n1518 ;
  buffer buf_n1520( .i (n1409), .o (n1520) );
  assign n1521 = n231 & n1520 ;
  buffer buf_n1522( .i (n230), .o (n1522) );
  buffer buf_n1523( .i (n943), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  assign n1525 = ~n1522 & n1524 ;
  assign n1526 = n1521 | n1525 ;
  assign n1527 = ~n700 & n1526 ;
  assign n1528 = n1519 | n1527 ;
  buffer buf_n1529( .i (n1528), .o (n1529) );
  assign n1530 = n1512 & n1529 ;
  assign n1531 = n1502 & n1530 ;
  assign n1532 = n1470 & n1531 ;
  assign n1533 = n1447 & n1532 ;
  buffer buf_n1534( .i (n1533), .o (n1534) );
  buffer buf_n1535( .i (n1534), .o (n1535) );
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n420( .i (G124), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  assign n1540 = n426 & n1152 ;
  assign n1541 = G97 & ~n426 ;
  assign n1542 = n1540 | n1541 ;
  buffer buf_n1543( .i (n1542), .o (n1543) );
  assign n1561 = n744 & n1543 ;
  buffer buf_n1562( .i (n1561), .o (n1562) );
  assign n1566 = n744 | n1543 ;
  buffer buf_n1567( .i (n1566), .o (n1567) );
  assign n1570 = ~n1562 & n1567 ;
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  assign n1579 = n259 & n424 ;
  assign n1580 = G110 & ~n424 ;
  assign n1581 = n1579 | n1580 ;
  buffer buf_n1582( .i (n1581), .o (n1582) );
  assign n1605 = n644 & n1582 ;
  buffer buf_n1606( .i (n1605), .o (n1606) );
  assign n1619 = n644 | n1582 ;
  buffer buf_n1620( .i (n1619), .o (n1620) );
  assign n1629 = ~n1606 & n1620 ;
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  assign n1647 = n235 & n424 ;
  buffer buf_n1648( .i (n423), .o (n1648) );
  assign n1649 = G108 & ~n1648 ;
  assign n1650 = n1647 | n1649 ;
  buffer buf_n1651( .i (n1650), .o (n1651) );
  assign n1674 = n701 | n1651 ;
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  assign n1684 = n701 & n1651 ;
  buffer buf_n1685( .i (n1684), .o (n1685) );
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  assign n1702 = n1677 & ~n1687 ;
  buffer buf_n1703( .i (n1702), .o (n1703) );
  assign n1718 = n1632 & n1703 ;
  buffer buf_n1719( .i (n1718), .o (n1719) );
  assign n1722 = n212 & n425 ;
  assign n1723 = G106 & ~n425 ;
  assign n1724 = n1722 | n1723 ;
  buffer buf_n1725( .i (n1724), .o (n1725) );
  assign n1747 = n682 & n1725 ;
  buffer buf_n1748( .i (n1747), .o (n1748) );
  assign n1749 = n682 | n1725 ;
  buffer buf_n1750( .i (n1749), .o (n1750) );
  assign n1753 = ~n1748 & n1750 ;
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  assign n1770 = n193 & n426 ;
  buffer buf_n1771( .i (n425), .o (n1771) );
  assign n1772 = G104 & ~n1771 ;
  assign n1773 = n1770 | n1772 ;
  buffer buf_n1774( .i (n1773), .o (n1774) );
  assign n1795 = n664 | n1774 ;
  buffer buf_n1796( .i (n1795), .o (n1796) );
  assign n1801 = n664 & n1774 ;
  buffer buf_n1802( .i (n1801), .o (n1802) );
  assign n1808 = n1796 & ~n1802 ;
  buffer buf_n1809( .i (n1808), .o (n1809) );
  assign n1824 = n1755 & n1809 ;
  buffer buf_n1825( .i (n1824), .o (n1825) );
  assign n1834 = n1719 & n1825 ;
  buffer buf_n1835( .i (n1834), .o (n1835) );
  assign n1845 = n1575 & n1835 ;
  buffer buf_n1846( .i (n1845), .o (n1846) );
  buffer buf_n1847( .i (n1846), .o (n1847) );
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n1849( .i (n1848), .o (n1849) );
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1850), .o (n1851) );
  buffer buf_n1852( .i (n1851), .o (n1852) );
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  assign n1855 = n423 & n1047 ;
  assign n1856 = G89 & ~n423 ;
  assign n1857 = n1855 | n1856 ;
  buffer buf_n1858( .i (n1857), .o (n1858) );
  assign n1879 = n762 & n1858 ;
  buffer buf_n1880( .i (n1879), .o (n1880) );
  assign n1900 = n762 | n1858 ;
  buffer buf_n1901( .i (n1900), .o (n1901) );
  assign n1920 = ~n1880 & n1901 ;
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  buffer buf_n1930( .i (n1929), .o (n1930) );
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n1934( .i (n1933), .o (n1934) );
  buffer buf_n1935( .i (n1934), .o (n1935) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1940( .i (n422), .o (n1940) );
  assign n1941 = n1072 & n1940 ;
  assign n1942 = G91 & ~n1940 ;
  assign n1943 = n1941 | n1942 ;
  buffer buf_n1944( .i (n1943), .o (n1944) );
  assign n1968 = n775 & n1944 ;
  buffer buf_n1969( .i (n1968), .o (n1969) );
  assign n1986 = n775 | n1944 ;
  buffer buf_n1987( .i (n1986), .o (n1987) );
  assign n1996 = ~n1969 & n1987 ;
  buffer buf_n1997( .i (n1996), .o (n1997) );
  buffer buf_n1998( .i (n1997), .o (n1998) );
  buffer buf_n1999( .i (n1998), .o (n1999) );
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n2001( .i (n2000), .o (n2001) );
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n2003), .o (n2004) );
  buffer buf_n2005( .i (n2004), .o (n2005) );
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n2007( .i (n2006), .o (n2007) );
  buffer buf_n2008( .i (n2007), .o (n2008) );
  buffer buf_n2009( .i (n2008), .o (n2009) );
  buffer buf_n2010( .i (n2009), .o (n2010) );
  assign n2014 = n420 & n1097 ;
  assign n2015 = G93 & ~n420 ;
  assign n2016 = n2014 | n2015 ;
  buffer buf_n2017( .i (n2016), .o (n2017) );
  assign n2044 = n795 & n2017 ;
  buffer buf_n2045( .i (n2044), .o (n2045) );
  assign n2049 = n795 | n2017 ;
  buffer buf_n2050( .i (n2049), .o (n2050) );
  assign n2052 = ~n2045 & n2050 ;
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  assign n2073 = n421 & n1125 ;
  assign n2074 = G95 & ~n421 ;
  assign n2075 = n2073 | n2074 ;
  buffer buf_n2076( .i (n2075), .o (n2076) );
  assign n2099 = n722 & n2076 ;
  buffer buf_n2100( .i (n2099), .o (n2100) );
  assign n2118 = n722 | n2076 ;
  buffer buf_n2119( .i (n2118), .o (n2119) );
  assign n2137 = ~n2100 & n2119 ;
  buffer buf_n2138( .i (n2137), .o (n2138) );
  assign n2157 = n2054 & n2138 ;
  buffer buf_n2158( .i (n2157), .o (n2158) );
  buffer buf_n2159( .i (n2158), .o (n2159) );
  buffer buf_n2160( .i (n2159), .o (n2160) );
  buffer buf_n2161( .i (n2160), .o (n2161) );
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n2163( .i (n2162), .o (n2163) );
  buffer buf_n2164( .i (n2163), .o (n2164) );
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n2166( .i (n2165), .o (n2166) );
  buffer buf_n2167( .i (n2166), .o (n2167) );
  buffer buf_n2168( .i (n2167), .o (n2168) );
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  buffer buf_n2171( .i (n2170), .o (n2171) );
  assign n2172 = n2010 & n2171 ;
  buffer buf_n2173( .i (n2172), .o (n2173) );
  assign n2174 = n1936 & n2173 ;
  buffer buf_n2175( .i (n2174), .o (n2175) );
  assign n2176 = n1854 & n2175 ;
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n2177), .o (n2178) );
  buffer buf_n2179( .i (n2178), .o (n2179) );
  buffer buf_n2180( .i (n2179), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  buffer buf_n2182( .i (n2181), .o (n2182) );
  buffer buf_n2183( .i (n2182), .o (n2183) );
  buffer buf_n2184( .i (n2183), .o (n2184) );
  buffer buf_n2185( .i (n2184), .o (n2185) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  buffer buf_n2187( .i (n2186), .o (n2187) );
  buffer buf_n398( .i (G123), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  assign n2188 = n403 | n444 ;
  buffer buf_n2189( .i (n2188), .o (n2189) );
  assign n2204 = n839 & n2189 ;
  buffer buf_n2205( .i (n2204), .o (n2205) );
  assign n2214 = n839 | n2189 ;
  buffer buf_n2215( .i (n2214), .o (n2215) );
  assign n2224 = ~n2205 & n2215 ;
  buffer buf_n2225( .i (n2224), .o (n2225) );
  assign n2235 = n398 & n530 ;
  assign n2236 = ~n398 & n553 ;
  assign n2237 = n2235 | n2236 ;
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  assign n2257 = n872 | n2240 ;
  buffer buf_n2258( .i (n2257), .o (n2258) );
  assign n2273 = n400 & n589 ;
  assign n2274 = ~n400 & n607 ;
  assign n2275 = n2273 | n2274 ;
  buffer buf_n2276( .i (n2275), .o (n2276) );
  assign n2296 = n870 & n2238 ;
  buffer buf_n2297( .i (n2296), .o (n2297) );
  assign n2314 = n2276 | n2297 ;
  buffer buf_n2315( .i (n2314), .o (n2315) );
  assign n2320 = n2258 & ~n2315 ;
  buffer buf_n2321( .i (n2320), .o (n2321) );
  assign n2336 = n400 & n475 ;
  buffer buf_n2337( .i (n399), .o (n2337) );
  assign n2338 = n496 & ~n2337 ;
  assign n2339 = n2336 | n2338 ;
  buffer buf_n2340( .i (n2339), .o (n2340) );
  assign n2357 = n852 & n2340 ;
  buffer buf_n2358( .i (n2357), .o (n2358) );
  assign n2361 = n852 | n2340 ;
  buffer buf_n2362( .i (n2361), .o (n2362) );
  assign n2364 = ~n2358 & n2362 ;
  buffer buf_n2365( .i (n2364), .o (n2365) );
  assign n2379 = n2321 & n2365 ;
  buffer buf_n2380( .i (n2379), .o (n2380) );
  assign n2385 = n2225 & n2380 ;
  buffer buf_n2386( .i (n2385), .o (n2386) );
  buffer buf_n2387( .i (n2386), .o (n2387) );
  buffer buf_n2388( .i (n2387), .o (n2388) );
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2391( .i (n2390), .o (n2391) );
  buffer buf_n2392( .i (n2391), .o (n2392) );
  buffer buf_n2393( .i (n2392), .o (n2393) );
  buffer buf_n2394( .i (n2393), .o (n2394) );
  buffer buf_n2395( .i (n2394), .o (n2395) );
  buffer buf_n2396( .i (n2395), .o (n2396) );
  buffer buf_n2397( .i (n2396), .o (n2397) );
  buffer buf_n2398( .i (n2397), .o (n2398) );
  buffer buf_n2399( .i (n2398), .o (n2399) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  assign n2400 = n349 & n407 ;
  assign n2401 = G118 & ~n407 ;
  assign n2402 = n2400 | n2401 ;
  buffer buf_n2403( .i (n2402), .o (n2403) );
  buffer buf_n2404( .i (n2403), .o (n2404) );
  assign n2407 = n819 & n2404 ;
  buffer buf_n2408( .i (n2407), .o (n2408) );
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n2405( .i (n2404), .o (n2405) );
  assign n2414 = n820 | n2405 ;
  buffer buf_n2415( .i (n2414), .o (n2415) );
  assign n2419 = ~n2409 & n2415 ;
  buffer buf_n2420( .i (n2419), .o (n2420) );
  assign n2425 = n363 & n405 ;
  assign n2426 = G120 & ~n405 ;
  assign n2427 = n2425 | n2426 ;
  buffer buf_n2428( .i (n2427), .o (n2428) );
  assign n2443 = n821 & n2428 ;
  buffer buf_n2444( .i (n2443), .o (n2444) );
  assign n2452 = n821 | n2428 ;
  buffer buf_n2453( .i (n2452), .o (n2453) );
  assign n2461 = ~n2444 & n2453 ;
  buffer buf_n2462( .i (n2461), .o (n2462) );
  buffer buf_n2463( .i (n2462), .o (n2463) );
  buffer buf_n2464( .i (n2463), .o (n2464) );
  buffer buf_n2465( .i (n2464), .o (n2465) );
  buffer buf_n2466( .i (n2465), .o (n2466) );
  assign n2471 = n2420 & n2466 ;
  buffer buf_n2472( .i (n2471), .o (n2472) );
  buffer buf_n2473( .i (n2472), .o (n2473) );
  buffer buf_n2474( .i (n2473), .o (n2474) );
  buffer buf_n2475( .i (n2474), .o (n2475) );
  buffer buf_n2476( .i (n2475), .o (n2476) );
  buffer buf_n2477( .i (n2476), .o (n2477) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  assign n2478 = n288 & n409 ;
  assign n2479 = n313 & ~n409 ;
  assign n2480 = n2478 | n2479 ;
  buffer buf_n2481( .i (n2480), .o (n2481) );
  buffer buf_n2482( .i (n2481), .o (n2482) );
  buffer buf_n2483( .i (n2482), .o (n2483) );
  buffer buf_n2484( .i (n2483), .o (n2484) );
  buffer buf_n2485( .i (n2484), .o (n2485) );
  buffer buf_n2486( .i (n2485), .o (n2486) );
  buffer buf_n2487( .i (n2486), .o (n2487) );
  buffer buf_n2488( .i (n2487), .o (n2488) );
  buffer buf_n2489( .i (n2488), .o (n2489) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  assign n2496 = n345 & n417 ;
  assign n2497 = G116 & ~n417 ;
  assign n2498 = n2496 | n2497 ;
  buffer buf_n2499( .i (n2498), .o (n2499) );
  assign n2502 = n2489 | n2499 ;
  buffer buf_n2503( .i (n2502), .o (n2503) );
  assign n2504 = G122 | n401 ;
  buffer buf_n2505( .i (n2504), .o (n2505) );
  assign n2522 = ~n379 & n402 ;
  assign n2523 = n2505 & ~n2522 ;
  buffer buf_n2524( .i (n2523), .o (n2524) );
  assign n2539 = n824 & n2524 ;
  buffer buf_n2540( .i (n2539), .o (n2540) );
  assign n2548 = n824 | n2524 ;
  buffer buf_n2549( .i (n2548), .o (n2549) );
  assign n2556 = ~n2540 & n2549 ;
  buffer buf_n2557( .i (n2556), .o (n2557) );
  buffer buf_n2558( .i (n2557), .o (n2558) );
  buffer buf_n2559( .i (n2558), .o (n2559) );
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  buffer buf_n2563( .i (n2562), .o (n2563) );
  buffer buf_n2564( .i (n2563), .o (n2564) );
  buffer buf_n2565( .i (n2564), .o (n2565) );
  buffer buf_n2566( .i (n2565), .o (n2566) );
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n2568( .i (n2567), .o (n2568) );
  buffer buf_n2569( .i (n2568), .o (n2569) );
  buffer buf_n2570( .i (n2569), .o (n2570) );
  assign n2571 = ~n2503 & n2570 ;
  assign n2572 = n2477 & n2571 ;
  assign n2573 = n2399 & n2572 ;
  buffer buf_n2574( .i (n2573), .o (n2574) );
  buffer buf_n2575( .i (n2574), .o (n2575) );
  buffer buf_n2576( .i (n2575), .o (n2576) );
  buffer buf_n2577( .i (n2576), .o (n2577) );
  buffer buf_n2578( .i (n2577), .o (n2578) );
  buffer buf_n2579( .i (n2578), .o (n2579) );
  buffer buf_n2580( .i (n2579), .o (n2580) );
  buffer buf_n2581( .i (n2580), .o (n2581) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  assign n2582 = n299 | n348 ;
  assign n2583 = n299 & n348 ;
  assign n2584 = n2582 & ~n2583 ;
  buffer buf_n2585( .i (n2584), .o (n2585) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  assign n2586 = n362 & ~n378 ;
  assign n2587 = ~n362 & n378 ;
  assign n2588 = n2586 | n2587 ;
  buffer buf_n2589( .i (n2588), .o (n2589) );
  assign n2590 = ~n2585 & n2589 ;
  assign n2591 = n2585 & ~n2589 ;
  assign n2592 = n2590 | n2591 ;
  buffer buf_n2593( .i (n2592), .o (n2593) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n641( .i (G132), .o (n641) );
  assign n2594 = n606 & ~n641 ;
  assign n2595 = ~n606 & n641 ;
  assign n2596 = n2594 | n2595 ;
  buffer buf_n2597( .i (n2596), .o (n2597) );
  assign n2598 = n397 & ~n2597 ;
  assign n2599 = ~n397 & n2597 ;
  assign n2600 = n2598 | n2599 ;
  buffer buf_n2601( .i (n2600), .o (n2601) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  assign n2602 = n495 & ~n552 ;
  assign n2603 = ~n495 & n552 ;
  assign n2604 = n2602 | n2603 ;
  buffer buf_n2605( .i (n2604), .o (n2605) );
  assign n2606 = n2601 & ~n2605 ;
  assign n2607 = ~n2601 & n2605 ;
  assign n2608 = n2606 | n2607 ;
  buffer buf_n2609( .i (n2608), .o (n2609) );
  assign n2610 = n2593 | n2609 ;
  assign n2611 = n2593 & n2609 ;
  assign n2612 = n2610 & ~n2611 ;
  buffer buf_n2613( .i (n2612), .o (n2613) );
  buffer buf_n2614( .i (n2613), .o (n2614) );
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  inverter inv_n2617( .i (n2616), .o (n2617) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n1095( .i (n1094), .o (n1095) );
  buffer buf_n1096( .i (n1095), .o (n1096) );
  assign n2618 = n1071 | n1096 ;
  assign n2619 = n1071 & n1096 ;
  assign n2620 = n2618 & ~n2619 ;
  buffer buf_n2621( .i (n2620), .o (n2621) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  assign n2622 = n1124 & ~n1151 ;
  assign n2623 = ~n1124 & n1151 ;
  assign n2624 = n2622 | n2623 ;
  buffer buf_n2625( .i (n2624), .o (n2625) );
  assign n2626 = ~n2621 & n2625 ;
  assign n2627 = n2621 & ~n2625 ;
  assign n2628 = n2626 | n2627 ;
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n210), .o (n2630) );
  buffer buf_n2631( .i (n1169), .o (n2631) );
  assign n2632 = n2630 | n2631 ;
  assign n2633 = n2630 & n2631 ;
  assign n2634 = n2632 & ~n2633 ;
  buffer buf_n2635( .i (n2634), .o (n2635) );
  buffer buf_n286( .i (G111), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n2636( .i (n278), .o (n2636) );
  assign n2637 = ~n287 & n2636 ;
  assign n2638 = n287 & ~n2636 ;
  assign n2639 = n2637 | n2638 ;
  buffer buf_n2640( .i (n2639), .o (n2640) );
  assign n2641 = n2635 | n2640 ;
  assign n2642 = n2635 & n2640 ;
  assign n2643 = n2641 & ~n2642 ;
  buffer buf_n2644( .i (n2643), .o (n2644) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  assign n2645 = n234 & ~n258 ;
  assign n2646 = ~n234 & n258 ;
  assign n2647 = n2645 | n2646 ;
  buffer buf_n2648( .i (n2647), .o (n2648) );
  assign n2649 = n2644 & ~n2648 ;
  assign n2650 = ~n2644 & n2648 ;
  assign n2651 = n2649 | n2650 ;
  buffer buf_n2652( .i (n2651), .o (n2652) );
  assign n2653 = n2629 & n2652 ;
  assign n2654 = n2629 | n2652 ;
  assign n2655 = ~n2653 & n2654 ;
  buffer buf_n2656( .i (n2655), .o (n2656) );
  buffer buf_n2657( .i (n2656), .o (n2657) );
  buffer buf_n2658( .i (n2657), .o (n2658) );
  inverter inv_n2659( .i (n2658), .o (n2659) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  assign n2660 = n1606 & n1675 ;
  buffer buf_n2661( .i (n2660), .o (n2661) );
  assign n2667 = n1686 | n1748 ;
  assign n2668 = n2661 | n2667 ;
  assign n2669 = n1752 & n2668 ;
  buffer buf_n2670( .i (n2669), .o (n2670) );
  assign n2681 = n1571 & n1809 ;
  assign n2682 = n2670 & n2681 ;
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  assign n2683 = n1569 & n1804 ;
  assign n2684 = n1565 | n2683 ;
  assign n2685 = n2682 | n2684 ;
  buffer buf_n2686( .i (n2685), .o (n2686) );
  buffer buf_n2687( .i (n2686), .o (n2687) );
  buffer buf_n2688( .i (n2687), .o (n2688) );
  buffer buf_n2689( .i (n2688), .o (n2689) );
  buffer buf_n2690( .i (n2689), .o (n2690) );
  buffer buf_n2691( .i (n2690), .o (n2691) );
  buffer buf_n2692( .i (n2691), .o (n2692) );
  buffer buf_n2693( .i (n2692), .o (n2693) );
  buffer buf_n2694( .i (n2693), .o (n2694) );
  buffer buf_n2695( .i (n2694), .o (n2695) );
  buffer buf_n2696( .i (n2695), .o (n2696) );
  assign n2697 = n2175 & n2696 ;
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  buffer buf_n1888( .i (n1887), .o (n1888) );
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1907( .i (n1906), .o (n1907) );
  buffer buf_n1908( .i (n1907), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n1915( .i (n1914), .o (n1915) );
  buffer buf_n1916( .i (n1915), .o (n1916) );
  buffer buf_n1917( .i (n1916), .o (n1917) );
  buffer buf_n1918( .i (n1917), .o (n1918) );
  buffer buf_n1919( .i (n1918), .o (n1919) );
  buffer buf_n1970( .i (n1969), .o (n1970) );
  buffer buf_n1971( .i (n1970), .o (n1971) );
  buffer buf_n1972( .i (n1971), .o (n1972) );
  buffer buf_n1973( .i (n1972), .o (n1973) );
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  buffer buf_n1983( .i (n1982), .o (n1983) );
  buffer buf_n1984( .i (n1983), .o (n1984) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n1988( .i (n1987), .o (n1988) );
  buffer buf_n1989( .i (n1988), .o (n1989) );
  buffer buf_n1990( .i (n1989), .o (n1990) );
  buffer buf_n1991( .i (n1990), .o (n1991) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  assign n2698 = n2051 & n2100 ;
  buffer buf_n2699( .i (n2698), .o (n2699) );
  assign n2705 = n2048 | n2699 ;
  buffer buf_n2706( .i (n2705), .o (n2706) );
  buffer buf_n2707( .i (n2706), .o (n2707) );
  buffer buf_n2708( .i (n2707), .o (n2708) );
  assign n2721 = n1991 & n2708 ;
  buffer buf_n2722( .i (n2721), .o (n2722) );
  buffer buf_n2723( .i (n2722), .o (n2723) );
  buffer buf_n2724( .i (n2723), .o (n2724) );
  buffer buf_n2725( .i (n2724), .o (n2725) );
  buffer buf_n2726( .i (n2725), .o (n2726) );
  buffer buf_n2727( .i (n2726), .o (n2727) );
  buffer buf_n2728( .i (n2727), .o (n2728) );
  buffer buf_n2729( .i (n2728), .o (n2729) );
  buffer buf_n2730( .i (n2729), .o (n2730) );
  buffer buf_n2731( .i (n2730), .o (n2731) );
  buffer buf_n2732( .i (n2731), .o (n2732) );
  assign n2733 = n1985 | n2732 ;
  buffer buf_n2734( .i (n2733), .o (n2734) );
  assign n2735 = n1919 & n2734 ;
  assign n2736 = n1899 | n2735 ;
  assign n2737 = n2697 | n2736 ;
  buffer buf_n2738( .i (n2737), .o (n2738) );
  buffer buf_n2739( .i (n2738), .o (n2739) );
  buffer buf_n2740( .i (n2739), .o (n2740) );
  buffer buf_n2741( .i (n2740), .o (n2741) );
  buffer buf_n2742( .i (n2741), .o (n2742) );
  buffer buf_n2743( .i (n2742), .o (n2743) );
  buffer buf_n2744( .i (n2743), .o (n2744) );
  buffer buf_n2745( .i (n2744), .o (n2745) );
  buffer buf_n2746( .i (n2745), .o (n2746) );
  buffer buf_n2747( .i (n2746), .o (n2747) );
  assign n2748 = ~n2489 & n2499 ;
  buffer buf_n2749( .i (n2748), .o (n2749) );
  buffer buf_n2750( .i (n2749), .o (n2750) );
  buffer buf_n2751( .i (n2750), .o (n2751) );
  buffer buf_n2752( .i (n2751), .o (n2752) );
  buffer buf_n2753( .i (n2752), .o (n2753) );
  buffer buf_n2754( .i (n2753), .o (n2754) );
  buffer buf_n2755( .i (n2754), .o (n2755) );
  buffer buf_n2756( .i (n2755), .o (n2756) );
  buffer buf_n2757( .i (n2756), .o (n2757) );
  buffer buf_n2758( .i (n2757), .o (n2758) );
  buffer buf_n2759( .i (n2758), .o (n2759) );
  inverter inv_n2760( .i (n2759), .o (n2760) );
  buffer buf_n976( .i (G176), .o (n976) );
  buffer buf_n982( .i (G177), .o (n982) );
  assign n2761 = n976 & ~n982 ;
  buffer buf_n2762( .i (n2761), .o (n2762) );
  buffer buf_n2763( .i (n2762), .o (n2763) );
  buffer buf_n2764( .i (n2763), .o (n2764) );
  buffer buf_n2765( .i (n2764), .o (n2765) );
  assign n2772 = G60 & n2765 ;
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n999( .i (G21), .o (n999) );
  buffer buf_n2277( .i (n2276), .o (n2277) );
  buffer buf_n2278( .i (n2277), .o (n2278) );
  buffer buf_n2279( .i (n2278), .o (n2279) );
  buffer buf_n2280( .i (n2279), .o (n2280) );
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n2289( .i (n2288), .o (n2289) );
  buffer buf_n2290( .i (n2289), .o (n2290) );
  buffer buf_n2291( .i (n2290), .o (n2291) );
  buffer buf_n2292( .i (n2291), .o (n2292) );
  buffer buf_n2293( .i (n2292), .o (n2293) );
  buffer buf_n2294( .i (n2293), .o (n2294) );
  assign n2773 = ~n999 & n2294 ;
  assign n2774 = n999 & ~n2294 ;
  assign n2775 = n2773 | n2774 ;
  buffer buf_n2776( .i (n2775), .o (n2776) );
  assign n2777 = ~n980 & n2776 ;
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  assign n2778 = n979 & ~n1361 ;
  assign n2779 = n986 & ~n2778 ;
  assign n2780 = ~n2777 & n2779 ;
  assign n2781 = n2772 | n2780 ;
  buffer buf_n2782( .i (n2781), .o (n2782) );
  buffer buf_n2783( .i (n2782), .o (n2783) );
  buffer buf_n2784( .i (n2783), .o (n2784) );
  buffer buf_n2785( .i (n2784), .o (n2785) );
  buffer buf_n2786( .i (n2785), .o (n2786) );
  inverter inv_n2787( .i (n2786), .o (n2787) );
  assign n2788 = G58 & n2764 ;
  buffer buf_n2322( .i (n2321), .o (n2322) );
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2325( .i (n2324), .o (n2325) );
  buffer buf_n2326( .i (n2325), .o (n2326) );
  buffer buf_n2327( .i (n2326), .o (n2327) );
  buffer buf_n2328( .i (n2327), .o (n2328) );
  buffer buf_n2329( .i (n2328), .o (n2329) );
  buffer buf_n2330( .i (n2329), .o (n2330) );
  buffer buf_n2331( .i (n2330), .o (n2331) );
  buffer buf_n2332( .i (n2331), .o (n2332) );
  buffer buf_n2333( .i (n2332), .o (n2333) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n2335( .i (n2334), .o (n2335) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  buffer buf_n2265( .i (n2264), .o (n2265) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  buffer buf_n2269( .i (n2268), .o (n2269) );
  buffer buf_n2270( .i (n2269), .o (n2270) );
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  buffer buf_n2307( .i (n2306), .o (n2307) );
  buffer buf_n2308( .i (n2307), .o (n2308) );
  buffer buf_n2309( .i (n2308), .o (n2309) );
  buffer buf_n2310( .i (n2309), .o (n2310) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  assign n2789 = n2272 & ~n2313 ;
  assign n2790 = n2293 & ~n2789 ;
  assign n2791 = n2335 | n2790 ;
  buffer buf_n2792( .i (n2791), .o (n2792) );
  assign n2795 = n979 | n2792 ;
  assign n2796 = n978 & n1304 ;
  assign n2797 = n985 & ~n2796 ;
  assign n2798 = n2795 & n2797 ;
  assign n2799 = n2788 | n2798 ;
  buffer buf_n2800( .i (n2799), .o (n2800) );
  buffer buf_n2801( .i (n2800), .o (n2801) );
  buffer buf_n2802( .i (n2801), .o (n2802) );
  buffer buf_n2803( .i (n2802), .o (n2803) );
  buffer buf_n2804( .i (n2803), .o (n2804) );
  buffer buf_n2805( .i (n2804), .o (n2805) );
  inverter inv_n2806( .i (n2805), .o (n2806) );
  assign n2807 = G48 & n2765 ;
  buffer buf_n990( .i (G2), .o (n990) );
  buffer buf_n1633( .i (n1632), .o (n1633) );
  buffer buf_n1634( .i (n1633), .o (n1634) );
  buffer buf_n1635( .i (n1634), .o (n1635) );
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n1637( .i (n1636), .o (n1637) );
  buffer buf_n1638( .i (n1637), .o (n1638) );
  assign n2808 = n990 & n1638 ;
  buffer buf_n2809( .i (n2808), .o (n2809) );
  buffer buf_n2810( .i (n2809), .o (n2810) );
  buffer buf_n2811( .i (n2810), .o (n2811) );
  buffer buf_n2812( .i (n2811), .o (n2812) );
  buffer buf_n2813( .i (n2812), .o (n2813) );
  buffer buf_n2814( .i (n2813), .o (n2814) );
  buffer buf_n2815( .i (n2814), .o (n2815) );
  buffer buf_n2816( .i (n2815), .o (n2816) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  assign n2817 = n998 | n1646 ;
  assign n2818 = ~n2816 & n2817 ;
  buffer buf_n2819( .i (n2818), .o (n2819) );
  assign n2820 = n980 | n2819 ;
  assign n2821 = n979 & n1457 ;
  assign n2822 = n986 & ~n2821 ;
  assign n2823 = n2820 & n2822 ;
  assign n2824 = n2807 | n2823 ;
  buffer buf_n2825( .i (n2824), .o (n2825) );
  buffer buf_n2826( .i (n2825), .o (n2826) );
  buffer buf_n2827( .i (n2826), .o (n2827) );
  buffer buf_n2828( .i (n2827), .o (n2828) );
  buffer buf_n2829( .i (n2828), .o (n2829) );
  inverter inv_n2830( .i (n2829), .o (n2830) );
  buffer buf_n2490( .i (n2489), .o (n2490) );
  buffer buf_n2500( .i (n2499), .o (n2500) );
  assign n2831 = n2490 & n2500 ;
  assign n2832 = n2503 & ~n2831 ;
  buffer buf_n2833( .i (n2832), .o (n2833) );
  buffer buf_n2834( .i (n2833), .o (n2834) );
  buffer buf_n2835( .i (n2834), .o (n2835) );
  buffer buf_n2836( .i (n2835), .o (n2836) );
  buffer buf_n2837( .i (n2836), .o (n2837) );
  buffer buf_n2838( .i (n2837), .o (n2838) );
  buffer buf_n2839( .i (n2838), .o (n2839) );
  buffer buf_n2840( .i (n2839), .o (n2840) );
  buffer buf_n2841( .i (n2840), .o (n2841) );
  buffer buf_n2842( .i (n2841), .o (n2842) );
  buffer buf_n964( .i (G173), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  assign n2843 = n967 | n2827 ;
  buffer buf_n960( .i (G172), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  assign n2844 = n966 & ~n2783 ;
  assign n2845 = n963 & ~n2844 ;
  assign n2846 = n2843 & n2845 ;
  buffer buf_n1006( .i (G3), .o (n1006) );
  assign n2847 = ~n960 & n964 ;
  buffer buf_n2848( .i (n2847), .o (n2848) );
  buffer buf_n2849( .i (n2848), .o (n2849) );
  assign n2850 = n1006 & n2849 ;
  buffer buf_n1000( .i (G22), .o (n1000) );
  assign n2851 = n960 | n964 ;
  buffer buf_n2852( .i (n2851), .o (n2852) );
  buffer buf_n2853( .i (n2852), .o (n2853) );
  assign n2854 = n1000 & ~n2853 ;
  assign n2855 = n2850 | n2854 ;
  assign n2856 = n2846 | n2855 ;
  assign n2857 = G19 & n2764 ;
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2206( .i (n2205), .o (n2206) );
  buffer buf_n2207( .i (n2206), .o (n2207) );
  buffer buf_n2359( .i (n2358), .o (n2359) );
  buffer buf_n2360( .i (n2359), .o (n2360) );
  buffer buf_n2363( .i (n2362), .o (n2363) );
  assign n2858 = n2300 & n2363 ;
  assign n2859 = n2360 | n2858 ;
  buffer buf_n2860( .i (n2859), .o (n2860) );
  assign n2865 = n2207 | n2860 ;
  assign n2866 = n2218 & n2865 ;
  assign n2867 = n2386 | n2866 ;
  buffer buf_n2868( .i (n2867), .o (n2868) );
  buffer buf_n2869( .i (n2868), .o (n2869) );
  buffer buf_n2870( .i (n2869), .o (n2870) );
  buffer buf_n2871( .i (n2870), .o (n2871) );
  buffer buf_n2872( .i (n2871), .o (n2872) );
  buffer buf_n2873( .i (n2872), .o (n2873) );
  buffer buf_n2874( .i (n2873), .o (n2874) );
  buffer buf_n2875( .i (n2874), .o (n2875) );
  assign n2876 = n2568 | n2875 ;
  assign n2877 = n2568 & n2875 ;
  assign n2878 = n2876 & ~n2877 ;
  buffer buf_n2879( .i (n2878), .o (n2879) );
  buffer buf_n2885( .i (n978), .o (n2885) );
  assign n2886 = n2879 & ~n2885 ;
  assign n2887 = n978 & n1379 ;
  assign n2888 = n985 & ~n2887 ;
  assign n2889 = ~n2886 & n2888 ;
  assign n2890 = n2857 | n2889 ;
  buffer buf_n2891( .i (n2890), .o (n2891) );
  buffer buf_n2892( .i (n2891), .o (n2892) );
  buffer buf_n2893( .i (n2892), .o (n2893) );
  buffer buf_n2894( .i (n2893), .o (n2894) );
  buffer buf_n2895( .i (n2894), .o (n2895) );
  buffer buf_n2896( .i (n2895), .o (n2896) );
  inverter inv_n2897( .i (n2896), .o (n2897) );
  assign n2898 = G59 & n2762 ;
  buffer buf_n2226( .i (n2225), .o (n2226) );
  buffer buf_n2227( .i (n2226), .o (n2227) );
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  buffer buf_n2231( .i (n2230), .o (n2231) );
  buffer buf_n2232( .i (n2231), .o (n2232) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  buffer buf_n2381( .i (n2380), .o (n2381) );
  buffer buf_n2382( .i (n2381), .o (n2382) );
  buffer buf_n2383( .i (n2382), .o (n2383) );
  buffer buf_n2384( .i (n2383), .o (n2384) );
  buffer buf_n2861( .i (n2860), .o (n2861) );
  buffer buf_n2862( .i (n2861), .o (n2862) );
  buffer buf_n2863( .i (n2862), .o (n2863) );
  buffer buf_n2864( .i (n2863), .o (n2864) );
  assign n2899 = n2384 | n2864 ;
  buffer buf_n2900( .i (n2899), .o (n2900) );
  buffer buf_n2901( .i (n2900), .o (n2901) );
  buffer buf_n2902( .i (n2901), .o (n2902) );
  buffer buf_n2903( .i (n2902), .o (n2903) );
  assign n2904 = ~n2234 & n2903 ;
  assign n2905 = n2234 & ~n2903 ;
  assign n2906 = n2904 | n2905 ;
  buffer buf_n2907( .i (n2906), .o (n2907) );
  assign n2914 = ~n977 & n2907 ;
  assign n2915 = n976 & n1365 ;
  assign n2916 = n983 & ~n2915 ;
  assign n2917 = ~n2914 & n2916 ;
  assign n2918 = n2898 | n2917 ;
  buffer buf_n2919( .i (n2918), .o (n2919) );
  buffer buf_n2920( .i (n2919), .o (n2920) );
  buffer buf_n2921( .i (n2920), .o (n2921) );
  buffer buf_n2922( .i (n2921), .o (n2922) );
  buffer buf_n2923( .i (n2922), .o (n2923) );
  buffer buf_n2924( .i (n2923), .o (n2924) );
  buffer buf_n2925( .i (n2924), .o (n2925) );
  buffer buf_n2926( .i (n2925), .o (n2926) );
  inverter inv_n2927( .i (n2926), .o (n2927) );
  assign n2928 = G50 & n2764 ;
  buffer buf_n2366( .i (n2365), .o (n2366) );
  buffer buf_n2367( .i (n2366), .o (n2367) );
  buffer buf_n2368( .i (n2367), .o (n2368) );
  buffer buf_n2369( .i (n2368), .o (n2369) );
  buffer buf_n2370( .i (n2369), .o (n2370) );
  buffer buf_n2371( .i (n2370), .o (n2371) );
  buffer buf_n2372( .i (n2371), .o (n2372) );
  buffer buf_n2373( .i (n2372), .o (n2373) );
  buffer buf_n2374( .i (n2373), .o (n2374) );
  buffer buf_n2375( .i (n2374), .o (n2375) );
  buffer buf_n2376( .i (n2375), .o (n2376) );
  buffer buf_n2377( .i (n2376), .o (n2377) );
  buffer buf_n2378( .i (n2377), .o (n2378) );
  assign n2929 = n2312 | n2332 ;
  buffer buf_n2930( .i (n2929), .o (n2930) );
  assign n2931 = n2378 | n2930 ;
  assign n2932 = n2378 & n2930 ;
  assign n2933 = n2931 & ~n2932 ;
  buffer buf_n2934( .i (n2933), .o (n2934) );
  assign n2938 = ~n2885 & n2934 ;
  buffer buf_n2939( .i (n977), .o (n2939) );
  assign n2940 = n1392 & n2939 ;
  assign n2941 = n985 & ~n2940 ;
  assign n2942 = ~n2938 & n2941 ;
  assign n2943 = n2928 | n2942 ;
  buffer buf_n2944( .i (n2943), .o (n2944) );
  buffer buf_n2945( .i (n2944), .o (n2945) );
  buffer buf_n2946( .i (n2945), .o (n2946) );
  buffer buf_n2947( .i (n2946), .o (n2947) );
  buffer buf_n2948( .i (n2947), .o (n2948) );
  buffer buf_n2949( .i (n2948), .o (n2949) );
  inverter inv_n2950( .i (n2949), .o (n2950) );
  buffer buf_n968( .i (G174), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  assign n2951 = n971 | n2827 ;
  buffer buf_n972( .i (G175), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  assign n2952 = n970 & ~n2783 ;
  assign n2953 = n975 & ~n2952 ;
  assign n2954 = n2951 & n2953 ;
  assign n2955 = n968 & ~n972 ;
  buffer buf_n2956( .i (n2955), .o (n2956) );
  buffer buf_n2957( .i (n2956), .o (n2957) );
  assign n2958 = n1006 & n2957 ;
  assign n2959 = n968 | n972 ;
  buffer buf_n2960( .i (n2959), .o (n2960) );
  buffer buf_n2961( .i (n2960), .o (n2961) );
  assign n2962 = n1000 & ~n2961 ;
  assign n2963 = n2958 | n2962 ;
  assign n2964 = n2954 | n2963 ;
  assign n2965 = G53 & n2765 ;
  assign n2966 = n990 & n1846 ;
  buffer buf_n2967( .i (n2966), .o (n2967) );
  buffer buf_n2968( .i (n2967), .o (n2968) );
  buffer buf_n2969( .i (n2968), .o (n2969) );
  buffer buf_n2970( .i (n2969), .o (n2970) );
  buffer buf_n2971( .i (n2970), .o (n2971) );
  buffer buf_n2972( .i (n2971), .o (n2972) );
  buffer buf_n2973( .i (n2972), .o (n2973) );
  buffer buf_n2974( .i (n2973), .o (n2974) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  assign n2975 = n997 & n1844 ;
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n2671( .i (n2670), .o (n2671) );
  assign n2976 = n1800 & n2671 ;
  assign n2977 = n1807 | n2976 ;
  buffer buf_n2978( .i (n2977), .o (n2978) );
  buffer buf_n2979( .i (n2978), .o (n2979) );
  buffer buf_n2980( .i (n2979), .o (n2980) );
  assign n2981 = ~n1578 & n2980 ;
  assign n2982 = n1578 & ~n2980 ;
  assign n2983 = n2981 | n2982 ;
  buffer buf_n2984( .i (n2983), .o (n2984) );
  buffer buf_n2985( .i (n2984), .o (n2985) );
  buffer buf_n2986( .i (n2985), .o (n2986) );
  buffer buf_n2987( .i (n2986), .o (n2987) );
  buffer buf_n2988( .i (n2987), .o (n2988) );
  assign n2989 = n2975 | n2988 ;
  assign n2990 = ~n2974 & n2989 ;
  buffer buf_n2991( .i (n2990), .o (n2991) );
  assign n2995 = ~n980 & n2991 ;
  assign n2996 = n1468 & n2885 ;
  assign n2997 = n986 & ~n2996 ;
  assign n2998 = ~n2995 & n2997 ;
  assign n2999 = n2965 | n2998 ;
  buffer buf_n3000( .i (n2999), .o (n3000) );
  buffer buf_n3001( .i (n3000), .o (n3001) );
  buffer buf_n3002( .i (n3001), .o (n3002) );
  buffer buf_n3003( .i (n3002), .o (n3003) );
  buffer buf_n3004( .i (n3003), .o (n3004) );
  inverter inv_n3005( .i (n3004), .o (n3005) );
  buffer buf_n3006( .i (n2763), .o (n3006) );
  buffer buf_n3007( .i (n3006), .o (n3007) );
  assign n3008 = G57 & n3007 ;
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  buffer buf_n1813( .i (n1812), .o (n1813) );
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  buffer buf_n1821( .i (n1820), .o (n1821) );
  buffer buf_n1822( .i (n1821), .o (n1822) );
  buffer buf_n1823( .i (n1822), .o (n1823) );
  buffer buf_n2672( .i (n2671), .o (n2672) );
  buffer buf_n2673( .i (n2672), .o (n2673) );
  buffer buf_n2674( .i (n2673), .o (n2674) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  assign n3009 = n1721 & n1759 ;
  assign n3010 = n2674 | n3009 ;
  buffer buf_n3011( .i (n3010), .o (n3011) );
  buffer buf_n3012( .i (n3011), .o (n3012) );
  buffer buf_n3013( .i (n3012), .o (n3013) );
  buffer buf_n3014( .i (n3013), .o (n3014) );
  buffer buf_n3015( .i (n3014), .o (n3015) );
  buffer buf_n3016( .i (n3015), .o (n3016) );
  buffer buf_n2675( .i (n2674), .o (n2675) );
  buffer buf_n2676( .i (n2675), .o (n2676) );
  buffer buf_n2677( .i (n2676), .o (n2677) );
  buffer buf_n2678( .i (n2677), .o (n2678) );
  buffer buf_n2679( .i (n2678), .o (n2679) );
  buffer buf_n2680( .i (n2679), .o (n2680) );
  assign n3017 = n995 | n2680 ;
  assign n3018 = n3016 & n3017 ;
  buffer buf_n3019( .i (n3018), .o (n3019) );
  assign n3020 = ~n1823 & n3019 ;
  assign n3021 = n1823 & ~n3019 ;
  assign n3022 = n3020 | n3021 ;
  buffer buf_n3023( .i (n3022), .o (n3023) );
  buffer buf_n3025( .i (n2885), .o (n3025) );
  assign n3026 = n3023 & ~n3025 ;
  buffer buf_n3027( .i (n2939), .o (n3027) );
  assign n3028 = n1512 & n3027 ;
  buffer buf_n3029( .i (n984), .o (n3029) );
  buffer buf_n3030( .i (n3029), .o (n3030) );
  assign n3031 = ~n3028 & n3030 ;
  assign n3032 = ~n3026 & n3031 ;
  assign n3033 = n3008 | n3032 ;
  buffer buf_n3034( .i (n3033), .o (n3034) );
  buffer buf_n3035( .i (n3034), .o (n3035) );
  buffer buf_n3036( .i (n3035), .o (n3036) );
  buffer buf_n3037( .i (n3036), .o (n3037) );
  buffer buf_n3038( .i (n3037), .o (n3038) );
  inverter inv_n3039( .i (n3038), .o (n3039) );
  assign n3040 = G56 & n3007 ;
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  assign n3041 = n1618 | n2809 ;
  buffer buf_n3042( .i (n3041), .o (n3042) );
  assign n3047 = n1713 & n3042 ;
  buffer buf_n3048( .i (n3047), .o (n3048) );
  assign n3052 = n1701 | n3048 ;
  buffer buf_n3053( .i (n3052), .o (n3053) );
  assign n3054 = n1769 | n3053 ;
  assign n3055 = n1769 & n3053 ;
  assign n3056 = n3054 & ~n3055 ;
  buffer buf_n3057( .i (n3056), .o (n3057) );
  assign n3060 = ~n3025 & n3057 ;
  assign n3061 = n1529 & n3027 ;
  assign n3062 = n3030 & ~n3061 ;
  assign n3063 = ~n3060 & n3062 ;
  assign n3064 = n3040 | n3063 ;
  buffer buf_n3065( .i (n3064), .o (n3065) );
  buffer buf_n3066( .i (n3065), .o (n3066) );
  buffer buf_n3067( .i (n3066), .o (n3067) );
  buffer buf_n3068( .i (n3067), .o (n3068) );
  buffer buf_n3069( .i (n3068), .o (n3069) );
  inverter inv_n3070( .i (n3069), .o (n3070) );
  assign n3071 = G55 & n3007 ;
  buffer buf_n3049( .i (n3048), .o (n3049) );
  buffer buf_n3050( .i (n3049), .o (n3050) );
  buffer buf_n3051( .i (n3050), .o (n3051) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n3043( .i (n3042), .o (n3043) );
  buffer buf_n3044( .i (n3043), .o (n3044) );
  buffer buf_n3045( .i (n3044), .o (n3045) );
  buffer buf_n3046( .i (n3045), .o (n3046) );
  assign n3072 = n1717 | n3046 ;
  assign n3073 = ~n3051 & n3072 ;
  buffer buf_n3074( .i (n3073), .o (n3074) );
  assign n3075 = ~n3025 & n3074 ;
  assign n3076 = n1481 & n3027 ;
  assign n3077 = n3030 & ~n3076 ;
  assign n3078 = ~n3075 & n3077 ;
  assign n3079 = n3071 | n3078 ;
  buffer buf_n3080( .i (n3079), .o (n3080) );
  buffer buf_n3081( .i (n3080), .o (n3081) );
  buffer buf_n3082( .i (n3081), .o (n3082) );
  buffer buf_n3083( .i (n3082), .o (n3083) );
  buffer buf_n3084( .i (n3083), .o (n3084) );
  inverter inv_n3085( .i (n3084), .o (n3085) );
  buffer buf_n2406( .i (n2405), .o (n2406) );
  assign n3086 = n2406 & n2482 ;
  assign n3087 = n2406 | n2482 ;
  assign n3088 = ~n3086 & n3087 ;
  buffer buf_n3089( .i (n3088), .o (n3089) );
  buffer buf_n3090( .i (n3089), .o (n3090) );
  buffer buf_n3091( .i (n3090), .o (n3091) );
  buffer buf_n3092( .i (n3091), .o (n3092) );
  buffer buf_n3093( .i (n3092), .o (n3093) );
  buffer buf_n3094( .i (n3093), .o (n3094) );
  buffer buf_n3095( .i (n3094), .o (n3095) );
  buffer buf_n3096( .i (n3095), .o (n3096) );
  buffer buf_n3097( .i (n3096), .o (n3097) );
  buffer buf_n3098( .i (n3097), .o (n3098) );
  buffer buf_n2429( .i (n2428), .o (n2429) );
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  buffer buf_n2432( .i (n2431), .o (n2432) );
  buffer buf_n2433( .i (n2432), .o (n2433) );
  buffer buf_n2434( .i (n2433), .o (n2434) );
  buffer buf_n2435( .i (n2434), .o (n2435) );
  buffer buf_n2436( .i (n2435), .o (n2436) );
  buffer buf_n2437( .i (n2436), .o (n2437) );
  buffer buf_n2438( .i (n2437), .o (n2438) );
  buffer buf_n2439( .i (n2438), .o (n2439) );
  buffer buf_n2440( .i (n2439), .o (n2440) );
  buffer buf_n2441( .i (n2440), .o (n2441) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  buffer buf_n2501( .i (n2500), .o (n2501) );
  assign n3099 = n2442 & n2501 ;
  assign n3100 = n2442 | n2501 ;
  assign n3101 = ~n3099 & n3100 ;
  buffer buf_n3102( .i (n3101), .o (n3102) );
  assign n3103 = ~n3098 & n3102 ;
  assign n3104 = n3098 & ~n3102 ;
  assign n3105 = n3103 | n3104 ;
  buffer buf_n3106( .i (n3105), .o (n3106) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  assign n3107 = n419 & n643 ;
  assign n3108 = G133 & ~n419 ;
  assign n3109 = n3107 | n3108 ;
  buffer buf_n3110( .i (n3109), .o (n3110) );
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  buffer buf_n2250( .i (n2249), .o (n2250) );
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n2341( .i (n2340), .o (n2341) );
  buffer buf_n2342( .i (n2341), .o (n2342) );
  buffer buf_n2343( .i (n2342), .o (n2343) );
  buffer buf_n2344( .i (n2343), .o (n2344) );
  buffer buf_n2345( .i (n2344), .o (n2345) );
  buffer buf_n2346( .i (n2345), .o (n2346) );
  buffer buf_n2347( .i (n2346), .o (n2347) );
  buffer buf_n2348( .i (n2347), .o (n2348) );
  buffer buf_n2349( .i (n2348), .o (n2349) );
  buffer buf_n2350( .i (n2349), .o (n2350) );
  buffer buf_n2351( .i (n2350), .o (n2351) );
  buffer buf_n2352( .i (n2351), .o (n2352) );
  buffer buf_n2353( .i (n2352), .o (n2353) );
  buffer buf_n2354( .i (n2353), .o (n2354) );
  buffer buf_n2355( .i (n2354), .o (n2355) );
  buffer buf_n2356( .i (n2355), .o (n2356) );
  assign n3111 = n2256 | n2356 ;
  assign n3112 = n2256 & n2356 ;
  assign n3113 = n3111 & ~n3112 ;
  buffer buf_n3114( .i (n3113), .o (n3114) );
  assign n3115 = n3110 | n3114 ;
  assign n3116 = n3110 & n3114 ;
  assign n3117 = n3115 & ~n3116 ;
  buffer buf_n3118( .i (n3117), .o (n3118) );
  buffer buf_n2295( .i (n2294), .o (n2295) );
  buffer buf_n2190( .i (n2189), .o (n2190) );
  buffer buf_n2191( .i (n2190), .o (n2191) );
  buffer buf_n2192( .i (n2191), .o (n2192) );
  buffer buf_n2193( .i (n2192), .o (n2193) );
  buffer buf_n2194( .i (n2193), .o (n2194) );
  buffer buf_n2195( .i (n2194), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  buffer buf_n2197( .i (n2196), .o (n2197) );
  buffer buf_n2198( .i (n2197), .o (n2198) );
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n2200( .i (n2199), .o (n2200) );
  buffer buf_n2201( .i (n2200), .o (n2201) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  buffer buf_n2203( .i (n2202), .o (n2203) );
  buffer buf_n2525( .i (n2524), .o (n2525) );
  buffer buf_n2526( .i (n2525), .o (n2526) );
  buffer buf_n2527( .i (n2526), .o (n2527) );
  buffer buf_n2528( .i (n2527), .o (n2528) );
  buffer buf_n2529( .i (n2528), .o (n2529) );
  buffer buf_n2530( .i (n2529), .o (n2530) );
  buffer buf_n2531( .i (n2530), .o (n2531) );
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n2532), .o (n2533) );
  buffer buf_n2534( .i (n2533), .o (n2534) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  buffer buf_n2536( .i (n2535), .o (n2536) );
  buffer buf_n2537( .i (n2536), .o (n2537) );
  buffer buf_n2538( .i (n2537), .o (n2538) );
  assign n3119 = n2203 & n2538 ;
  buffer buf_n2506( .i (n2505), .o (n2506) );
  buffer buf_n2507( .i (n2506), .o (n2507) );
  buffer buf_n2508( .i (n2507), .o (n2508) );
  buffer buf_n2509( .i (n2508), .o (n2509) );
  buffer buf_n2510( .i (n2509), .o (n2510) );
  buffer buf_n2511( .i (n2510), .o (n2511) );
  buffer buf_n2512( .i (n2511), .o (n2512) );
  buffer buf_n2513( .i (n2512), .o (n2513) );
  buffer buf_n2514( .i (n2513), .o (n2514) );
  buffer buf_n2515( .i (n2514), .o (n2515) );
  buffer buf_n2516( .i (n2515), .o (n2516) );
  buffer buf_n2517( .i (n2516), .o (n2517) );
  buffer buf_n2518( .i (n2517), .o (n2518) );
  buffer buf_n2519( .i (n2518), .o (n2519) );
  buffer buf_n2520( .i (n2519), .o (n2520) );
  buffer buf_n2521( .i (n2520), .o (n2521) );
  assign n3120 = n460 | n2521 ;
  assign n3121 = ~n3119 & n3120 ;
  buffer buf_n3122( .i (n3121), .o (n3122) );
  assign n3123 = ~n2295 & n3122 ;
  assign n3124 = n2295 & ~n3122 ;
  assign n3125 = n3123 | n3124 ;
  buffer buf_n3126( .i (n3125), .o (n3126) );
  assign n3127 = n3118 & ~n3126 ;
  assign n3128 = ~n3118 & n3126 ;
  assign n3129 = n3127 | n3128 ;
  buffer buf_n3130( .i (n3129), .o (n3130) );
  assign n3131 = ~n3106 & n3130 ;
  assign n3132 = n3106 & ~n3130 ;
  assign n3133 = n3131 | n3132 ;
  buffer buf_n3134( .i (n3133), .o (n3134) );
  buffer buf_n3135( .i (n3134), .o (n3135) );
  inverter inv_n3136( .i (n3135), .o (n3136) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  assign n3137 = n1746 & n1794 ;
  assign n3138 = n1746 | n1794 ;
  assign n3139 = ~n3137 & n3138 ;
  buffer buf_n3140( .i (n3139), .o (n3140) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  buffer buf_n1658( .i (n1657), .o (n1658) );
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  assign n3141 = ~n1604 & n1673 ;
  assign n3142 = n1604 & ~n1673 ;
  assign n3143 = n3141 | n3142 ;
  buffer buf_n3144( .i (n3143), .o (n3144) );
  assign n3145 = n3140 | n3144 ;
  assign n3146 = n3140 & n3144 ;
  assign n3147 = n3145 & ~n3146 ;
  buffer buf_n3148( .i (n3147), .o (n3148) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  buffer buf_n1954( .i (n1953), .o (n1954) );
  buffer buf_n1955( .i (n1954), .o (n1955) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  buffer buf_n1960( .i (n1959), .o (n1960) );
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1966( .i (n1965), .o (n1966) );
  buffer buf_n1967( .i (n1966), .o (n1967) );
  buffer buf_n2018( .i (n2017), .o (n2018) );
  buffer buf_n2019( .i (n2018), .o (n2019) );
  buffer buf_n2020( .i (n2019), .o (n2020) );
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2028( .i (n2027), .o (n2028) );
  buffer buf_n2029( .i (n2028), .o (n2029) );
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n2031( .i (n2030), .o (n2031) );
  buffer buf_n2032( .i (n2031), .o (n2032) );
  buffer buf_n2033( .i (n2032), .o (n2033) );
  buffer buf_n2034( .i (n2033), .o (n2034) );
  buffer buf_n2035( .i (n2034), .o (n2035) );
  buffer buf_n2036( .i (n2035), .o (n2036) );
  buffer buf_n2037( .i (n2036), .o (n2037) );
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  assign n3149 = n1967 & n2043 ;
  assign n3150 = n1967 | n2043 ;
  assign n3151 = ~n3149 & n3150 ;
  buffer buf_n3152( .i (n3151), .o (n3152) );
  buffer buf_n2077( .i (n2076), .o (n2077) );
  buffer buf_n2078( .i (n2077), .o (n2078) );
  buffer buf_n2079( .i (n2078), .o (n2079) );
  buffer buf_n2080( .i (n2079), .o (n2080) );
  buffer buf_n2081( .i (n2080), .o (n2081) );
  buffer buf_n2082( .i (n2081), .o (n2082) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2089( .i (n2088), .o (n2089) );
  buffer buf_n2090( .i (n2089), .o (n2090) );
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  assign n3153 = n286 & n443 ;
  assign n3154 = G112 & ~n443 ;
  assign n3155 = n3153 | n3154 ;
  buffer buf_n3156( .i (n3155), .o (n3156) );
  assign n3157 = n2098 & ~n3156 ;
  assign n3158 = ~n2098 & n3156 ;
  assign n3159 = n3157 | n3158 ;
  buffer buf_n3160( .i (n3159), .o (n3160) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n1556( .i (n1555), .o (n1556) );
  buffer buf_n1557( .i (n1556), .o (n1557) );
  buffer buf_n1558( .i (n1557), .o (n1558) );
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  buffer buf_n1872( .i (n1871), .o (n1872) );
  buffer buf_n1873( .i (n1872), .o (n1873) );
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  assign n3161 = ~n1560 & n1878 ;
  assign n3162 = n1560 & ~n1878 ;
  assign n3163 = n3161 | n3162 ;
  buffer buf_n3164( .i (n3163), .o (n3164) );
  assign n3165 = ~n3160 & n3164 ;
  assign n3166 = n3160 & ~n3164 ;
  assign n3167 = n3165 | n3166 ;
  buffer buf_n3168( .i (n3167), .o (n3168) );
  assign n3169 = ~n3152 & n3168 ;
  assign n3170 = n3152 & ~n3168 ;
  assign n3171 = n3169 | n3170 ;
  buffer buf_n3172( .i (n3171), .o (n3172) );
  assign n3173 = ~n3148 & n3172 ;
  assign n3174 = n3148 & ~n3172 ;
  assign n3175 = n3173 | n3174 ;
  buffer buf_n3176( .i (n3175), .o (n3176) );
  inverter inv_n3177( .i (n3176), .o (n3177) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  assign n3178 = n2690 | n2967 ;
  buffer buf_n3179( .i (n3178), .o (n3179) );
  buffer buf_n3180( .i (n3179), .o (n3180) );
  buffer buf_n3181( .i (n3180), .o (n3181) );
  assign n3183 = n2173 & n3181 ;
  assign n3184 = n2734 | n3183 ;
  buffer buf_n3185( .i (n3184), .o (n3185) );
  assign n3186 = n1939 | n3185 ;
  assign n3187 = n1939 & n3185 ;
  assign n3188 = n3186 & ~n3187 ;
  buffer buf_n3189( .i (n3188), .o (n3189) );
  buffer buf_n3190( .i (n3189), .o (n3190) );
  buffer buf_n3191( .i (n3190), .o (n3191) );
  buffer buf_n3192( .i (n3191), .o (n3192) );
  buffer buf_n3193( .i (n3192), .o (n3193) );
  buffer buf_n2139( .i (n2138), .o (n2139) );
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n2143( .i (n2142), .o (n2143) );
  buffer buf_n2144( .i (n2143), .o (n2144) );
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  buffer buf_n2152( .i (n2151), .o (n2152) );
  buffer buf_n2153( .i (n2152), .o (n2153) );
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n2155( .i (n2154), .o (n2155) );
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n3182( .i (n3181), .o (n3182) );
  assign n3194 = n2156 | n3182 ;
  assign n3195 = n2156 & n3182 ;
  assign n3196 = n3194 & ~n3195 ;
  buffer buf_n3197( .i (n3196), .o (n3197) );
  buffer buf_n3198( .i (n3197), .o (n3198) );
  buffer buf_n3199( .i (n3198), .o (n3199) );
  buffer buf_n3200( .i (n3199), .o (n3200) );
  buffer buf_n3201( .i (n3200), .o (n3201) );
  buffer buf_n3202( .i (n3201), .o (n3202) );
  buffer buf_n2992( .i (n2991), .o (n2992) );
  buffer buf_n2993( .i (n2992), .o (n2993) );
  buffer buf_n2994( .i (n2993), .o (n2994) );
  buffer buf_n3058( .i (n3057), .o (n3058) );
  buffer buf_n3059( .i (n3058), .o (n3059) );
  buffer buf_n3024( .i (n3023), .o (n3024) );
  assign n3203 = ~n2819 & n3074 ;
  assign n3204 = n3024 & n3203 ;
  assign n3205 = n3059 & n3204 ;
  assign n3206 = n2994 & n3205 ;
  assign n3207 = ~n3202 & n3206 ;
  assign n3208 = n3193 & n3207 ;
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n2012( .i (n2011), .o (n2012) );
  buffer buf_n2013( .i (n2012), .o (n2013) );
  buffer buf_n2709( .i (n2708), .o (n2709) );
  buffer buf_n2710( .i (n2709), .o (n2710) );
  buffer buf_n2711( .i (n2710), .o (n2711) );
  buffer buf_n2712( .i (n2711), .o (n2712) );
  buffer buf_n2713( .i (n2712), .o (n2713) );
  buffer buf_n2714( .i (n2713), .o (n2714) );
  buffer buf_n2715( .i (n2714), .o (n2715) );
  buffer buf_n2716( .i (n2715), .o (n2716) );
  buffer buf_n2717( .i (n2716), .o (n2717) );
  buffer buf_n2718( .i (n2717), .o (n2718) );
  buffer buf_n2719( .i (n2718), .o (n2719) );
  buffer buf_n2720( .i (n2719), .o (n2720) );
  assign n3209 = n2171 & n3179 ;
  assign n3210 = n2720 | n3209 ;
  buffer buf_n3211( .i (n3210), .o (n3211) );
  assign n3212 = ~n2013 & n3211 ;
  assign n3213 = n2013 & ~n3211 ;
  assign n3214 = n3212 | n3213 ;
  buffer buf_n3215( .i (n3214), .o (n3215) );
  buffer buf_n3216( .i (n3215), .o (n3216) );
  buffer buf_n3217( .i (n3216), .o (n3217) );
  buffer buf_n3218( .i (n3217), .o (n3218) );
  buffer buf_n3219( .i (n3218), .o (n3219) );
  buffer buf_n3220( .i (n3219), .o (n3220) );
  buffer buf_n3221( .i (n3220), .o (n3221) );
  buffer buf_n2055( .i (n2054), .o (n2055) );
  buffer buf_n2056( .i (n2055), .o (n2056) );
  buffer buf_n2057( .i (n2056), .o (n2057) );
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  buffer buf_n2064( .i (n2063), .o (n2064) );
  buffer buf_n2065( .i (n2064), .o (n2065) );
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n2120( .i (n2119), .o (n2120) );
  buffer buf_n2121( .i (n2120), .o (n2121) );
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  buffer buf_n2129( .i (n2128), .o (n2129) );
  buffer buf_n2130( .i (n2129), .o (n2130) );
  buffer buf_n2131( .i (n2130), .o (n2131) );
  buffer buf_n2132( .i (n2131), .o (n2132) );
  buffer buf_n2133( .i (n2132), .o (n2133) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  assign n3222 = n2136 & n3179 ;
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n2102( .i (n2101), .o (n2102) );
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  buffer buf_n2111( .i (n2110), .o (n2111) );
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  assign n3223 = n2117 | n3179 ;
  assign n3224 = ~n3222 & n3223 ;
  buffer buf_n3225( .i (n3224), .o (n3225) );
  assign n3226 = n2072 | n3225 ;
  assign n3227 = n2072 & n3225 ;
  assign n3228 = n3226 & ~n3227 ;
  buffer buf_n3229( .i (n3228), .o (n3229) );
  buffer buf_n3230( .i (n3229), .o (n3230) );
  buffer buf_n3231( .i (n3230), .o (n3231) );
  buffer buf_n3232( .i (n3231), .o (n3232) );
  buffer buf_n3233( .i (n3232), .o (n3233) );
  buffer buf_n3234( .i (n3233), .o (n3234) );
  buffer buf_n3235( .i (n3234), .o (n3235) );
  assign n3236 = n3221 & ~n3235 ;
  assign n3237 = n3208 & n3236 ;
  buffer buf_n3238( .i (n3237), .o (n3238) );
  buffer buf_n3239( .i (n3238), .o (n3239) );
  buffer buf_n2421( .i (n2420), .o (n2421) );
  buffer buf_n2422( .i (n2421), .o (n2422) );
  buffer buf_n2423( .i (n2422), .o (n2423) );
  buffer buf_n2424( .i (n2423), .o (n2424) );
  buffer buf_n2454( .i (n2453), .o (n2454) );
  buffer buf_n2455( .i (n2454), .o (n2455) );
  buffer buf_n2456( .i (n2455), .o (n2456) );
  buffer buf_n2457( .i (n2456), .o (n2457) );
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n2460( .i (n2459), .o (n2460) );
  buffer buf_n2541( .i (n2540), .o (n2541) );
  buffer buf_n2542( .i (n2541), .o (n2542) );
  buffer buf_n2543( .i (n2542), .o (n2543) );
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  buffer buf_n2551( .i (n2550), .o (n2551) );
  buffer buf_n2552( .i (n2551), .o (n2552) );
  buffer buf_n2553( .i (n2552), .o (n2553) );
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2555( .i (n2554), .o (n2555) );
  assign n3240 = n2555 & n2868 ;
  assign n3241 = n2547 | n3240 ;
  buffer buf_n3242( .i (n3241), .o (n3242) );
  buffer buf_n3243( .i (n3242), .o (n3243) );
  assign n3247 = n2460 & n3243 ;
  buffer buf_n2445( .i (n2444), .o (n2445) );
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n2448( .i (n2447), .o (n2448) );
  buffer buf_n2449( .i (n2448), .o (n2449) );
  buffer buf_n2450( .i (n2449), .o (n2450) );
  buffer buf_n2451( .i (n2450), .o (n2451) );
  assign n3248 = n2451 | n3243 ;
  assign n3249 = ~n3247 & n3248 ;
  buffer buf_n3250( .i (n3249), .o (n3250) );
  assign n3251 = n2424 & n3250 ;
  assign n3252 = n2424 | n3250 ;
  assign n3253 = ~n3251 & n3252 ;
  buffer buf_n3254( .i (n3253), .o (n3254) );
  buffer buf_n3255( .i (n3254), .o (n3255) );
  buffer buf_n3256( .i (n3255), .o (n3256) );
  buffer buf_n3257( .i (n3256), .o (n3257) );
  buffer buf_n3258( .i (n3257), .o (n3258) );
  buffer buf_n3259( .i (n3258), .o (n3259) );
  buffer buf_n3260( .i (n3259), .o (n3260) );
  buffer buf_n3261( .i (n3260), .o (n3261) );
  buffer buf_n3262( .i (n3261), .o (n3262) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  buffer buf_n2411( .i (n2410), .o (n2411) );
  buffer buf_n2412( .i (n2411), .o (n2412) );
  buffer buf_n2413( .i (n2412), .o (n2413) );
  buffer buf_n2416( .i (n2415), .o (n2416) );
  buffer buf_n2417( .i (n2416), .o (n2417) );
  buffer buf_n2418( .i (n2417), .o (n2418) );
  assign n3263 = n2418 & n2451 ;
  assign n3264 = n2413 | n3263 ;
  buffer buf_n3244( .i (n3243), .o (n3244) );
  assign n3265 = n2472 & n3244 ;
  assign n3266 = n3264 | n3265 ;
  buffer buf_n3267( .i (n3266), .o (n3267) );
  assign n3268 = n2500 | n3267 ;
  assign n3269 = n2500 & n3267 ;
  assign n3270 = n3268 & ~n3269 ;
  buffer buf_n3271( .i (n3270), .o (n3271) );
  buffer buf_n3272( .i (n3271), .o (n3272) );
  buffer buf_n3273( .i (n3272), .o (n3273) );
  buffer buf_n3274( .i (n3273), .o (n3274) );
  buffer buf_n3275( .i (n3274), .o (n3275) );
  buffer buf_n3276( .i (n3275), .o (n3276) );
  buffer buf_n3277( .i (n3276), .o (n3277) );
  buffer buf_n2467( .i (n2466), .o (n2467) );
  buffer buf_n2468( .i (n2467), .o (n2468) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  buffer buf_n2470( .i (n2469), .o (n2470) );
  buffer buf_n3245( .i (n3244), .o (n3245) );
  buffer buf_n3246( .i (n3245), .o (n3246) );
  assign n3278 = n2470 & n3246 ;
  assign n3279 = n2470 | n3246 ;
  assign n3280 = ~n3278 & n3279 ;
  buffer buf_n3281( .i (n3280), .o (n3281) );
  buffer buf_n3282( .i (n3281), .o (n3282) );
  buffer buf_n3283( .i (n3282), .o (n3283) );
  buffer buf_n3284( .i (n3283), .o (n3284) );
  buffer buf_n3285( .i (n3284), .o (n3285) );
  buffer buf_n3286( .i (n3285), .o (n3286) );
  buffer buf_n3287( .i (n3286), .o (n3287) );
  buffer buf_n2880( .i (n2879), .o (n2880) );
  buffer buf_n2881( .i (n2880), .o (n2881) );
  buffer buf_n2882( .i (n2881), .o (n2882) );
  buffer buf_n2883( .i (n2882), .o (n2883) );
  buffer buf_n2884( .i (n2883), .o (n2884) );
  buffer buf_n2908( .i (n2907), .o (n2908) );
  buffer buf_n2909( .i (n2908), .o (n2909) );
  buffer buf_n2910( .i (n2909), .o (n2910) );
  buffer buf_n2911( .i (n2910), .o (n2911) );
  buffer buf_n2912( .i (n2911), .o (n2912) );
  buffer buf_n2913( .i (n2912), .o (n2913) );
  buffer buf_n2935( .i (n2934), .o (n2935) );
  buffer buf_n2936( .i (n2935), .o (n2936) );
  buffer buf_n2937( .i (n2936), .o (n2937) );
  buffer buf_n2793( .i (n2792), .o (n2793) );
  buffer buf_n2794( .i (n2793), .o (n2794) );
  assign n3288 = n2776 & n2833 ;
  assign n3289 = ~n2794 & n3288 ;
  assign n3290 = n2937 & n3289 ;
  assign n3291 = n2913 & n3290 ;
  assign n3292 = n2884 & n3291 ;
  assign n3293 = ~n3287 & n3292 ;
  assign n3294 = ~n3277 & n3293 ;
  assign n3295 = ~n3262 & n3294 ;
  buffer buf_n3296( .i (n3295), .o (n3296) );
  buffer buf_n920( .i (G158), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  assign n3297 = n923 | n2826 ;
  buffer buf_n924( .i (G159), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  assign n3298 = n922 & ~n2782 ;
  assign n3299 = n927 & ~n3298 ;
  assign n3300 = n3297 & n3299 ;
  buffer buf_n1040( .i (G81), .o (n1040) );
  assign n3301 = n920 | n924 ;
  buffer buf_n3302( .i (n3301), .o (n3302) );
  buffer buf_n3303( .i (n3302), .o (n3303) );
  assign n3304 = n1040 & ~n3303 ;
  buffer buf_n1039( .i (G80), .o (n1039) );
  assign n3305 = n920 & ~n924 ;
  buffer buf_n3306( .i (n3305), .o (n3306) );
  buffer buf_n3307( .i (n3306), .o (n3307) );
  assign n3308 = n1039 & n3307 ;
  assign n3309 = n3304 | n3308 ;
  assign n3310 = n3300 | n3309 ;
  assign n3311 = n1022 & n3310 ;
  buffer buf_n929( .i (G160), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  assign n3312 = n932 | n2826 ;
  buffer buf_n933( .i (G161), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  assign n3313 = n931 & ~n2782 ;
  assign n3314 = n936 & ~n3313 ;
  assign n3315 = n3312 & n3314 ;
  assign n3316 = n929 | n933 ;
  buffer buf_n3317( .i (n3316), .o (n3317) );
  buffer buf_n3318( .i (n3317), .o (n3318) );
  assign n3319 = n1040 & ~n3318 ;
  assign n3320 = n929 & ~n933 ;
  buffer buf_n3321( .i (n3320), .o (n3321) );
  buffer buf_n3322( .i (n3321), .o (n3322) );
  assign n3323 = n1039 & n3322 ;
  assign n3324 = n3319 | n3323 ;
  assign n3325 = n3315 | n3324 ;
  assign n3326 = n1022 & n3325 ;
  assign n3327 = n967 | n3002 ;
  assign n3328 = n966 & ~n2893 ;
  assign n3329 = n963 & ~n3328 ;
  assign n3330 = n3327 & n3329 ;
  buffer buf_n928( .i (G16), .o (n928) );
  assign n3331 = n928 & n2849 ;
  buffer buf_n721( .i (G14), .o (n721) );
  assign n3332 = n721 & ~n2853 ;
  assign n3333 = n3331 | n3332 ;
  assign n3334 = n3330 | n3333 ;
  assign n3335 = n967 | n3036 ;
  assign n3336 = n966 & ~n2923 ;
  assign n3337 = n963 & ~n3336 ;
  assign n3338 = n3335 & n3337 ;
  buffer buf_n1018( .i (G6), .o (n1018) );
  assign n3339 = n1018 & ~n2853 ;
  buffer buf_n1005( .i (G27), .o (n1005) );
  assign n3340 = n1005 & n2849 ;
  assign n3341 = n3339 | n3340 ;
  assign n3342 = n3338 | n3341 ;
  assign n3343 = n967 | n3067 ;
  buffer buf_n3344( .i (n965), .o (n3344) );
  assign n3345 = ~n2946 & n3344 ;
  assign n3346 = n963 & ~n3345 ;
  assign n3347 = n3343 & n3346 ;
  buffer buf_n1004( .i (G26), .o (n1004) );
  assign n3348 = n1004 & n2849 ;
  buffer buf_n1013( .i (G5), .o (n1013) );
  assign n3349 = n1013 & ~n2853 ;
  assign n3350 = n3348 | n3349 ;
  assign n3351 = n3347 | n3350 ;
  buffer buf_n3352( .i (n3344), .o (n3352) );
  assign n3353 = n3082 | n3352 ;
  assign n3354 = ~n2802 & n3344 ;
  buffer buf_n3355( .i (n962), .o (n3355) );
  assign n3356 = ~n3354 & n3355 ;
  assign n3357 = n3353 & n3356 ;
  buffer buf_n1002( .i (G24), .o (n1002) );
  buffer buf_n3358( .i (n2848), .o (n3358) );
  assign n3359 = n1002 & n3358 ;
  buffer buf_n1003( .i (G25), .o (n1003) );
  buffer buf_n3360( .i (n2852), .o (n3360) );
  assign n3361 = n1003 & ~n3360 ;
  assign n3362 = n3359 | n3361 ;
  assign n3363 = n3357 | n3362 ;
  assign n3364 = n971 | n3002 ;
  assign n3365 = n970 & ~n2893 ;
  assign n3366 = n975 & ~n3365 ;
  assign n3367 = n3364 & n3366 ;
  assign n3368 = n721 & ~n2961 ;
  assign n3369 = n928 & n2957 ;
  assign n3370 = n3368 | n3369 ;
  assign n3371 = n3367 | n3370 ;
  assign n3372 = n971 | n3036 ;
  assign n3373 = n970 & ~n2923 ;
  assign n3374 = n975 & ~n3373 ;
  assign n3375 = n3372 & n3374 ;
  assign n3376 = n1005 & n2957 ;
  assign n3377 = n1018 & ~n2961 ;
  assign n3378 = n3376 | n3377 ;
  assign n3379 = n3375 | n3378 ;
  assign n3380 = n971 | n3067 ;
  buffer buf_n3381( .i (n969), .o (n3381) );
  assign n3382 = ~n2946 & n3381 ;
  assign n3383 = n975 & ~n3382 ;
  assign n3384 = n3380 & n3383 ;
  assign n3385 = n1013 & ~n2961 ;
  assign n3386 = n1004 & n2957 ;
  assign n3387 = n3385 | n3386 ;
  assign n3388 = n3384 | n3387 ;
  buffer buf_n3389( .i (n3381), .o (n3389) );
  assign n3390 = n3082 | n3389 ;
  assign n3391 = ~n2802 & n3381 ;
  buffer buf_n3392( .i (n974), .o (n3392) );
  assign n3393 = ~n3391 & n3392 ;
  assign n3394 = n3390 & n3393 ;
  buffer buf_n3395( .i (n2956), .o (n3395) );
  assign n3396 = n1002 & n3395 ;
  buffer buf_n3397( .i (n2960), .o (n3397) );
  assign n3398 = n1003 & ~n3397 ;
  assign n3399 = n3396 | n3398 ;
  assign n3400 = n3394 | n3399 ;
  assign n3401 = n923 | n3001 ;
  assign n3402 = n922 & ~n2892 ;
  assign n3403 = n927 & ~n3402 ;
  assign n3404 = n3401 & n3403 ;
  buffer buf_n1035( .i (G76), .o (n1035) );
  assign n3405 = n1035 & ~n3303 ;
  buffer buf_n1045( .i (G86), .o (n1045) );
  assign n3406 = n1045 & n3307 ;
  assign n3407 = n3405 | n3406 ;
  assign n3408 = n3404 | n3407 ;
  assign n3409 = n1022 & n3408 ;
  assign n3410 = n923 | n3081 ;
  assign n3411 = n922 & ~n2801 ;
  assign n3412 = n927 & ~n3411 ;
  assign n3413 = n3410 & n3412 ;
  buffer buf_n1031( .i (G72), .o (n1031) );
  assign n3414 = n1031 & ~n3303 ;
  buffer buf_n1041( .i (G82), .o (n1041) );
  assign n3415 = n1041 & n3307 ;
  assign n3416 = n3414 | n3415 ;
  assign n3417 = n3413 | n3416 ;
  buffer buf_n3418( .i (n1021), .o (n3418) );
  assign n3419 = n3417 & n3418 ;
  assign n3420 = n923 | n3066 ;
  buffer buf_n3421( .i (n921), .o (n3421) );
  assign n3422 = ~n2945 & n3421 ;
  assign n3423 = n927 & ~n3422 ;
  assign n3424 = n3420 & n3423 ;
  buffer buf_n1029( .i (G70), .o (n1029) );
  assign n3425 = n1029 & ~n3303 ;
  buffer buf_n1030( .i (G71), .o (n1030) );
  assign n3426 = n1030 & n3307 ;
  assign n3427 = n3425 | n3426 ;
  assign n3428 = n3424 | n3427 ;
  assign n3429 = n3418 & n3428 ;
  buffer buf_n3430( .i (n3421), .o (n3430) );
  assign n3431 = n3035 | n3430 ;
  assign n3432 = ~n2922 & n3421 ;
  buffer buf_n3433( .i (n926), .o (n3433) );
  assign n3434 = ~n3432 & n3433 ;
  assign n3435 = n3431 & n3434 ;
  buffer buf_n1027( .i (G68), .o (n1027) );
  buffer buf_n3436( .i (n3302), .o (n3436) );
  assign n3437 = n1027 & ~n3436 ;
  buffer buf_n1028( .i (G69), .o (n1028) );
  buffer buf_n3438( .i (n3306), .o (n3438) );
  assign n3439 = n1028 & n3438 ;
  assign n3440 = n3437 | n3439 ;
  assign n3441 = n3435 | n3440 ;
  assign n3442 = n3418 & n3441 ;
  assign n3443 = n932 | n3001 ;
  assign n3444 = n931 & ~n2892 ;
  assign n3445 = n936 & ~n3444 ;
  assign n3446 = n3443 & n3445 ;
  assign n3447 = n1035 & ~n3318 ;
  assign n3448 = n1045 & n3322 ;
  assign n3449 = n3447 | n3448 ;
  assign n3450 = n3446 | n3449 ;
  assign n3451 = n3418 & n3450 ;
  assign n3452 = n932 | n3081 ;
  assign n3453 = n931 & ~n2801 ;
  assign n3454 = n936 & ~n3453 ;
  assign n3455 = n3452 & n3454 ;
  assign n3456 = n1031 & ~n3318 ;
  assign n3457 = n1041 & n3322 ;
  assign n3458 = n3456 | n3457 ;
  assign n3459 = n3455 | n3458 ;
  buffer buf_n3460( .i (n1021), .o (n3460) );
  assign n3461 = n3459 & n3460 ;
  assign n3462 = n932 | n3066 ;
  buffer buf_n3463( .i (n930), .o (n3463) );
  assign n3464 = ~n2945 & n3463 ;
  assign n3465 = n936 & ~n3464 ;
  assign n3466 = n3462 & n3465 ;
  assign n3467 = n1029 & ~n3318 ;
  assign n3468 = n1030 & n3322 ;
  assign n3469 = n3467 | n3468 ;
  assign n3470 = n3466 | n3469 ;
  assign n3471 = n3460 & n3470 ;
  buffer buf_n3472( .i (n3463), .o (n3472) );
  assign n3473 = n3035 | n3472 ;
  assign n3474 = ~n2922 & n3463 ;
  buffer buf_n3475( .i (n935), .o (n3475) );
  assign n3476 = ~n3474 & n3475 ;
  assign n3477 = n3473 & n3476 ;
  buffer buf_n3478( .i (n3317), .o (n3478) );
  assign n3479 = n1027 & ~n3478 ;
  buffer buf_n3480( .i (n3321), .o (n3480) );
  assign n3481 = n1028 & n3480 ;
  assign n3482 = n3479 | n3481 ;
  assign n3483 = n3477 | n3482 ;
  assign n3484 = n3460 & n3483 ;
  buffer buf_n958( .i (G171), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n956( .i (G170), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  assign n3485 = n957 & n2838 ;
  buffer buf_n1019( .i (G61), .o (n1019) );
  buffer buf_n2491( .i (n2490), .o (n2491) );
  buffer buf_n2492( .i (n2491), .o (n2492) );
  buffer buf_n2493( .i (n2492), .o (n2493) );
  buffer buf_n2494( .i (n2493), .o (n2494) );
  buffer buf_n2495( .i (n2494), .o (n2495) );
  assign n3486 = ~n1019 & n2495 ;
  assign n3487 = n1019 & ~n2495 ;
  assign n3488 = n3486 | n3487 ;
  buffer buf_n3489( .i (n3488), .o (n3489) );
  assign n3492 = n957 | n3489 ;
  assign n3493 = ~n3485 & n3492 ;
  assign n3494 = n959 & ~n3493 ;
  assign n3495 = G178 & G62 ;
  buffer buf_n1014( .i (G54), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  assign n3496 = n956 & ~n1017 ;
  buffer buf_n1309( .i (n1308), .o (n1309) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  assign n3497 = n956 | n1323 ;
  assign n3498 = ~n3496 & n3497 ;
  assign n3499 = n958 | n3498 ;
  assign n3500 = ~n3495 & n3499 ;
  assign n3501 = ~n3494 & n3500 ;
  buffer buf_n3490( .i (n3489), .o (n3490) );
  buffer buf_n3491( .i (n3490), .o (n3491) );
  assign n3502 = n2840 & n3491 ;
  assign n3503 = n2840 | n3491 ;
  assign n3504 = n3502 | ~n3503 ;
  assign n3505 = n1014 & n3007 ;
  assign n3506 = n2833 & ~n3025 ;
  assign n3507 = ~n1318 & n3027 ;
  assign n3508 = n3030 & ~n3507 ;
  assign n3509 = ~n3506 & n3508 ;
  assign n3510 = n3505 | n3509 ;
  buffer buf_n3511( .i (n3510), .o (n3511) );
  buffer buf_n3512( .i (n3511), .o (n3512) );
  buffer buf_n3513( .i (n3512), .o (n3513) );
  buffer buf_n3514( .i (n3513), .o (n3514) );
  buffer buf_n3515( .i (n3514), .o (n3515) );
  inverter inv_n3516( .i (n3515), .o (n3516) );
  buffer buf_n3517( .i (n3006), .o (n3517) );
  assign n3518 = G52 & n3517 ;
  buffer buf_n3519( .i (n2939), .o (n3519) );
  buffer buf_n3520( .i (n3519), .o (n3520) );
  assign n3521 = n3271 | n3520 ;
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  assign n3522 = ~n1337 & n3519 ;
  buffer buf_n3523( .i (n3029), .o (n3523) );
  assign n3524 = ~n3522 & n3523 ;
  assign n3525 = n3521 & n3524 ;
  assign n3526 = n3518 | n3525 ;
  buffer buf_n3527( .i (n3526), .o (n3527) );
  buffer buf_n3528( .i (n3527), .o (n3528) );
  buffer buf_n3529( .i (n3528), .o (n3529) );
  buffer buf_n3530( .i (n3529), .o (n3530) );
  buffer buf_n3531( .i (n3530), .o (n3531) );
  inverter inv_n3532( .i (n3531), .o (n3532) );
  assign n3533 = G47 & n3006 ;
  assign n3534 = n3254 | n3519 ;
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  assign n3535 = n1262 & n2939 ;
  assign n3536 = n3029 & ~n3535 ;
  assign n3537 = n3534 & n3536 ;
  assign n3538 = n3533 | n3537 ;
  buffer buf_n3539( .i (n3538), .o (n3539) );
  buffer buf_n3540( .i (n3539), .o (n3540) );
  buffer buf_n3541( .i (n3540), .o (n3541) );
  buffer buf_n3542( .i (n3541), .o (n3542) );
  buffer buf_n3543( .i (n3542), .o (n3543) );
  buffer buf_n3544( .i (n3543), .o (n3544) );
  inverter inv_n3545( .i (n3544), .o (n3545) );
  assign n3546 = G43 & n3006 ;
  assign n3547 = n3281 | n3519 ;
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n3548( .i (n977), .o (n3548) );
  assign n3549 = n1282 & n3548 ;
  assign n3550 = n3029 & ~n3549 ;
  assign n3551 = n3547 & n3550 ;
  assign n3552 = n3546 | n3551 ;
  buffer buf_n3553( .i (n3552), .o (n3553) );
  buffer buf_n3554( .i (n3553), .o (n3554) );
  buffer buf_n3555( .i (n3554), .o (n3555) );
  buffer buf_n3556( .i (n3555), .o (n3556) );
  buffer buf_n3557( .i (n3556), .o (n3557) );
  buffer buf_n3558( .i (n3557), .o (n3558) );
  inverter inv_n3559( .i (n3558), .o (n3559) );
  assign n3560 = n900 & n1175 ;
  assign n3561 = n1195 & n3560 ;
  assign n3562 = n1184 & n3561 ;
  assign n3563 = ~n2613 & n3562 ;
  assign n3564 = ~n2656 & n3563 ;
  assign n3565 = ~n3134 & n3564 ;
  assign n3566 = ~n3176 & n3565 ;
  buffer buf_n2766( .i (n2765), .o (n2766) );
  assign n3567 = G46 & n2766 ;
  buffer buf_n981( .i (n980), .o (n981) );
  assign n3568 = ~n981 & n3189 ;
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  assign n3569 = n1501 & n3520 ;
  assign n3570 = n987 & ~n3569 ;
  assign n3571 = ~n3568 & n3570 ;
  assign n3572 = n3567 | n3571 ;
  buffer buf_n3573( .i (n3572), .o (n3573) );
  buffer buf_n3574( .i (n3573), .o (n3574) );
  buffer buf_n3575( .i (n3574), .o (n3575) );
  buffer buf_n3576( .i (n3575), .o (n3576) );
  inverter inv_n3577( .i (n3576), .o (n3577) );
  buffer buf_n3578( .i (n2763), .o (n3578) );
  assign n3579 = G45 & n3578 ;
  buffer buf_n3580( .i (n3548), .o (n3580) );
  assign n3581 = n3215 & ~n3580 ;
  assign n3582 = n1430 & n3548 ;
  buffer buf_n3583( .i (n984), .o (n3583) );
  assign n3584 = ~n3582 & n3583 ;
  assign n3585 = ~n3581 & n3584 ;
  assign n3586 = n3579 | n3585 ;
  buffer buf_n3587( .i (n3586), .o (n3587) );
  buffer buf_n3588( .i (n3587), .o (n3588) );
  buffer buf_n3589( .i (n3588), .o (n3589) );
  buffer buf_n3590( .i (n3589), .o (n3590) );
  buffer buf_n3591( .i (n3590), .o (n3591) );
  buffer buf_n3592( .i (n3591), .o (n3592) );
  inverter inv_n3593( .i (n3592), .o (n3593) );
  assign n3594 = G20 & n3578 ;
  assign n3595 = n3229 | n3580 ;
  assign n3596 = n1443 & n3548 ;
  assign n3597 = n3583 & ~n3596 ;
  assign n3598 = n3595 & n3597 ;
  assign n3599 = n3594 | n3598 ;
  buffer buf_n3600( .i (n3599), .o (n3600) );
  buffer buf_n3601( .i (n3600), .o (n3601) );
  buffer buf_n3602( .i (n3601), .o (n3602) );
  buffer buf_n3603( .i (n3602), .o (n3603) );
  buffer buf_n3604( .i (n3603), .o (n3604) );
  buffer buf_n3605( .i (n3604), .o (n3605) );
  inverter inv_n3606( .i (n3605), .o (n3606) );
  assign n3607 = G44 & n3578 ;
  assign n3608 = n3197 | n3580 ;
  buffer buf_n3609( .i (n976), .o (n3609) );
  buffer buf_n3610( .i (n3609), .o (n3610) );
  assign n3611 = n1416 & n3610 ;
  assign n3612 = n3583 & ~n3611 ;
  assign n3613 = n3608 & n3612 ;
  assign n3614 = n3607 | n3613 ;
  buffer buf_n3615( .i (n3614), .o (n3615) );
  buffer buf_n3616( .i (n3615), .o (n3616) );
  buffer buf_n3617( .i (n3616), .o (n3617) );
  buffer buf_n3618( .i (n3617), .o (n3618) );
  buffer buf_n3619( .i (n3618), .o (n3619) );
  buffer buf_n3620( .i (n3619), .o (n3620) );
  inverter inv_n3621( .i (n3620), .o (n3621) );
  assign n3622 = n3389 | n3574 ;
  assign n3623 = n3381 & ~n3512 ;
  assign n3624 = n3392 & ~n3623 ;
  assign n3625 = n3622 & n3624 ;
  buffer buf_n1011( .i (G41), .o (n1011) );
  assign n3626 = n1011 & ~n3397 ;
  buffer buf_n1012( .i (G42), .o (n1012) );
  assign n3627 = n1012 & n3395 ;
  assign n3628 = n3626 | n3627 ;
  assign n3629 = n3625 | n3628 ;
  assign n3630 = n3352 | n3574 ;
  assign n3631 = n3344 & ~n3512 ;
  assign n3632 = n3355 & ~n3631 ;
  assign n3633 = n3630 & n3632 ;
  assign n3634 = n1011 & ~n3360 ;
  assign n3635 = n1012 & n3358 ;
  assign n3636 = n3634 | n3635 ;
  assign n3637 = n3633 | n3636 ;
  assign n3638 = n3352 & ~n3529 ;
  buffer buf_n3639( .i (n965), .o (n3639) );
  assign n3640 = n3589 | n3639 ;
  assign n3641 = n3355 & n3640 ;
  assign n3642 = ~n3638 & n3641 ;
  buffer buf_n955( .i (G17), .o (n955) );
  assign n3643 = n955 & n3358 ;
  buffer buf_n989( .i (G18), .o (n989) );
  assign n3644 = n989 & ~n3360 ;
  assign n3645 = n3643 | n3644 ;
  assign n3646 = n3642 | n3645 ;
  assign n3647 = n3352 & ~n3542 ;
  assign n3648 = n3602 | n3639 ;
  assign n3649 = n3355 & n3648 ;
  assign n3650 = ~n3647 & n3649 ;
  buffer buf_n1008( .i (G39), .o (n1008) );
  assign n3651 = n1008 & n3358 ;
  buffer buf_n1010( .i (G40), .o (n1010) );
  assign n3652 = n1010 & ~n3360 ;
  assign n3653 = n3651 | n3652 ;
  assign n3654 = n3650 | n3653 ;
  buffer buf_n3655( .i (n3639), .o (n3655) );
  assign n3656 = ~n3556 & n3655 ;
  assign n3657 = n3617 | n3639 ;
  buffer buf_n3658( .i (n962), .o (n3658) );
  assign n3659 = n3657 & n3658 ;
  assign n3660 = ~n3656 & n3659 ;
  buffer buf_n1007( .i (G36), .o (n1007) );
  buffer buf_n3661( .i (n2848), .o (n3661) );
  assign n3662 = n1007 & n3661 ;
  buffer buf_n869( .i (G15), .o (n869) );
  buffer buf_n3663( .i (n2852), .o (n3663) );
  assign n3664 = n869 & ~n3663 ;
  assign n3665 = n3662 | n3664 ;
  assign n3666 = n3660 | n3665 ;
  assign n3667 = n3389 | n3590 ;
  buffer buf_n3668( .i (n969), .o (n3668) );
  assign n3669 = ~n3528 & n3668 ;
  assign n3670 = n3392 & ~n3669 ;
  assign n3671 = n3667 & n3670 ;
  assign n3672 = n955 & n3395 ;
  assign n3673 = n989 & ~n3397 ;
  assign n3674 = n3672 | n3673 ;
  assign n3675 = n3671 | n3674 ;
  assign n3676 = n3389 | n3603 ;
  assign n3677 = ~n3541 & n3668 ;
  assign n3678 = n3392 & ~n3677 ;
  assign n3679 = n3676 & n3678 ;
  assign n3680 = n1008 & n3395 ;
  assign n3681 = n1010 & ~n3397 ;
  assign n3682 = n3680 | n3681 ;
  assign n3683 = n3679 | n3682 ;
  buffer buf_n3684( .i (n3668), .o (n3684) );
  assign n3685 = n3618 | n3684 ;
  assign n3686 = ~n3555 & n3668 ;
  buffer buf_n3687( .i (n974), .o (n3687) );
  assign n3688 = ~n3686 & n3687 ;
  assign n3689 = n3685 & n3688 ;
  buffer buf_n3690( .i (n2956), .o (n3690) );
  assign n3691 = n1007 & n3690 ;
  buffer buf_n3692( .i (n2960), .o (n3692) );
  assign n3693 = n869 & ~n3692 ;
  assign n3694 = n3691 | n3693 ;
  assign n3695 = n3689 | n3694 ;
  assign n3696 = n3430 & ~n3555 ;
  assign n3697 = n3421 | n3616 ;
  assign n3698 = n3433 & n3697 ;
  assign n3699 = ~n3696 & n3698 ;
  buffer buf_n1036( .i (G77), .o (n1036) );
  assign n3700 = n1036 & ~n3436 ;
  buffer buf_n1046( .i (G87), .o (n1046) );
  assign n3701 = n1046 & n3438 ;
  assign n3702 = n3700 | n3701 ;
  assign n3703 = n3699 | n3702 ;
  assign n3704 = n3460 & n3703 ;
  assign n3705 = n3430 & ~n3541 ;
  buffer buf_n3706( .i (n921), .o (n3706) );
  assign n3707 = n3601 | n3706 ;
  assign n3708 = n3433 & n3707 ;
  assign n3709 = ~n3705 & n3708 ;
  buffer buf_n1034( .i (G75), .o (n1034) );
  assign n3710 = n1034 & ~n3436 ;
  buffer buf_n1044( .i (G85), .o (n1044) );
  assign n3711 = n1044 & n3438 ;
  assign n3712 = n3710 | n3711 ;
  assign n3713 = n3709 | n3712 ;
  buffer buf_n3714( .i (n1021), .o (n3714) );
  assign n3715 = n3713 & n3714 ;
  assign n3716 = n3430 & ~n3528 ;
  assign n3717 = n3588 | n3706 ;
  assign n3718 = n3433 & n3717 ;
  assign n3719 = ~n3716 & n3718 ;
  buffer buf_n1043( .i (G84), .o (n1043) );
  assign n3720 = n1043 & n3438 ;
  buffer buf_n1033( .i (G74), .o (n1033) );
  assign n3721 = n1033 & ~n3436 ;
  assign n3722 = n3720 | n3721 ;
  assign n3723 = n3719 | n3722 ;
  assign n3724 = n3714 & n3723 ;
  buffer buf_n3725( .i (n3706), .o (n3725) );
  assign n3726 = n3573 | n3725 ;
  assign n3727 = ~n3511 & n3706 ;
  buffer buf_n3728( .i (n926), .o (n3728) );
  assign n3729 = ~n3727 & n3728 ;
  assign n3730 = n3726 & n3729 ;
  buffer buf_n1032( .i (G73), .o (n1032) );
  buffer buf_n3731( .i (n3302), .o (n3731) );
  assign n3732 = n1032 & ~n3731 ;
  buffer buf_n1042( .i (G83), .o (n1042) );
  buffer buf_n3733( .i (n3306), .o (n3733) );
  assign n3734 = n1042 & n3733 ;
  assign n3735 = n3732 | n3734 ;
  assign n3736 = n3730 | n3735 ;
  assign n3737 = n3714 & n3736 ;
  assign n3738 = n3472 | n3617 ;
  assign n3739 = n3463 & ~n3554 ;
  assign n3740 = n3475 & ~n3739 ;
  assign n3741 = n3738 & n3740 ;
  assign n3742 = n1036 & ~n3478 ;
  assign n3743 = n1046 & n3480 ;
  assign n3744 = n3742 | n3743 ;
  assign n3745 = n3741 | n3744 ;
  assign n3746 = n3714 & n3745 ;
  assign n3747 = n3472 | n3602 ;
  buffer buf_n3748( .i (n930), .o (n3748) );
  assign n3749 = ~n3540 & n3748 ;
  assign n3750 = n3475 & ~n3749 ;
  assign n3751 = n3747 & n3750 ;
  assign n3752 = n1044 & n3480 ;
  assign n3753 = n1034 & ~n3478 ;
  assign n3754 = n3752 | n3753 ;
  assign n3755 = n3751 | n3754 ;
  buffer buf_n3756( .i (n1020), .o (n3756) );
  buffer buf_n3757( .i (n3756), .o (n3757) );
  assign n3758 = n3755 & n3757 ;
  assign n3759 = n3472 & ~n3528 ;
  assign n3760 = n3588 | n3748 ;
  assign n3761 = n3475 & n3760 ;
  assign n3762 = ~n3759 & n3761 ;
  assign n3763 = n1033 & ~n3478 ;
  assign n3764 = n1043 & n3480 ;
  assign n3765 = n3763 | n3764 ;
  assign n3766 = n3762 | n3765 ;
  assign n3767 = n3757 & n3766 ;
  buffer buf_n3768( .i (n3748), .o (n3768) );
  assign n3769 = n3573 | n3768 ;
  assign n3770 = ~n3511 & n3748 ;
  buffer buf_n3771( .i (n935), .o (n3771) );
  assign n3772 = ~n3770 & n3771 ;
  assign n3773 = n3769 & n3772 ;
  buffer buf_n3774( .i (n3317), .o (n3774) );
  assign n3775 = n1032 & ~n3774 ;
  buffer buf_n3776( .i (n3321), .o (n3776) );
  assign n3777 = n1042 & n3776 ;
  assign n3778 = n3775 | n3777 ;
  assign n3779 = n3773 | n3778 ;
  assign n3780 = n3757 & n3779 ;
  assign n3781 = ~n818 & n2403 ;
  buffer buf_n3782( .i (n3781), .o (n3782) );
  buffer buf_n3783( .i (n3782), .o (n3783) );
  assign n3784 = n2447 & ~n3783 ;
  assign n3785 = n819 & ~n2454 ;
  assign n3786 = n3782 | n3785 ;
  assign n3787 = n2405 & ~n2462 ;
  assign n3788 = n3786 & ~n3787 ;
  assign n3789 = n3784 | n3788 ;
  buffer buf_n3790( .i (n3789), .o (n3790) );
  assign n3791 = n3089 & n3790 ;
  assign n3792 = n3089 | n3790 ;
  assign n3793 = ~n3791 & n3792 ;
  assign n3794 = n3244 & ~n3793 ;
  assign n3795 = ~n2408 & n2447 ;
  assign n3796 = n2415 & ~n3795 ;
  buffer buf_n3797( .i (n3796), .o (n3797) );
  assign n3798 = ~n2456 & n2482 ;
  buffer buf_n3799( .i (n2481), .o (n3799) );
  assign n3800 = n2456 & ~n3799 ;
  assign n3801 = n3798 | n3800 ;
  buffer buf_n3802( .i (n3801), .o (n3802) );
  assign n3803 = n3797 & n3802 ;
  assign n3804 = n3797 | n3802 ;
  assign n3805 = ~n3803 & n3804 ;
  assign n3806 = n3244 | n3805 ;
  assign n3807 = ~n3794 & n3806 ;
  buffer buf_n3808( .i (n3807), .o (n3808) );
  buffer buf_n3809( .i (n3808), .o (n3809) );
  buffer buf_n2208( .i (n2207), .o (n2208) );
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n2211( .i (n2210), .o (n2211) );
  buffer buf_n2212( .i (n2211), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  assign n3810 = n2213 & ~n2900 ;
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n2221( .i (n2220), .o (n2221) );
  buffer buf_n2222( .i (n2221), .o (n2222) );
  buffer buf_n2223( .i (n2222), .o (n2223) );
  assign n3811 = ~n2223 & n2900 ;
  assign n3812 = n3810 | n3811 ;
  buffer buf_n3813( .i (n3812), .o (n3813) );
  buffer buf_n937( .i (G162), .o (n937) );
  assign n3814 = n937 & n2281 ;
  assign n3815 = n2262 & n3814 ;
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  assign n3816 = n937 | n2261 ;
  assign n3817 = n2319 & n3816 ;
  assign n3818 = ~n3815 & n3817 ;
  buffer buf_n3819( .i (n3818), .o (n3819) );
  assign n3820 = ~n2225 & n2557 ;
  assign n3821 = n2225 & ~n2557 ;
  assign n3822 = n3820 | n3821 ;
  buffer buf_n3823( .i (n3822), .o (n3823) );
  assign n3824 = n3819 & n3823 ;
  assign n3825 = n3819 | n3823 ;
  assign n3826 = ~n3824 & n3825 ;
  buffer buf_n3827( .i (n3826), .o (n3827) );
  assign n3828 = ~n2373 & n3827 ;
  assign n3829 = n2373 & ~n3827 ;
  assign n3830 = n3828 | n3829 ;
  buffer buf_n3831( .i (n3830), .o (n3831) );
  assign n3832 = n3813 & ~n3831 ;
  assign n3833 = ~n3813 & n3831 ;
  assign n3834 = n3832 | n3833 ;
  buffer buf_n3835( .i (n3834), .o (n3835) );
  buffer buf_n3836( .i (n3835), .o (n3836) );
  assign n3837 = n3809 | n3836 ;
  assign n3838 = n3808 & n3835 ;
  assign n3839 = n3610 | n3838 ;
  assign n3840 = n3837 & ~n3839 ;
  assign n3841 = ~n842 & n1172 ;
  buffer buf_n3842( .i (n181), .o (n3842) );
  assign n3843 = n842 & ~n3842 ;
  assign n3844 = n3841 | n3843 ;
  buffer buf_n3845( .i (n3844), .o (n3845) );
  assign n3846 = ~n1349 & n3845 ;
  assign n3847 = n1349 & ~n3845 ;
  assign n3848 = n3846 | n3847 ;
  buffer buf_n3849( .i (n3848), .o (n3849) );
  assign n3850 = n183 | n386 ;
  assign n3851 = ~n187 & n386 ;
  assign n3852 = n3850 & ~n3851 ;
  assign n3853 = n830 & ~n3852 ;
  assign n3854 = n191 & n386 ;
  buffer buf_n3855( .i (n385), .o (n3855) );
  assign n3856 = n1173 & ~n3855 ;
  assign n3857 = n3854 | n3856 ;
  assign n3858 = ~n830 & n3857 ;
  assign n3859 = n3853 | n3858 ;
  buffer buf_n3860( .i (n3859), .o (n3860) );
  assign n3861 = n3849 | n3860 ;
  assign n3862 = n3849 & n3860 ;
  assign n3863 = n3861 & ~n3862 ;
  buffer buf_n3864( .i (n3863), .o (n3864) );
  assign n3865 = n183 | n541 ;
  assign n3866 = ~n187 & n541 ;
  assign n3867 = n3865 & ~n3866 ;
  assign n3868 = n880 & ~n3867 ;
  assign n3869 = n191 & n541 ;
  buffer buf_n3870( .i (n540), .o (n3870) );
  assign n3871 = n1173 & ~n3870 ;
  assign n3872 = n3869 | n3871 ;
  assign n3873 = ~n880 & n3872 ;
  assign n3874 = n3868 | n3873 ;
  buffer buf_n3875( .i (n3874), .o (n3875) );
  assign n3876 = n183 | n484 ;
  assign n3877 = ~n187 & n484 ;
  assign n3878 = n3876 & ~n3877 ;
  assign n3879 = n860 & ~n3878 ;
  assign n3880 = n191 & n484 ;
  buffer buf_n3881( .i (n483), .o (n3881) );
  assign n3882 = n1173 & ~n3881 ;
  assign n3883 = n3880 | n3882 ;
  assign n3884 = ~n860 & n3883 ;
  assign n3885 = n3879 | n3884 ;
  buffer buf_n3886( .i (n3885), .o (n3886) );
  assign n3887 = n3875 | n3886 ;
  assign n3888 = n3875 & n3886 ;
  assign n3889 = n3887 & ~n3888 ;
  buffer buf_n3890( .i (n3889), .o (n3890) );
  assign n3891 = n3864 | n3890 ;
  assign n3892 = n3864 & n3890 ;
  assign n3893 = n3891 & ~n3892 ;
  buffer buf_n3894( .i (n3893), .o (n3894) );
  buffer buf_n3895( .i (n3894), .o (n3895) );
  assign n3896 = n1254 | n1274 ;
  assign n3897 = ~n1284 & n3896 ;
  buffer buf_n3898( .i (n3897), .o (n3898) );
  assign n3899 = ~n1309 & n1328 ;
  assign n3900 = n1339 | n3899 ;
  buffer buf_n3901( .i (n3900), .o (n3901) );
  assign n3902 = n3898 | n3901 ;
  assign n3903 = n3898 & n3901 ;
  assign n3904 = n3902 & ~n3903 ;
  buffer buf_n3905( .i (n3904), .o (n3905) );
  buffer buf_n3906( .i (n3905), .o (n3906) );
  assign n3907 = n3895 | n3906 ;
  assign n3908 = n3894 & n3905 ;
  assign n3909 = n3609 & ~n3908 ;
  assign n3910 = n3907 & n3909 ;
  assign n3911 = n3583 & ~n3910 ;
  assign n3912 = ~n3840 & n3911 ;
  buffer buf_n3913( .i (n3912), .o (n3913) );
  buffer buf_n3914( .i (n3913), .o (n3914) );
  buffer buf_n3915( .i (n3914), .o (n3915) );
  buffer buf_n3916( .i (n3915), .o (n3916) );
  buffer buf_n3917( .i (n3916), .o (n3917) );
  buffer buf_n3918( .i (n3917), .o (n3918) );
  buffer buf_n3919( .i (n3918), .o (n3919) );
  buffer buf_n2767( .i (n2766), .o (n2767) );
  buffer buf_n2768( .i (n2767), .o (n2768) );
  buffer buf_n2769( .i (n2768), .o (n2769) );
  buffer buf_n2770( .i (n2769), .o (n2770) );
  buffer buf_n2771( .i (n2770), .o (n2771) );
  assign n3920 = ~G51 & n2771 ;
  assign n3921 = ~n3919 & ~n3920 ;
  assign n3922 = n1636 & n1693 ;
  assign n3923 = n1633 | n1704 ;
  assign n3924 = ~n1719 & n3923 ;
  buffer buf_n3925( .i (n3924), .o (n3925) );
  buffer buf_n2662( .i (n2661), .o (n2662) );
  buffer buf_n2663( .i (n2662), .o (n2663) );
  buffer buf_n2664( .i (n2663), .o (n2664) );
  buffer buf_n2665( .i (n2664), .o (n2665) );
  buffer buf_n2666( .i (n2665), .o (n2666) );
  assign n3926 = n1612 | n1691 ;
  assign n3927 = ~n2666 & n3926 ;
  assign n3928 = n3925 | n3927 ;
  assign n3929 = ~n3922 & n3928 ;
  buffer buf_n3930( .i (n3929), .o (n3930) );
  assign n3931 = n2676 & ~n3930 ;
  assign n3932 = ~n2676 & n3930 ;
  assign n3933 = n3931 | n3932 ;
  buffer buf_n3934( .i (n3933), .o (n3934) );
  buffer buf_n3935( .i (n3934), .o (n3935) );
  assign n3936 = n2985 | n3935 ;
  buffer buf_n916( .i (G157), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  assign n3937 = n2984 & n3934 ;
  assign n3938 = n919 | n3937 ;
  assign n3939 = n3936 & ~n3938 ;
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  assign n3940 = n1628 & n1683 ;
  assign n3941 = n1628 | n1693 ;
  assign n3942 = ~n3940 & n3941 ;
  buffer buf_n3943( .i (n3942), .o (n3943) );
  assign n3944 = n3011 & ~n3943 ;
  assign n3945 = ~n3011 & n3943 ;
  assign n3946 = n3944 | n3945 ;
  buffer buf_n3947( .i (n3946), .o (n3947) );
  buffer buf_n3948( .i (n3947), .o (n3948) );
  assign n3949 = n1575 | n3925 ;
  assign n3950 = n1575 & n3925 ;
  assign n3951 = n3949 & ~n3950 ;
  buffer buf_n3952( .i (n3951), .o (n3952) );
  assign n3953 = n1836 | n2978 ;
  buffer buf_n3954( .i (n3953), .o (n3954) );
  assign n3955 = n3952 & ~n3954 ;
  assign n3956 = ~n3952 & n3954 ;
  assign n3957 = n3955 | n3956 ;
  buffer buf_n3958( .i (n3957), .o (n3958) );
  buffer buf_n3959( .i (n3958), .o (n3959) );
  assign n3960 = n3948 & n3959 ;
  assign n3961 = n3947 | n3958 ;
  assign n3962 = n919 & n3961 ;
  assign n3963 = ~n3960 & n3962 ;
  assign n3964 = n3939 | n3963 ;
  buffer buf_n3965( .i (n3964), .o (n3965) );
  buffer buf_n3966( .i (n3965), .o (n3966) );
  buffer buf_n1992( .i (n1991), .o (n1992) );
  buffer buf_n1993( .i (n1992), .o (n1993) );
  buffer buf_n1994( .i (n1993), .o (n1994) );
  buffer buf_n1995( .i (n1994), .o (n1995) );
  assign n3967 = n2158 | n2706 ;
  buffer buf_n3968( .i (n3967), .o (n3968) );
  buffer buf_n3969( .i (n3968), .o (n3969) );
  buffer buf_n3970( .i (n3969), .o (n3970) );
  buffer buf_n3971( .i (n3970), .o (n3971) );
  assign n3972 = ~n1976 & n3971 ;
  assign n3973 = n1995 & ~n3972 ;
  buffer buf_n3974( .i (n3973), .o (n3974) );
  assign n3975 = n1921 | n2056 ;
  assign n3976 = n1921 & n2056 ;
  assign n3977 = n3975 & ~n3976 ;
  buffer buf_n3978( .i (n3977), .o (n3978) );
  buffer buf_n3979( .i (n3978), .o (n3979) );
  buffer buf_n3980( .i (n3979), .o (n3980) );
  buffer buf_n2700( .i (n2699), .o (n2700) );
  buffer buf_n2701( .i (n2700), .o (n2701) );
  buffer buf_n2702( .i (n2701), .o (n2702) );
  buffer buf_n2703( .i (n2702), .o (n2703) );
  buffer buf_n2704( .i (n2703), .o (n2704) );
  assign n3981 = n2106 | n3968 ;
  assign n3982 = ~n2704 & n3981 ;
  buffer buf_n3983( .i (n3982), .o (n3983) );
  assign n3984 = n3980 & n3983 ;
  assign n3985 = n3980 | n3983 ;
  assign n3986 = ~n3984 & n3985 ;
  buffer buf_n3987( .i (n3986), .o (n3987) );
  assign n3988 = n3974 & n3987 ;
  assign n3989 = n3974 | n3987 ;
  assign n3990 = ~n3988 & n3989 ;
  buffer buf_n3991( .i (n3990), .o (n3991) );
  assign n3992 = n2690 & n3991 ;
  assign n3993 = n1974 | n2709 ;
  assign n3994 = ~n2722 & n3993 ;
  buffer buf_n3995( .i (n3994), .o (n3995) );
  buffer buf_n3996( .i (n3995), .o (n3996) );
  assign n3997 = ~n1997 & n2123 ;
  assign n3998 = n1997 & ~n2123 ;
  assign n3999 = n3997 | n3998 ;
  buffer buf_n4000( .i (n3999), .o (n4000) );
  assign n4001 = n3978 & ~n4000 ;
  assign n4002 = ~n3978 & n4000 ;
  assign n4003 = n4001 | n4002 ;
  buffer buf_n4004( .i (n4003), .o (n4004) );
  buffer buf_n4005( .i (n4004), .o (n4005) );
  assign n4006 = n3996 | n4005 ;
  assign n4007 = n3995 & n4004 ;
  assign n4008 = n2686 | n4007 ;
  assign n4009 = n4006 & ~n4008 ;
  buffer buf_n4010( .i (n4009), .o (n4010) );
  buffer buf_n4011( .i (n4010), .o (n4011) );
  assign n4012 = n916 | n4011 ;
  assign n4013 = n3992 | n4012 ;
  assign n4014 = n1847 | n2689 ;
  assign n4015 = n3991 & n4014 ;
  assign n4016 = ~n1847 & n4010 ;
  assign n4017 = n916 & ~n4016 ;
  assign n4018 = ~n4015 & n4017 ;
  assign n4019 = n4013 & ~n4018 ;
  buffer buf_n4020( .i (n4019), .o (n4020) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  buffer buf_n1828( .i (n1827), .o (n1828) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  assign n4021 = n1764 | n1818 ;
  assign n4022 = ~n1833 & n4021 ;
  buffer buf_n4023( .i (n4022), .o (n4023) );
  assign n4024 = n4020 & ~n4023 ;
  assign n4025 = ~n4020 & n4023 ;
  assign n4026 = n4024 | n4025 ;
  buffer buf_n4027( .i (n4026), .o (n4027) );
  buffer buf_n4028( .i (n4027), .o (n4028) );
  assign n4029 = ~n3966 & n4028 ;
  assign n4030 = n3965 & ~n4027 ;
  assign n4031 = n3580 | n4030 ;
  assign n4032 = n4029 | n4031 ;
  assign n4033 = n184 | n1085 ;
  assign n4034 = ~n188 & n1085 ;
  assign n4035 = n4033 & ~n4034 ;
  assign n4036 = n787 & ~n4035 ;
  assign n4037 = n192 & n1085 ;
  buffer buf_n4038( .i (n1084), .o (n4038) );
  assign n4039 = n1174 & ~n4038 ;
  assign n4040 = n4037 | n4039 ;
  assign n4041 = ~n787 & n4040 ;
  assign n4042 = n4036 | n4041 ;
  buffer buf_n4043( .i (n4042), .o (n4043) );
  assign n4044 = n184 | n1113 ;
  assign n4045 = ~n188 & n1113 ;
  assign n4046 = n4044 & ~n4045 ;
  assign n4047 = n810 & ~n4046 ;
  assign n4048 = n192 & n1113 ;
  buffer buf_n4049( .i (n1112), .o (n4049) );
  assign n4050 = n1174 & ~n4049 ;
  assign n4051 = n4048 | n4050 ;
  assign n4052 = ~n810 & n4051 ;
  assign n4053 = n4047 | n4052 ;
  buffer buf_n4054( .i (n4053), .o (n4054) );
  assign n4055 = n4043 & ~n4054 ;
  assign n4056 = ~n4043 & n4054 ;
  assign n4057 = n4055 | n4056 ;
  buffer buf_n4058( .i (n4057), .o (n4058) );
  buffer buf_n4059( .i (n3842), .o (n4059) );
  buffer buf_n4060( .i (n4059), .o (n4060) );
  assign n4061 = n1140 | n4060 ;
  buffer buf_n4062( .i (n185), .o (n4062) );
  buffer buf_n4063( .i (n4062), .o (n4063) );
  buffer buf_n4064( .i (n4063), .o (n4064) );
  assign n4065 = n1140 & ~n4064 ;
  assign n4066 = n4061 & ~n4065 ;
  assign n4067 = n736 & ~n4066 ;
  buffer buf_n4068( .i (n190), .o (n4068) );
  buffer buf_n4069( .i (n4068), .o (n4069) );
  assign n4070 = n1140 & n4069 ;
  buffer buf_n4071( .i (n1139), .o (n4071) );
  buffer buf_n4072( .i (n1171), .o (n4072) );
  buffer buf_n4073( .i (n4072), .o (n4073) );
  buffer buf_n4074( .i (n4073), .o (n4074) );
  assign n4075 = ~n4071 & n4074 ;
  assign n4076 = n4070 | n4075 ;
  assign n4077 = ~n736 & n4076 ;
  assign n4078 = n4067 | n4077 ;
  buffer buf_n4079( .i (n4078), .o (n4079) );
  assign n4080 = n1492 & n4079 ;
  assign n4081 = n1492 | n4079 ;
  assign n4082 = ~n4080 & n4081 ;
  buffer buf_n4083( .i (n4082), .o (n4083) );
  assign n4084 = ~n4058 & n4083 ;
  assign n4085 = n4058 & ~n4083 ;
  assign n4086 = n4084 | n4085 ;
  buffer buf_n4087( .i (n4086), .o (n4087) );
  buffer buf_n4088( .i (n4087), .o (n4088) );
  assign n4089 = n247 | n4060 ;
  assign n4090 = n247 & ~n4064 ;
  assign n4091 = n4089 & ~n4090 ;
  assign n4092 = n712 & ~n4091 ;
  assign n4093 = n247 & n4069 ;
  buffer buf_n4094( .i (n246), .o (n4094) );
  assign n4095 = n4074 & ~n4094 ;
  assign n4096 = n4093 | n4095 ;
  assign n4097 = ~n712 & n4096 ;
  assign n4098 = n4092 | n4097 ;
  buffer buf_n4099( .i (n4098), .o (n4099) );
  assign n4100 = n223 | n4060 ;
  assign n4101 = n223 & ~n4064 ;
  assign n4102 = n4100 & ~n4101 ;
  assign n4103 = n692 & ~n4102 ;
  assign n4104 = n223 & n4069 ;
  buffer buf_n4105( .i (n222), .o (n4105) );
  assign n4106 = n4074 & ~n4105 ;
  assign n4107 = n4104 | n4106 ;
  assign n4108 = ~n692 & n4107 ;
  assign n4109 = n4103 | n4108 ;
  buffer buf_n4110( .i (n4109), .o (n4110) );
  assign n4111 = n4099 & n4110 ;
  assign n4112 = n4099 | n4110 ;
  assign n4113 = ~n4111 & n4112 ;
  buffer buf_n4114( .i (n4113), .o (n4114) );
  assign n4115 = n1162 | n4060 ;
  assign n4116 = n1162 & ~n4064 ;
  assign n4117 = n4115 & ~n4116 ;
  assign n4118 = n753 & ~n4117 ;
  assign n4119 = n1162 & n4069 ;
  buffer buf_n4120( .i (n1161), .o (n4120) );
  assign n4121 = n4074 & ~n4120 ;
  assign n4122 = n4119 | n4121 ;
  assign n4123 = ~n753 & n4122 ;
  assign n4124 = n4118 | n4123 ;
  buffer buf_n4125( .i (n4124), .o (n4125) );
  assign n4126 = n181 | n268 ;
  assign n4127 = ~n185 & n268 ;
  assign n4128 = n4126 & ~n4127 ;
  assign n4129 = n652 & ~n4128 ;
  assign n4130 = n189 & n268 ;
  buffer buf_n4131( .i (n267), .o (n4131) );
  assign n4132 = n1171 & ~n4131 ;
  assign n4133 = n4130 | n4132 ;
  assign n4134 = ~n652 & n4133 ;
  assign n4135 = n4129 | n4134 ;
  buffer buf_n4136( .i (n4135), .o (n4136) );
  assign n4137 = n181 | n200 ;
  assign n4138 = ~n185 & n200 ;
  assign n4139 = n4137 & ~n4138 ;
  assign n4140 = n670 & ~n4139 ;
  assign n4141 = n189 & n200 ;
  buffer buf_n4142( .i (n199), .o (n4142) );
  assign n4143 = n1171 & ~n4142 ;
  assign n4144 = n4141 | n4143 ;
  assign n4145 = ~n670 & n4144 ;
  assign n4146 = n4140 | n4145 ;
  buffer buf_n4147( .i (n4146), .o (n4147) );
  assign n4148 = n4136 & n4147 ;
  assign n4149 = n4136 | n4147 ;
  assign n4150 = ~n4148 & n4149 ;
  buffer buf_n4151( .i (n4150), .o (n4151) );
  assign n4152 = n4125 & ~n4151 ;
  assign n4153 = ~n4125 & n4151 ;
  assign n4154 = n4152 | n4153 ;
  buffer buf_n4155( .i (n4154), .o (n4155) );
  assign n4156 = ~n4114 & n4155 ;
  assign n4157 = n4114 & ~n4155 ;
  assign n4158 = n4156 | n4157 ;
  buffer buf_n4159( .i (n4158), .o (n4159) );
  buffer buf_n4160( .i (n4159), .o (n4160) );
  assign n4161 = ~n4088 & n4160 ;
  assign n4162 = n4087 & ~n4159 ;
  assign n4163 = n3610 & ~n4162 ;
  assign n4164 = ~n4161 & n4163 ;
  assign n4165 = n3523 & ~n4164 ;
  assign n4166 = n4032 & n4165 ;
  buffer buf_n4167( .i (n4166), .o (n4167) );
  buffer buf_n4168( .i (n4167), .o (n4168) );
  buffer buf_n4169( .i (n4168), .o (n4169) );
  buffer buf_n4170( .i (n4169), .o (n4170) );
  buffer buf_n4171( .i (n4170), .o (n4171) );
  buffer buf_n4172( .i (n4171), .o (n4172) );
  assign n4173 = ~G49 & n2771 ;
  assign n4174 = ~n4172 & ~n4173 ;
  buffer buf_n988( .i (n987), .o (n988) );
  assign n4175 = G38 & ~n988 ;
  assign n4176 = n4167 | n4175 ;
  buffer buf_n4177( .i (n4176), .o (n4177) );
  buffer buf_n4178( .i (n4177), .o (n4178) );
  assign n4179 = n3655 | n4178 ;
  assign n4180 = G37 & ~n987 ;
  assign n4181 = n3913 | n4180 ;
  buffer buf_n4182( .i (n4181), .o (n4182) );
  buffer buf_n4183( .i (n4182), .o (n4183) );
  buffer buf_n4184( .i (n965), .o (n4184) );
  assign n4185 = ~n4183 & n4184 ;
  assign n4186 = n3658 & ~n4185 ;
  assign n4187 = n4179 & n4186 ;
  buffer buf_n1001( .i (G23), .o (n1001) );
  assign n4188 = n1001 & ~n3663 ;
  buffer buf_n1009( .i (G4), .o (n1009) );
  assign n4189 = n1009 & n3661 ;
  assign n4190 = n4188 | n4189 ;
  assign n4191 = n4187 | n4190 ;
  assign n4192 = n3684 | n4178 ;
  buffer buf_n4193( .i (n969), .o (n4193) );
  assign n4194 = ~n4183 & n4193 ;
  assign n4195 = n3687 & ~n4194 ;
  assign n4196 = n4192 & n4195 ;
  assign n4197 = n1001 & ~n3692 ;
  assign n4198 = n1009 & n3690 ;
  assign n4199 = n4197 | n4198 ;
  assign n4200 = n4196 | n4199 ;
  assign n4201 = n3725 | n4177 ;
  buffer buf_n4202( .i (n921), .o (n4202) );
  assign n4203 = ~n4182 & n4202 ;
  assign n4204 = n3728 & ~n4203 ;
  assign n4205 = n4201 & n4204 ;
  buffer buf_n1038( .i (G79), .o (n1038) );
  assign n4206 = n1038 & ~n3731 ;
  buffer buf_n1037( .i (G78), .o (n1037) );
  assign n4207 = n1037 & n3733 ;
  assign n4208 = n4206 | n4207 ;
  assign n4209 = n4205 | n4208 ;
  assign n4210 = ~n3757 | ~n4209 ;
  assign n4211 = n3768 | n4177 ;
  buffer buf_n4212( .i (n930), .o (n4212) );
  assign n4213 = ~n4182 & n4212 ;
  assign n4214 = n3771 & ~n4213 ;
  assign n4215 = n4211 & n4214 ;
  assign n4216 = n1038 & ~n3774 ;
  assign n4217 = n1037 & n3776 ;
  assign n4218 = n4216 | n4217 ;
  assign n4219 = n4215 | n4218 ;
  buffer buf_n4220( .i (n3756), .o (n4220) );
  assign n4221 = ~n4219 | ~n4220 ;
  assign G5193 = n1026 ;
  assign G5194 = n312 ;
  assign G5195 = n942 ;
  assign G5196 = n889 ;
  assign G5197 = n529 ;
  assign G5198 = n640 ;
  assign G5199 = n1189 ;
  assign G5200 = n891 ;
  assign G5201 = n889 ;
  assign G5202 = n889 ;
  assign G5203 = n474 ;
  assign G5204 = n588 ;
  assign G5205 = n1190 ;
  assign G5206 = n1182 ;
  assign G5207 = n899 ;
  assign G5208 = n915 ;
  assign G5209 = n907 ;
  assign G5210 = n1191 ;
  assign G5211 = n1192 ;
  assign G5212 = n1193 ;
  assign G5213 = n1201 ;
  assign G5214 = n1023 ;
  assign G5215 = n4222 ;
  assign G5216 = n180 ;
  assign G5217 = n4223 ;
  assign G5218 = n337 ;
  assign G5219 = n4223 ;
  assign G5220 = n1208 ;
  assign G5221 = n1207 ;
  assign G5222 = n4224 ;
  assign G5223 = n4224 ;
  assign G5224 = n4224 ;
  assign G5225 = n4224 ;
  assign G5226 = n4225 ;
  assign G5227 = n4225 ;
  assign G5228 = n1212 ;
  assign G5229 = n1217 ;
  assign G5230 = n1217 ;
  assign G5231 = n1218 ;
  assign G5232 = n1223 ;
  assign G5233 = n1229 ;
  assign G5234 = n1236 ;
  assign G5235 = n1242 ;
  assign G5236 = n1403 ;
  assign G5237 = n1539 ;
  assign G5238 = n2187 ;
  assign G5239 = n2581 ;
  assign G5240 = n2581 ;
  assign G5241 = n2187 ;
  assign G5242 = n2617 ;
  assign G5243 = n2659 ;
  assign G5244 = n2747 ;
  assign G5245 = n2760 ;
  assign G5246 = n2747 ;
  assign G5247 = n2760 ;
  assign G5248 = n2787 ;
  assign G5249 = n2806 ;
  assign G5250 = n2830 ;
  assign G5251 = n2842 ;
  assign G5252 = n2856 ;
  assign G5253 = n2897 ;
  assign G5254 = n2927 ;
  assign G5255 = n2950 ;
  assign G5256 = n2964 ;
  assign G5257 = n3005 ;
  assign G5258 = n3039 ;
  assign G5259 = n3070 ;
  assign G5260 = n3085 ;
  assign G5261 = n3136 ;
  assign G5262 = n3177 ;
  assign G5263 = n3239 ;
  assign G5264 = n3296 ;
  assign G5265 = n3311 ;
  assign G5266 = n3326 ;
  assign G5267 = n3334 ;
  assign G5268 = n3342 ;
  assign G5269 = n3351 ;
  assign G5270 = n3363 ;
  assign G5271 = n3371 ;
  assign G5272 = n3379 ;
  assign G5273 = n3388 ;
  assign G5274 = n3400 ;
  assign G5275 = n3409 ;
  assign G5276 = n3419 ;
  assign G5277 = n3429 ;
  assign G5278 = n3442 ;
  assign G5279 = n3451 ;
  assign G5280 = n3461 ;
  assign G5281 = n3471 ;
  assign G5282 = n3484 ;
  assign G5283 = n3501 ;
  assign G5284 = n3504 ;
  assign G5285 = n3516 ;
  assign G5286 = n3532 ;
  assign G5287 = n3545 ;
  assign G5288 = n3559 ;
  assign G5289 = n3566 ;
  assign G5290 = n3577 ;
  assign G5291 = n3593 ;
  assign G5292 = n3606 ;
  assign G5293 = n3621 ;
  assign G5294 = n3629 ;
  assign G5295 = n3637 ;
  assign G5296 = n3646 ;
  assign G5297 = n3654 ;
  assign G5298 = n3666 ;
  assign G5299 = n3675 ;
  assign G5300 = n3683 ;
  assign G5301 = n3695 ;
  assign G5302 = n3704 ;
  assign G5303 = n3715 ;
  assign G5304 = n3724 ;
  assign G5305 = n3737 ;
  assign G5306 = n3746 ;
  assign G5307 = n3758 ;
  assign G5308 = n3767 ;
  assign G5309 = n3780 ;
  assign G5310 = n3921 ;
  assign G5311 = n4174 ;
  assign G5312 = n4191 ;
  assign G5313 = n4200 ;
  assign G5314 = n4210 ;
  assign G5315 = n4221 ;
endmodule
