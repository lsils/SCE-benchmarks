module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 ;
  buffer buf_n418( .i (x13), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n515( .i (x16), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n549( .i (x17), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n450( .i (x14), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n603( .i (x19), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n580( .i (x18), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n630( .i (x20), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n676( .i (x22), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n652( .i (x21), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n697( .i (x23), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n720( .i (x24), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n763( .i (x26), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  assign n841 = n710 & ~n776 ;
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  assign n847 = ( n714 & ~n737 ) | ( n714 & n844 ) | ( ~n737 & n844 ) ;
  assign n848 = ~n670 & n847 ;
  assign n849 = ( n649 & ~n695 ) | ( n649 & n848 ) | ( ~n695 & n848 ) ;
  assign n850 = ~n650 & n849 ;
  assign n851 = ~n601 & n850 ;
  assign n852 = ~n625 & n851 ;
  assign n853 = n473 & n852 ;
  assign n854 = ( n539 & n573 ) | ( n539 & n853 ) | ( n573 & n853 ) ;
  assign n855 = ~n574 & n854 ;
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n351( .i (x11), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n93( .i (x2), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  assign n858 = n119 & n444 ;
  assign n859 = ( n378 & ~n856 ) | ( n378 & n858 ) | ( ~n856 & n858 ) ;
  assign n860 = n857 & n859 ;
  buffer buf_n861( .i (n860), .o (n861) );
  assign n862 = ( n448 & ~n545 ) | ( n448 & n861 ) | ( ~n545 & n861 ) ;
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  assign n863 = n381 & ~n861 ;
  assign n864 = ( n449 & ~n862 ) | ( n449 & n863 ) | ( ~n862 & n863 ) ;
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n384( .i (x12), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n156( .i (x4), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n482( .i (x15), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  assign n867 = ~n188 & n514 ;
  assign n868 = ( n417 & n865 ) | ( n417 & n867 ) | ( n865 & n867 ) ;
  assign n869 = ~n866 & n868 ;
  assign n870 = ~n676 & n763 ;
  assign n871 = ( n653 & n698 ) | ( n653 & n870 ) | ( n698 & n870 ) ;
  assign n872 = ~n654 & n871 ;
  assign n873 = ~n606 & n872 ;
  assign n874 = ( n584 & ~n634 ) | ( n584 & n873 ) | ( ~n634 & n873 ) ;
  assign n875 = ~n585 & n874 ;
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  assign n878 = n419 & n451 ;
  assign n879 = ( n484 & n551 ) | ( n484 & n878 ) | ( n551 & n878 ) ;
  assign n880 = ~n552 & n879 ;
  assign n881 = n388 & n880 ;
  assign n882 = ( n98 & n356 ) | ( n98 & n881 ) | ( n356 & n881 ) ;
  assign n883 = ~n99 & n882 ;
  assign n884 = ( n522 & ~n876 ) | ( n522 & n883 ) | ( ~n876 & n883 ) ;
  assign n885 = n389 | n455 ;
  assign n886 = n356 | n487 ;
  assign n887 = ( ~n390 & n885 ) | ( ~n390 & n886 ) | ( n885 & n886 ) ;
  assign n888 = n522 & ~n887 ;
  assign n889 = ( n877 & n884 ) | ( n877 & n888 ) | ( n884 & n888 ) ;
  assign n890 = ~n165 & n889 ;
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n122( .i (x3), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n742( .i (x25), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  assign n916 = ( n104 & n753 ) | ( n104 & n774 ) | ( n753 & n774 ) ;
  buffer buf_n917( .i (n916), .o (n917) );
  assign n918 = n733 | n917 ;
  assign n919 = n666 & ~n918 ;
  assign n920 = ( n691 & n712 ) | ( n691 & n919 ) | ( n712 & n919 ) ;
  assign n921 = ~n713 & n920 ;
  assign n922 = ~n620 & n921 ;
  assign n923 = ( n598 & ~n648 ) | ( n598 & n922 ) | ( ~n648 & n922 ) ;
  assign n924 = ~n599 & n923 ;
  assign n925 = ~n569 & n924 ;
  assign n926 = ( ~n405 & n503 ) | ( ~n405 & n925 ) | ( n503 & n925 ) ;
  assign n927 = n406 & ~n926 ;
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  assign n930 = ~n404 & n502 ;
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  assign n937 = ( ~n117 & n928 ) | ( ~n117 & n933 ) | ( n928 & n933 ) ;
  assign n938 = n929 | n937 ;
  assign n939 = n541 & ~n938 ;
  assign n940 = n445 & ~n939 ;
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  assign n941 = n445 | n936 ;
  assign n942 = ~n940 & n941 ;
  assign n943 = n380 & ~n942 ;
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  assign n944 = n508 & n541 ;
  assign n945 = n410 | n444 ;
  assign n946 = ( n509 & ~n944 ) | ( n509 & n945 ) | ( ~n944 & n945 ) ;
  assign n947 = n121 & ~n946 ;
  assign n948 = n380 | n947 ;
  assign n949 = ~n943 & n948 ;
  assign n950 = n481 & ~n949 ;
  assign n951 = ( ~n407 & n441 ) | ( ~n407 & n505 ) | ( n441 & n505 ) ;
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  assign n956 = ~n507 & n952 ;
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  assign n959 = ( n411 & n542 ) | ( n411 & n957 ) | ( n542 & n957 ) ;
  assign n960 = ( n955 & n958 ) | ( n955 & n959 ) | ( n958 & n959 ) ;
  assign n961 = ~n409 & n540 ;
  assign n962 = ~n508 & n961 ;
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  assign n965 = n121 | n963 ;
  assign n966 = ( n960 & n964 ) | ( n960 & n965 ) | ( n964 & n965 ) ;
  assign n967 = ~n381 & n966 ;
  assign n968 = n481 | n967 ;
  assign n969 = ~n950 & n968 ;
  assign n970 = n155 & n969 ;
  assign n971 = ~n190 & n970 ;
  assign n972 = n440 & n537 ;
  buffer buf_n973( .i (n972), .o (n973) );
  assign n974 = n506 & n973 ;
  buffer buf_n975( .i (n974), .o (n975) );
  assign n982 = ~n699 & n765 ;
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  assign n994 = n690 | n993 ;
  assign n995 = ~n709 & n732 ;
  buffer buf_n996( .i (n995), .o (n996) );
  assign n998 = ( n690 & n993 ) | ( n690 & n996 ) | ( n993 & n996 ) ;
  assign n999 = n994 & ~n998 ;
  buffer buf_n293( .i (x9), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  assign n1000 = ~n305 & n709 ;
  assign n1001 = ~n689 & n1000 ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  assign n1004 = n757 & ~n1002 ;
  assign n1005 = ( n999 & n1003 ) | ( n999 & ~n1004 ) | ( n1003 & ~n1004 ) ;
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  assign n1008 = ( n111 & n670 ) | ( n111 & n1006 ) | ( n670 & n1006 ) ;
  assign n1009 = n303 & ~n686 ;
  assign n1010 = n303 | n730 ;
  assign n1011 = ( n774 & n1009 ) | ( n774 & n1010 ) | ( n1009 & n1010 ) ;
  assign n1012 = n105 & ~n1011 ;
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  assign n1015 = n690 | n1013 ;
  assign n1016 = ( ~n735 & n1014 ) | ( ~n735 & n1015 ) | ( n1014 & n1015 ) ;
  assign n1017 = n713 & n1016 ;
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  assign n1018 = n688 & n775 ;
  assign n1019 = ( n689 & ~n755 ) | ( n689 & n1018 ) | ( ~n755 & n1018 ) ;
  assign n1020 = ( n307 & n734 ) | ( n307 & n1019 ) | ( n734 & n1019 ) ;
  assign n1021 = ( ~n105 & n688 ) | ( ~n105 & n775 ) | ( n688 & n775 ) ;
  assign n1022 = n917 & ~n1021 ;
  assign n1023 = n734 & n1022 ;
  assign n1024 = ( ~n308 & n1020 ) | ( ~n308 & n1023 ) | ( n1020 & n1023 ) ;
  assign n1025 = n713 | n1024 ;
  assign n1026 = ( ~n714 & n1017 ) | ( ~n714 & n1025 ) | ( n1017 & n1025 ) ;
  assign n1027 = ~n670 & n1026 ;
  assign n1028 = ( n1007 & ~n1008 ) | ( n1007 & n1027 ) | ( ~n1008 & n1027 ) ;
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n777( .i (n776), .o (n777) );
  assign n1031 = ~n307 & n777 ;
  assign n1032 = ~n757 & n1031 ;
  assign n1033 = n109 & n1032 ;
  buffer buf_n778( .i (n777), .o (n778) );
  assign n1034 = n710 & n755 ;
  assign n1035 = n777 & n1034 ;
  assign n1036 = ( n778 & n842 ) | ( n778 & ~n1035 ) | ( n842 & ~n1035 ) ;
  assign n1037 = ~n109 & n1036 ;
  assign n1038 = ( n669 & n1033 ) | ( n669 & ~n1037 ) | ( n1033 & ~n1037 ) ;
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  assign n1041 = ( n695 & n739 ) | ( n695 & n1039 ) | ( n739 & n1039 ) ;
  assign n1042 = n94 | n764 ;
  buffer buf_n1043( .i (n1042), .o (n1043) );
  assign n1061 = n655 | n1043 ;
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n1076( .i (n712), .o (n1076) );
  assign n1077 = n758 & ~n1076 ;
  assign n1078 = ( n737 & ~n1074 ) | ( n737 & n1077 ) | ( ~n1074 & n1077 ) ;
  assign n1079 = n1075 & n1078 ;
  assign n1080 = ~n695 & n1079 ;
  assign n1081 = ( n1040 & ~n1041 ) | ( n1040 & n1080 ) | ( ~n1041 & n1080 ) ;
  assign n1082 = ~n1029 & n1081 ;
  buffer buf_n651( .i (n650), .o (n651) );
  assign n1083 = n624 | n651 ;
  assign n1084 = ( n1030 & n1082 ) | ( n1030 & ~n1083 ) | ( n1082 & ~n1083 ) ;
  buffer buf_n602( .i (n601), .o (n602) );
  assign n1085 = n472 & ~n602 ;
  assign n1086 = ( n572 & n1084 ) | ( n572 & n1085 ) | ( n1084 & n1085 ) ;
  assign n1087 = ~n573 & n1086 ;
  assign n1088 = n376 & n1087 ;
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  assign n1089 = n318 & ~n376 ;
  assign n1090 = ( n975 & ~n1088 ) | ( n975 & n1089 ) | ( ~n1088 & n1089 ) ;
  buffer buf_n218( .i (x6), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (x7), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  assign n1091 = ~n369 & n533 ;
  buffer buf_n1092( .i (n1091), .o (n1092) );
  assign n1095 = ( n433 & n465 ) | ( n433 & n530 ) | ( n465 & n530 ) ;
  buffer buf_n1096( .i (n1095), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  assign n1098 = ~n652 & n742 ;
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  assign n1102 = n96 & n655 ;
  assign n1103 = ( n724 & n1101 ) | ( n724 & ~n1102 ) | ( n1101 & ~n1102 ) ;
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  assign n1106 = n769 & ~n1104 ;
  assign n1107 = n655 & n745 ;
  assign n1108 = n724 & n1107 ;
  buffer buf_n1109( .i (n1108), .o (n1109) );
  assign n1121 = ~n722 & n744 ;
  assign n1122 = ~n653 & n764 ;
  assign n1123 = n744 | n1122 ;
  assign n1124 = ~n1121 & n1123 ;
  assign n1125 = ( ~n97 & n519 ) | ( ~n97 & n1124 ) | ( n519 & n1124 ) ;
  assign n1126 = n721 & n764 ;
  assign n1127 = ( ~n722 & n1099 ) | ( ~n722 & n1126 ) | ( n1099 & n1126 ) ;
  buffer buf_n1128( .i (n1127), .o (n1128) );
  assign n1131 = ( n97 & n519 ) | ( n97 & n1128 ) | ( n519 & n1128 ) ;
  assign n1132 = n1125 & n1131 ;
  assign n1133 = n1109 | n1132 ;
  assign n1134 = ( n1105 & n1106 ) | ( n1105 & ~n1133 ) | ( n1106 & ~n1133 ) ;
  assign n1135 = n98 & ~n725 ;
  assign n1136 = n658 & n1135 ;
  buffer buf_n1137( .i (n1136), .o (n1137) );
  assign n1138 = ( n705 & n1134 ) | ( n705 & ~n1137 ) | ( n1134 & ~n1137 ) ;
  assign n1139 = n744 & n765 ;
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  assign n1155 = ( ~n657 & n725 ) | ( ~n657 & n1062 ) | ( n725 & n1062 ) ;
  assign n1156 = n1142 & n1155 ;
  assign n1157 = ( n1064 & ~n1143 ) | ( n1064 & n1156 ) | ( ~n1143 & n1156 ) ;
  assign n1158 = ( n705 & n1137 ) | ( n705 & ~n1157 ) | ( n1137 & ~n1157 ) ;
  assign n1159 = n1138 & ~n1158 ;
  buffer buf_n1160( .i (n1159), .o (n1160) );
  buffer buf_n1161( .i (n1160), .o (n1161) );
  assign n1162 = ( n641 & n687 ) | ( n641 & ~n1160 ) | ( n687 & ~n1160 ) ;
  assign n1163 = n96 & ~n766 ;
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  assign n1177 = n725 & ~n1164 ;
  assign n1178 = ( n748 & ~n1165 ) | ( n748 & n1177 ) | ( ~n1165 & n1177 ) ;
  assign n1179 = n704 & ~n1178 ;
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n1181( .i (n1180), .o (n1181) );
  assign n1182 = ( n661 & ~n685 ) | ( n661 & n1180 ) | ( ~n685 & n1180 ) ;
  buffer buf_n1183( .i (n743), .o (n1183) );
  assign n1184 = ( n699 & ~n722 ) | ( n699 & n1183 ) | ( ~n722 & n1183 ) ;
  buffer buf_n1185( .i (n1184), .o (n1185) );
  assign n1186 = n746 & ~n1185 ;
  assign n1187 = ( n724 & n983 ) | ( n724 & n1185 ) | ( n983 & n1185 ) ;
  assign n1188 = ( n702 & n1186 ) | ( n702 & ~n1187 ) | ( n1186 & ~n1187 ) ;
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  assign n1191 = ( n100 & ~n683 ) | ( n100 & n1189 ) | ( ~n683 & n1189 ) ;
  buffer buf_n1192( .i (n723), .o (n1192) );
  assign n1193 = n767 | n1192 ;
  assign n1194 = ( ~n702 & n747 ) | ( ~n702 & n1193 ) | ( n747 & n1193 ) ;
  assign n1195 = n703 | n1194 ;
  assign n1196 = n100 | n1195 ;
  assign n1197 = ( ~n1190 & n1191 ) | ( ~n1190 & n1196 ) | ( n1191 & n1196 ) ;
  assign n1198 = n661 | n1197 ;
  assign n1199 = ( ~n1181 & n1182 ) | ( ~n1181 & n1198 ) | ( n1182 & n1198 ) ;
  assign n1200 = n641 | n1199 ;
  assign n1201 = ( n1161 & n1162 ) | ( n1161 & n1200 ) | ( n1162 & n1200 ) ;
  assign n1202 = n593 | n1201 ;
  assign n1203 = ( ~n563 & n617 ) | ( ~n563 & n1202 ) | ( n617 & n1202 ) ;
  assign n1204 = n564 | n1203 ;
  assign n1205 = ( ~n434 & n531 ) | ( ~n434 & n1204 ) | ( n531 & n1204 ) ;
  assign n1206 = n1096 & n1205 ;
  assign n1207 = ( ~n468 & n1097 ) | ( ~n468 & n1206 ) | ( n1097 & n1206 ) ;
  assign n1208 = n370 & ~n1207 ;
  assign n1209 = ( n502 & n1092 ) | ( n502 & ~n1208 ) | ( n1092 & ~n1208 ) ;
  assign n1210 = n264 & ~n1209 ;
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  assign n1213 = n745 & ~n766 ;
  assign n1214 = ( n767 & n1192 ) | ( n767 & ~n1213 ) | ( n1192 & ~n1213 ) ;
  assign n1215 = n657 & n1214 ;
  assign n1216 = n765 & ~n1183 ;
  assign n1217 = ( n723 & n766 ) | ( n723 & n1216 ) | ( n766 & n1216 ) ;
  assign n1218 = n97 & n1217 ;
  assign n1219 = n657 | n1218 ;
  assign n1220 = ~n1215 & n1219 ;
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  assign n1223 = n705 & n1221 ;
  buffer buf_n1224( .i (n656), .o (n1224) );
  assign n1225 = ~n768 & n1224 ;
  assign n1226 = ( n99 & n726 ) | ( n99 & n1225 ) | ( n726 & n1225 ) ;
  assign n1227 = ~n727 & n1226 ;
  buffer buf_n1228( .i (n654), .o (n1228) );
  assign n1229 = n723 & n1228 ;
  assign n1230 = ( n656 & ~n1140 ) | ( n656 & n1229 ) | ( ~n1140 & n1229 ) ;
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  assign n1233 = ( ~n99 & n703 ) | ( ~n99 & n1231 ) | ( n703 & n1231 ) ;
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1234( .i (n98), .o (n1234) );
  assign n1235 = n1130 & ~n1234 ;
  assign n1236 = ( ~n1232 & n1233 ) | ( ~n1232 & n1235 ) | ( n1233 & n1235 ) ;
  assign n1237 = n1227 | n1236 ;
  assign n1238 = ( n1222 & ~n1223 ) | ( n1222 & n1237 ) | ( ~n1223 & n1237 ) ;
  assign n1239 = ~n686 & n1238 ;
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  assign n1242 = ( ~n100 & n727 ) | ( ~n100 & n770 ) | ( n727 & n770 ) ;
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  assign n1245 = n102 & n1243 ;
  assign n1246 = ( n752 & n1244 ) | ( n752 & n1245 ) | ( n1244 & n1245 ) ;
  assign n1247 = n745 | n1043 ;
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  assign n1263 = ( n702 & n1141 ) | ( n702 & n1248 ) | ( n1141 & n1248 ) ;
  assign n1264 = n726 & n1263 ;
  assign n1265 = ( ~n727 & n1250 ) | ( ~n727 & n1264 ) | ( n1250 & n1264 ) ;
  assign n1266 = n684 & ~n1265 ;
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  assign n1269 = n707 | n1267 ;
  assign n1270 = ( ~n1246 & n1268 ) | ( ~n1246 & n1269 ) | ( n1268 & n1269 ) ;
  assign n1271 = n1240 | n1270 ;
  assign n1272 = ( ~n665 & n1241 ) | ( ~n665 & n1271 ) | ( n1241 & n1271 ) ;
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  assign n1275 = n593 | n643 ;
  buffer buf_n1276( .i (n1275), .o (n1276) );
  assign n1288 = ( n618 & n1273 ) | ( n618 & n1276 ) | ( n1273 & n1276 ) ;
  assign n1289 = n1274 & ~n1288 ;
  assign n1290 = n499 & n1289 ;
  assign n1291 = ( n533 & n567 ) | ( n533 & n1290 ) | ( n567 & n1290 ) ;
  assign n1292 = ~n568 & n1291 ;
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  assign n1295 = n371 & n470 ;
  assign n1296 = ( n439 & ~n1293 ) | ( n439 & n1295 ) | ( ~n1293 & n1295 ) ;
  assign n1297 = n1294 & n1296 ;
  assign n1298 = n1211 | n1297 ;
  assign n1299 = ( n242 & n1212 ) | ( n242 & n1298 ) | ( n1212 & n1298 ) ;
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n191( .i (x5), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  assign n1302 = n217 | n1300 ;
  assign n1303 = ( ~n1090 & n1301 ) | ( ~n1090 & n1302 ) | ( n1301 & n1302 ) ;
  assign n1304 = ( n469 & ~n501 ) | ( n469 & n534 ) | ( ~n501 & n534 ) ;
  assign n1305 = ( ~n437 & n469 ) | ( ~n437 & n501 ) | ( n469 & n501 ) ;
  assign n1306 = ~n1304 & n1305 ;
  assign n1307 = n211 & ~n371 ;
  assign n1308 = ( n314 & n1306 ) | ( n314 & n1307 ) | ( n1306 & n1307 ) ;
  assign n1309 = ~n315 & n1308 ;
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  assign n1313 = n472 & ~n504 ;
  assign n1314 = ~n538 & n1313 ;
  assign n1315 = ( n267 & n1310 ) | ( n267 & n1314 ) | ( n1310 & n1314 ) ;
  assign n1316 = n443 & ~n1315 ;
  assign n1317 = ( n444 & n1312 ) | ( n444 & ~n1316 ) | ( n1312 & ~n1316 ) ;
  buffer buf_n1318( .i (n1317), .o (n1318) );
  assign n1319 = ( n412 & n1303 ) | ( n412 & n1318 ) | ( n1303 & n1318 ) ;
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  assign n1320 = ( n370 & ~n501 ) | ( n370 & n534 ) | ( ~n501 & n534 ) ;
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  assign n1323 = ( n472 & n1094 ) | ( n472 & ~n1322 ) | ( n1094 & ~n1322 ) ;
  assign n1324 = n214 & n1323 ;
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  assign n1327 = ( n241 & n473 ) | ( n241 & n538 ) | ( n473 & n538 ) ;
  assign n1328 = n266 & n473 ;
  assign n1329 = ( ~n539 & n1327 ) | ( ~n539 & n1328 ) | ( n1327 & n1328 ) ;
  assign n1330 = n1325 | n1329 ;
  assign n1331 = ( ~n377 & n1326 ) | ( ~n377 & n1330 ) | ( n1326 & n1330 ) ;
  assign n1332 = ( ~n313 & n371 ) | ( ~n313 & n535 ) | ( n371 & n535 ) ;
  buffer buf_n1333( .i (n370), .o (n1333) );
  assign n1334 = ( n313 & ~n438 ) | ( n313 & n1333 ) | ( ~n438 & n1333 ) ;
  assign n1335 = n1332 & ~n1334 ;
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n471), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  assign n1340 = ( ~n214 & n1336 ) | ( ~n214 & n1339 ) | ( n1336 & n1339 ) ;
  assign n1341 = ( ~n438 & n502 ) | ( ~n438 & n535 ) | ( n502 & n535 ) ;
  assign n1342 = ~n1321 & n1341 ;
  buffer buf_n274( .i (x8), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  assign n1343 = n368 & ~n499 ;
  assign n1344 = ( n292 & n436 ) | ( n292 & n1343 ) | ( n436 & n1343 ) ;
  assign n1345 = ~n437 & n1344 ;
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  assign n1348 = n264 | n1346 ;
  assign n1349 = ( n1342 & n1347 ) | ( n1342 & n1348 ) | ( n1347 & n1348 ) ;
  assign n1350 = ~n1339 & n1349 ;
  assign n1351 = ( n1337 & ~n1340 ) | ( n1337 & n1350 ) | ( ~n1340 & n1350 ) ;
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n443), .o (n1354) );
  assign n1355 = n1352 | n1354 ;
  assign n1356 = ( n1331 & n1353 ) | ( n1331 & n1355 ) | ( n1353 & n1355 ) ;
  assign n1357 = ( ~n412 & n1318 ) | ( ~n412 & n1356 ) | ( n1318 & n1356 ) ;
  assign n1358 = n1319 | n1357 ;
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n319( .i (x10), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  assign n1361 = ( n187 & ~n350 ) | ( n187 & n1359 ) | ( ~n350 & n1359 ) ;
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n780( .i (x27), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (x28), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  assign n1362 = n272 & n840 ;
  assign n1363 = ( n273 & n810 ) | ( n273 & n1362 ) | ( n810 & n1362 ) ;
  assign n1364 = n350 & n1363 ;
  assign n1365 = ( n1360 & ~n1361 ) | ( n1360 & n1364 ) | ( ~n1361 & n1364 ) ;
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n30( .i (x0), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  assign n1368 = n471 & n503 ;
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  assign n1371 = ~n729 & n1252 ;
  assign n1372 = ( n1146 & n1253 ) | ( n1146 & n1371 ) | ( n1253 & n1371 ) ;
  assign n1373 = n687 & ~n1372 ;
  assign n1374 = ~n709 & n1373 ;
  assign n1375 = ~n643 & n1374 ;
  assign n1376 = ( n617 & ~n666 ) | ( n617 & n1375 ) | ( ~n666 & n1375 ) ;
  assign n1377 = ~n618 & n1376 ;
  assign n1378 = n530 & ~n595 ;
  assign n1379 = ( n565 & n1377 ) | ( n565 & n1378 ) | ( n1377 & n1378 ) ;
  assign n1380 = ~n566 & n1379 ;
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  assign n1383 = n367 & n434 ;
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  assign n1386 = ( n403 & ~n1381 ) | ( n403 & n1385 ) | ( ~n1381 & n1385 ) ;
  assign n1387 = n1382 & n1386 ;
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n997( .i (n996), .o (n997) );
  assign n1390 = n691 & n997 ;
  assign n1391 = ~n646 & n1390 ;
  assign n1392 = ( n620 & ~n669 ) | ( n620 & n1391 ) | ( ~n669 & n1391 ) ;
  assign n1393 = ~n621 & n1392 ;
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  assign n1396 = n530 & ~n564 ;
  assign n1397 = ~n596 & n1396 ;
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  assign n1400 = ( n402 & n1384 ) | ( n402 & ~n1398 ) | ( n1384 & ~n1398 ) ;
  assign n1401 = n1399 & n1400 ;
  assign n1402 = ( n313 & n1394 ) | ( n313 & ~n1401 ) | ( n1394 & ~n1401 ) ;
  assign n1403 = n401 | n532 ;
  assign n1404 = ( ~n369 & n436 ) | ( ~n369 & n1403 ) | ( n436 & n1403 ) ;
  buffer buf_n1405( .i (n369), .o (n1405) );
  assign n1406 = n1404 | n1405 ;
  buffer buf_n1407( .i (n312), .o (n1407) );
  assign n1408 = n1406 | n1407 ;
  assign n1409 = ( ~n1395 & n1402 ) | ( ~n1395 & n1408 ) | ( n1402 & n1408 ) ;
  assign n1410 = n1388 | n1409 ;
  assign n1411 = ( n1369 & n1389 ) | ( n1369 & ~n1410 ) | ( n1389 & ~n1410 ) ;
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  assign n1415 = ( ~n442 & n973 ) | ( ~n442 & n1370 ) | ( n973 & n1370 ) ;
  assign n1416 = ( n409 & ~n1412 ) | ( n409 & n1415 ) | ( ~n1412 & n1415 ) ;
  assign n1417 = n377 & n1416 ;
  assign n1418 = ( n378 & n1414 ) | ( n378 & ~n1417 ) | ( n1414 & ~n1417 ) ;
  assign n1419 = n58 & n1418 ;
  assign n1420 = ~n185 & n1419 ;
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n59( .i (x1), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  assign n1426 = ( ~n411 & n477 ) | ( ~n411 & n509 ) | ( n477 & n509 ) ;
  assign n1427 = n543 & ~n1426 ;
  assign n1428 = ( n413 & ~n544 ) | ( n413 & n1427 ) | ( ~n544 & n1427 ) ;
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  assign n1431 = ~n447 & n544 ;
  assign n1432 = n479 | n511 ;
  assign n1433 = ( n448 & n1431 ) | ( n448 & ~n1432 ) | ( n1431 & ~n1432 ) ;
  assign n1434 = ( n144 & n373 ) | ( n144 & n931 ) | ( n373 & n931 ) ;
  assign n1435 = ~n145 & n1434 ;
  buffer buf_n1436( .i (n1435), .o (n1436) );
  assign n1437 = ( n507 & n540 ) | ( n507 & ~n1436 ) | ( n540 & ~n1436 ) ;
  assign n1438 = n376 & ~n1436 ;
  assign n1439 = ( ~n541 & n1437 ) | ( ~n541 & n1438 ) | ( n1437 & n1438 ) ;
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  assign n1442 = ( ~n446 & n478 ) | ( ~n446 & n1440 ) | ( n478 & n1440 ) ;
  assign n1443 = n685 & ~n706 ;
  assign n1444 = ~n773 & n1443 ;
  assign n1445 = ~n132 & n662 ;
  assign n1446 = ( n104 & n1444 ) | ( n104 & n1445 ) | ( n1444 & n1445 ) ;
  assign n1447 = ~n105 & n1446 ;
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n689), .o (n1451) );
  assign n1452 = ( n666 & ~n1448 ) | ( n666 & n1451 ) | ( ~n1448 & n1451 ) ;
  assign n1453 = n712 & n1452 ;
  assign n1454 = ( n1076 & n1450 ) | ( n1076 & ~n1453 ) | ( n1450 & ~n1453 ) ;
  buffer buf_n1455( .i (n1454), .o (n1455) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  assign n1457 = ( n648 & n738 ) | ( n648 & n1455 ) | ( n738 & n1455 ) ;
  assign n1458 = n703 | n748 ;
  buffer buf_n1459( .i (n726), .o (n1459) );
  assign n1460 = n1458 | n1459 ;
  assign n1461 = n684 & ~n1460 ;
  assign n1462 = ( n131 & n661 ) | ( n131 & n1461 ) | ( n661 & n1461 ) ;
  assign n1463 = ~n132 & n1462 ;
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n708), .o (n1467) );
  assign n1468 = ( ~n688 & n1464 ) | ( ~n688 & n1467 ) | ( n1464 & n1467 ) ;
  assign n1469 = n733 & ~n1468 ;
  assign n1470 = ( n734 & n1466 ) | ( n734 & ~n1469 ) | ( n1466 & ~n1469 ) ;
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n779( .i (n778), .o (n779) );
  assign n1473 = ~n779 & n1471 ;
  assign n1474 = ( ~n110 & n1472 ) | ( ~n110 & n1473 ) | ( n1472 & n1473 ) ;
  assign n1475 = ~n648 & n1474 ;
  assign n1476 = ( n1456 & ~n1457 ) | ( n1456 & n1475 ) | ( ~n1457 & n1475 ) ;
  assign n1477 = ~n600 & n1476 ;
  assign n1478 = ( n570 & ~n624 ) | ( n570 & n1477 ) | ( ~n624 & n1477 ) ;
  assign n1479 = ~n571 & n1478 ;
  assign n1480 = n407 & ~n1479 ;
  assign n1481 = n145 | n407 ;
  assign n1482 = ( ~n506 & n1480 ) | ( ~n506 & n1481 ) | ( n1480 & n1481 ) ;
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n375), .o (n1485) );
  assign n1486 = n540 & n1485 ;
  assign n1487 = ( n1354 & n1483 ) | ( n1354 & n1486 ) | ( n1483 & n1486 ) ;
  assign n1488 = ~n1484 & n1487 ;
  assign n1489 = n478 & n1488 ;
  assign n1490 = ( ~n1441 & n1442 ) | ( ~n1441 & n1489 ) | ( n1442 & n1489 ) ;
  buffer buf_n1491( .i (n1490), .o (n1491) );
  assign n1492 = ( ~n1429 & n1433 ) | ( ~n1429 & n1491 ) | ( n1433 & n1491 ) ;
  buffer buf_n382( .i (n381), .o (n382) );
  assign n1493 = n382 & ~n1491 ;
  assign n1494 = ( n1430 & n1492 ) | ( n1430 & ~n1493 ) | ( n1492 & ~n1493 ) ;
  assign n1495 = n92 & n1494 ;
  assign n1496 = ~n190 & n1495 ;
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  assign n1497 = ( n382 & ~n415 ) | ( n382 & n481 ) | ( ~n415 & n481 ) ;
  assign n1498 = ~n547 & n1497 ;
  assign n1499 = ( ~n417 & n548 ) | ( ~n417 & n1498 ) | ( n548 & n1498 ) ;
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  assign n1500 = n415 & ~n980 ;
  assign n1501 = ( n383 & ~n981 ) | ( n383 & n1500 ) | ( ~n981 & n1500 ) ;
  assign n1502 = ( ~n184 & n379 ) | ( ~n184 & n478 ) | ( n379 & n478 ) ;
  assign n1503 = n413 & n1502 ;
  assign n1504 = ( n186 & n414 ) | ( n186 & ~n1503 ) | ( n414 & ~n1503 ) ;
  assign n1505 = ( ~n449 & n513 ) | ( ~n449 & n1504 ) | ( n513 & n1504 ) ;
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n759( .i (n758), .o (n759) );
  assign n1506 = n779 | n843 ;
  assign n1507 = n759 | n1506 ;
  assign n1508 = ( ~n715 & n845 ) | ( ~n715 & n1507 ) | ( n845 & n1507 ) ;
  assign n1509 = ( n739 & n846 ) | ( n739 & n1508 ) | ( n846 & n1508 ) ;
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  assign n1512 = ~n114 & n1510 ;
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n1513( .i (n694), .o (n1513) );
  assign n1514 = ( n716 & n739 ) | ( n716 & n1513 ) | ( n739 & n1513 ) ;
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  assign n1515 = ~n1262 & n1513 ;
  assign n1516 = ( ~n717 & n1514 ) | ( ~n717 & n1515 ) | ( n1514 & n1515 ) ;
  assign n1517 = ~n107 & n711 ;
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  assign n1520 = n736 & ~n1518 ;
  assign n1521 = ( n693 & ~n1519 ) | ( n693 & n1520 ) | ( ~n1519 & n1520 ) ;
  buffer buf_n1522( .i (n1521), .o (n1522) );
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  assign n1524 = n761 & ~n1522 ;
  assign n1525 = ( ~n110 & n693 ) | ( ~n110 & n714 ) | ( n693 & n714 ) ;
  buffer buf_n1526( .i (n1076), .o (n1526) );
  assign n1527 = ~n737 & n1526 ;
  assign n1528 = ( ~n694 & n1525 ) | ( ~n694 & n1527 ) | ( n1525 & n1527 ) ;
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1529( .i (n736), .o (n1529) );
  assign n1530 = n1153 | n1529 ;
  assign n1531 = n110 | n693 ;
  assign n1532 = ( ~n1154 & n1530 ) | ( ~n1154 & n1531 ) | ( n1530 & n1531 ) ;
  assign n1533 = ~n1528 & n1532 ;
  assign n1534 = ( n1523 & n1524 ) | ( n1523 & n1533 ) | ( n1524 & n1533 ) ;
  assign n1535 = ~n1516 & n1534 ;
  assign n1536 = ( ~n1511 & n1512 ) | ( ~n1511 & n1535 ) | ( n1512 & n1535 ) ;
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  assign n1537 = ( n1120 & ~n1153 ) | ( n1120 & n1529 ) | ( ~n1153 & n1529 ) ;
  assign n1538 = n1120 | n1526 ;
  assign n1539 = ( n1154 & n1537 ) | ( n1154 & n1538 ) | ( n1537 & n1538 ) ;
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n696( .i (n695), .o (n696) );
  assign n1542 = ( n113 & n696 ) | ( n113 & n1540 ) | ( n696 & n1540 ) ;
  assign n1543 = n106 & n755 ;
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  assign n1546 = n778 & ~n1544 ;
  assign n1547 = ( n736 & ~n1545 ) | ( n736 & n1546 ) | ( ~n1545 & n1546 ) ;
  buffer buf_n1548( .i (n1547), .o (n1548) );
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1550( .i (n669), .o (n1550) );
  assign n1551 = ( ~n715 & n1548 ) | ( ~n715 & n1550 ) | ( n1548 & n1550 ) ;
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1552( .i (n109), .o (n1552) );
  assign n1553 = ( n1176 & ~n1529 ) | ( n1176 & n1552 ) | ( ~n1529 & n1552 ) ;
  assign n1554 = n1550 & n1553 ;
  assign n1555 = ( ~n1549 & n1551 ) | ( ~n1549 & n1554 ) | ( n1551 & n1554 ) ;
  assign n1556 = ~n696 & n1555 ;
  assign n1557 = ( n1541 & ~n1542 ) | ( n1541 & n1556 ) | ( ~n1542 & n1556 ) ;
  buffer buf_n1558( .i (n1557), .o (n1558) );
  assign n1559 = ( n675 & n1536 ) | ( n675 & ~n1558 ) | ( n1536 & ~n1558 ) ;
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n1560 = n1059 & ~n1513 ;
  assign n1561 = ( n762 & n1060 ) | ( n762 & n1560 ) | ( n1060 & n1560 ) ;
  assign n1562 = n741 | n1561 ;
  assign n1563 = n719 | n1562 ;
  assign n1564 = ( n675 & n1558 ) | ( n675 & ~n1563 ) | ( n1558 & ~n1563 ) ;
  assign n1565 = n1559 & ~n1564 ;
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  assign n1568 = ( n629 & n1287 ) | ( n629 & ~n1566 ) | ( n1287 & ~n1566 ) ;
  assign n1569 = n1567 | n1568 ;
  assign n1570 = n379 & ~n1569 ;
  assign n1571 = ( n479 & n578 ) | ( n479 & n1570 ) | ( n578 & n1570 ) ;
  assign n1572 = ~n579 & n1571 ;
  assign n1573 = ( n449 & ~n513 ) | ( n449 & n1572 ) | ( ~n513 & n1572 ) ;
  assign n1574 = n1505 | n1573 ;
  assign n1575 = n1501 | n1574 ;
  assign n1576 = n1499 | n1575 ;
  assign y0 = n869 ;
  assign y1 = n915 ;
  assign y2 = n971 ;
  assign y3 = n1367 ;
  assign y4 = n1425 ;
  assign y5 = n1496 ;
  assign y6 = n1576 ;
endmodule
