module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 ;
  wire n2 , n3 , n4 , n5 , n7 , n8 , n10 , n11 , n12 , n13 , n15 , n16 , n17 , n18 , n20 , n21 , n22 , n24 , n25 , n26 , n27 , n28 , n30 , n31 , n32 , n34 , n35 , n36 , n37 , n38 , n40 , n41 , n42 , n43 , n44 , n46 , n47 , n49 , n50 , n51 , n53 , n54 , n56 , n57 , n58 , n60 , n61 , n62 , n63 , n65 , n66 , n67 , n68 , n69 , n70 , n72 , n73 , n74 , n75 , n76 , n77 , n79 , n80 , n81 , n82 , n83 , n89 , n90 , n92 , n93 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n178 , n179 , n180 , n181 , n183 , n184 , n185 , n186 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n212 , n214 , n215 , n216 , n217 , n218 , n219 , n221 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n341 , n342 , n343 , n344 , n345 , n346 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n392 , n393 , n394 , n395 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n407 , n408 , n410 , n411 , n413 , n414 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n427 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 ;
  buffer buf_n72( .i (x15), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n24( .i (x5), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n34( .i (x7), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  assign n432 = n28 & n38 ;
  assign n433 = n77 & n432 ;
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n79( .i (x16), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n30( .i (x6), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  assign n446 = n26 & n32 ;
  buffer buf_n447( .i (n446), .o (n447) );
  assign n448 = n83 & n447 ;
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  assign n462 = n38 & n447 ;
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  assign n476 = x17 & x18 ;
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n7( .i (x1), .o (n7) );
  assign n495 = n2 & n7 ;
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n10( .i (x2), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n15( .i (x3), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  assign n500 = n13 & n18 ;
  buffer buf_n501( .i (n500), .o (n501) );
  assign n502 = n499 & n501 ;
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n20( .i (x4), .o (n20) );
  assign n515 = n2 & n20 ;
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  assign n520 = n501 & n519 ;
  buffer buf_n521( .i (n520), .o (n521) );
  assign n522 = ~n464 & n521 ;
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n49( .i (x10), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  assign n533 = n72 & n79 ;
  buffer buf_n534( .i (n533), .o (n534) );
  assign n535 = n51 & n534 ;
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  assign n551 = n32 & n51 ;
  assign n552 = n82 & n551 ;
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  assign n567 = n34 & n49 ;
  buffer buf_n568( .i (n567), .o (n568) );
  assign n569 = n32 & n568 ;
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n92( .i (x22), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  assign n585 = x19 | x20 ;
  buffer buf_n586( .i (n585), .o (n586) );
  assign n587 = n93 & n586 ;
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  assign n604 = n464 & n521 ;
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n40( .i (x8), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  assign n615 = n44 & n518 ;
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n53( .i (x11), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n46( .i (x9), .o (n46) );
  assign n629 = n10 & n46 ;
  assign n630 = n54 & n629 ;
  buffer buf_n631( .i (n630), .o (n631) );
  assign n632 = n497 & n631 ;
  assign n633 = n28 & n632 ;
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n65( .i (x14), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  assign n647 = n51 & n496 ;
  assign n648 = n631 & n647 ;
  buffer buf_n649( .i (n648), .o (n649) );
  assign n651 = n70 & n649 ;
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n89( .i (x21), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  assign n664 = n90 & n586 ;
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n123( .i (x26), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n95( .i (x23), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n115( .i (x25), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n135( .i (x27), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  assign n681 = ( ~n101 & n121 ) | ( ~n101 & n141 ) | ( n121 & n141 ) ;
  assign n682 = ( n101 & n121 ) | ( n101 & n141 ) | ( n121 & n141 ) ;
  assign n683 = ( n102 & n681 ) | ( n102 & ~n682 ) | ( n681 & ~n682 ) ;
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n153( .i (x29), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n170( .i (x31), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n162( .i (x30), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n178( .i (x32), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n105( .i (x24), .o (n105) );
  buffer buf_n144( .i (x28), .o (n144) );
  assign n685 = n105 | n144 ;
  assign n686 = n105 & n144 ;
  assign n687 = n685 & ~n686 ;
  buffer buf_n688( .i (n687), .o (n688) );
  assign n689 = ( ~n165 & n181 ) | ( ~n165 & n688 ) | ( n181 & n688 ) ;
  assign n690 = ( n165 & n181 ) | ( n165 & n688 ) | ( n181 & n688 ) ;
  assign n691 = ( n166 & n689 ) | ( n166 & ~n690 ) | ( n689 & ~n690 ) ;
  buffer buf_n692( .i (n691), .o (n692) );
  assign n693 = ( n159 & ~n176 ) | ( n159 & n692 ) | ( ~n176 & n692 ) ;
  assign n694 = ( n159 & n176 ) | ( n159 & ~n692 ) | ( n176 & ~n692 ) ;
  assign n695 = ( ~n160 & n693 ) | ( ~n160 & n694 ) | ( n693 & n694 ) ;
  buffer buf_n696( .i (n695), .o (n696) );
  assign n697 = ( n132 & ~n684 ) | ( n132 & n696 ) | ( ~n684 & n696 ) ;
  assign n698 = ( n132 & n684 ) | ( n132 & ~n696 ) | ( n684 & ~n696 ) ;
  assign n699 = ( ~n133 & n697 ) | ( ~n133 & n698 ) | ( n697 & n698 ) ;
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n223( .i (x40), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n258( .i (x42), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n241( .i (x41), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n316( .i (x46), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  assign n707 = ( ~n172 & n243 ) | ( ~n172 & n318 ) | ( n243 & n318 ) ;
  assign n708 = ( n172 & n243 ) | ( n172 & n318 ) | ( n243 & n318 ) ;
  assign n709 = ( n173 & n707 ) | ( n173 & ~n708 ) | ( n707 & ~n708 ) ;
  buffer buf_n710( .i (n709), .o (n710) );
  assign n711 = ( n228 & ~n263 ) | ( n228 & n710 ) | ( ~n263 & n710 ) ;
  assign n712 = ( n228 & n263 ) | ( n228 & ~n710 ) | ( n263 & ~n710 ) ;
  assign n713 = ( ~n229 & n711 ) | ( ~n229 & n712 ) | ( n711 & n712 ) ;
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n287( .i (x44), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n341( .i (x48), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n272( .i (x43), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n302( .i (x45), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n330( .i (x47), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  assign n715 = ( ~n274 & n304 ) | ( ~n274 & n332 ) | ( n304 & n332 ) ;
  assign n716 = ( n274 & n304 ) | ( n274 & n332 ) | ( n304 & n332 ) ;
  assign n717 = ( n275 & n715 ) | ( n275 & ~n716 ) | ( n715 & ~n716 ) ;
  buffer buf_n718( .i (n717), .o (n718) );
  assign n719 = ( n292 & ~n346 ) | ( n292 & n718 ) | ( ~n346 & n718 ) ;
  assign n720 = ( n292 & n346 ) | ( n292 & ~n718 ) | ( n346 & ~n718 ) ;
  assign n721 = ( ~n293 & n719 ) | ( ~n293 & n720 ) | ( n719 & n720 ) ;
  buffer buf_n722( .i (n721), .o (n722) );
  assign n723 = n714 | n722 ;
  assign n724 = n714 & n722 ;
  assign n725 = n723 & ~n724 ;
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n60( .i (x13), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n56( .i (x12), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  assign n734 = n36 & n58 ;
  assign n735 = n63 & n734 ;
  buffer buf_n736( .i (n735), .o (n736) );
  assign n737 = n649 & n736 ;
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n348( .i (x49), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  assign n745 = n158 & n353 ;
  buffer buf_n407( .i (x54), .o (n407) );
  buffer buf_n427( .i (x58), .o (n427) );
  assign n746 = n407 & n427 ;
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  assign n752 = n745 | n751 ;
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  assign n755 = n338 | n753 ;
  assign n756 = ( n740 & n754 ) | ( n740 & n755 ) | ( n754 & n755 ) ;
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  assign n757 = n74 & n568 ;
  assign n758 = n15 & n40 ;
  buffer buf_n759( .i (n758), .o (n759) );
  assign n761 = n496 & n759 ;
  assign n762 = ~n757 & n761 ;
  buffer buf_n221( .i (x39), .o (n221) );
  assign n763 = n49 & n221 ;
  buffer buf_n764( .i (n763), .o (n764) );
  assign n767 = ( n17 & n36 ) | ( n17 & ~n764 ) | ( n36 & ~n764 ) ;
  assign n768 = n16 & n35 ;
  assign n769 = ( n16 & n35 ) | ( n16 & n41 ) | ( n35 & n41 ) ;
  assign n770 = ( n516 & n768 ) | ( n516 & n769 ) | ( n768 & n769 ) ;
  assign n771 = ~n767 & n770 ;
  assign n772 = n762 | n771 ;
  buffer buf_n773( .i (n772), .o (n773) );
  assign n775 = n168 & n773 ;
  buffer buf_n429( .i (x59), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  assign n776 = n25 & ~n430 ;
  assign n777 = n534 & n776 ;
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n47( .i (n46), .o (n47) );
  assign n779 = n41 & n47 ;
  assign n780 = n516 & n779 ;
  buffer buf_n781( .i (n780), .o (n781) );
  assign n784 = n778 & n781 ;
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n214( .i (x38), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n5( .i (n4), .o (n5) );
  assign n787 = n4 & n764 ;
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  assign n788 = n22 & n759 ;
  assign n789 = ( n5 & n787 ) | ( n5 & ~n788 ) | ( n787 & ~n788 ) ;
  buffer buf_n790( .i (n789), .o (n790) );
  assign n792 = n219 & ~n790 ;
  assign n793 = n785 | n792 ;
  assign n794 = n775 | n793 ;
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n376( .i (x51), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  assign n796 = n337 & ~n383 ;
  buffer buf_n416( .i (x57), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  assign n797 = n337 & ~n423 ;
  buffer buf_n358( .i (x50), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  assign n798 = ( n337 & n365 ) | ( n337 & n423 ) | ( n365 & n423 ) ;
  assign n799 = ( ~n796 & n797 ) | ( ~n796 & n798 ) | ( n797 & n798 ) ;
  assign n800 = n795 | n799 ;
  buffer buf_n397( .i (x53), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  assign n801 = n381 | n402 ;
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n336), .o (n803) );
  assign n804 = n802 | n803 ;
  buffer buf_n392( .i (x52), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  assign n805 = n395 | n400 ;
  buffer buf_n806( .i (n805), .o (n806) );
  assign n814 = n335 & ~n806 ;
  buffer buf_n815( .i (n814), .o (n815) );
  assign n816 = ( n365 & n423 ) | ( n365 & ~n815 ) | ( n423 & ~n815 ) ;
  buffer buf_n817( .i (n422), .o (n817) );
  assign n818 = n815 | n817 ;
  assign n819 = ( n804 & n816 ) | ( n804 & ~n818 ) | ( n816 & ~n818 ) ;
  assign n820 = n795 & ~n819 ;
  assign n821 = ( n756 & n800 ) | ( n756 & ~n820 ) | ( n800 & ~n820 ) ;
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n774( .i (n773), .o (n774) );
  assign n829 = n142 & n774 ;
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n188( .i (x34), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n791( .i (n790), .o (n791) );
  assign n830 = n194 & ~n791 ;
  assign n831 = n786 | n830 ;
  assign n832 = n829 | n831 ;
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  assign n837 = ~n298 & n834 ;
  assign n838 = n298 & ~n834 ;
  assign n839 = n837 | n838 ;
  buffer buf_n840( .i (n839), .o (n840) );
  assign n842 = n390 & n840 ;
  assign n843 = n290 & n395 ;
  assign n844 = n401 | n843 ;
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  assign n850 = n833 & n849 ;
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  assign n851 = n130 & n355 ;
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  assign n854 = n296 | n852 ;
  assign n855 = ( n741 & n853 ) | ( n741 & n854 ) | ( n853 & n854 ) ;
  assign n856 = n850 | n855 ;
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  assign n860 = n842 | n859 ;
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  assign n861 = ( n339 & n425 ) | ( n339 & n795 ) | ( n425 & n795 ) ;
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  assign n865 = n151 & n774 ;
  buffer buf_n196( .i (x35), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  assign n866 = n202 & ~n791 ;
  assign n867 = n786 | n866 ;
  assign n868 = n865 | n867 ;
  buffer buf_n869( .i (n868), .o (n869) );
  assign n872 = ( n312 & n326 ) | ( n312 & n869 ) | ( n326 & n869 ) ;
  assign n873 = n160 & n774 ;
  buffer buf_n204( .i (x36), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  assign n874 = n210 & ~n791 ;
  assign n875 = n786 | n874 ;
  assign n876 = n873 | n875 ;
  buffer buf_n877( .i (n876), .o (n877) );
  assign n880 = ( n312 & n869 ) | ( n312 & n877 ) | ( n869 & n877 ) ;
  assign n881 = ( n862 & n872 ) | ( n862 & n880 ) | ( n872 & n880 ) ;
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  assign n885 = n841 | n884 ;
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  assign n886 = ( ~n373 & n841 ) | ( ~n373 & n884 ) | ( n841 & n884 ) ;
  assign n887 = ( n860 & n885 ) | ( n860 & ~n886 ) | ( n885 & ~n886 ) ;
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  assign n889 = ( n328 & n863 ) | ( n328 & n879 ) | ( n863 & n879 ) ;
  buffer buf_n890( .i (n889), .o (n890) );
  assign n891 = n372 & n890 ;
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  assign n892 = n314 | n871 ;
  buffer buf_n893( .i (n892), .o (n893) );
  assign n894 = n314 & n871 ;
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  assign n895 = n742 | n812 ;
  buffer buf_n896( .i (n895), .o (n896) );
  assign n897 = n894 & ~n896 ;
  assign n898 = n893 & ~n897 ;
  assign n899 = n891 | n898 ;
  assign n900 = n890 & n893 ;
  assign n901 = n307 | n402 ;
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  assign n907 = n741 & n905 ;
  assign n908 = ( n870 & n906 ) | ( n870 & n907 ) | ( n906 & n907 ) ;
  assign n909 = n388 | n908 ;
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  assign n912 = n372 | n910 ;
  assign n913 = ( ~n900 & n911 ) | ( ~n900 & n912 ) | ( n911 & n912 ) ;
  assign n914 = n899 & n913 ;
  assign n915 = n139 & n352 ;
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n410( .i (x55), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  assign n916 = n408 & n411 ;
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  assign n920 = n915 | n919 ;
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  assign n932 = n914 | n931 ;
  buffer buf_n864( .i (n863), .o (n864) );
  assign n933 = n371 & n864 ;
  buffer buf_n934( .i (n933), .o (n934) );
  assign n935 = n327 | n878 ;
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  assign n938 = n328 & n879 ;
  assign n939 = ~n896 & n938 ;
  assign n940 = n937 & ~n939 ;
  assign n941 = n934 | n940 ;
  assign n942 = n864 & n936 ;
  assign n943 = n372 & ~n942 ;
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  assign n944 = n324 | n405 ;
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  assign n947 = n741 & n945 ;
  assign n948 = ( n878 & n946 ) | ( n878 & n947 ) | ( n946 & n947 ) ;
  assign n949 = n388 | n948 ;
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  assign n952 = n943 | n951 ;
  assign n953 = n941 & n952 ;
  assign n954 = n148 & n352 ;
  buffer buf_n413( .i (x56), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  assign n955 = n408 & n414 ;
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  assign n959 = n954 | n958 ;
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  assign n971 = n953 | n970 ;
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  assign n972 = n102 & n774 ;
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n183( .i (x33), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  assign n973 = n8 & n184 ;
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n760( .i (n759), .o (n760) );
  assign n978 = n517 & n760 ;
  assign n979 = n778 & n978 ;
  buffer buf_n980( .i (n979), .o (n980) );
  assign n982 = n977 | n980 ;
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  assign n983 = n192 & ~n766 ;
  buffer buf_n984( .i (n983), .o (n984) );
  assign n985 = n783 & n984 ;
  assign n986 = n982 | n985 ;
  assign n987 = n972 | n986 ;
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n995( .i (n773), .o (n995) );
  assign n996 = n112 & n995 ;
  buffer buf_n185( .i (n184), .o (n185) );
  assign n997 = n42 & n185 ;
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  assign n1001 = n980 | n1000 ;
  assign n1002 = n200 & ~n766 ;
  buffer buf_n1003( .i (n1002), .o (n1003) );
  assign n1004 = n783 & n1003 ;
  assign n1005 = n1001 | n1004 ;
  assign n1006 = n996 | n1005 ;
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  assign n1013 = n121 & n773 ;
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n186( .i (n185), .o (n186) );
  assign n1016 = n18 & n186 ;
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  assign n1020 = n981 | n1019 ;
  assign n1021 = n208 & ~n766 ;
  buffer buf_n1022( .i (n1021), .o (n1022) );
  assign n1023 = n783 & n1022 ;
  buffer buf_n1024( .i (n1023), .o (n1024) );
  assign n1025 = n1020 | n1024 ;
  assign n1026 = n1015 | n1025 ;
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1028( .i (n1027), .o (n1028) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  assign n1029 = n130 & n995 ;
  buffer buf_n212( .i (x37), .o (n212) );
  assign n1030 = n183 & n212 ;
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  assign n1036 = n980 | n1035 ;
  assign n1037 = n218 & ~n766 ;
  assign n1038 = n782 & n1037 ;
  buffer buf_n1039( .i (n1038), .o (n1039) );
  assign n1040 = n1036 | n1039 ;
  assign n1041 = n1029 | n1040 ;
  buffer buf_n1042( .i (n1041), .o (n1042) );
  assign n1045 = ( n282 & n297 ) | ( n282 & n1042 ) | ( n297 & n1042 ) ;
  buffer buf_n1046( .i (n1045), .o (n1046) );
  assign n1048 = ( n270 & n1028 ) | ( n270 & n1046 ) | ( n1028 & n1046 ) ;
  assign n1049 = ( n282 & n833 ) | ( n282 & n1042 ) | ( n833 & n1042 ) ;
  buffer buf_n1050( .i (n1049), .o (n1050) );
  assign n1052 = ( n270 & n1028 ) | ( n270 & n1050 ) | ( n1028 & n1050 ) ;
  assign n1053 = ( n882 & n1048 ) | ( n882 & n1052 ) | ( n1048 & n1052 ) ;
  buffer buf_n1054( .i (n1053), .o (n1054) );
  assign n1056 = ( n256 & n1012 ) | ( n256 & n1054 ) | ( n1012 & n1054 ) ;
  assign n1057 = ( n239 & n994 ) | ( n239 & n1056 ) | ( n994 & n1056 ) ;
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  assign n1059 = ~n813 & n1044 ;
  assign n1060 = n388 | n1044 ;
  assign n1061 = ( n744 & ~n1059 ) | ( n744 & n1060 ) | ( ~n1059 & n1060 ) ;
  assign n1062 = n121 & n354 ;
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  assign n1066 = ~n279 & n802 ;
  assign n1067 = n1063 | n1066 ;
  buffer buf_n1068( .i (n1067), .o (n1068) );
  assign n1069 = ( n1042 & n1065 ) | ( n1042 & n1068 ) | ( n1065 & n1068 ) ;
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  assign n1073 = n285 | n1071 ;
  assign n1074 = ( n1061 & n1072 ) | ( n1061 & n1073 ) | ( n1072 & n1073 ) ;
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  assign n1076 = ( n300 & n836 ) | ( n300 & n882 ) | ( n836 & n882 ) ;
  buffer buf_n1077( .i (n1076), .o (n1077) );
  assign n1078 = ~n284 & n1044 ;
  assign n1079 = n284 & ~n1044 ;
  assign n1080 = n1078 | n1079 ;
  buffer buf_n1081( .i (n1080), .o (n1081) );
  assign n1082 = n1077 & n1081 ;
  assign n1083 = ( n373 & n1077 ) | ( n373 & n1081 ) | ( n1077 & n1081 ) ;
  assign n1084 = ( n1075 & ~n1082 ) | ( n1075 & n1083 ) | ( ~n1082 & n1083 ) ;
  buffer buf_n1085( .i (n1084), .o (n1085) );
  assign n1086 = ~n233 & n988 ;
  assign n1087 = n233 & ~n988 ;
  assign n1088 = n1086 | n1087 ;
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n431( .i (n430), .o (n431) );
  assign n1091 = n350 & n431 ;
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  assign n1095 = n227 | n1092 ;
  assign n1096 = ( n736 & n1093 ) | ( n736 & n1095 ) | ( n1093 & n1095 ) ;
  assign n1097 = ( n650 & n1094 ) | ( n650 & n1096 ) | ( n1094 & n1096 ) ;
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  assign n1101 = n225 & n394 ;
  assign n1102 = n400 | n1101 ;
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  assign n1107 = n1098 | n1106 ;
  buffer buf_n1108( .i (n1107), .o (n1108) );
  assign n1109 = ( n988 & n1100 ) | ( n988 & n1108 ) | ( n1100 & n1108 ) ;
  buffer buf_n1110( .i (n1109), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n387), .o (n1112) );
  assign n1113 = n1110 | n1112 ;
  assign n1114 = ( n1089 & n1111 ) | ( n1089 & n1113 ) | ( n1111 & n1113 ) ;
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  assign n1117 = n255 & n1090 ;
  assign n1118 = n1011 & n1090 ;
  assign n1119 = ( n1054 & n1117 ) | ( n1054 & n1118 ) | ( n1117 & n1118 ) ;
  buffer buf_n1120( .i (n371), .o (n1120) );
  assign n1121 = ( n255 & n1090 ) | ( n255 & n1120 ) | ( n1090 & n1120 ) ;
  assign n1122 = ( n1011 & n1090 ) | ( n1011 & n1120 ) | ( n1090 & n1120 ) ;
  assign n1123 = ( n1054 & n1121 ) | ( n1054 & n1122 ) | ( n1121 & n1122 ) ;
  assign n1124 = ( n1116 & ~n1119 ) | ( n1116 & n1123 ) | ( ~n1119 & n1123 ) ;
  buffer buf_n1125( .i (n1124), .o (n1125) );
  assign n1126 = ~n251 & n1007 ;
  assign n1127 = n251 & ~n1007 ;
  assign n1128 = n1126 | n1127 ;
  buffer buf_n1129( .i (n1128), .o (n1129) );
  assign n1133 = n389 & n1129 ;
  assign n1134 = n244 & n395 ;
  assign n1135 = n401 | n1134 ;
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  assign n1143 = n1009 & n1142 ;
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n356( .i (n355), .o (n356) );
  assign n1144 = n103 & n356 ;
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  assign n1147 = n251 | n1145 ;
  assign n1148 = ( n742 & n1146 ) | ( n742 & n1147 ) | ( n1146 & n1147 ) ;
  buffer buf_n1149( .i (n1148), .o (n1149) );
  assign n1150 = n1143 | n1149 ;
  assign n1151 = n1133 | n1150 ;
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  assign n1154 = n1055 & n1132 ;
  buffer buf_n374( .i (n373), .o (n374) );
  assign n1155 = ( n374 & n1055 ) | ( n374 & n1132 ) | ( n1055 & n1132 ) ;
  assign n1156 = ( n1153 & ~n1154 ) | ( n1153 & n1155 ) | ( ~n1154 & n1155 ) ;
  assign n1157 = ~n269 & n1027 ;
  assign n1158 = n269 & ~n1027 ;
  assign n1159 = n1157 | n1158 ;
  buffer buf_n1160( .i (n1159), .o (n1160) );
  assign n1162 = n390 & n1160 ;
  assign n1163 = n261 & n395 ;
  assign n1164 = n401 | n1163 ;
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  assign n1171 = n1027 & n1170 ;
  buffer buf_n113( .i (n112), .o (n113) );
  assign n1172 = n113 & n356 ;
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  assign n1175 = n268 | n1173 ;
  assign n1176 = ( n742 & n1174 ) | ( n742 & n1175 ) | ( n1174 & n1175 ) ;
  assign n1177 = n1171 | n1176 ;
  buffer buf_n1178( .i (n1177), .o (n1178) );
  buffer buf_n1179( .i (n1178), .o (n1179) );
  assign n1180 = n1162 | n1179 ;
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  assign n1181 = ( n882 & n1047 ) | ( n882 & n1051 ) | ( n1047 & n1051 ) ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  assign n1183 = n1161 & n1182 ;
  assign n1184 = ( n373 & n1161 ) | ( n373 & n1182 ) | ( n1161 & n1182 ) ;
  assign n1185 = ( n1180 & ~n1183 ) | ( n1180 & n1184 ) | ( ~n1183 & n1184 ) ;
  buffer buf_n1186( .i (n1185), .o (n1186) );
  assign y0 = n445 ;
  assign y1 = n461 ;
  assign y2 = n475 ;
  assign y3 = n494 ;
  assign y4 = n514 ;
  assign y5 = ~n532 ;
  assign y6 = ~n550 ;
  assign y7 = ~n566 ;
  assign y8 = ~n584 ;
  assign y9 = n603 ;
  assign y10 = ~n614 ;
  assign y11 = n628 ;
  assign y12 = n646 ;
  assign y13 = n663 ;
  assign y14 = n680 ;
  assign y15 = n706 ;
  assign y16 = n733 ;
  assign y17 = n828 ;
  assign y18 = n888 ;
  assign y19 = n932 ;
  assign y20 = n971 ;
  assign y21 = n1058 ;
  assign y22 = n1085 ;
  assign y23 = n1125 ;
  assign y24 = n1156 ;
  assign y25 = n1186 ;
endmodule
