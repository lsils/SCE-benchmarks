module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n13 , n14 , n15 , n16 , n17 , n19 , n20 , n22 , n23 , n24 , n25 , n27 , n28 , n29 , n30 , n31 , n32 , n34 , n35 , n36 , n37 , n38 , n40 , n41 , n42 , n43 , n45 , n46 , n47 , n48 , n50 , n51 , n52 , n54 , n55 , n56 , n57 , n58 , n60 , n61 , n62 , n63 , n64 , n66 , n67 , n69 , n70 , n72 , n74 , n75 , n76 , n78 , n79 , n80 , n82 , n83 , n84 , n86 , n87 , n88 , n89 , n90 , n91 , n93 , n94 , n95 , n96 , n97 , n98 , n100 , n101 , n103 , n105 , n106 , n107 , n109 , n110 , n111 , n113 , n115 , n116 , n117 , n118 , n119 , n120 , n122 , n124 , n125 , n126 , n127 , n128 , n130 , n131 , n132 , n133 , n135 , n136 , n137 , n138 , n139 , n141 , n142 , n143 , n144 , n145 , n147 , n148 , n149 , n150 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 ;
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n152( .i (x31), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n109( .i (x22), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n147( .i (x30), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  assign n168 = n111 & n149 ;
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n13( .i (x1), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n135( .i (x28), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  assign n170 = n15 & n137 ;
  buffer buf_n171( .i (n170), .o (n171) );
  assign n172 = n169 & n171 ;
  buffer buf_n173( .i (n172), .o (n173) );
  assign n174 = ~n158 & n173 ;
  buffer buf_n78( .i (x15), .o (n78) );
  buffer buf_n82( .i (x16), .o (n82) );
  assign n175 = n78 | n82 ;
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  assign n179 = n156 & ~n178 ;
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  assign n182 = ( ~n9 & n174 ) | ( ~n9 & n181 ) | ( n174 & n181 ) ;
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n160( .i (x32), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n27( .i (x4), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  assign n186 = n7 | n32 ;
  buffer buf_n187( .i (n186), .o (n187) );
  assign n188 = n167 & ~n187 ;
  buffer buf_n141( .i (x29), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  assign n189 = n145 & n171 ;
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n115( .i (x24), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  assign n191 = ~n7 & n120 ;
  assign n192 = n190 & n191 ;
  buffer buf_n193( .i (n192), .o (n193) );
  assign n197 = n167 & n187 ;
  assign n198 = ( n188 & n193 ) | ( n188 & ~n197 ) | ( n193 & ~n197 ) ;
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  assign n201 = n2 | n135 ;
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n22( .i (x3), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n150( .i (n149), .o (n150) );
  assign n206 = n25 & ~n150 ;
  buffer buf_n207( .i (n206), .o (n207) );
  assign n208 = ~n205 & n207 ;
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n138( .i (n137), .o (n138) );
  assign n214 = n138 | n150 ;
  buffer buf_n215( .i (n214), .o (n215) );
  assign n216 = n25 & n144 ;
  buffer buf_n217( .i (n216), .o (n217) );
  assign n218 = ~n215 & n217 ;
  buffer buf_n219( .i (n218), .o (n219) );
  assign n220 = n9 | n219 ;
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n66( .i (x11), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n69( .i (x12), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  assign n224 = ~n67 & n70 ;
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n54( .i (x9), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n100( .i (x19), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  assign n227 = ~n70 & n101 ;
  assign n228 = n56 & ~n227 ;
  buffer buf_n105( .i (x21), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  assign n229 = n67 & n106 ;
  assign n230 = n143 & n229 ;
  assign n231 = ~n228 & n230 ;
  assign n232 = n226 | n231 ;
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  assign n234 = n66 & n69 ;
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  assign n238 = n58 | n237 ;
  buffer buf_n60( .i (x10), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  assign n239 = n62 & n149 ;
  assign n240 = ~n203 & n239 ;
  buffer buf_n241( .i (n240), .o (n241) );
  assign n242 = n238 & n241 ;
  assign n243 = n233 & n242 ;
  buffer buf_n244( .i (n243), .o (n244) );
  assign n246 = n149 & ~n202 ;
  buffer buf_n247( .i (n246), .o (n247) );
  assign n248 = n55 & n101 ;
  buffer buf_n103( .i (x20), .o (n103) );
  assign n249 = n103 & n141 ;
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = n248 & n250 ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n253 = n247 & n252 ;
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n107( .i (n106), .o (n107) );
  assign n261 = ~n62 & n107 ;
  assign n262 = ~n225 & n261 ;
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  assign n265 = n254 & n264 ;
  buffer buf_n266( .i (n265), .o (n266) );
  assign n267 = n244 | n266 ;
  buffer buf_n268( .i (n267), .o (n268) );
  assign n255 = n60 & n69 ;
  buffer buf_n256( .i (n255), .o (n256) );
  assign n269 = n66 & ~n69 ;
  buffer buf_n270( .i (n269), .o (n270) );
  assign n271 = n256 | n270 ;
  buffer buf_n272( .i (n271), .o (n272) );
  assign n273 = n58 | n272 ;
  assign n274 = n241 & ~n273 ;
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  assign n257 = n107 | n256 ;
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  assign n278 = n254 & n260 ;
  assign n279 = n54 | n60 ;
  buffer buf_n280( .i (n279), .o (n280) );
  assign n281 = n270 & ~n280 ;
  buffer buf_n282( .i (n281), .o (n282) );
  assign n283 = n247 & n282 ;
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  assign n286 = ~n237 & n272 ;
  buffer buf_n287( .i (n286), .o (n287) );
  assign n288 = ~n284 & n287 ;
  assign n289 = ( n278 & n285 ) | ( n278 & ~n288 ) | ( n285 & ~n288 ) ;
  buffer buf_n290( .i (n289), .o (n290) );
  assign n292 = n277 | n290 ;
  assign n293 = n268 | n292 ;
  buffer buf_n86( .i (x17), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n93( .i (x18), .o (n93) );
  assign n294 = n82 | n93 ;
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = n88 & ~n295 ;
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n74( .i (x14), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  assign n299 = ~n76 & n80 ;
  buffer buf_n300( .i (n299), .o (n300) );
  assign n301 = n297 & n300 ;
  buffer buf_n302( .i (n301), .o (n302) );
  assign n303 = n80 & ~n295 ;
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n40( .i (x6), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n45( .i (x7), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  assign n307 = ~n42 & n47 ;
  assign n308 = ~n89 & n307 ;
  assign n309 = n304 & n308 ;
  buffer buf_n310( .i (n309), .o (n310) );
  assign n312 = n302 | n310 ;
  buffer buf_n313( .i (n312), .o (n313) );
  assign n315 = n88 & ~n176 ;
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  assign n319 = n42 | n95 ;
  buffer buf_n320( .i (n319), .o (n320) );
  assign n321 = n316 & ~n320 ;
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  assign n325 = n313 | n324 ;
  buffer buf_n139( .i (n138), .o (n139) );
  assign n326 = ~n3 & n14 ;
  buffer buf_n113( .i (x23), .o (n113) );
  assign n327 = n113 & n147 ;
  buffer buf_n328( .i (n327), .o (n328) );
  assign n329 = n326 & n328 ;
  buffer buf_n330( .i (n329), .o (n330) );
  assign n332 = n139 & n330 ;
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  assign n335 = n302 | n333 ;
  assign n336 = ( n275 & n334 ) | ( n275 & n335 ) | ( n334 & n335 ) ;
  buffer buf_n337( .i (n336), .o (n337) );
  assign n338 = n325 & n337 ;
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n96( .i (n95), .o (n96) );
  assign n340 = n89 | n96 ;
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n50( .i (x8), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  assign n343 = ~n42 & n52 ;
  buffer buf_n344( .i (n343), .o (n344) );
  assign n346 = n320 & ~n344 ;
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  assign n348 = ~n91 & n341 ;
  assign n349 = ( n342 & ~n347 ) | ( n342 & n348 ) | ( ~n347 & n348 ) ;
  assign n350 = n235 & ~n280 ;
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n331( .i (n330), .o (n331) );
  assign n354 = n139 | n178 ;
  assign n355 = n331 & ~n354 ;
  assign n356 = n353 & n355 ;
  assign n357 = ~n349 & n356 ;
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  assign n359 = ~n80 & n84 ;
  buffer buf_n360( .i (n359), .o (n360) );
  assign n361 = ~n89 & n96 ;
  assign n362 = n360 & n361 ;
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  assign n367 = n333 & n363 ;
  assign n368 = ( n275 & n364 ) | ( n275 & n367 ) | ( n364 & n367 ) ;
  buffer buf_n369( .i (n368), .o (n369) );
  assign n370 = n358 | n369 ;
  assign n371 = n322 & n333 ;
  assign n372 = ( n275 & n323 ) | ( n275 & n371 ) | ( n323 & n371 ) ;
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  assign n375 = n370 | n374 ;
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  assign n376 = n139 | n351 ;
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  assign n378 = n17 & n169 ;
  assign n379 = ~n341 & n378 ;
  assign n380 = n377 & n379 ;
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  assign n383 = n80 & n84 ;
  assign n384 = n5 | n383 ;
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  assign n390 = ( n11 & n382 ) | ( n11 & n389 ) | ( n382 & n389 ) ;
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  assign n391 = ~n8 & n173 ;
  buffer buf_n392( .i (n391), .o (n392) );
  assign n394 = n365 & n392 ;
  assign n395 = ( n277 & n366 ) | ( n277 & n394 ) | ( n366 & n394 ) ;
  assign n396 = n390 | n395 ;
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  assign n397 = n173 & n306 ;
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  assign n400 = n276 & n313 ;
  assign n401 = n399 | n400 ;
  buffer buf_n345( .i (n344), .o (n345) );
  assign n402 = n205 | n345 ;
  assign n403 = n386 & n402 ;
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  assign n406 = ( n11 & n382 ) | ( n11 & n405 ) | ( n382 & n405 ) ;
  assign n407 = n401 | n406 ;
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n393( .i (n392), .o (n393) );
  assign n408 = n324 & n392 ;
  assign n409 = ( n314 & n393 ) | ( n314 & n408 ) | ( n393 & n408 ) ;
  buffer buf_n48( .i (n47), .o (n48) );
  assign n410 = n5 & n48 ;
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  assign n416 = n302 | n412 ;
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  assign n419 = ( n277 & n415 ) | ( n277 & n418 ) | ( n415 & n418 ) ;
  assign n420 = n409 | n419 ;
  buffer buf_n43( .i (n42), .o (n43) );
  assign n421 = n52 & n84 ;
  assign n422 = n43 | n421 ;
  buffer buf_n423( .i (n422), .o (n423) );
  assign n424 = n204 | n360 ;
  assign n425 = n423 & ~n424 ;
  assign n426 = n48 & ~n138 ;
  assign n427 = ~n178 & n426 ;
  buffer buf_n428( .i (n427), .o (n428) );
  assign n429 = n425 | n428 ;
  buffer buf_n430( .i (n429), .o (n430) );
  assign n431 = n381 & n430 ;
  assign n432 = n415 | n431 ;
  assign n433 = n276 | n392 ;
  buffer buf_n311( .i (n310), .o (n311) );
  assign n434 = n311 | n364 ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n436 = n433 & n435 ;
  assign n437 = n432 | n436 ;
  assign n438 = n4 & ~n47 ;
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  assign n444 = n98 & n331 ;
  assign n445 = n318 & n444 ;
  buffer buf_n446( .i (n445), .o (n446) );
  assign n447 = n377 | n441 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = ( n443 & n446 ) | ( n443 & n448 ) | ( n446 & n448 ) ;
  assign n450 = n369 | n449 ;
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n298( .i (n297), .o (n298) );
  assign n452 = n298 | n317 ;
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  assign n456 = n337 & n455 ;
  buffer buf_n457( .i (n41), .o (n457) );
  assign n458 = n52 | n457 ;
  buffer buf_n459( .i (n458), .o (n459) );
  assign n460 = ~n439 & n459 ;
  assign n461 = ( n352 & n440 ) | ( n352 & ~n460 ) | ( n440 & ~n460 ) ;
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  assign n464 = ( n443 & n446 ) | ( n443 & n463 ) | ( n446 & n463 ) ;
  assign n465 = n373 | n464 ;
  assign n466 = n456 | n465 ;
  buffer buf_n122( .i (x25), .o (n122) );
  assign n467 = n115 | n122 ;
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  assign n472 = n7 | n471 ;
  assign n473 = ( n8 & n190 ) | ( n8 & n472 ) | ( n190 & n472 ) ;
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n72( .i (x13), .o (n72) );
  assign n478 = n72 & ~n109 ;
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  assign n486 = n193 & n485 ;
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  assign n489 = n139 & n169 ;
  buffer buf_n34( .i (x5), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  assign n490 = ~n6 & n38 ;
  buffer buf_n491( .i (n6), .o (n491) );
  assign n492 = ( n489 & n490 ) | ( n489 & ~n491 ) | ( n490 & ~n491 ) ;
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  assign n498 = n10 | n276 ;
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n124( .i (x26), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n130( .i (x27), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  assign n500 = n24 & ~n132 ;
  buffer buf_n501( .i (n500), .o (n501) );
  assign n502 = n128 & ~n501 ;
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  assign n508 = n499 | n507 ;
  buffer buf_n133( .i (n132), .o (n133) );
  assign n509 = ~n25 & n133 ;
  buffer buf_n510( .i (n509), .o (n510) );
  assign n511 = n128 & n501 ;
  assign n512 = n510 | n511 ;
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  assign n517 = n499 | n516 ;
  buffer buf_n291( .i (n290), .o (n291) );
  assign n518 = n268 | n291 ;
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n19( .i (x2), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  assign n519 = n20 | n23 ;
  buffer buf_n520( .i (n519), .o (n520) );
  assign n521 = n144 | n520 ;
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  assign n524 = n215 | n217 ;
  assign n525 = n523 & ~n524 ;
  assign n526 = n9 | n525 ;
  assign n527 = n266 | n526 ;
  assign n528 = n245 | n527 ;
  buffer buf_n529( .i (n528), .o (n529) );
  assign n530 = n212 | n291 ;
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  assign n531 = n64 & n237 ;
  buffer buf_n532( .i (n531), .o (n532) );
  assign n533 = n254 & n532 ;
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  assign y0 = n185 ;
  assign y1 = n200 ;
  assign y2 = n213 ;
  assign y3 = n223 ;
  assign y4 = n293 ;
  assign y5 = n339 ;
  assign y6 = n375 ;
  assign y7 = n396 ;
  assign y8 = n407 ;
  assign y9 = n420 ;
  assign y10 = n437 ;
  assign y11 = n451 ;
  assign y12 = n466 ;
  assign y13 = n477 ;
  assign y14 = n488 ;
  assign y15 = n196 ;
  assign y16 = n497 ;
  assign y17 = n508 ;
  assign y18 = n517 ;
  assign y19 = n518 ;
  assign y20 = n529 ;
  assign y21 = n530 ;
  assign y22 = n537 ;
endmodule
