module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 ;
  buffer buf_n66( .i (x2), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n124( .i (x4), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n94( .i (x3), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n154( .i (x5), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n212( .i (x7), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n240( .i (x8), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  assign n268 = n220 & ~n248 ;
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  assign n286 = ~n168 & n273 ;
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = ~n118 & n295 ;
  assign n297 = ( n91 & ~n149 ) | ( n91 & n296 ) | ( ~n149 & n296 ) ;
  assign n298 = ~n92 & n297 ;
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n10( .i (x0), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n38( .i (x1), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  assign n301 = n46 | n74 ;
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  assign n317 = n113 | n311 ;
  buffer buf_n318( .i (n317), .o (n318) );
  assign n319 = n31 & n318 ;
  assign n320 = n31 | n318 ;
  assign n321 = ~n319 & n320 ;
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  assign n324 = n218 | n246 ;
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  assign n342 = ( ~n222 & n269 ) | ( ~n222 & n327 ) | ( n269 & n327 ) ;
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  assign n362 = ~n130 & n160 ;
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  assign n380 = ~n113 & n374 ;
  buffer buf_n381( .i (n380), .o (n381) );
  assign n388 = ~n31 & n381 ;
  assign n389 = ~n314 & n388 ;
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  assign n390 = ~n103 & n133 ;
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  assign n405 = ~n83 & n397 ;
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n30), .o (n409) );
  assign n410 = n408 & ~n409 ;
  assign n411 = ~n60 & n410 ;
  assign n412 = ( n354 & n389 ) | ( n354 & n411 ) | ( n389 & n411 ) ;
  assign n413 = ~n322 & n412 ;
  assign n414 = ( n323 & n356 ) | ( n323 & n413 ) | ( n356 & n413 ) ;
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  assign n418 = ( n37 & n65 ) | ( n37 & ~n415 ) | ( n65 & ~n415 ) ;
  assign n419 = n299 & n418 ;
  assign n420 = ( n300 & n417 ) | ( n300 & ~n419 ) | ( n417 & ~n419 ) ;
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  assign n422 = n77 & n105 ;
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  assign n436 = ~n103 & n163 ;
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  assign n448 = n162 | n248 ;
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  assign n461 = n84 & n457 ;
  assign n462 = ( n429 & n445 ) | ( n429 & ~n461 ) | ( n445 & ~n461 ) ;
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  assign n465 = n58 | n232 ;
  assign n466 = ( n145 & n463 ) | ( n145 & n465 ) | ( n463 & n465 ) ;
  assign n467 = n464 & ~n466 ;
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  assign n470 = ( n76 & ~n164 ) | ( n76 & n222 ) | ( ~n164 & n222 ) ;
  buffer buf_n471( .i (n470), .o (n471) );
  assign n479 = ( ~n136 & n224 ) | ( ~n136 & n471 ) | ( n224 & n471 ) ;
  buffer buf_n480( .i (n479), .o (n480) );
  assign n483 = n226 & ~n480 ;
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  assign n486 = n482 | n484 ;
  assign n487 = ( ~n229 & n485 ) | ( ~n229 & n486 ) | ( n485 & n486 ) ;
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n182( .i (x6), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  assign n490 = ~n193 & n251 ;
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  assign n507 = ( n57 & ~n488 ) | ( n57 & n497 ) | ( ~n488 & n497 ) ;
  assign n508 = n489 & n507 ;
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  assign n511 = ~n167 & n195 ;
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  assign n524 = n79 | n137 ;
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  assign n532 = n516 & ~n529 ;
  assign n533 = ( n58 & ~n337 ) | ( n58 & n532 ) | ( ~n337 & n532 ) ;
  assign n534 = ~n59 & n533 ;
  assign n535 = ~n50 & n78 ;
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  assign n547 = n193 | n328 ;
  buffer buf_n548( .i (n547), .o (n548) );
  assign n556 = n167 & ~n548 ;
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  assign n562 = n107 & ~n137 ;
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  assign n574 = n561 & n567 ;
  assign n575 = n542 & n574 ;
  buffer buf_n576( .i (n575), .o (n576) );
  assign n577 = ( ~n509 & n534 ) | ( ~n509 & n576 ) | ( n534 & n576 ) ;
  assign n578 = n116 & ~n576 ;
  assign n579 = ( n510 & n577 ) | ( n510 & ~n578 ) | ( n577 & ~n578 ) ;
  assign n580 = n75 | n103 ;
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  assign n593 = n140 & ~n170 ;
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  assign n603 = n222 & n250 ;
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  assign n614 = n58 & n612 ;
  assign n615 = ( n591 & n597 ) | ( n591 & n614 ) | ( n597 & n614 ) ;
  assign n616 = ~n592 & n615 ;
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  assign n617 = ( n49 & n77 ) | ( n49 & ~n223 ) | ( n77 & ~n223 ) ;
  buffer buf_n618( .i (n617), .o (n618) );
  assign n629 = n225 | n618 ;
  assign n630 = ~n49 & n105 ;
  buffer buf_n631( .i (n630), .o (n631) );
  assign n639 = ( ~n79 & n618 ) | ( ~n79 & n631 ) | ( n618 & n631 ) ;
  assign n640 = ( ~n52 & n629 ) | ( ~n52 & n639 ) | ( n629 & n639 ) ;
  assign n641 = n255 & n640 ;
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  assign n644 = ( n81 & n109 ) | ( n81 & ~n227 ) | ( n109 & ~n227 ) ;
  assign n645 = ( n81 & n109 ) | ( n81 & n255 ) | ( n109 & n255 ) ;
  assign n646 = n644 & ~n645 ;
  assign n647 = n642 | n646 ;
  assign n648 = ( ~n56 & n643 ) | ( ~n56 & n647 ) | ( n643 & n647 ) ;
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  assign n652 = n135 & ~n223 ;
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  assign n663 = n51 & n225 ;
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n256( .i (n255), .o (n256) );
  assign n669 = ~n140 & n256 ;
  buffer buf_n670( .i (n669), .o (n670) );
  assign n673 = n56 & ~n670 ;
  assign n674 = ( n659 & n668 ) | ( n659 & ~n673 ) | ( n668 & ~n673 ) ;
  assign n675 = ( ~n86 & n649 ) | ( ~n86 & n674 ) | ( n649 & n674 ) ;
  assign n676 = n115 | n675 ;
  assign n677 = ( ~n116 & n651 ) | ( ~n116 & n676 ) | ( n651 & n676 ) ;
  assign n678 = n616 | n677 ;
  assign n679 = ( ~n468 & n579 ) | ( ~n468 & n678 ) | ( n579 & n678 ) ;
  assign n680 = n469 | n679 ;
  assign n681 = ~n36 & n680 ;
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  assign n684 = n106 | n136 ;
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  assign n697 = n522 & ~n696 ;
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  assign n698 = n87 & n401 ;
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  assign n701 = n23 & ~n51 ;
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  assign n712 = ~n587 & n704 ;
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  assign n723 = ( n433 & ~n699 ) | ( n433 & n717 ) | ( ~n699 & n717 ) ;
  assign n724 = ~n22 & n50 ;
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  assign n736 = n717 | n734 ;
  assign n737 = ( n700 & n723 ) | ( n700 & n736 ) | ( n723 & n736 ) ;
  buffer buf_n738( .i (n737), .o (n738) );
  assign n739 = ( ~n386 & n697 ) | ( ~n386 & n738 ) | ( n697 & n738 ) ;
  assign n740 = n49 & n77 ;
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  assign n752 = ~n26 & n744 ;
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  assign n763 = n738 | n761 ;
  assign n764 = ( n387 & n739 ) | ( n387 & n763 ) | ( n739 & n763 ) ;
  assign n765 = n682 | n764 ;
  assign n766 = ( n360 & n683 ) | ( n360 & n765 ) | ( n683 & n765 ) ;
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  assign n768 = ( n130 & n160 ) | ( n130 & ~n188 ) | ( n160 & ~n188 ) ;
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  assign n785 = ( ~n117 & n205 ) | ( ~n117 & n784 ) | ( n205 & n784 ) ;
  assign n786 = ( n117 & ~n147 ) | ( n117 & n784 ) | ( ~n147 & n784 ) ;
  assign n787 = n785 | n786 ;
  assign n788 = n91 & ~n787 ;
  assign n789 = ( n36 & n64 ) | ( n36 & n788 ) | ( n64 & n788 ) ;
  assign n790 = ~n37 & n789 ;
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  assign n793 = n133 & n163 ;
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  assign n809 = n112 & n801 ;
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  assign n819 = n22 & ~n106 ;
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n828( .i (n48), .o (n828) );
  assign n829 = ~n105 & n828 ;
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  assign n841 = ( n725 & n820 ) | ( n725 & ~n831 ) | ( n820 & ~n831 ) ;
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  assign n850 = ( n383 & ~n403 ) | ( n383 & n849 ) | ( ~n403 & n849 ) ;
  assign n851 = n734 | n849 ;
  assign n852 = ( n404 & n850 ) | ( n404 & n851 ) | ( n850 & n851 ) ;
  assign n853 = ~n91 & n852 ;
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n762( .i (n761), .o (n762) );
  assign n856 = n762 | n854 ;
  assign n857 = ( n818 & n855 ) | ( n818 & n856 ) | ( n855 & n856 ) ;
  buffer buf_n858( .i (n102), .o (n858) );
  assign n859 = ~n221 & n858 ;
  buffer buf_n860( .i (n859), .o (n860) );
  assign n866 = n162 & ~n220 ;
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  assign n880 = ( n437 & n860 ) | ( n437 & ~n868 ) | ( n860 & ~n868 ) ;
  buffer buf_n881( .i (n880), .o (n881) );
  assign n886 = n253 & n881 ;
  assign n887 = n80 & ~n886 ;
  assign n888 = n164 | n327 ;
  buffer buf_n889( .i (n888), .o (n889) );
  assign n896 = n106 & ~n889 ;
  assign n897 = n79 | n896 ;
  buffer buf_n898( .i (n897), .o (n898) );
  assign n904 = ~n887 & n898 ;
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  assign n907 = ( ~n141 & n199 ) | ( ~n141 & n905 ) | ( n199 & n905 ) ;
  assign n908 = n196 & n440 ;
  assign n909 = ( n81 & n607 ) | ( n81 & n908 ) | ( n607 & n908 ) ;
  assign n910 = ~n82 & n909 ;
  assign n911 = n141 & n910 ;
  assign n912 = ( n906 & ~n907 ) | ( n906 & n911 ) | ( ~n907 & n911 ) ;
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  assign n916 = n83 & ~n688 ;
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  assign n921 = ~n223 & n251 ;
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  assign n935 = ( n913 & n918 ) | ( n913 & n929 ) | ( n918 & n929 ) ;
  assign n936 = n518 & ~n935 ;
  assign n937 = ( n519 & n915 ) | ( n519 & ~n936 ) | ( n915 & ~n936 ) ;
  assign n938 = n61 & ~n937 ;
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n939( .i (n104), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  assign n941 = ( n194 & n252 ) | ( n194 & n940 ) | ( n252 & n940 ) ;
  buffer buf_n942( .i (n941), .o (n942) );
  assign n948 = ( ~n226 & n254 ) | ( ~n226 & n942 ) | ( n254 & n942 ) ;
  buffer buf_n949( .i (n948), .o (n949) );
  assign n952 = n256 & ~n949 ;
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  assign n955 = n951 | n953 ;
  assign n956 = ( ~n259 & n954 ) | ( ~n259 & n955 ) | ( n954 & n955 ) ;
  buffer buf_n957( .i (n80), .o (n957) );
  assign n958 = ~n169 & n957 ;
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  assign n965 = n84 & ~n960 ;
  buffer buf_n966( .i (n965), .o (n966) );
  assign n967 = n956 & n966 ;
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  assign n968 = ( n101 & n189 ) | ( n101 & ~n219 ) | ( n189 & ~n219 ) ;
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  assign n980 = ~n947 & n979 ;
  assign n981 = ( ~n962 & n966 ) | ( ~n962 & n980 ) | ( n966 & n980 ) ;
  assign n982 = ( ~n175 & n967 ) | ( ~n175 & n981 ) | ( n967 & n981 ) ;
  assign n983 = ~n146 & n982 ;
  assign n984 = n61 | n983 ;
  assign n985 = ~n938 & n984 ;
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  assign n988 = ( ~n52 & n168 ) | ( ~n52 & n226 ) | ( n168 & n226 ) ;
  assign n989 = ( n169 & n957 ) | ( n169 & n988 ) | ( n957 & n988 ) ;
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  assign n993 = ( n55 & ~n83 ) | ( n55 & n990 ) | ( ~n83 & n990 ) ;
  assign n994 = ~n230 & n993 ;
  assign n995 = ( ~n173 & n992 ) | ( ~n173 & n994 ) | ( n992 & n994 ) ;
  assign n996 = n144 | n995 ;
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  assign n997 = ~n163 & n221 ;
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  assign n1008 = n747 & n1006 ;
  assign n1009 = n144 & ~n1008 ;
  assign n1010 = n996 & ~n1009 ;
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  assign n1013 = ( n117 & ~n263 ) | ( n117 & n1011 ) | ( ~n263 & n1011 ) ;
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  assign n1014 = n167 & ~n330 ;
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  assign n1022 = ( n59 & ~n531 ) | ( n59 & n1021 ) | ( ~n531 & n1021 ) ;
  assign n1023 = ~n60 & n1022 ;
  buffer buf_n1024( .i (n116), .o (n1024) );
  assign n1025 = n1023 & ~n1024 ;
  assign n1026 = ( n1012 & ~n1013 ) | ( n1012 & n1025 ) | ( ~n1013 & n1025 ) ;
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  assign n1027 = ( n50 & n136 ) | ( n50 & ~n252 ) | ( n136 & ~n252 ) ;
  buffer buf_n1028( .i (n1027), .o (n1028) );
  assign n1033 = ( n80 & n254 ) | ( n80 & n1028 ) | ( n254 & n1028 ) ;
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  assign n1038 = ( n54 & n140 ) | ( n54 & n1034 ) | ( n140 & n1034 ) ;
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  assign n1041 = n1032 & ~n1039 ;
  assign n1042 = ( n1037 & ~n1040 ) | ( n1037 & n1041 ) | ( ~n1040 & n1041 ) ;
  assign n1043 = n114 | n1042 ;
  assign n1044 = n134 & n250 ;
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  assign n1052 = ( n84 & n142 ) | ( n84 & n1051 ) | ( n142 & n1051 ) ;
  assign n1053 = ~n57 & n1052 ;
  assign n1054 = n114 & ~n1053 ;
  assign n1055 = n1043 & ~n1054 ;
  assign n1056 = n107 & n137 ;
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  assign n1066 = ( n85 & ~n259 ) | ( n85 & n311 ) | ( ~n259 & n311 ) ;
  assign n1067 = ( n85 & n259 ) | ( n85 & ~n311 ) | ( n259 & ~n311 ) ;
  assign n1068 = ( ~n86 & n1066 ) | ( ~n86 & n1067 ) | ( n1066 & n1067 ) ;
  assign n1069 = ( n115 & n145 ) | ( n115 & n1068 ) | ( n145 & n1068 ) ;
  assign n1070 = ( n1055 & ~n1064 ) | ( n1055 & n1069 ) | ( ~n1064 & n1069 ) ;
  assign n1071 = n235 | n1070 ;
  buffer buf_n1072( .i (n82), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  assign n1074 = ( n56 & n112 ) | ( n56 & ~n1073 ) | ( n112 & ~n1073 ) ;
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n57), .o (n1076) );
  assign n1077 = ~n1075 & n1076 ;
  buffer buf_n1078( .i (n78), .o (n1078) );
  buffer buf_n1079( .i (n1078), .o (n1079) );
  assign n1080 = n138 & n1079 ;
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  assign n1088 = ( ~n114 & n1075 ) | ( ~n114 & n1085 ) | ( n1075 & n1085 ) ;
  assign n1089 = ( n87 & ~n1077 ) | ( n87 & n1088 ) | ( ~n1077 & n1088 ) ;
  assign n1090 = n262 & ~n1089 ;
  assign n1091 = n235 & ~n1090 ;
  assign n1092 = n1071 & ~n1091 ;
  assign n1093 = ( ~n35 & n1026 ) | ( ~n35 & n1092 ) | ( n1026 & n1092 ) ;
  assign n1094 = ~n986 & n1093 ;
  assign n1095 = ( ~n37 & n987 ) | ( ~n37 & n1094 ) | ( n987 & n1094 ) ;
  buffer buf_n1096( .i (n1095), .o (n1096) );
  assign n1097 = ( ~n791 & n857 ) | ( ~n791 & n1096 ) | ( n857 & n1096 ) ;
  assign n1098 = n360 | n1096 ;
  assign n1099 = ( n792 & n1097 ) | ( n792 & n1098 ) | ( n1097 & n1098 ) ;
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n1100( .i (n221), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  assign n1102 = ( n165 & n939 ) | ( n165 & ~n1101 ) | ( n939 & ~n1101 ) ;
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  assign n1108 = n168 & ~n1104 ;
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  assign n1111 = ( ~n228 & n256 ) | ( ~n228 & n1109 ) | ( n256 & n1109 ) ;
  assign n1112 = ( ~n1107 & n1110 ) | ( ~n1107 & n1111 ) | ( n1110 & n1111 ) ;
  assign n1113 = n1073 & n1112 ;
  assign n1114 = ( n102 & ~n220 ) | ( n102 & n248 ) | ( ~n220 & n248 ) ;
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  assign n1125 = ( ~n165 & n251 ) | ( ~n165 & n1116 ) | ( n251 & n1116 ) ;
  buffer buf_n1126( .i (n1125), .o (n1126) );
  assign n1129 = n253 & ~n1126 ;
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  assign n1132 = n1128 | n1130 ;
  buffer buf_n1133( .i (n255), .o (n1133) );
  assign n1134 = ( n1131 & n1132 ) | ( n1131 & ~n1133 ) | ( n1132 & ~n1133 ) ;
  buffer buf_n1135( .i (n1134), .o (n1135) );
  assign n1136 = n1073 | n1135 ;
  assign n1137 = ( ~n85 & n1113 ) | ( ~n85 & n1136 ) | ( n1113 & n1136 ) ;
  assign n1138 = n1076 & ~n1137 ;
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  assign n1139 = n170 & n275 ;
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  assign n1143 = n72 & ~n100 ;
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  assign n1156 = n1141 & n1155 ;
  assign n1157 = n1076 | n1156 ;
  assign n1158 = ~n1138 & n1157 ;
  assign n1159 = n146 & ~n1158 ;
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  assign n1160 = ( n165 & n939 ) | ( n165 & n1101 ) | ( n939 & n1101 ) ;
  buffer buf_n1161( .i (n1160), .o (n1161) );
  buffer buf_n1162( .i (n1161), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  assign n1168 = ( n111 & n257 ) | ( n111 & ~n1165 ) | ( n257 & ~n1165 ) ;
  assign n1169 = ( ~n225 & n253 ) | ( ~n225 & n1161 ) | ( n253 & n1161 ) ;
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  assign n1174 = ~n1168 & n1173 ;
  buffer buf_n1175( .i (n1073), .o (n1175) );
  assign n1176 = ~n1174 & n1175 ;
  assign n1177 = n903 & ~n1176 ;
  assign n1178 = ~n59 & n1177 ;
  assign n1179 = n146 | n1178 ;
  assign n1180 = ~n1159 & n1179 ;
  assign n1181 = n206 & ~n1180 ;
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  assign n1182 = n135 | n1101 ;
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1189( .i (n135), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  assign n1191 = ( n653 & n1183 ) | ( n653 & ~n1190 ) | ( n1183 & ~n1190 ) ;
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1203( .i (n254), .o (n1203) );
  assign n1204 = n1192 | n1203 ;
  assign n1205 = n170 | n1204 ;
  assign n1206 = n1072 & n1205 ;
  buffer buf_n1207( .i (n166), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  assign n1209 = n606 & n1208 ;
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1220( .i (n139), .o (n1220) );
  assign n1221 = n1210 & n1220 ;
  assign n1222 = n1072 | n1221 ;
  assign n1223 = ~n1206 & n1222 ;
  assign n1224 = n113 & n1223 ;
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  assign n1227 = n292 | n1225 ;
  assign n1228 = ( n920 & n1226 ) | ( n920 & n1227 ) | ( n1226 & n1227 ) ;
  assign n1229 = n61 & n1228 ;
  assign n1230 = n206 | n1229 ;
  assign n1231 = ~n1181 & n1230 ;
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  assign n1234 = n37 & n1232 ;
  assign n1235 = n196 & n273 ;
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  assign n1247 = n378 & n717 ;
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  assign n1250 = n1246 & n1249 ;
  assign n1251 = n563 & n957 ;
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1253( .i (n1252), .o (n1253) );
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  assign n1256 = n26 & n54 ;
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1260( .i (n55), .o (n1260) );
  assign n1261 = ~n1257 & n1260 ;
  buffer buf_n1262( .i (n1261), .o (n1262) );
  assign n1263 = n1255 & n1262 ;
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  assign n1264 = ( n407 & ~n1259 ) | ( n407 & n1262 ) | ( ~n1259 & n1262 ) ;
  assign n1265 = ( n409 & n1263 ) | ( n409 & n1264 ) | ( n1263 & n1264 ) ;
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  assign n1270 = ~n356 & n1268 ;
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  assign n1271 = ( n112 & ~n172 ) | ( n112 & n258 ) | ( ~n172 & n258 ) ;
  assign n1272 = n1124 & ~n1271 ;
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n219), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  assign n1277 = ( ~n249 & n858 ) | ( ~n249 & n1276 ) | ( n858 & n1276 ) ;
  assign n1278 = ( n134 & ~n250 ) | ( n134 & n1277 ) | ( ~n250 & n1277 ) ;
  buffer buf_n1279( .i (n1278), .o (n1279) );
  assign n1282 = n252 & n1279 ;
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  assign n1285 = n1281 & ~n1283 ;
  assign n1286 = ( n1203 & ~n1284 ) | ( n1203 & n1285 ) | ( ~n1284 & n1285 ) ;
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  assign n1289 = ( ~n171 & n1072 ) | ( ~n171 & n1287 ) | ( n1072 & n1287 ) ;
  assign n1290 = n139 & n274 ;
  assign n1291 = ~n586 & n1290 ;
  assign n1292 = ~n171 & n1291 ;
  assign n1293 = ( ~n1288 & n1289 ) | ( ~n1288 & n1292 ) | ( n1289 & n1292 ) ;
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  assign n1297 = ( n86 & n144 ) | ( n86 & ~n1294 ) | ( n144 & ~n1294 ) ;
  assign n1298 = n1273 & n1297 ;
  assign n1299 = ( n1274 & n1296 ) | ( n1274 & ~n1298 ) | ( n1296 & ~n1298 ) ;
  buffer buf_n1300( .i (n60), .o (n1300) );
  assign n1301 = ( ~n33 & n1299 ) | ( ~n33 & n1300 ) | ( n1299 & n1300 ) ;
  assign n1302 = n922 & n1207 ;
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  assign n1310 = ~n1078 & n1190 ;
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  assign n1318 = n141 & ~n1313 ;
  buffer buf_n1319( .i (n1318), .o (n1319) );
  assign n1320 = n1307 & n1319 ;
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  assign n1321 = ( n290 & ~n1315 ) | ( n290 & n1319 ) | ( ~n1315 & n1319 ) ;
  buffer buf_n1322( .i (n1175), .o (n1322) );
  assign n1323 = ( n1320 & n1321 ) | ( n1320 & ~n1322 ) | ( n1321 & ~n1322 ) ;
  assign n1324 = n115 | n1323 ;
  buffer buf_n1325( .i (n249), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  assign n1328 = ( n224 & n1189 ) | ( n224 & n1327 ) | ( n1189 & n1327 ) ;
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1334( .i (n1327), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  assign n1336 = ( n1208 & n1329 ) | ( n1208 & ~n1335 ) | ( n1329 & ~n1335 ) ;
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  assign n1341 = ( n228 & n1220 ) | ( n228 & n1337 ) | ( n1220 & n1337 ) ;
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  assign n1344 = ~n1333 & n1342 ;
  assign n1345 = ( ~n1340 & n1343 ) | ( ~n1340 & n1344 ) | ( n1343 & n1344 ) ;
  assign n1346 = ~n1322 & n1345 ;
  buffer buf_n1347( .i (n111), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  assign n1351 = ~n1346 & n1350 ;
  assign n1352 = n1324 & ~n1351 ;
  assign n1353 = ( n33 & n1300 ) | ( n33 & ~n1352 ) | ( n1300 & ~n1352 ) ;
  assign n1354 = n1301 & ~n1353 ;
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  assign n1355 = ( n110 & n1133 ) | ( n110 & n1186 ) | ( n1133 & n1186 ) ;
  buffer buf_n1356( .i (n1355), .o (n1356) );
  assign n1357 = n230 & ~n1356 ;
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  assign n1358 = ( ~n142 & n1188 ) | ( ~n142 & n1356 ) | ( n1188 & n1356 ) ;
  assign n1359 = ( ~n231 & n1357 ) | ( ~n231 & n1358 ) | ( n1357 & n1358 ) ;
  assign n1360 = ( ~n1076 & n1322 ) | ( ~n1076 & n1359 ) | ( n1322 & n1359 ) ;
  assign n1361 = ~n940 & n1327 ;
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  assign n1371 = ( ~n142 & n230 ) | ( ~n142 & n1366 ) | ( n230 & n1366 ) ;
  buffer buf_n1372( .i (n1220), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  assign n1374 = ( ~n258 & n1366 ) | ( ~n258 & n1373 ) | ( n1366 & n1373 ) ;
  assign n1375 = ( n1348 & n1371 ) | ( n1348 & n1374 ) | ( n1371 & n1374 ) ;
  buffer buf_n1376( .i (n1260), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  assign n1378 = ( n1322 & ~n1375 ) | ( n1322 & n1377 ) | ( ~n1375 & n1377 ) ;
  assign n1379 = n1360 & ~n1378 ;
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  assign n1382 = n1079 | n1335 ;
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1386( .i (n1385), .o (n1386) );
  assign n1389 = ( n143 & ~n231 ) | ( n143 & n1386 ) | ( ~n231 & n1386 ) ;
  assign n1390 = ( n143 & n1175 ) | ( n143 & ~n1386 ) | ( n1175 & ~n1386 ) ;
  assign n1391 = ( n260 & ~n1389 ) | ( n260 & n1390 ) | ( ~n1389 & n1390 ) ;
  buffer buf_n1392( .i (n1377), .o (n1392) );
  assign n1393 = ( ~n1350 & n1391 ) | ( ~n1350 & n1392 ) | ( n1391 & n1392 ) ;
  buffer buf_n1394( .i (n1175), .o (n1394) );
  assign n1395 = ( n337 & n530 ) | ( n337 & ~n1394 ) | ( n530 & ~n1394 ) ;
  assign n1396 = ( n1350 & n1392 ) | ( n1350 & ~n1395 ) | ( n1392 & ~n1395 ) ;
  assign n1397 = n1393 & n1396 ;
  buffer buf_n930( .i (n929), .o (n930) );
  assign n1398 = n26 & ~n308 ;
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  assign n1407 = ~n690 & n1400 ;
  buffer buf_n1408( .i (n1407), .o (n1408) );
  assign n1412 = n930 & n1408 ;
  buffer buf_n1413( .i (n1412), .o (n1413) );
  assign n1414 = ( ~n1380 & n1397 ) | ( ~n1380 & n1413 ) | ( n1397 & n1413 ) ;
  assign n1415 = n33 & ~n1413 ;
  assign n1416 = ( n1381 & n1414 ) | ( n1381 & ~n1415 ) | ( n1414 & ~n1415 ) ;
  assign n1417 = n1354 | n1416 ;
  assign n1418 = ( n1269 & ~n1270 ) | ( n1269 & n1417 ) | ( ~n1270 & n1417 ) ;
  assign n1419 = n1250 | n1418 ;
  assign n1420 = ( n1233 & ~n1234 ) | ( n1233 & n1419 ) | ( ~n1234 & n1419 ) ;
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  assign n1423 = n132 & ~n190 ;
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1434( .i (n1433), .o (n1434) );
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n207( .i (n206), .o (n207) );
  assign n1445 = ~n171 & n609 ;
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  assign n1450 = ( n166 & ~n940 ) | ( n166 & n1327 ) | ( ~n940 & n1327 ) ;
  buffer buf_n1451( .i (n1450), .o (n1451) );
  assign n1452 = ( n138 & ~n1335 ) | ( n138 & n1451 ) | ( ~n1335 & n1451 ) ;
  assign n1453 = ( n138 & n1208 ) | ( n138 & ~n1451 ) | ( n1208 & ~n1451 ) ;
  assign n1454 = n1452 & ~n1453 ;
  buffer buf_n1455( .i (n1454), .o (n1455) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  assign n1457 = ( ~n55 & n229 ) | ( ~n55 & n1455 ) | ( n229 & n1455 ) ;
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n1458( .i (n1190), .o (n1458) );
  assign n1459 = n632 & n1458 ;
  assign n1460 = ( n169 & n1203 ) | ( n169 & n1459 ) | ( n1203 & n1459 ) ;
  assign n1461 = ~n1133 & n1460 ;
  assign n1462 = ~n229 & n1461 ;
  assign n1463 = ( n1456 & ~n1457 ) | ( n1456 & n1462 ) | ( ~n1457 & n1462 ) ;
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n568( .i (n567), .o (n568) );
  assign n1467 = ( n568 & ~n1377 ) | ( n568 & n1464 ) | ( ~n1377 & n1464 ) ;
  assign n1468 = n1448 & ~n1467 ;
  assign n1469 = ( n1449 & n1466 ) | ( n1449 & ~n1468 ) | ( n1466 & ~n1468 ) ;
  assign n1470 = n89 & ~n1469 ;
  assign n1471 = ( n110 & n228 ) | ( n110 & n1220 ) | ( n228 & n1220 ) ;
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1326), .o (n1475) );
  assign n1476 = ( n940 & n1189 ) | ( n940 & ~n1475 ) | ( n1189 & ~n1475 ) ;
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  assign n1484 = n1474 & ~n1483 ;
  assign n1485 = n175 & n1484 ;
  buffer buf_n1486( .i (n1392), .o (n1486) );
  assign n1487 = n1485 & ~n1486 ;
  assign n1488 = n89 | n1487 ;
  assign n1489 = ~n1470 & n1488 ;
  assign n1490 = ( ~n35 & n207 ) | ( ~n35 & n1489 ) | ( n207 & n1489 ) ;
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  assign n1491 = ~n51 & n1190 ;
  buffer buf_n1492( .i (n1491), .o (n1492) );
  assign n1497 = n139 & ~n1492 ;
  buffer buf_n1498( .i (n1497), .o (n1498) );
  assign n1499 = n885 & n1498 ;
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1500( .i (n164), .o (n1500) );
  assign n1501 = n1101 | n1500 ;
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  assign n1514 = ( n1494 & ~n1498 ) | ( n1494 & n1506 ) | ( ~n1498 & n1506 ) ;
  assign n1515 = ( n1260 & ~n1499 ) | ( n1260 & n1514 ) | ( ~n1499 & n1514 ) ;
  buffer buf_n1516( .i (n82), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1518( .i (n1517), .o (n1518) );
  assign n1519 = n1515 & ~n1518 ;
  buffer buf_n1520( .i (n162), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  assign n1522 = ( n48 & n104 ) | ( n48 & n1521 ) | ( n104 & n1521 ) ;
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1528( .i (n939), .o (n1528) );
  assign n1529 = ( n224 & n1523 ) | ( n224 & ~n1528 ) | ( n1523 & ~n1528 ) ;
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  assign n1534 = ( n52 & n1208 ) | ( n52 & n1530 ) | ( n1208 & n1530 ) ;
  buffer buf_n1535( .i (n1534), .o (n1535) );
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  assign n1537 = n1527 & ~n1535 ;
  assign n1538 = ( n1533 & ~n1536 ) | ( n1533 & n1537 ) | ( ~n1536 & n1537 ) ;
  assign n1539 = ~n1373 & n1538 ;
  assign n1540 = n1518 & ~n1539 ;
  assign n1541 = n1519 | n1540 ;
  assign n1542 = n261 | n1541 ;
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  assign n1545 = ~n110 & n1210 ;
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n145), .o (n1551) );
  assign n1552 = n1550 & ~n1551 ;
  assign n1553 = n1543 & ~n1552 ;
  assign n1554 = ( n62 & n1544 ) | ( n62 & n1553 ) | ( n1544 & n1553 ) ;
  assign n1555 = ( n35 & n207 ) | ( n35 & n1554 ) | ( n207 & n1554 ) ;
  assign n1556 = n1490 & ~n1555 ;
  buffer buf_n1557( .i (n1556), .o (n1557) );
  buffer buf_n1558( .i (n1557), .o (n1558) );
  assign n1559 = n166 | n1528 ;
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  assign n1566 = n143 | n1565 ;
  buffer buf_n1567( .i (n1566), .o (n1567) );
  assign n1570 = n23 & n1078 ;
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  assign n1578 = n29 & ~n1575 ;
  buffer buf_n1579( .i (n1578), .o (n1579) );
  assign n1580 = ~n1567 & n1579 ;
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  assign n1581 = ( n811 & ~n1577 ) | ( n811 & n1579 ) | ( ~n1577 & n1579 ) ;
  assign n1582 = ( n88 & n1580 ) | ( n88 & n1581 ) | ( n1580 & n1581 ) ;
  assign n1583 = n1300 | n1582 ;
  buffer buf_n1584( .i (n1207), .o (n1584) );
  assign n1585 = ( n1079 & n1458 ) | ( n1079 & ~n1584 ) | ( n1458 & ~n1584 ) ;
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  assign n1592 = n172 | n1588 ;
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  assign n1595 = ( n1349 & n1394 ) | ( n1349 & ~n1593 ) | ( n1394 & ~n1593 ) ;
  assign n1596 = ( n1591 & n1594 ) | ( n1591 & ~n1595 ) | ( n1594 & ~n1595 ) ;
  assign n1597 = n32 | n1596 ;
  assign n1598 = n1300 & n1597 ;
  assign n1599 = n1583 & ~n1598 ;
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  assign n1602 = ~n238 & n1600 ;
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  assign n1603 = n759 & ~n1513 ;
  assign n1604 = ~n696 & n1603 ;
  buffer buf_n1605( .i (n134), .o (n1605) );
  buffer buf_n1606( .i (n1100), .o (n1606) );
  assign n1607 = n1605 & n1606 ;
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n1613( .i (n1612), .o (n1613) );
  assign n1616 = ( n257 & ~n1313 ) | ( n257 & n1372 ) | ( ~n1313 & n1372 ) ;
  buffer buf_n1617( .i (n227), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  assign n1619 = ( ~n257 & n1313 ) | ( ~n257 & n1618 ) | ( n1313 & n1618 ) ;
  assign n1620 = ( ~n1613 & n1616 ) | ( ~n1613 & n1619 ) | ( n1616 & n1619 ) ;
  assign n1621 = n173 & n1620 ;
  buffer buf_n1622( .i (n1606), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  assign n1625 = ( ~n1079 & n1335 ) | ( ~n1079 & n1624 ) | ( n1335 & n1624 ) ;
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  assign n1631 = ~n1617 & n1626 ;
  assign n1632 = ( n1516 & n1627 ) | ( n1516 & n1631 ) | ( n1627 & n1631 ) ;
  assign n1633 = n1373 & n1632 ;
  assign n1634 = n173 | n1633 ;
  assign n1635 = ~n1621 & n1634 ;
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  assign n1636 = ( n368 & n653 ) | ( n368 & ~n870 ) | ( n653 & ~n870 ) ;
  buffer buf_n1637( .i (n1636), .o (n1637) );
  assign n1640 = ( n957 & n1203 ) | ( n957 & n1637 ) | ( n1203 & n1637 ) ;
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1133), .o (n1642) );
  assign n1643 = ( n27 & n1641 ) | ( n27 & ~n1642 ) | ( n1641 & ~n1642 ) ;
  assign n1644 = ( n27 & n1516 ) | ( n27 & ~n1641 ) | ( n1516 & ~n1641 ) ;
  assign n1645 = n1643 & ~n1644 ;
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  assign n1648 = n30 & ~n1646 ;
  assign n1649 = ( n1635 & n1647 ) | ( n1635 & ~n1648 ) | ( n1647 & ~n1648 ) ;
  buffer buf_n1650( .i (n1350), .o (n1650) );
  assign n1651 = n1649 | n1650 ;
  assign n1652 = n527 & n1642 ;
  assign n1653 = ( n610 & n658 ) | ( n610 & ~n1652 ) | ( n658 & ~n1652 ) ;
  buffer buf_n1654( .i (n172), .o (n1654) );
  assign n1655 = n1653 | n1654 ;
  assign n1656 = n335 | n528 ;
  assign n1657 = n1654 & n1656 ;
  assign n1658 = n1655 & ~n1657 ;
  assign n1659 = ~n409 & n1658 ;
  assign n1660 = n1650 & ~n1659 ;
  assign n1661 = n1651 & ~n1660 ;
  assign n1662 = n62 | n1661 ;
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  assign n1663 = n919 & ~n1309 ;
  buffer buf_n1664( .i (n133), .o (n1664) );
  assign n1665 = ( ~n76 & n1521 ) | ( ~n76 & n1664 ) | ( n1521 & n1664 ) ;
  buffer buf_n1666( .i (n1665), .o (n1666) );
  assign n1672 = ( n78 & ~n1622 ) | ( n78 & n1666 ) | ( ~n1622 & n1666 ) ;
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  assign n1677 = ( n1458 & n1584 ) | ( n1458 & n1673 ) | ( n1584 & n1673 ) ;
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  assign n1680 = ~n1670 & n1678 ;
  assign n1681 = ( ~n1676 & n1679 ) | ( ~n1676 & n1680 ) | ( n1679 & n1680 ) ;
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n258), .o (n1684) );
  assign n1685 = ( ~n1348 & n1682 ) | ( ~n1348 & n1684 ) | ( n1682 & n1684 ) ;
  assign n1686 = ~n581 & n1605 ;
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  assign n1694 = ~n1507 & n1692 ;
  assign n1695 = ~n1684 & n1694 ;
  assign n1696 = ( n1683 & ~n1685 ) | ( n1683 & n1695 ) | ( ~n1685 & n1695 ) ;
  assign n1697 = ~n1082 & n1516 ;
  buffer buf_n1698( .i (n1697), .o (n1698) );
  assign n1699 = n1446 & n1698 ;
  assign n1700 = ( n1019 & ~n1084 ) | ( n1019 & n1698 ) | ( ~n1084 & n1698 ) ;
  buffer buf_n1701( .i (n1373), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  assign n1703 = ( n1699 & n1700 ) | ( n1699 & n1702 ) | ( n1700 & n1702 ) ;
  assign n1704 = n1696 | n1703 ;
  assign n1705 = ( n920 & ~n1663 ) | ( n920 & n1704 ) | ( ~n1663 & n1704 ) ;
  buffer buf_n1706( .i (n32), .o (n1706) );
  assign n1707 = n1705 & ~n1706 ;
  assign n1708 = n62 & ~n1707 ;
  assign n1709 = n1662 & ~n1708 ;
  assign n1710 = n1604 | n1709 ;
  assign n1711 = ( n1601 & ~n1602 ) | ( n1601 & n1710 ) | ( ~n1602 & n1710 ) ;
  assign n1712 = n132 | n190 ;
  buffer buf_n1713( .i (n1712), .o (n1713) );
  assign n1732 = ( n1424 & ~n1664 ) | ( n1424 & n1713 ) | ( ~n1664 & n1713 ) ;
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1078), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  assign n1747 = n1642 & ~n1746 ;
  buffer buf_n1748( .i (n1747), .o (n1748) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  assign n1751 = ( n1349 & n1741 ) | ( n1349 & ~n1749 ) | ( n1741 & ~n1749 ) ;
  assign n1752 = n1742 & ~n1751 ;
  assign n1753 = n1486 | n1752 ;
  assign n1754 = n194 | n1475 ;
  buffer buf_n1755( .i (n1754), .o (n1755) );
  assign n1763 = n1458 & ~n1755 ;
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  assign n1770 = n431 & n1769 ;
  assign n1771 = n1486 & ~n1770 ;
  assign n1772 = n1753 & ~n1771 ;
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n871( .i (n870), .o (n871) );
  assign n1775 = ( n871 & n1503 ) | ( n871 & ~n1584 ) | ( n1503 & ~n1584 ) ;
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n34), .o (n1786) );
  assign n1787 = ( n1773 & ~n1785 ) | ( n1773 & n1786 ) | ( ~n1785 & n1786 ) ;
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  assign n1788 = n260 & n400 ;
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  assign n1791 = ( n205 & n1404 ) | ( n205 & n1790 ) | ( n1404 & n1790 ) ;
  assign n1792 = ~n206 & n1791 ;
  assign n1793 = n1785 & n1792 ;
  assign n1794 = ( n1774 & ~n1787 ) | ( n1774 & n1793 ) | ( ~n1787 & n1793 ) ;
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  assign n1795 = ~n130 & n188 ;
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  buffer buf_n1813( .i (n1812), .o (n1813) );
  assign n1814 = n934 & n1813 ;
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n1815( .i (n1334), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  assign n1817 = ( n53 & n1744 ) | ( n53 & ~n1816 ) | ( n1744 & ~n1816 ) ;
  assign n1818 = n621 & ~n1817 ;
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  buffer buf_n1821( .i (n1820), .o (n1821) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  assign n1822 = ( n277 & ~n310 ) | ( n277 & n1819 ) | ( ~n310 & n1819 ) ;
  assign n1823 = n1348 & ~n1822 ;
  assign n1824 = ( n1349 & n1821 ) | ( n1349 & ~n1823 ) | ( n1821 & ~n1823 ) ;
  buffer buf_n1825( .i (n1189), .o (n1825) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1827( .i (n1826), .o (n1827) );
  assign n1828 = n197 & n1827 ;
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  assign n1834 = n201 & ~n1831 ;
  buffer buf_n1835( .i (n1834), .o (n1835) );
  assign n1836 = n1824 & n1835 ;
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  assign n1837 = ( n108 & n1743 ) | ( n108 & ~n1815 ) | ( n1743 & ~n1815 ) ;
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n109), .o (n1842) );
  assign n1843 = n1838 & ~n1842 ;
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  assign n1846 = ( n1260 & n1517 ) | ( n1260 & ~n1844 ) | ( n1517 & ~n1844 ) ;
  assign n1847 = ( n1841 & n1845 ) | ( n1841 & ~n1846 ) | ( n1845 & ~n1846 ) ;
  assign n1848 = n231 | n1820 ;
  assign n1849 = ( n1821 & n1847 ) | ( n1821 & n1848 ) | ( n1847 & n1848 ) ;
  assign n1850 = ( ~n1833 & n1835 ) | ( ~n1833 & n1849 ) | ( n1835 & n1849 ) ;
  assign n1851 = ( n1551 & n1836 ) | ( n1551 & n1850 ) | ( n1836 & n1850 ) ;
  assign n1852 = ~n1706 & n1851 ;
  buffer buf_n1853( .i (n1852), .o (n1853) );
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  assign n1855 = n719 | n1853 ;
  assign n1856 = ( n1814 & n1854 ) | ( n1814 & n1855 ) | ( n1854 & n1855 ) ;
  assign n1857 = n1794 | n1856 ;
  assign n1858 = ( ~n1557 & n1711 ) | ( ~n1557 & n1857 ) | ( n1711 & n1857 ) ;
  assign n1859 = n1558 | n1858 ;
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  assign n1860 = ( n76 & n1100 ) | ( n76 & ~n1325 ) | ( n1100 & ~n1325 ) ;
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  buffer buf_n1872( .i (n1871), .o (n1872) );
  assign n1873 = ( n1100 & n1325 ) | ( n1100 & n1521 ) | ( n1325 & n1521 ) ;
  buffer buf_n1874( .i (n1873), .o (n1874) );
  buffer buf_n1875( .i (n1874), .o (n1875) );
  buffer buf_n1876( .i (n1875), .o (n1876) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  buffer buf_n1878( .i (n1877), .o (n1878) );
  buffer buf_n1879( .i (n1878), .o (n1879) );
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  assign n1886 = ~n1872 & n1885 ;
  buffer buf_n1887( .i (n1584), .o (n1887) );
  buffer buf_n1888( .i (n1887), .o (n1888) );
  buffer buf_n1889( .i (n1888), .o (n1889) );
  buffer buf_n1890( .i (n1889), .o (n1890) );
  assign n1891 = ( n349 & n1517 ) | ( n349 & n1890 ) | ( n1517 & n1890 ) ;
  buffer buf_n1892( .i (n1891), .o (n1892) );
  assign n1893 = ( n30 & ~n174 ) | ( n30 & n1892 ) | ( ~n174 & n1892 ) ;
  buffer buf_n1894( .i (n29), .o (n1894) );
  assign n1895 = ( n1394 & ~n1892 ) | ( n1394 & n1894 ) | ( ~n1892 & n1894 ) ;
  assign n1896 = n1893 & ~n1895 ;
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  assign n1899 = n1706 & ~n1897 ;
  assign n1900 = ( n1886 & n1898 ) | ( n1886 & ~n1899 ) | ( n1898 & ~n1899 ) ;
  assign n1901 = n63 | n1900 ;
  assign n1902 = ( n1618 & ~n1627 ) | ( n1618 & n1889 ) | ( ~n1627 & n1889 ) ;
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1907( .i (n1906), .o (n1907) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1908( .i (n1618), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  assign n1910 = ( n1684 & n1903 ) | ( n1684 & ~n1909 ) | ( n1903 & ~n1909 ) ;
  assign n1911 = n1630 & n1910 ;
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n176( .i (n175), .o (n176) );
  assign n1914 = n176 & ~n1912 ;
  assign n1915 = ( n1907 & n1913 ) | ( n1907 & ~n1914 ) | ( n1913 & ~n1914 ) ;
  assign n1916 = ~n34 & n1915 ;
  assign n1917 = n63 & ~n1916 ;
  assign n1918 = n1901 & ~n1917 ;
  assign n1919 = n121 | n1918 ;
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  assign n1920 = ( n53 & n1744 ) | ( n53 & n1816 ) | ( n1744 & n1816 ) ;
  buffer buf_n1921( .i (n1920), .o (n1921) );
  assign n1926 = ( n1618 & ~n1642 ) | ( n1618 & n1921 ) | ( ~n1642 & n1921 ) ;
  buffer buf_n1927( .i (n1926), .o (n1927) );
  buffer buf_n1928( .i (n1927), .o (n1928) );
  buffer buf_n1929( .i (n1928), .o (n1929) );
  buffer buf_n1930( .i (n1929), .o (n1930) );
  assign n1931 = ( n1376 & n1518 ) | ( n1376 & n1927 ) | ( n1518 & n1927 ) ;
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1925( .i (n1924), .o (n1925) );
  assign n1934 = n1925 & ~n1932 ;
  assign n1935 = ( n1930 & ~n1933 ) | ( n1930 & n1934 ) | ( ~n1933 & n1934 ) ;
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n828), .o (n1938) );
  buffer buf_n1939( .i (n75), .o (n1939) );
  buffer buf_n1940( .i (n1939), .o (n1940) );
  buffer buf_n1941( .i (n1940), .o (n1941) );
  assign n1942 = n1938 & ~n1941 ;
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  assign n1954 = n1936 | n1953 ;
  assign n1955 = ( n1219 & n1937 ) | ( n1219 & n1954 ) | ( n1937 & n1954 ) ;
  assign n1956 = ~n36 & n1955 ;
  assign n1957 = n121 & ~n1956 ;
  assign n1958 = n1919 & ~n1957 ;
  assign n1959 = ( n153 & ~n211 ) | ( n153 & n1958 ) | ( ~n211 & n1958 ) ;
  assign n1960 = ( ~n1444 & n1859 ) | ( ~n1444 & n1959 ) | ( n1859 & n1959 ) ;
  buffer buf_n177( .i (n176), .o (n177) );
  assign n1961 = ( n27 & ~n1372 ) | ( n27 & n1889 ) | ( ~n1372 & n1889 ) ;
  assign n1962 = ( ~n1347 & n1890 ) | ( ~n1347 & n1961 ) | ( n1890 & n1961 ) ;
  buffer buf_n1963( .i (n1962), .o (n1963) );
  assign n1966 = n174 & ~n1963 ;
  buffer buf_n1967( .i (n1966), .o (n1967) );
  buffer buf_n1968( .i (n1967), .o (n1968) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  assign n1969 = n1965 | n1967 ;
  assign n1970 = ( ~n177 & n1968 ) | ( ~n177 & n1969 ) | ( n1968 & n1969 ) ;
  assign n1971 = n90 | n1970 ;
  buffer buf_n1972( .i (n1827), .o (n1972) );
  assign n1973 = ( n1842 & n1888 ) | ( n1842 & ~n1972 ) | ( n1888 & ~n1972 ) ;
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  assign n1978 = n203 | n1977 ;
  assign n1979 = ( ~n175 & n203 ) | ( ~n175 & n1977 ) | ( n203 & n1977 ) ;
  assign n1980 = ( n176 & ~n1978 ) | ( n176 & n1979 ) | ( ~n1978 & n1979 ) ;
  assign n1981 = ~n1706 & n1980 ;
  assign n1982 = n90 & ~n1981 ;
  assign n1983 = n1971 & ~n1982 ;
  assign n1984 = n64 | n1983 ;
  buffer buf_n1985( .i (n108), .o (n1985) );
  assign n1986 = ( ~n1744 & n1887 ) | ( ~n1744 & n1985 ) | ( n1887 & n1985 ) ;
  buffer buf_n1987( .i (n1986), .o (n1987) );
  assign n1992 = ( ~n1372 & n1746 ) | ( ~n1372 & n1987 ) | ( n1746 & n1987 ) ;
  buffer buf_n1993( .i (n1992), .o (n1993) );
  buffer buf_n1994( .i (n1993), .o (n1994) );
  buffer buf_n1995( .i (n1994), .o (n1995) );
  buffer buf_n1996( .i (n1995), .o (n1996) );
  buffer buf_n1997( .i (n1347), .o (n1997) );
  assign n1998 = ( n1654 & n1993 ) | ( n1654 & n1997 ) | ( n1993 & n1997 ) ;
  buffer buf_n1999( .i (n1998), .o (n1999) );
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n1988( .i (n1987), .o (n1988) );
  buffer buf_n1989( .i (n1988), .o (n1989) );
  buffer buf_n1990( .i (n1989), .o (n1990) );
  buffer buf_n1991( .i (n1990), .o (n1991) );
  assign n2001 = ~n1991 & n1999 ;
  assign n2002 = ( ~n1996 & n2000 ) | ( ~n1996 & n2001 ) | ( n2000 & n2001 ) ;
  assign n2003 = n205 & ~n2002 ;
  buffer buf_n2004( .i (n1941), .o (n2004) );
  assign n2005 = ~n1825 & n2004 ;
  buffer buf_n2006( .i (n2005), .o (n2006) );
  buffer buf_n2007( .i (n2006), .o (n2007) );
  buffer buf_n2008( .i (n2007), .o (n2008) );
  buffer buf_n2009( .i (n2008), .o (n2009) );
  buffer buf_n2010( .i (n2009), .o (n2010) );
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n2012( .i (n2011), .o (n2012) );
  buffer buf_n2016( .i (n1702), .o (n2016) );
  assign n2017 = ( ~n401 & n2012 ) | ( ~n401 & n2016 ) | ( n2012 & n2016 ) ;
  assign n2018 = n176 | n2017 ;
  buffer buf_n2019( .i (n204), .o (n2019) );
  assign n2020 = n2018 & ~n2019 ;
  assign n2021 = n2003 | n2020 ;
  assign n2022 = n1786 | n2021 ;
  assign n2023 = n64 & n2022 ;
  assign n2024 = n1984 & ~n2023 ;
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  assign n2027 = n360 & n2025 ;
  assign n2028 = ~n200 & n1778 ;
  buffer buf_n2029( .i (n1972), .o (n2029) );
  assign n2030 = ~n1082 & n2029 ;
  buffer buf_n2031( .i (n2030), .o (n2031) );
  assign n2032 = n2028 & n2031 ;
  assign n2033 = ~n191 & n1276 ;
  buffer buf_n2034( .i (n2033), .o (n2034) );
  assign n2051 = ~n1500 & n2034 ;
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  buffer buf_n2055( .i (n2054), .o (n2055) );
  buffer buf_n2056( .i (n2055), .o (n2056) );
  buffer buf_n2057( .i (n2056), .o (n2057) );
  assign n2059 = n196 & n871 ;
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  assign n2063 = n2057 | n2062 ;
  assign n2064 = ( ~n1084 & n2031 ) | ( ~n1084 & n2063 ) | ( n2031 & n2063 ) ;
  assign n2065 = ( n1394 & n2032 ) | ( n1394 & n2064 ) | ( n2032 & n2064 ) ;
  assign n2066 = n1392 & ~n2065 ;
  buffer buf_n2067( .i (n1276), .o (n2067) );
  assign n2068 = ( n1521 & n1664 ) | ( n1521 & ~n2067 ) | ( n1664 & ~n2067 ) ;
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n2073( .i (n2072), .o (n2073) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n2075( .i (n2074), .o (n2075) );
  buffer buf_n2076( .i (n2075), .o (n2076) );
  assign n2077 = n1972 & ~n2073 ;
  buffer buf_n2078( .i (n2077), .o (n2078) );
  buffer buf_n2079( .i (n2078), .o (n2079) );
  assign n2080 = ( n200 & n1890 ) | ( n200 & n2078 ) | ( n1890 & n2078 ) ;
  assign n2081 = ( ~n2076 & n2079 ) | ( ~n2076 & n2080 ) | ( n2079 & n2080 ) ;
  buffer buf_n2082( .i (n1518), .o (n2082) );
  assign n2083 = n2081 & ~n2082 ;
  buffer buf_n2084( .i (n1377), .o (n2084) );
  assign n2085 = n2083 | n2084 ;
  assign n2086 = ~n2066 & n2085 ;
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  assign n2089 = ( n34 & ~n118 ) | ( n34 & n2087 ) | ( ~n118 & n2087 ) ;
  assign n2090 = n193 | n1606 ;
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n2099( .i (n2098), .o (n2099) );
  buffer buf_n2100( .i (n2099), .o (n2100) );
  assign n2104 = ~n591 & n597 ;
  assign n2105 = ( n1486 & ~n2100 ) | ( n1486 & n2104 ) | ( ~n2100 & n2104 ) ;
  buffer buf_n2106( .i (n2084), .o (n2106) );
  buffer buf_n2107( .i (n2106), .o (n2107) );
  assign n2108 = n2105 & ~n2107 ;
  buffer buf_n2109( .i (n32), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  assign n2111 = n2108 & ~n2110 ;
  assign n2112 = ( n2088 & ~n2089 ) | ( n2088 & n2111 ) | ( ~n2089 & n2111 ) ;
  buffer buf_n2113( .i (n2112), .o (n2113) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  assign n2115 = n192 & n2067 ;
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n2118( .i (n2117), .o (n2118) );
  buffer buf_n2119( .i (n2118), .o (n2119) );
  buffer buf_n2120( .i (n2119), .o (n2120) );
  buffer buf_n2121( .i (n2120), .o (n2121) );
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  buffer buf_n2129( .i (n2128), .o (n2129) );
  assign n2130 = n719 & n2129 ;
  assign n2131 = n602 & n2130 ;
  buffer buf_n2132( .i (n195), .o (n2132) );
  assign n2133 = n923 & n2132 ;
  buffer buf_n2134( .i (n2133), .o (n2134) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  buffer buf_n2137( .i (n2136), .o (n2137) );
  buffer buf_n2138( .i (n2137), .o (n2138) );
  buffer buf_n2139( .i (n2138), .o (n2139) );
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n2143( .i (n2142), .o (n2143) );
  buffer buf_n633( .i (n632), .o (n633) );
  assign n2144 = ~n44 & n160 ;
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2147( .i (n2146), .o (n2147) );
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  buffer buf_n2152( .i (n2151), .o (n2152) );
  assign n2159 = ( n633 & n1151 ) | ( n633 & ~n2152 ) | ( n1151 & ~n2152 ) ;
  assign n2160 = ( n1152 & ~n1745 ) | ( n1152 & n2159 ) | ( ~n1745 & n2159 ) ;
  assign n2161 = ~n2029 & n2160 ;
  assign n2162 = ~n28 & n2161 ;
  buffer buf_n2163( .i (n2162), .o (n2163) );
  buffer buf_n2164( .i (n2163), .o (n2164) );
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n2166( .i (n1997), .o (n2166) );
  assign n2167 = ( n803 & n2163 ) | ( n803 & ~n2166 ) | ( n2163 & ~n2166 ) ;
  assign n2168 = n1402 & ~n2167 ;
  assign n2169 = ( n1403 & n2165 ) | ( n1403 & ~n2168 ) | ( n2165 & ~n2168 ) ;
  buffer buf_n2170( .i (n2169), .o (n2170) );
  buffer buf_n2171( .i (n2170), .o (n2171) );
  assign n2172 = ~n192 & n269 ;
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n2175( .i (n2174), .o (n2175) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n2177), .o (n2178) );
  buffer buf_n2179( .i (n2178), .o (n2179) );
  buffer buf_n2180( .i (n2179), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  buffer buf_n2182( .i (n2181), .o (n2182) );
  buffer buf_n2183( .i (n2182), .o (n2183) );
  buffer buf_n2184( .i (n2183), .o (n2184) );
  buffer buf_n2185( .i (n2184), .o (n2185) );
  assign n2186 = n2170 & n2185 ;
  assign n2187 = ( n2143 & n2171 ) | ( n2143 & n2186 ) | ( n2171 & n2186 ) ;
  buffer buf_n2188( .i (n161), .o (n2188) );
  assign n2189 = n190 | n2188 ;
  buffer buf_n2190( .i (n2189), .o (n2190) );
  buffer buf_n2191( .i (n2190), .o (n2191) );
  buffer buf_n2192( .i (n2191), .o (n2192) );
  buffer buf_n2193( .i (n2192), .o (n2193) );
  buffer buf_n2194( .i (n2193), .o (n2194) );
  buffer buf_n2195( .i (n2194), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  buffer buf_n2197( .i (n2196), .o (n2197) );
  buffer buf_n2198( .i (n2197), .o (n2198) );
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n2200( .i (n2199), .o (n2200) );
  buffer buf_n2201( .i (n2200), .o (n2201) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  buffer buf_n2203( .i (n2202), .o (n2203) );
  assign n2205 = ( n195 & n1334 ) | ( n195 & n2004 ) | ( n1334 & n2004 ) ;
  buffer buf_n2206( .i (n1500), .o (n2206) );
  assign n2207 = n1475 & n2206 ;
  buffer buf_n2208( .i (n2207), .o (n2208) );
  assign n2214 = ( ~n2132 & n2205 ) | ( ~n2132 & n2208 ) | ( n2205 & n2208 ) ;
  buffer buf_n2215( .i (n2214), .o (n2215) );
  buffer buf_n2216( .i (n2215), .o (n2216) );
  assign n2217 = ( ~n72 & n188 ) | ( ~n72 & n218 ) | ( n188 & n218 ) ;
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n2221( .i (n2220), .o (n2221) );
  assign n2222 = n74 & n2218 ;
  buffer buf_n2223( .i (n2222), .o (n2223) );
  buffer buf_n2224( .i (n2223), .o (n2224) );
  buffer buf_n2225( .i (n1520), .o (n2225) );
  assign n2226 = ( n192 & ~n2223 ) | ( n192 & n2225 ) | ( ~n2223 & n2225 ) ;
  assign n2227 = ( n2221 & n2224 ) | ( n2221 & ~n2226 ) | ( n2224 & ~n2226 ) ;
  buffer buf_n2228( .i (n1605), .o (n2228) );
  assign n2229 = ( ~n1475 & n2227 ) | ( ~n1475 & n2228 ) | ( n2227 & n2228 ) ;
  buffer buf_n2230( .i (n159), .o (n2230) );
  buffer buf_n2231( .i (n187), .o (n2231) );
  assign n2232 = n2230 & n2231 ;
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2234( .i (n2233), .o (n2234) );
  buffer buf_n2235( .i (n2234), .o (n2235) );
  assign n2252 = n189 & ~n219 ;
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  assign n2264 = ( ~n1939 & n2235 ) | ( ~n1939 & n2254 ) | ( n2235 & n2254 ) ;
  assign n2265 = ( ~n1939 & n2067 ) | ( ~n1939 & n2235 ) | ( n2067 & n2235 ) ;
  assign n2266 = ( n1606 & n2264 ) | ( n1606 & ~n2265 ) | ( n2264 & ~n2265 ) ;
  buffer buf_n2267( .i (n1326), .o (n2267) );
  assign n2268 = ( n2228 & ~n2266 ) | ( n2228 & n2267 ) | ( ~n2266 & n2267 ) ;
  assign n2269 = n2229 & ~n2268 ;
  buffer buf_n2270( .i (n2269), .o (n2270) );
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  assign n2273 = ( n227 & n1827 ) | ( n227 & ~n2270 ) | ( n1827 & ~n2270 ) ;
  assign n2274 = n2215 & n2273 ;
  assign n2275 = ( n2216 & n2272 ) | ( n2216 & ~n2274 ) | ( n2272 & ~n2274 ) ;
  assign n2276 = ( ~n28 & n1347 ) | ( ~n28 & n2275 ) | ( n1347 & n2275 ) ;
  buffer buf_n2277( .i (n218), .o (n2277) );
  assign n2278 = ( n161 & n247 ) | ( n161 & ~n2277 ) | ( n247 & ~n2277 ) ;
  buffer buf_n2279( .i (n2278), .o (n2279) );
  assign n2288 = ( n75 & n1276 ) | ( n75 & n2279 ) | ( n1276 & n2279 ) ;
  buffer buf_n2289( .i (n2288), .o (n2289) );
  buffer buf_n2290( .i (n2289), .o (n2290) );
  buffer buf_n2291( .i (n2290), .o (n2291) );
  buffer buf_n2280( .i (n2279), .o (n2280) );
  buffer buf_n2281( .i (n2280), .o (n2281) );
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2292( .i (n2067), .o (n2292) );
  assign n2293 = ( n1326 & ~n2289 ) | ( n1326 & n2292 ) | ( ~n2289 & n2292 ) ;
  assign n2294 = n2282 & n2293 ;
  assign n2295 = ( n2004 & ~n2291 ) | ( n2004 & n2294 ) | ( ~n2291 & n2294 ) ;
  assign n2296 = n2132 | n2295 ;
  assign n2297 = ~n246 & n2230 ;
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  assign n2308 = ( n449 & ~n2225 ) | ( n449 & n2300 ) | ( ~n2225 & n2300 ) ;
  buffer buf_n2309( .i (n2308), .o (n2309) );
  assign n2324 = n1622 & n2309 ;
  assign n2325 = n2004 & n2324 ;
  assign n2326 = n2132 & ~n2325 ;
  assign n2327 = n2296 & ~n2326 ;
  assign n2328 = n1972 | n2327 ;
  buffer buf_n2329( .i (n189), .o (n2329) );
  buffer buf_n2330( .i (n247), .o (n2330) );
  assign n2331 = ( n2188 & n2329 ) | ( n2188 & ~n2330 ) | ( n2329 & ~n2330 ) ;
  buffer buf_n2332( .i (n2331), .o (n2332) );
  assign n2336 = ( n1939 & ~n2225 ) | ( n1939 & n2332 ) | ( ~n2225 & n2332 ) ;
  buffer buf_n2337( .i (n2336), .o (n2337) );
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  buffer buf_n2333( .i (n2332), .o (n2333) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n2335( .i (n2334), .o (n2335) );
  assign n2340 = ( n2206 & n2267 ) | ( n2206 & n2337 ) | ( n2267 & n2337 ) ;
  assign n2341 = n2335 & ~n2340 ;
  assign n2342 = ( n1743 & ~n2339 ) | ( n1743 & n2341 ) | ( ~n2339 & n2341 ) ;
  buffer buf_n2343( .i (n1624), .o (n2343) );
  assign n2344 = n2342 & n2343 ;
  buffer buf_n2345( .i (n1827), .o (n2345) );
  assign n2346 = ~n2344 & n2345 ;
  assign n2347 = n2328 & ~n2346 ;
  buffer buf_n2348( .i (n111), .o (n2348) );
  assign n2349 = ( n28 & ~n2347 ) | ( n28 & n2348 ) | ( ~n2347 & n2348 ) ;
  assign n2350 = n2276 & ~n2349 ;
  buffer buf_n2351( .i (n2350), .o (n2351) );
  buffer buf_n2352( .i (n2351), .o (n2352) );
  buffer buf_n2353( .i (n2352), .o (n2353) );
  assign n2354 = n685 | n1743 ;
  buffer buf_n2355( .i (n2354), .o (n2355) );
  buffer buf_n2356( .i (n2355), .o (n2356) );
  buffer buf_n2357( .i (n2356), .o (n2357) );
  buffer buf_n2358( .i (n2357), .o (n2358) );
  buffer buf_n2359( .i (n2358), .o (n2359) );
  assign n2360 = n1894 & ~n2359 ;
  assign n2361 = ( n930 & n2351 ) | ( n930 & n2360 ) | ( n2351 & n2360 ) ;
  assign n2362 = n2202 | n2361 ;
  assign n2363 = ( ~n2203 & n2353 ) | ( ~n2203 & n2362 ) | ( n2353 & n2362 ) ;
  buffer buf_n2364( .i (n2107), .o (n2364) );
  assign n2365 = n2363 | n2364 ;
  buffer buf_n2366( .i (n132), .o (n2366) );
  assign n2367 = ( n191 & ~n1520 ) | ( n191 & n2366 ) | ( ~n1520 & n2366 ) ;
  buffer buf_n2368( .i (n2367), .o (n2368) );
  assign n2374 = ( n1500 & ~n2292 ) | ( n1500 & n2368 ) | ( ~n2292 & n2368 ) ;
  buffer buf_n2375( .i (n2374), .o (n2375) );
  buffer buf_n2376( .i (n2375), .o (n2376) );
  buffer buf_n2377( .i (n2376), .o (n2377) );
  buffer buf_n2378( .i (n2377), .o (n2378) );
  buffer buf_n2379( .i (n194), .o (n2379) );
  assign n2380 = ( n1825 & n2375 ) | ( n1825 & n2379 ) | ( n2375 & n2379 ) ;
  buffer buf_n2381( .i (n2380), .o (n2381) );
  buffer buf_n2382( .i (n2381), .o (n2382) );
  buffer buf_n2369( .i (n2368), .o (n2369) );
  buffer buf_n2370( .i (n2369), .o (n2370) );
  buffer buf_n2371( .i (n2370), .o (n2371) );
  buffer buf_n2372( .i (n2371), .o (n2372) );
  assign n2383 = n2372 & ~n2381 ;
  assign n2384 = ( n2378 & ~n2382 ) | ( n2378 & n2383 ) | ( ~n2382 & n2383 ) ;
  buffer buf_n2385( .i (n1842), .o (n2385) );
  assign n2386 = n2384 & n2385 ;
  buffer buf_n2387( .i (n191), .o (n2387) );
  assign n2388 = ( n1664 & n2225 ) | ( n1664 & n2387 ) | ( n2225 & n2387 ) ;
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2391( .i (n2390), .o (n2391) );
  buffer buf_n2392( .i (n2391), .o (n2392) );
  buffer buf_n2393( .i (n2392), .o (n2393) );
  buffer buf_n2236( .i (n2235), .o (n2236) );
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  buffer buf_n2394( .i (n1826), .o (n2394) );
  assign n2395 = ( n2240 & ~n2343 ) | ( n2240 & n2394 ) | ( ~n2343 & n2394 ) ;
  assign n2396 = n2393 & ~n2395 ;
  assign n2397 = n2385 | n2396 ;
  assign n2398 = ( ~n2348 & n2386 ) | ( ~n2348 & n2397 ) | ( n2386 & n2397 ) ;
  assign n2399 = n1684 | n2398 ;
  buffer buf_n2400( .i (n2387), .o (n2400) );
  buffer buf_n2401( .i (n2400), .o (n2401) );
  assign n2402 = ( n1622 & ~n2389 ) | ( n1622 & n2401 ) | ( ~n2389 & n2401 ) ;
  buffer buf_n2403( .i (n2402), .o (n2403) );
  buffer buf_n2404( .i (n2403), .o (n2404) );
  buffer buf_n2405( .i (n2404), .o (n2405) );
  buffer buf_n2406( .i (n2405), .o (n2406) );
  buffer buf_n2407( .i (n1207), .o (n2407) );
  assign n2408 = ( n1826 & ~n2403 ) | ( n1826 & n2407 ) | ( ~n2403 & n2407 ) ;
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  assign n2411 = ~n2393 & n2409 ;
  assign n2412 = ( n2406 & n2410 ) | ( n2406 & n2411 ) | ( n2410 & n2411 ) ;
  assign n2413 = ~n2348 & n2412 ;
  buffer buf_n2414( .i (n1816), .o (n2414) );
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n2416( .i (n2415), .o (n2416) );
  buffer buf_n2417( .i (n2416), .o (n2417) );
  assign n2418 = ~n2413 & n2417 ;
  assign n2419 = n2399 & ~n2418 ;
  assign n2420 = n1059 & n1746 ;
  buffer buf_n2421( .i (n2420), .o (n2421) );
  assign n2426 = n287 & ~n2355 ;
  buffer buf_n2427( .i (n2426), .o (n2427) );
  buffer buf_n2428( .i (n2427), .o (n2428) );
  assign n2429 = n1306 | n2427 ;
  assign n2430 = ( n2421 & n2428 ) | ( n2421 & n2429 ) | ( n2428 & n2429 ) ;
  buffer buf_n2431( .i (n2430), .o (n2431) );
  assign n2432 = ( n87 & n2419 ) | ( n87 & n2431 ) | ( n2419 & n2431 ) ;
  buffer buf_n2433( .i (n2366), .o (n2433) );
  assign n2434 = ( ~n104 & n2387 ) | ( ~n104 & n2433 ) | ( n2387 & n2433 ) ;
  buffer buf_n2435( .i (n2434), .o (n2435) );
  buffer buf_n2440( .i (n2292), .o (n2440) );
  assign n2441 = ( n2228 & ~n2435 ) | ( n2228 & n2440 ) | ( ~n2435 & n2440 ) ;
  buffer buf_n2442( .i (n2441), .o (n2442) );
  buffer buf_n2443( .i (n2442), .o (n2443) );
  buffer buf_n2444( .i (n2443), .o (n2444) );
  buffer buf_n2445( .i (n2444), .o (n2445) );
  buffer buf_n2446( .i (n2379), .o (n2446) );
  assign n2447 = ( n108 & n2442 ) | ( n108 & ~n2446 ) | ( n2442 & ~n2446 ) ;
  buffer buf_n2448( .i (n2447), .o (n2448) );
  buffer buf_n2449( .i (n2448), .o (n2449) );
  buffer buf_n2436( .i (n2435), .o (n2436) );
  buffer buf_n2437( .i (n2436), .o (n2437) );
  buffer buf_n2438( .i (n2437), .o (n2438) );
  buffer buf_n2439( .i (n2438), .o (n2439) );
  assign n2450 = n2439 & n2448 ;
  assign n2451 = ( ~n2445 & n2449 ) | ( ~n2445 & n2450 ) | ( n2449 & n2450 ) ;
  assign n2452 = n2416 | n2451 ;
  assign n2453 = ( n563 & n1985 ) | ( n563 & n2343 ) | ( n1985 & n2343 ) ;
  assign n2454 = ( n563 & ~n1985 ) | ( n563 & n2343 ) | ( ~n1985 & n2343 ) ;
  assign n2455 = ( n1842 & ~n2453 ) | ( n1842 & n2454 ) | ( ~n2453 & n2454 ) ;
  assign n2456 = n199 & n2455 ;
  assign n2457 = n2416 & ~n2456 ;
  assign n2458 = n2452 & ~n2457 ;
  assign n2459 = n1528 & ~n2206 ;
  buffer buf_n2460( .i (n2459), .o (n2460) );
  buffer buf_n2461( .i (n2460), .o (n2461) );
  buffer buf_n2462( .i (n2461), .o (n2462) );
  assign n2468 = ( n2177 & n2345 ) | ( n2177 & n2462 ) | ( n2345 & n2462 ) ;
  assign n2469 = ~n2029 & n2468 ;
  buffer buf_n2470( .i (n2469), .o (n2470) );
  buffer buf_n2471( .i (n2470), .o (n2471) );
  assign n2472 = n1654 | n2470 ;
  assign n2473 = ( n2458 & n2471 ) | ( n2458 & n2472 ) | ( n2471 & n2472 ) ;
  buffer buf_n2474( .i (n2082), .o (n2474) );
  assign n2475 = ( n2431 & n2473 ) | ( n2431 & ~n2474 ) | ( n2473 & ~n2474 ) ;
  assign n2476 = n2432 | n2475 ;
  assign n2477 = ~n2109 & n2476 ;
  assign n2478 = n2364 & ~n2477 ;
  assign n2479 = n2365 & ~n2478 ;
  assign n2480 = n2187 | n2479 ;
  assign n2481 = ( ~n2113 & n2131 ) | ( ~n2113 & n2480 ) | ( n2131 & n2480 ) ;
  assign n2482 = n2114 | n2481 ;
  assign n2483 = ( n200 & n1517 ) | ( n200 & ~n2416 ) | ( n1517 & ~n2416 ) ;
  buffer buf_n2484( .i (n2483), .o (n2484) );
  assign n2485 = ( n1702 & ~n2082 ) | ( n1702 & n2484 ) | ( ~n2082 & n2484 ) ;
  assign n2486 = ( n260 & ~n1702 ) | ( n260 & n2484 ) | ( ~n1702 & n2484 ) ;
  assign n2487 = n2485 & n2486 ;
  buffer buf_n2488( .i (n2487), .o (n2488) );
  buffer buf_n2489( .i (n2488), .o (n2489) );
  buffer buf_n2490( .i (n1325), .o (n2490) );
  assign n2491 = n1605 & ~n2490 ;
  buffer buf_n2492( .i (n2491), .o (n2492) );
  buffer buf_n2500( .i (n1941), .o (n2500) );
  assign n2501 = ( n23 & n2492 ) | ( n23 & n2500 ) | ( n2492 & n2500 ) ;
  buffer buf_n2502( .i (n2501), .o (n2502) );
  buffer buf_n2503( .i (n2502), .o (n2503) );
  buffer buf_n2504( .i (n2503), .o (n2504) );
  buffer buf_n2505( .i (n2500), .o (n2505) );
  buffer buf_n2506( .i (n2505), .o (n2506) );
  assign n2507 = ( n2394 & ~n2502 ) | ( n2394 & n2506 ) | ( ~n2502 & n2506 ) ;
  buffer buf_n2508( .i (n25), .o (n2508) );
  assign n2509 = ( ~n2414 & n2507 ) | ( ~n2414 & n2508 ) | ( n2507 & n2508 ) ;
  assign n2510 = ~n2504 & n2509 ;
  buffer buf_n2511( .i (n2510), .o (n2511) );
  buffer buf_n2512( .i (n2511), .o (n2512) );
  buffer buf_n2513( .i (n1890), .o (n2513) );
  assign n2514 = ( n201 & n2511 ) | ( n201 & ~n2513 ) | ( n2511 & ~n2513 ) ;
  assign n2515 = ~n2206 & n2267 ;
  buffer buf_n2516( .i (n2515), .o (n2516) );
  buffer buf_n2517( .i (n2516), .o (n2517) );
  buffer buf_n2518( .i (n2517), .o (n2518) );
  assign n2523 = n2345 & n2518 ;
  buffer buf_n2524( .i (n2508), .o (n2524) );
  assign n2525 = ( n1746 & n2523 ) | ( n1746 & n2524 ) | ( n2523 & n2524 ) ;
  buffer buf_n2526( .i (n2524), .o (n2526) );
  assign n2527 = n2525 & ~n2526 ;
  assign n2528 = ~n201 & n2527 ;
  assign n2529 = ( n2512 & ~n2514 ) | ( n2512 & n2528 ) | ( ~n2514 & n2528 ) ;
  buffer buf_n2530( .i (n2529), .o (n2530) );
  buffer buf_n2531( .i (n2530), .o (n2531) );
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n409), .o (n2533) );
  buffer buf_n2534( .i (n174), .o (n2534) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  assign n2536 = ( ~n2530 & n2533 ) | ( ~n2530 & n2535 ) | ( n2533 & n2535 ) ;
  assign n2537 = n2488 & n2536 ;
  assign n2538 = ( n2489 & n2532 ) | ( n2489 & ~n2537 ) | ( n2532 & ~n2537 ) ;
  assign n2539 = n119 | n2538 ;
  buffer buf_n2540( .i (n1520), .o (n2540) );
  buffer buf_n2541( .i (n2540), .o (n2541) );
  assign n2542 = ( ~n1940 & n2400 ) | ( ~n1940 & n2541 ) | ( n2400 & n2541 ) ;
  buffer buf_n2543( .i (n2542), .o (n2543) );
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2552( .i (n1745), .o (n2552) );
  assign n2553 = ( n2029 & n2547 ) | ( n2029 & n2552 ) | ( n2547 & n2552 ) ;
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2555( .i (n2554), .o (n2555) );
  buffer buf_n2556( .i (n2555), .o (n2556) );
  buffer buf_n2557( .i (n2556), .o (n2557) );
  buffer buf_n2558( .i (n199), .o (n2558) );
  buffer buf_n2559( .i (n2558), .o (n2559) );
  assign n2560 = ( n2513 & n2554 ) | ( n2513 & n2559 ) | ( n2554 & n2559 ) ;
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  buffer buf_n2550( .i (n2549), .o (n2550) );
  buffer buf_n2551( .i (n2550), .o (n2551) );
  assign n2563 = n2551 & ~n2561 ;
  assign n2564 = ( n2557 & ~n2562 ) | ( n2557 & n2563 ) | ( ~n2562 & n2563 ) ;
  assign n2565 = ~n263 & n2564 ;
  assign n2566 = ~n2110 & n2565 ;
  assign n2567 = n119 & ~n2566 ;
  assign n2568 = n2539 & ~n2567 ;
  assign n2569 = n65 | n2568 ;
  buffer buf_n178( .i (n177), .o (n178) );
  assign n2570 = n1745 & ~n2414 ;
  buffer buf_n2571( .i (n2570), .o (n2571) );
  buffer buf_n2574( .i (n2552), .o (n2574) );
  assign n2575 = ~n2571 & n2574 ;
  buffer buf_n2576( .i (n2575), .o (n2576) );
  buffer buf_n2577( .i (n1701), .o (n2577) );
  assign n2578 = n2576 & n2577 ;
  buffer buf_n2572( .i (n2571), .o (n2572) );
  buffer buf_n2573( .i (n2572), .o (n2573) );
  assign n2579 = ( n202 & ~n2573 ) | ( n202 & n2576 ) | ( ~n2573 & n2576 ) ;
  assign n2580 = ( ~n261 & n2578 ) | ( ~n261 & n2579 ) | ( n2578 & n2579 ) ;
  assign n2581 = n1650 & n2580 ;
  buffer buf_n2582( .i (n131), .o (n2582) );
  assign n2583 = ( n74 & n2330 ) | ( n74 & n2582 ) | ( n2330 & n2582 ) ;
  buffer buf_n2584( .i (n2583), .o (n2584) );
  buffer buf_n2585( .i (n2584), .o (n2585) );
  buffer buf_n2586( .i (n2585), .o (n2586) );
  buffer buf_n2587( .i (n2586), .o (n2587) );
  buffer buf_n2588( .i (n2587), .o (n2588) );
  buffer buf_n2589( .i (n2588), .o (n2589) );
  buffer buf_n2590( .i (n2589), .o (n2590) );
  assign n2591 = ( ~n198 & n2345 ) | ( ~n198 & n2590 ) | ( n2345 & n2590 ) ;
  buffer buf_n2592( .i (n2591), .o (n2592) );
  buffer buf_n2595( .i (n2394), .o (n2595) );
  buffer buf_n2596( .i (n2595), .o (n2596) );
  buffer buf_n2597( .i (n2596), .o (n2597) );
  assign n2598 = ~n2592 & n2597 ;
  buffer buf_n2599( .i (n2598), .o (n2599) );
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2593( .i (n2592), .o (n2593) );
  buffer buf_n2594( .i (n2593), .o (n2594) );
  assign n2601 = n2594 | n2599 ;
  assign n2602 = ( ~n2016 & n2600 ) | ( ~n2016 & n2601 ) | ( n2600 & n2601 ) ;
  assign n2603 = n1650 | n2602 ;
  assign n2604 = ( ~n1024 & n2581 ) | ( ~n1024 & n2603 ) | ( n2581 & n2603 ) ;
  assign n2605 = n178 | n2604 ;
  buffer buf_n2422( .i (n2421), .o (n2422) );
  buffer buf_n2423( .i (n2422), .o (n2423) );
  buffer buf_n2424( .i (n2423), .o (n2424) );
  buffer buf_n2425( .i (n2424), .o (n2425) );
  assign n2606 = ~n2267 & n2401 ;
  buffer buf_n2607( .i (n2606), .o (n2607) );
  buffer buf_n2608( .i (n2607), .o (n2608) );
  buffer buf_n2609( .i (n2608), .o (n2609) );
  buffer buf_n2610( .i (n2609), .o (n2610) );
  buffer buf_n2611( .i (n2610), .o (n2611) );
  buffer buf_n2612( .i (n2611), .o (n2612) );
  buffer buf_n2613( .i (n2612), .o (n2613) );
  buffer buf_n2614( .i (n2613), .o (n2614) );
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2616( .i (n2615), .o (n2616) );
  assign n2617 = n2425 & n2616 ;
  assign n2618 = n178 & ~n2617 ;
  assign n2619 = n2605 & ~n2618 ;
  buffer buf_n2620( .i (n1786), .o (n2620) );
  assign n2621 = n2619 & ~n2620 ;
  assign n2622 = n65 & ~n2621 ;
  assign n2623 = n2569 & ~n2622 ;
  assign n2624 = n2482 | n2623 ;
  assign n2625 = ( n2026 & ~n2027 ) | ( n2026 & n2624 ) | ( ~n2027 & n2624 ) ;
  assign n2626 = n2292 & n2541 ;
  buffer buf_n2627( .i (n2626), .o (n2627) );
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  buffer buf_n2631( .i (n2630), .o (n2631) );
  buffer buf_n2632( .i (n2631), .o (n2632) );
  buffer buf_n2633( .i (n2632), .o (n2633) );
  buffer buf_n2634( .i (n2633), .o (n2634) );
  buffer buf_n2635( .i (n2634), .o (n2635) );
  buffer buf_n2636( .i (n2635), .o (n2636) );
  buffer buf_n2637( .i (n2636), .o (n2637) );
  assign n2638 = ( ~n177 & n403 ) | ( ~n177 & n2637 ) | ( n403 & n2637 ) ;
  assign n2639 = ~n2364 & n2638 ;
  buffer buf_n2640( .i (n90), .o (n2640) );
  assign n2641 = n2639 & ~n2640 ;
  assign n2642 = n2620 & n2641 ;
  buffer buf_n2643( .i (n54), .o (n2643) );
  buffer buf_n2644( .i (n1617), .o (n2644) );
  assign n2645 = ( n2552 & ~n2643 ) | ( n2552 & n2644 ) | ( ~n2643 & n2644 ) ;
  buffer buf_n2646( .i (n2645), .o (n2646) );
  buffer buf_n2647( .i (n2646), .o (n2647) );
  buffer buf_n2648( .i (n2647), .o (n2648) );
  buffer buf_n2649( .i (n2648), .o (n2649) );
  buffer buf_n2650( .i (n2574), .o (n2650) );
  assign n2651 = n2646 & ~n2650 ;
  buffer buf_n2652( .i (n2651), .o (n2652) );
  buffer buf_n2653( .i (n2652), .o (n2653) );
  assign n2654 = ( n2084 & ~n2534 ) | ( n2084 & n2652 ) | ( ~n2534 & n2652 ) ;
  assign n2655 = ( n2649 & n2653 ) | ( n2649 & n2654 ) | ( n2653 & n2654 ) ;
  assign n2656 = ( n147 & ~n1024 ) | ( n147 & n2655 ) | ( ~n1024 & n2655 ) ;
  assign n2657 = ( n1889 & ~n2552 ) | ( n1889 & n2643 ) | ( ~n2552 & n2643 ) ;
  buffer buf_n2658( .i (n2657), .o (n2658) );
  buffer buf_n2659( .i (n2658), .o (n2659) );
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2660), .o (n2661) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  assign n2662 = n478 & ~n2658 ;
  buffer buf_n2663( .i (n2662), .o (n2663) );
  buffer buf_n2664( .i (n2663), .o (n2664) );
  assign n2665 = n233 & ~n2663 ;
  assign n2666 = ( n2661 & n2664 ) | ( n2661 & ~n2665 ) | ( n2664 & ~n2665 ) ;
  assign n2667 = ( n147 & n1024 ) | ( n147 & n2666 ) | ( n1024 & n2666 ) ;
  assign n2668 = n2656 & ~n2667 ;
  assign n2669 = ( ~n796 & n870 ) | ( ~n796 & n1183 ) | ( n870 & n1183 ) ;
  buffer buf_n2670( .i (n2669), .o (n2670) );
  buffer buf_n2671( .i (n2670), .o (n2671) );
  buffer buf_n2672( .i (n2671), .o (n2672) );
  buffer buf_n2673( .i (n2672), .o (n2673) );
  buffer buf_n2674( .i (n2673), .o (n2674) );
  buffer buf_n2675( .i (n2674), .o (n2675) );
  buffer buf_n2676( .i (n2675), .o (n2676) );
  buffer buf_n2685( .i (n2166), .o (n2685) );
  assign n2686 = ( n2474 & ~n2676 ) | ( n2474 & n2685 ) | ( ~n2676 & n2685 ) ;
  buffer buf_n2687( .i (n2686), .o (n2687) );
  buffer buf_n2688( .i (n2685), .o (n2688) );
  buffer buf_n2689( .i (n2688), .o (n2689) );
  assign n2690 = ( n2107 & n2687 ) | ( n2107 & ~n2689 ) | ( n2687 & ~n2689 ) ;
  assign n2691 = ( n89 & n2107 ) | ( n89 & ~n2687 ) | ( n2107 & ~n2687 ) ;
  assign n2692 = n2690 & ~n2691 ;
  assign n2693 = n2668 | n2692 ;
  assign n2694 = ~n2620 & n2693 ;
  assign n2695 = n2642 | n2694 ;
  buffer buf_n2696( .i (n2695), .o (n2696) );
  buffer buf_n2697( .i (n2696), .o (n2697) );
  assign n2698 = ( n1755 & ~n2446 ) | ( n1755 & n2607 ) | ( ~n2446 & n2607 ) ;
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n2700( .i (n2699), .o (n2700) );
  buffer buf_n2701( .i (n2700), .o (n2701) );
  buffer buf_n2702( .i (n2701), .o (n2702) );
  buffer buf_n2703( .i (n2702), .o (n2703) );
  buffer buf_n2704( .i (n2703), .o (n2704) );
  buffer buf_n2705( .i (n2704), .o (n2705) );
  buffer buf_n2706( .i (n2705), .o (n2706) );
  buffer buf_n2707( .i (n2706), .o (n2707) );
  buffer buf_n2708( .i (n2707), .o (n2708) );
  buffer buf_n2709( .i (n2708), .o (n2709) );
  buffer buf_n2710( .i (n2709), .o (n2710) );
  buffer buf_n2711( .i (n2710), .o (n2711) );
  buffer buf_n2712( .i (n2711), .o (n2712) );
  assign n2714 = n2696 & n2712 ;
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n2715( .i (n2541), .o (n2715) );
  buffer buf_n2716( .i (n2715), .o (n2716) );
  assign n2717 = n1825 | n2716 ;
  buffer buf_n2718( .i (n2717), .o (n2718) );
  buffer buf_n2719( .i (n2718), .o (n2719) );
  buffer buf_n2720( .i (n2719), .o (n2720) );
  buffer buf_n2721( .i (n2720), .o (n2721) );
  buffer buf_n2722( .i (n2721), .o (n2722) );
  assign n2727 = ( n1997 & n2650 ) | ( n1997 & n2722 ) | ( n2650 & n2722 ) ;
  assign n2728 = ( n1985 & n2506 ) | ( n1985 & ~n2718 ) | ( n2506 & ~n2718 ) ;
  buffer buf_n2729( .i (n2728), .o (n2729) );
  buffer buf_n2730( .i (n2729), .o (n2730) );
  buffer buf_n2731( .i (n2730), .o (n2731) );
  assign n2732 = ( n1701 & n2513 ) | ( n1701 & n2731 ) | ( n2513 & n2731 ) ;
  assign n2733 = n2727 & ~n2732 ;
  assign n2734 = n2084 & n2733 ;
  buffer buf_n2735( .i (n1888), .o (n2735) );
  buffer buf_n2736( .i (n2735), .o (n2736) );
  assign n2737 = n2574 | n2736 ;
  buffer buf_n2738( .i (n2737), .o (n2738) );
  assign n2739 = ( n568 & n2082 ) | ( n568 & ~n2738 ) | ( n2082 & ~n2738 ) ;
  buffer buf_n2740( .i (n1376), .o (n2740) );
  buffer buf_n2741( .i (n2740), .o (n2741) );
  assign n2742 = n2739 | n2741 ;
  assign n2743 = ( ~n2106 & n2734 ) | ( ~n2106 & n2742 ) | ( n2734 & n2742 ) ;
  assign n2744 = ( n235 & ~n2109 ) | ( n235 & n2743 ) | ( ~n2109 & n2743 ) ;
  buffer buf_n2745( .i (n2506), .o (n2745) );
  buffer buf_n2746( .i (n2745), .o (n2746) );
  assign n2747 = n443 | n2746 ;
  buffer buf_n2748( .i (n2747), .o (n2748) );
  buffer buf_n2749( .i (n2748), .o (n2749) );
  assign n2750 = ( n444 & n2574 ) | ( n444 & ~n2597 ) | ( n2574 & ~n2597 ) ;
  assign n2751 = n2748 & ~n2750 ;
  buffer buf_n2752( .i (n2650), .o (n2752) );
  assign n2753 = ( n2749 & n2751 ) | ( n2749 & ~n2752 ) | ( n2751 & ~n2752 ) ;
  assign n2754 = n2741 | n2753 ;
  assign n2755 = n810 & n2752 ;
  assign n2756 = n2741 & ~n2755 ;
  assign n2757 = n2754 & ~n2756 ;
  buffer buf_n2758( .i (n234), .o (n2758) );
  assign n2759 = ( n2109 & ~n2757 ) | ( n2109 & n2758 ) | ( ~n2757 & n2758 ) ;
  assign n2760 = n2744 & ~n2759 ;
  buffer buf_n2761( .i (n1275), .o (n2761) );
  buffer buf_n2762( .i (n2761), .o (n2762) );
  assign n2763 = ~n2433 & n2762 ;
  buffer buf_n2764( .i (n2763), .o (n2764) );
  buffer buf_n2765( .i (n2764), .o (n2765) );
  buffer buf_n2766( .i (n2765), .o (n2766) );
  buffer buf_n2767( .i (n2766), .o (n2767) );
  buffer buf_n2768( .i (n2767), .o (n2768) );
  buffer buf_n2769( .i (n2768), .o (n2769) );
  buffer buf_n2770( .i (n2769), .o (n2770) );
  buffer buf_n2771( .i (n2770), .o (n2771) );
  buffer buf_n2772( .i (n2771), .o (n2772) );
  buffer buf_n2773( .i (n2772), .o (n2773) );
  buffer buf_n2774( .i (n2773), .o (n2774) );
  buffer buf_n2775( .i (n2774), .o (n2775) );
  buffer buf_n2776( .i (n2775), .o (n2776) );
  assign n2777 = n1888 & n2745 ;
  buffer buf_n2778( .i (n2777), .o (n2778) );
  buffer buf_n2779( .i (n2778), .o (n2779) );
  assign n2780 = ( ~n730 & n1997 ) | ( ~n730 & n2779 ) | ( n1997 & n2779 ) ;
  assign n2781 = n731 & n2780 ;
  buffer buf_n2782( .i (n107), .o (n2782) );
  buffer buf_n2783( .i (n2782), .o (n2783) );
  assign n2784 = n702 & ~n2783 ;
  buffer buf_n2785( .i (n2784), .o (n2785) );
  buffer buf_n2786( .i (n2785), .o (n2786) );
  buffer buf_n2787( .i (n2786), .o (n2787) );
  assign n2788 = ( ~n2513 & n2650 ) | ( ~n2513 & n2787 ) | ( n2650 & n2787 ) ;
  assign n2789 = ~n2752 & n2788 ;
  assign n2790 = n2781 | n2789 ;
  buffer buf_n2791( .i (n2790), .o (n2791) );
  buffer buf_n2792( .i (n2791), .o (n2792) );
  buffer buf_n2793( .i (n1551), .o (n2793) );
  assign n2794 = ( n2758 & n2791 ) | ( n2758 & ~n2793 ) | ( n2791 & ~n2793 ) ;
  assign n2795 = ( n2776 & n2792 ) | ( n2776 & ~n2794 ) | ( n2792 & ~n2794 ) ;
  assign n2796 = n2760 | n2795 ;
  buffer buf_n2797( .i (n2796), .o (n2797) );
  buffer buf_n2798( .i (n2797), .o (n2798) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  assign n2799 = ( ~n209 & n267 ) | ( ~n209 & n2797 ) | ( n267 & n2797 ) ;
  assign n2800 = ( n506 & n2798 ) | ( n506 & ~n2799 ) | ( n2798 & ~n2799 ) ;
  assign n2801 = ( n1528 & n1941 ) | ( n1528 & n2440 ) | ( n1941 & n2440 ) ;
  buffer buf_n2802( .i (n2801), .o (n2802) );
  assign n2808 = ( n1624 & ~n2407 ) | ( n1624 & n2802 ) | ( ~n2407 & n2802 ) ;
  buffer buf_n2809( .i (n2808), .o (n2809) );
  assign n2813 = n1617 & ~n2809 ;
  buffer buf_n2814( .i (n2813), .o (n2814) );
  buffer buf_n2815( .i (n2814), .o (n2815) );
  buffer buf_n2810( .i (n2809), .o (n2810) );
  buffer buf_n2811( .i (n2810), .o (n2811) );
  assign n2816 = n2811 | n2814 ;
  assign n2817 = ( ~n1909 & n2815 ) | ( ~n1909 & n2816 ) | ( n2815 & n2816 ) ;
  buffer buf_n2818( .i (n2817), .o (n2818) );
  buffer buf_n2819( .i (n2818), .o (n2819) );
  assign n2820 = ( n203 & n2741 ) | ( n203 & ~n2818 ) | ( n2741 & ~n2818 ) ;
  buffer buf_n2821( .i (n2348), .o (n2821) );
  assign n2822 = n541 & n2821 ;
  assign n2823 = ~n1509 & n2822 ;
  buffer buf_n2824( .i (n202), .o (n2824) );
  assign n2825 = n2823 & n2824 ;
  assign n2826 = ( n2819 & n2820 ) | ( n2819 & n2825 ) | ( n2820 & n2825 ) ;
  buffer buf_n2827( .i (n2826), .o (n2827) );
  buffer buf_n2828( .i (n2827), .o (n2828) );
  assign n2829 = n2201 | n2685 ;
  assign n2830 = ( n88 & n2106 ) | ( n88 & ~n2829 ) | ( n2106 & ~n2829 ) ;
  buffer buf_n2831( .i (n2106), .o (n2831) );
  assign n2832 = n2830 & ~n2831 ;
  assign n2833 = ~n2092 & n2407 ;
  buffer buf_n2834( .i (n2833), .o (n2834) );
  buffer buf_n2835( .i (n2834), .o (n2835) );
  buffer buf_n2836( .i (n2835), .o (n2836) );
  assign n2839 = ~n73 & n161 ;
  buffer buf_n2840( .i (n2839), .o (n2840) );
  assign n2849 = ( ~n858 & n2366 ) | ( ~n858 & n2840 ) | ( n2366 & n2840 ) ;
  buffer buf_n2850( .i (n2849), .o (n2850) );
  buffer buf_n2851( .i (n2850), .o (n2851) );
  buffer buf_n2852( .i (n2851), .o (n2852) );
  buffer buf_n2853( .i (n858), .o (n2853) );
  buffer buf_n2854( .i (n2853), .o (n2854) );
  assign n2855 = ( n1940 & n2850 ) | ( n1940 & n2854 ) | ( n2850 & n2854 ) ;
  assign n2856 = ( n2228 & n2715 ) | ( n2228 & ~n2855 ) | ( n2715 & ~n2855 ) ;
  assign n2857 = ~n2852 & n2856 ;
  assign n2858 = n1145 & n2366 ;
  buffer buf_n2859( .i (n2858), .o (n2859) );
  assign n2866 = n998 & n2859 ;
  buffer buf_n2867( .i (n2866), .o (n2867) );
  buffer buf_n2868( .i (n2867), .o (n2868) );
  assign n2869 = n1623 & ~n2867 ;
  assign n2870 = ( n2857 & n2868 ) | ( n2857 & ~n2869 ) | ( n2868 & ~n2869 ) ;
  assign n2871 = n197 & n2870 ;
  buffer buf_n2872( .i (n2871), .o (n2872) );
  buffer buf_n2873( .i (n2872), .o (n2873) );
  assign n2874 = n1252 | n2872 ;
  assign n2875 = ( n2836 & n2873 ) | ( n2836 & n2874 ) | ( n2873 & n2874 ) ;
  assign n2876 = n2417 & n2875 ;
  assign n2877 = n2230 & ~n2231 ;
  buffer buf_n2878( .i (n2877), .o (n2878) );
  assign n2887 = ( ~n363 & n1796 ) | ( ~n363 & n2878 ) | ( n1796 & n2878 ) ;
  buffer buf_n2888( .i (n73), .o (n2888) );
  buffer buf_n2889( .i (n2888), .o (n2889) );
  assign n2890 = ( n2761 & n2887 ) | ( n2761 & ~n2889 ) | ( n2887 & ~n2889 ) ;
  buffer buf_n2891( .i (n2890), .o (n2891) );
  buffer buf_n2892( .i (n2891), .o (n2892) );
  buffer buf_n2893( .i (n2892), .o (n2893) );
  buffer buf_n2894( .i (n2893), .o (n2894) );
  buffer buf_n2895( .i (n2762), .o (n2895) );
  assign n2896 = n2891 & ~n2895 ;
  buffer buf_n2897( .i (n2896), .o (n2897) );
  buffer buf_n2898( .i (n2897), .o (n2898) );
  buffer buf_n2899( .i (n2854), .o (n2899) );
  buffer buf_n2900( .i (n2899), .o (n2900) );
  assign n2901 = ( n2500 & n2897 ) | ( n2500 & n2900 ) | ( n2897 & n2900 ) ;
  assign n2902 = ( n2894 & n2898 ) | ( n2894 & n2901 ) | ( n2898 & n2901 ) ;
  buffer buf_n2903( .i (n2902), .o (n2903) );
  buffer buf_n2904( .i (n2903), .o (n2904) );
  buffer buf_n2905( .i (n2904), .o (n2905) );
  assign n2906 = ( n391 & n1940 ) | ( n391 & ~n2541 ) | ( n1940 & ~n2541 ) ;
  buffer buf_n2907( .i (n2906), .o (n2907) );
  buffer buf_n2908( .i (n2907), .o (n2908) );
  buffer buf_n2909( .i (n2908), .o (n2909) );
  buffer buf_n2910( .i (n102), .o (n2910) );
  buffer buf_n2911( .i (n2188), .o (n2911) );
  assign n2912 = ( n2889 & n2910 ) | ( n2889 & ~n2911 ) | ( n2910 & ~n2911 ) ;
  buffer buf_n2913( .i (n2912), .o (n2913) );
  buffer buf_n2914( .i (n2913), .o (n2914) );
  buffer buf_n2915( .i (n2914), .o (n2915) );
  buffer buf_n2916( .i (n2915), .o (n2916) );
  buffer buf_n2917( .i (n2433), .o (n2917) );
  buffer buf_n2918( .i (n2917), .o (n2918) );
  buffer buf_n2919( .i (n2918), .o (n2919) );
  assign n2920 = ( ~n2900 & n2907 ) | ( ~n2900 & n2919 ) | ( n2907 & n2919 ) ;
  assign n2921 = ( n394 & n2916 ) | ( n394 & ~n2920 ) | ( n2916 & ~n2920 ) ;
  assign n2922 = n2909 & ~n2921 ;
  assign n2923 = ( ~n198 & n2903 ) | ( ~n198 & n2922 ) | ( n2903 & n2922 ) ;
  assign n2924 = n2644 | n2923 ;
  assign n2925 = ( ~n1908 & n2905 ) | ( ~n1908 & n2924 ) | ( n2905 & n2924 ) ;
  assign n2926 = n2417 | n2925 ;
  buffer buf_n2927( .i (n2417), .o (n2927) );
  assign n2928 = ( n2876 & n2926 ) | ( n2876 & ~n2927 ) | ( n2926 & ~n2927 ) ;
  buffer buf_n2929( .i (n2740), .o (n2929) );
  assign n2930 = n2928 & n2929 ;
  assign n2931 = ~n2500 & n2900 ;
  buffer buf_n2932( .i (n2931), .o (n2932) );
  buffer buf_n2841( .i (n2840), .o (n2841) );
  buffer buf_n2842( .i (n2841), .o (n2842) );
  buffer buf_n2843( .i (n2842), .o (n2843) );
  buffer buf_n2844( .i (n2843), .o (n2844) );
  buffer buf_n2845( .i (n2844), .o (n2845) );
  assign n2939 = ( n1624 & n2505 ) | ( n1624 & n2845 ) | ( n2505 & n2845 ) ;
  buffer buf_n2940( .i (n1623), .o (n2940) );
  assign n2941 = ( n2782 & n2845 ) | ( n2782 & n2940 ) | ( n2845 & n2940 ) ;
  assign n2942 = ( n2932 & n2939 ) | ( n2932 & ~n2941 ) | ( n2939 & ~n2941 ) ;
  assign n2943 = ~n583 & n2052 ;
  buffer buf_n2944( .i (n2943), .o (n2944) );
  buffer buf_n2945( .i (n2944), .o (n2945) );
  assign n2946 = n197 | n2944 ;
  assign n2947 = ( n2942 & n2945 ) | ( n2942 & n2946 ) | ( n2945 & n2946 ) ;
  buffer buf_n2948( .i (n2947), .o (n2948) );
  buffer buf_n2949( .i (n2948), .o (n2949) );
  buffer buf_n2950( .i (n2415), .o (n2950) );
  assign n2951 = ( n2597 & n2948 ) | ( n2597 & ~n2950 ) | ( n2948 & ~n2950 ) ;
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  assign n2952 = ~n551 & n2745 ;
  assign n2953 = n443 & n2952 ;
  assign n2954 = ~n2597 & n2953 ;
  assign n2955 = ( n2949 & ~n2951 ) | ( n2949 & n2954 ) | ( ~n2951 & n2954 ) ;
  assign n2956 = ( ~n2280 & n2387 ) | ( ~n2280 & n2540 ) | ( n2387 & n2540 ) ;
  buffer buf_n2957( .i (n2956), .o (n2957) );
  buffer buf_n2958( .i (n2957), .o (n2958) );
  buffer buf_n2959( .i (n2958), .o (n2959) );
  buffer buf_n2960( .i (n2959), .o (n2960) );
  buffer buf_n2961( .i (n2490), .o (n2961) );
  assign n2962 = ( n2440 & n2957 ) | ( n2440 & ~n2961 ) | ( n2957 & ~n2961 ) ;
  buffer buf_n2963( .i (n2962), .o (n2963) );
  buffer buf_n2964( .i (n2963), .o (n2964) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  assign n2965 = n2284 & n2963 ;
  assign n2966 = ( ~n2960 & n2964 ) | ( ~n2960 & n2965 ) | ( n2964 & n2965 ) ;
  assign n2967 = n2745 & n2966 ;
  assign n2968 = ( n1334 & n1623 ) | ( n1334 & ~n2379 ) | ( n1623 & ~n2379 ) ;
  assign n2969 = ( n2407 & n2446 ) | ( n2407 & ~n2968 ) | ( n2446 & ~n2968 ) ;
  buffer buf_n2970( .i (n2446), .o (n2970) );
  assign n2971 = ( n2517 & n2969 ) | ( n2517 & ~n2970 ) | ( n2969 & ~n2970 ) ;
  buffer buf_n2972( .i (n2506), .o (n2972) );
  assign n2973 = n2971 | n2972 ;
  assign n2974 = ( ~n2746 & n2967 ) | ( ~n2746 & n2973 ) | ( n2967 & n2973 ) ;
  buffer buf_n2975( .i (n2385), .o (n2975) );
  buffer buf_n2976( .i (n2596), .o (n2976) );
  assign n2977 = ( n2974 & ~n2975 ) | ( n2974 & n2976 ) | ( ~n2975 & n2976 ) ;
  assign n2978 = ( n2401 & ~n2440 ) | ( n2401 & n2961 ) | ( ~n2440 & n2961 ) ;
  buffer buf_n2979( .i (n2978), .o (n2979) );
  assign n2980 = ( ~n1815 & n2505 ) | ( ~n1815 & n2979 ) | ( n2505 & n2979 ) ;
  buffer buf_n2981( .i (n2379), .o (n2981) );
  assign n2982 = ( n2505 & ~n2979 ) | ( n2505 & n2981 ) | ( ~n2979 & n2981 ) ;
  assign n2983 = n2980 & ~n2982 ;
  buffer buf_n2984( .i (n1887), .o (n2984) );
  assign n2985 = ~n2983 & n2984 ;
  buffer buf_n2986( .i (n2889), .o (n2986) );
  buffer buf_n2987( .i (n2986), .o (n2987) );
  buffer buf_n2988( .i (n2987), .o (n2988) );
  buffer buf_n2989( .i (n2988), .o (n2989) );
  buffer buf_n2990( .i (n2989), .o (n2990) );
  buffer buf_n2991( .i (n2990), .o (n2991) );
  assign n2992 = n607 & ~n2991 ;
  assign n2993 = n2984 | n2992 ;
  assign n2994 = ~n2985 & n2993 ;
  assign n2995 = ( n2975 & n2976 ) | ( n2975 & n2994 ) | ( n2976 & n2994 ) ;
  assign n2996 = n2977 & n2995 ;
  assign n2997 = n2955 | n2996 ;
  assign n2998 = ~n2929 & n2997 ;
  assign n2999 = n2930 | n2998 ;
  buffer buf_n3000( .i (n2999), .o (n3000) );
  assign n3001 = ( ~n2827 & n2832 ) | ( ~n2827 & n3000 ) | ( n2832 & n3000 ) ;
  buffer buf_n3002( .i (n2582), .o (n3002) );
  assign n3003 = n249 | n3002 ;
  buffer buf_n3004( .i (n3003), .o (n3004) );
  buffer buf_n3005( .i (n3004), .o (n3005) );
  buffer buf_n3006( .i (n3005), .o (n3006) );
  assign n3010 = ( n2492 & ~n2919 ) | ( n2492 & n3006 ) | ( ~n2919 & n3006 ) ;
  buffer buf_n3011( .i (n3010), .o (n3011) );
  buffer buf_n3012( .i (n3011), .o (n3012) );
  buffer buf_n3013( .i (n3012), .o (n3013) );
  buffer buf_n3014( .i (n3013), .o (n3014) );
  buffer buf_n3015( .i (n3014), .o (n3015) );
  buffer buf_n3016( .i (n3015), .o (n3016) );
  buffer buf_n3017( .i (n3016), .o (n3017) );
  buffer buf_n3018( .i (n3017), .o (n3018) );
  buffer buf_n3019( .i (n3018), .o (n3019) );
  buffer buf_n3020( .i (n3019), .o (n3020) );
  assign n3021 = n3000 | n3020 ;
  assign n3022 = ( n2828 & n3001 ) | ( n2828 & n3021 ) | ( n3001 & n3021 ) ;
  buffer buf_n3023( .i (n3022), .o (n3023) );
  buffer buf_n3024( .i (n3023), .o (n3024) );
  buffer buf_n3025( .i (n2620), .o (n3025) );
  assign n3026 = n3023 & n3025 ;
  assign n3027 = n604 & ~n2401 ;
  buffer buf_n3028( .i (n3027), .o (n3028) );
  buffer buf_n3029( .i (n3028), .o (n3029) );
  buffer buf_n3030( .i (n3029), .o (n3030) );
  buffer buf_n3031( .i (n3030), .o (n3031) );
  buffer buf_n3032( .i (n3031), .o (n3032) );
  buffer buf_n3033( .i (n3032), .o (n3033) );
  buffer buf_n3034( .i (n3033), .o (n3034) );
  buffer buf_n3035( .i (n3034), .o (n3035) );
  buffer buf_n3036( .i (n3035), .o (n3036) );
  buffer buf_n3037( .i (n3036), .o (n3037) );
  buffer buf_n3038( .i (n3037), .o (n3038) );
  buffer buf_n3039( .i (n3038), .o (n3039) );
  assign n3040 = n1248 & n3039 ;
  buffer buf_n3041( .i (n3040), .o (n3041) );
  assign n3042 = n22 & n2715 ;
  buffer buf_n3043( .i (n2400), .o (n3043) );
  buffer buf_n3044( .i (n3043), .o (n3044) );
  assign n3045 = ( n2900 & n3042 ) | ( n2900 & ~n3044 ) | ( n3042 & ~n3044 ) ;
  buffer buf_n3046( .i (n3045), .o (n3046) );
  buffer buf_n3047( .i (n3046), .o (n3047) );
  buffer buf_n3048( .i (n3047), .o (n3048) );
  assign n3049 = ( n25 & n2783 ) | ( n25 & ~n3046 ) | ( n2783 & ~n3046 ) ;
  assign n3050 = ( ~n198 & n2984 ) | ( ~n198 & n3049 ) | ( n2984 & n3049 ) ;
  assign n3051 = ~n3048 & n3050 ;
  assign n3052 = ~n1908 & n3051 ;
  assign n3053 = n1376 | n3052 ;
  assign n3054 = ( ~n1563 & n2121 ) | ( ~n1563 & n2385 ) | ( n2121 & n2385 ) ;
  assign n3055 = ~n2526 & n3054 ;
  buffer buf_n3056( .i (n2643), .o (n3056) );
  buffer buf_n3057( .i (n3056), .o (n3057) );
  assign n3058 = ~n3055 & n3057 ;
  assign n3059 = n3053 & ~n3058 ;
  assign n3060 = n2474 | n3059 ;
  buffer buf_n3061( .i (n2329), .o (n3061) );
  assign n3062 = ( n47 & n2911 ) | ( n47 & n3061 ) | ( n2911 & n3061 ) ;
  buffer buf_n3063( .i (n3062), .o (n3063) );
  buffer buf_n3064( .i (n3063), .o (n3064) );
  buffer buf_n3065( .i (n3064), .o (n3065) );
  buffer buf_n3070( .i (n1938), .o (n3070) );
  buffer buf_n3071( .i (n2899), .o (n3071) );
  assign n3072 = ( n3065 & ~n3070 ) | ( n3065 & n3071 ) | ( ~n3070 & n3071 ) ;
  buffer buf_n3073( .i (n3072), .o (n3073) );
  buffer buf_n3074( .i (n3073), .o (n3074) );
  buffer buf_n3075( .i (n3074), .o (n3075) );
  buffer buf_n3076( .i (n3075), .o (n3076) );
  assign n3077 = ( n1887 & n2970 ) | ( n1887 & n3073 ) | ( n2970 & n3073 ) ;
  buffer buf_n3078( .i (n3077), .o (n3078) );
  buffer buf_n3079( .i (n3078), .o (n3079) );
  buffer buf_n3066( .i (n3065), .o (n3066) );
  buffer buf_n3067( .i (n3066), .o (n3067) );
  buffer buf_n3068( .i (n3067), .o (n3068) );
  buffer buf_n3069( .i (n3068), .o (n3069) );
  assign n3080 = ~n3069 & n3078 ;
  assign n3081 = ( ~n3076 & n3079 ) | ( ~n3076 & n3080 ) | ( n3079 & n3080 ) ;
  assign n3082 = n1909 & n3081 ;
  assign n3083 = ~n1894 & n3082 ;
  assign n3084 = n2474 & ~n3083 ;
  assign n3085 = n3060 & ~n3084 ;
  assign n3086 = ~n2793 & n3085 ;
  buffer buf_n3087( .i (n3086), .o (n3087) );
  buffer buf_n3088( .i (n3087), .o (n3088) );
  buffer buf_n3089( .i (n2746), .o (n3089) );
  buffer buf_n3090( .i (n3089), .o (n3090) );
  assign n3091 = ( ~n1909 & n2559 ) | ( ~n1909 & n3090 ) | ( n2559 & n3090 ) ;
  buffer buf_n3092( .i (n3091), .o (n3092) );
  buffer buf_n3094( .i (n2736), .o (n3094) );
  buffer buf_n3095( .i (n3094), .o (n3095) );
  assign n3096 = ( n202 & n2752 ) | ( n202 & ~n3095 ) | ( n2752 & ~n3095 ) ;
  assign n3097 = ~n3092 & n3096 ;
  buffer buf_n3098( .i (n3097), .o (n3098) );
  buffer buf_n3099( .i (n3098), .o (n3099) );
  assign n3100 = n53 & n2394 ;
  buffer buf_n3101( .i (n3100), .o (n3101) );
  buffer buf_n3102( .i (n3101), .o (n3102) );
  buffer buf_n3103( .i (n3102), .o (n3103) );
  buffer buf_n3104( .i (n3103), .o (n3104) );
  buffer buf_n3105( .i (n3104), .o (n3105) );
  buffer buf_n3106( .i (n3105), .o (n3106) );
  buffer buf_n3107( .i (n3106), .o (n3107) );
  assign n3108 = ( n2689 & ~n3098 ) | ( n2689 & n3107 ) | ( ~n3098 & n3107 ) ;
  assign n3109 = n3099 & n3108 ;
  assign n3110 = n3087 | n3109 ;
  buffer buf_n3111( .i (n1786), .o (n3111) );
  assign n3112 = ( n3088 & n3110 ) | ( n3088 & ~n3111 ) | ( n3110 & ~n3111 ) ;
  assign n3113 = n3041 | n3112 ;
  assign n3114 = ( n3024 & ~n3026 ) | ( n3024 & n3113 ) | ( ~n3026 & n3113 ) ;
  assign n3115 = n2800 | n3114 ;
  assign n3116 = ( n2697 & ~n2714 ) | ( n2697 & n3115 ) | ( ~n2714 & n3115 ) ;
  buffer buf_n2713( .i (n2712), .o (n2713) );
  assign n3117 = n2961 & n3043 ;
  buffer buf_n3118( .i (n3117), .o (n3118) );
  buffer buf_n3119( .i (n3118), .o (n3119) );
  buffer buf_n3120( .i (n3119), .o (n3120) );
  buffer buf_n3121( .i (n3120), .o (n3121) );
  buffer buf_n3122( .i (n3121), .o (n3122) );
  buffer buf_n3123( .i (n3122), .o (n3123) );
  buffer buf_n3124( .i (n3123), .o (n3124) );
  buffer buf_n3125( .i (n3124), .o (n3125) );
  buffer buf_n3126( .i (n3125), .o (n3126) );
  buffer buf_n3127( .i (n3126), .o (n3127) );
  buffer buf_n3128( .i (n3127), .o (n3128) );
  buffer buf_n3129( .i (n3128), .o (n3129) );
  buffer buf_n3130( .i (n3129), .o (n3130) );
  buffer buf_n3131( .i (n3130), .o (n3131) );
  buffer buf_n2204( .i (n2203), .o (n2204) );
  buffer buf_n3132( .i (n3070), .o (n3132) );
  assign n3133 = ~n1826 & n3132 ;
  buffer buf_n3134( .i (n3133), .o (n3134) );
  buffer buf_n3135( .i (n3134), .o (n3135) );
  buffer buf_n3137( .i (n2783), .o (n3137) );
  buffer buf_n3138( .i (n3137), .o (n3138) );
  assign n3139 = n3135 & n3138 ;
  buffer buf_n3140( .i (n3132), .o (n3140) );
  buffer buf_n3141( .i (n3140), .o (n3141) );
  assign n3142 = ( n2972 & n3134 ) | ( n2972 & ~n3141 ) | ( n3134 & ~n3141 ) ;
  assign n3143 = ( n1946 & ~n3138 ) | ( n1946 & n3142 ) | ( ~n3138 & n3142 ) ;
  assign n3144 = ( n2975 & ~n3139 ) | ( n2975 & n3143 ) | ( ~n3139 & n3143 ) ;
  assign n3145 = ( n48 & ~n2433 ) | ( n48 & n2986 ) | ( ~n2433 & n2986 ) ;
  buffer buf_n3146( .i (n2540), .o (n3146) );
  assign n3147 = ( n828 & n3145 ) | ( n828 & ~n3146 ) | ( n3145 & ~n3146 ) ;
  buffer buf_n3148( .i (n3147), .o (n3148) );
  assign n3151 = n3070 & ~n3148 ;
  buffer buf_n3152( .i (n3151), .o (n3152) );
  buffer buf_n3153( .i (n3152), .o (n3153) );
  buffer buf_n3149( .i (n3148), .o (n3149) );
  buffer buf_n3150( .i (n3149), .o (n3150) );
  assign n3154 = n3150 | n3152 ;
  assign n3155 = ( ~n3141 & n3153 ) | ( ~n3141 & n3154 ) | ( n3153 & n3154 ) ;
  buffer buf_n3156( .i (n3155), .o (n3156) );
  buffer buf_n3157( .i (n3156), .o (n3157) );
  assign n3158 = n2736 & ~n3156 ;
  assign n3159 = ( n3144 & ~n3157 ) | ( n3144 & n3158 ) | ( ~n3157 & n3158 ) ;
  assign n3160 = n2927 & ~n3159 ;
  assign n3161 = ( n397 & ~n959 ) | ( n397 & n2729 ) | ( ~n959 & n2729 ) ;
  assign n3162 = n3056 | n3161 ;
  assign n3163 = n370 & n2783 ;
  buffer buf_n3164( .i (n3163), .o (n3164) );
  assign n3171 = n2746 & n3164 ;
  assign n3172 = n3056 & ~n3171 ;
  assign n3173 = n3162 & ~n3172 ;
  assign n3174 = n2927 | n3173 ;
  assign n3175 = ( ~n261 & n3160 ) | ( ~n261 & n3174 ) | ( n3160 & n3174 ) ;
  assign n3176 = ( n204 & ~n2533 ) | ( n204 & n3175 ) | ( ~n2533 & n3175 ) ;
  buffer buf_n3177( .i (n2972), .o (n3177) );
  assign n3178 = ( n2415 & n3138 ) | ( n2415 & ~n3177 ) | ( n3138 & ~n3177 ) ;
  assign n3179 = n1988 & ~n3178 ;
  buffer buf_n3180( .i (n3179), .o (n3180) );
  buffer buf_n3181( .i (n3180), .o (n3181) );
  assign n3182 = ( ~n423 & n2989 ) | ( ~n423 & n3071 ) | ( n2989 & n3071 ) ;
  buffer buf_n3183( .i (n2919), .o (n3183) );
  assign n3184 = ( n3132 & n3182 ) | ( n3132 & ~n3183 ) | ( n3182 & ~n3183 ) ;
  assign n3185 = ~n425 & n3184 ;
  assign n3186 = ( n2414 & ~n2984 ) | ( n2414 & n3185 ) | ( ~n2984 & n3185 ) ;
  buffer buf_n3187( .i (n101), .o (n3187) );
  assign n3188 = ( n46 & n2582 ) | ( n46 & n3187 ) | ( n2582 & n3187 ) ;
  buffer buf_n3189( .i (n3188), .o (n3189) );
  buffer buf_n3201( .i (n3002), .o (n3201) );
  assign n3202 = ( ~n2986 & n3189 ) | ( ~n2986 & n3201 ) | ( n3189 & n3201 ) ;
  buffer buf_n3203( .i (n3202), .o (n3203) );
  assign n3206 = n2918 & ~n3203 ;
  buffer buf_n3207( .i (n3206), .o (n3207) );
  buffer buf_n3208( .i (n3207), .o (n3208) );
  buffer buf_n3204( .i (n3203), .o (n3204) );
  buffer buf_n3205( .i (n3204), .o (n3205) );
  assign n3209 = n3205 | n3207 ;
  buffer buf_n3210( .i (n3183), .o (n3210) );
  assign n3211 = ( n3208 & n3209 ) | ( n3208 & ~n3210 ) | ( n3209 & ~n3210 ) ;
  buffer buf_n3212( .i (n2716), .o (n3212) );
  buffer buf_n3213( .i (n3212), .o (n3213) );
  buffer buf_n3214( .i (n3213), .o (n3214) );
  buffer buf_n3215( .i (n1816), .o (n3215) );
  assign n3216 = ( n3211 & n3214 ) | ( n3211 & n3215 ) | ( n3214 & n3215 ) ;
  assign n3217 = n3186 & n3216 ;
  buffer buf_n3218( .i (n3217), .o (n3218) );
  buffer buf_n3219( .i (n3218), .o (n3219) );
  buffer buf_n3220( .i (n3219), .o (n3220) );
  assign n3221 = ( ~n1701 & n3057 ) | ( ~n1701 & n3218 ) | ( n3057 & n3218 ) ;
  assign n3222 = n3180 & ~n3221 ;
  assign n3223 = ( n3181 & n3220 ) | ( n3181 & ~n3222 ) | ( n3220 & ~n3222 ) ;
  assign n3224 = ( n204 & n2533 ) | ( n204 & ~n3223 ) | ( n2533 & ~n3223 ) ;
  assign n3225 = n3176 & ~n3224 ;
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  assign n3226 = n1369 & ~n2016 ;
  assign n3227 = ( n1938 & ~n2918 ) | ( n1938 & n2961 ) | ( ~n2918 & n2961 ) ;
  buffer buf_n3228( .i (n3227), .o (n3228) );
  buffer buf_n3229( .i (n3228), .o (n3229) );
  buffer buf_n3230( .i (n3229), .o (n3230) );
  buffer buf_n3231( .i (n3230), .o (n3231) );
  assign n3232 = n1815 & ~n3228 ;
  buffer buf_n3233( .i (n3232), .o (n3233) );
  buffer buf_n3234( .i (n3233), .o (n3234) );
  assign n3235 = ( n2972 & n3141 ) | ( n2972 & n3233 ) | ( n3141 & n3233 ) ;
  assign n3236 = ( ~n3231 & n3234 ) | ( ~n3231 & n3235 ) | ( n3234 & n3235 ) ;
  assign n3237 = n2975 & n3236 ;
  assign n3238 = ~n29 & n3237 ;
  buffer buf_n3239( .i (n3238), .o (n3239) );
  buffer buf_n3240( .i (n3239), .o (n3240) );
  assign n3241 = n313 & ~n3239 ;
  assign n3242 = ( n3226 & n3240 ) | ( n3226 & ~n3241 ) | ( n3240 & ~n3241 ) ;
  assign n3243 = ( n177 & n2019 ) | ( n177 & ~n3242 ) | ( n2019 & ~n3242 ) ;
  assign n3244 = ( n2204 & n3225 ) | ( n2204 & ~n3243 ) | ( n3225 & ~n3243 ) ;
  assign n3245 = n237 & ~n3244 ;
  assign n3246 = ( n2716 & ~n2919 ) | ( n2716 & n3044 ) | ( ~n2919 & n3044 ) ;
  buffer buf_n3247( .i (n3246), .o (n3247) );
  buffer buf_n3248( .i (n3247), .o (n3248) );
  buffer buf_n3249( .i (n3248), .o (n3249) );
  buffer buf_n3250( .i (n3249), .o (n3250) );
  assign n3251 = n3210 & n3247 ;
  buffer buf_n3252( .i (n3251), .o (n3252) );
  buffer buf_n3253( .i (n3252), .o (n3253) );
  buffer buf_n3254( .i (n2970), .o (n3254) );
  buffer buf_n3255( .i (n3254), .o (n3255) );
  assign n3256 = ( n3138 & n3252 ) | ( n3138 & ~n3255 ) | ( n3252 & ~n3255 ) ;
  assign n3257 = ( n3250 & n3253 ) | ( n3250 & n3256 ) | ( n3253 & n3256 ) ;
  buffer buf_n3258( .i (n3257), .o (n3258) );
  buffer buf_n3259( .i (n3258), .o (n3259) );
  buffer buf_n3260( .i (n3090), .o (n3260) );
  assign n3261 = n3258 & ~n3260 ;
  buffer buf_n3262( .i (n2490), .o (n3262) );
  assign n3263 = ( n2715 & n2918 ) | ( n2715 & ~n3262 ) | ( n2918 & ~n3262 ) ;
  buffer buf_n3264( .i (n3263), .o (n3264) );
  buffer buf_n3265( .i (n3264), .o (n3265) );
  buffer buf_n3266( .i (n3265), .o (n3266) );
  buffer buf_n3268( .i (n3262), .o (n3268) );
  buffer buf_n3269( .i (n3268), .o (n3269) );
  assign n3270 = ( n2981 & ~n3212 ) | ( n2981 & n3269 ) | ( ~n3212 & n3269 ) ;
  assign n3271 = ~n3210 & n3270 ;
  assign n3272 = n3266 | n3271 ;
  buffer buf_n3273( .i (n3272), .o (n3273) );
  buffer buf_n3274( .i (n3273), .o (n3274) );
  buffer buf_n3275( .i (n3137), .o (n3275) );
  buffer buf_n3276( .i (n3275), .o (n3276) );
  assign n3277 = ( n3089 & ~n3273 ) | ( n3089 & n3276 ) | ( ~n3273 & n3276 ) ;
  assign n3278 = n1755 | n3212 ;
  buffer buf_n3279( .i (n3278), .o (n3279) );
  assign n3289 = n2595 & ~n3279 ;
  assign n3290 = n3177 & n3289 ;
  assign n3291 = ~n3276 & n3290 ;
  assign n3292 = ( n3274 & n3277 ) | ( n3274 & ~n3291 ) | ( n3277 & ~n3291 ) ;
  buffer buf_n2933( .i (n2932), .o (n2933) );
  buffer buf_n2934( .i (n2933), .o (n2934) );
  buffer buf_n2935( .i (n2934), .o (n2935) );
  assign n3293 = n2935 & ~n2976 ;
  assign n3294 = ~n2199 & n3293 ;
  assign n3295 = n3292 & ~n3294 ;
  assign n3296 = ( ~n3259 & n3261 ) | ( ~n3259 & n3295 ) | ( n3261 & n3295 ) ;
  buffer buf_n3297( .i (n2929), .o (n3297) );
  assign n3298 = ~n3296 & n3297 ;
  buffer buf_n2310( .i (n2309), .o (n2310) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  assign n3299 = ( n1311 & n2312 ) | ( n1311 & ~n2970 ) | ( n2312 & ~n2970 ) ;
  assign n3300 = ~n2313 & n3299 ;
  buffer buf_n3301( .i (n3300), .o (n3301) );
  buffer buf_n3302( .i (n3301), .o (n3302) );
  buffer buf_n3303( .i (n3302), .o (n3303) );
  assign n3304 = ( n2009 & n3122 ) | ( n2009 & n3301 ) | ( n3122 & n3301 ) ;
  assign n3305 = n3094 & ~n3304 ;
  assign n3306 = ( n3095 & n3303 ) | ( n3095 & ~n3305 ) | ( n3303 & ~n3305 ) ;
  assign n3307 = ( n2400 & n2490 ) | ( n2400 & n2917 ) | ( n2490 & n2917 ) ;
  buffer buf_n3308( .i (n3307), .o (n3308) );
  buffer buf_n3309( .i (n3308), .o (n3309) );
  buffer buf_n3310( .i (n3309), .o (n3310) );
  buffer buf_n3311( .i (n3269), .o (n3311) );
  assign n3312 = n3310 & n3311 ;
  assign n3313 = ( n2990 & n3183 ) | ( n2990 & n3309 ) | ( n3183 & n3309 ) ;
  assign n3314 = n3311 | n3313 ;
  assign n3315 = ~n3312 & n3314 ;
  assign n3316 = n3275 | n3315 ;
  buffer buf_n3317( .i (n2991), .o (n3317) );
  assign n3318 = n1049 & n3317 ;
  assign n3319 = n3275 & ~n3318 ;
  assign n3320 = n3316 & ~n3319 ;
  assign n3321 = n3094 | n3320 ;
  assign n3322 = ~n2357 & n3122 ;
  assign n3323 = n3094 & ~n3322 ;
  assign n3324 = n3321 & ~n3323 ;
  assign n3325 = n3306 | n3324 ;
  assign n3326 = ~n3297 & n3325 ;
  assign n3327 = n3298 | n3326 ;
  assign n3328 = ~n2110 & n3327 ;
  assign n3329 = n237 | n3328 ;
  assign n3330 = ~n3245 & n3329 ;
  assign n3331 = ( n21 & n2917 ) | ( n21 & n3146 ) | ( n2917 & n3146 ) ;
  buffer buf_n3332( .i (n3331), .o (n3332) );
  buffer buf_n3337( .i (n2917), .o (n3337) );
  buffer buf_n3338( .i (n3337), .o (n3338) );
  buffer buf_n3339( .i (n2895), .o (n3339) );
  buffer buf_n3340( .i (n3339), .o (n3340) );
  assign n3341 = ( ~n3332 & n3338 ) | ( ~n3332 & n3340 ) | ( n3338 & n3340 ) ;
  buffer buf_n3342( .i (n3341), .o (n3342) );
  buffer buf_n3343( .i (n3342), .o (n3343) );
  buffer buf_n3344( .i (n3343), .o (n3344) );
  buffer buf_n3345( .i (n3344), .o (n3345) );
  assign n3346 = ( n25 & n3213 ) | ( n25 & ~n3342 ) | ( n3213 & ~n3342 ) ;
  buffer buf_n3347( .i (n3346), .o (n3347) );
  buffer buf_n3348( .i (n3347), .o (n3348) );
  buffer buf_n3333( .i (n3332), .o (n3333) );
  buffer buf_n3334( .i (n3333), .o (n3334) );
  buffer buf_n3335( .i (n3334), .o (n3335) );
  buffer buf_n3336( .i (n3335), .o (n3336) );
  assign n3349 = ~n3336 & n3347 ;
  assign n3350 = ( n3345 & n3348 ) | ( n3345 & n3349 ) | ( n3348 & n3349 ) ;
  buffer buf_n3351( .i (n3350), .o (n3351) );
  buffer buf_n3352( .i (n3351), .o (n3352) );
  assign n3353 = n2740 & n3351 ;
  assign n3354 = ( n1776 & n2508 ) | ( n1776 & n2595 ) | ( n2508 & n2595 ) ;
  buffer buf_n3355( .i (n3354), .o (n3355) );
  assign n3356 = ( ~n2976 & n3056 ) | ( ~n2976 & n3355 ) | ( n3056 & n3355 ) ;
  buffer buf_n3357( .i (n2643), .o (n3357) );
  assign n3358 = ( n2526 & ~n3355 ) | ( n2526 & n3357 ) | ( ~n3355 & n3357 ) ;
  assign n3359 = n3356 & ~n3358 ;
  buffer buf_n3360( .i (n2596), .o (n3360) );
  assign n3361 = n729 & ~n3360 ;
  assign n3362 = ~n1508 & n3361 ;
  assign n3363 = n3359 | n3362 ;
  assign n3364 = ( n3352 & ~n3353 ) | ( n3352 & n3363 ) | ( ~n3353 & n3363 ) ;
  assign n3365 = n88 | n3364 ;
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n3366( .i (n2736), .o (n3366) );
  assign n3367 = ( ~n1614 & n3057 ) | ( ~n1614 & n3366 ) | ( n3057 & n3366 ) ;
  buffer buf_n3368( .i (n2940), .o (n3368) );
  assign n3369 = ( n3140 & ~n3213 ) | ( n3140 & n3368 ) | ( ~n3213 & n3368 ) ;
  buffer buf_n3370( .i (n3369), .o (n3370) );
  buffer buf_n3371( .i (n3370), .o (n3371) );
  buffer buf_n3372( .i (n3371), .o (n3372) );
  assign n3373 = n3057 & ~n3372 ;
  assign n3374 = n3367 & ~n3373 ;
  buffer buf_n3375( .i (n1894), .o (n3375) );
  assign n3376 = n3374 & ~n3375 ;
  buffer buf_n3377( .i (n3260), .o (n3377) );
  buffer buf_n3378( .i (n3377), .o (n3378) );
  assign n3379 = ~n3376 & n3378 ;
  assign n3380 = n3365 & ~n3379 ;
  assign n3381 = n118 | n3380 ;
  assign n3382 = n2735 & n2769 ;
  buffer buf_n3383( .i (n3382), .o (n3383) );
  assign n3387 = ~n3090 & n3383 ;
  assign n3388 = ( n596 & ~n3260 ) | ( n596 & n3387 ) | ( ~n3260 & n3387 ) ;
  assign n3389 = n2929 & ~n3388 ;
  buffer buf_n3390( .i (n2735), .o (n3390) );
  assign n3391 = ( n1908 & n3089 ) | ( n1908 & n3390 ) | ( n3089 & n3390 ) ;
  buffer buf_n3392( .i (n3360), .o (n3392) );
  assign n3393 = n3391 & n3392 ;
  assign n3394 = ( n530 & n2634 ) | ( n530 & ~n3393 ) | ( n2634 & ~n3393 ) ;
  buffer buf_n3395( .i (n2740), .o (n3395) );
  assign n3396 = n3394 | n3395 ;
  assign n3397 = ( ~n3297 & n3389 ) | ( ~n3297 & n3396 ) | ( n3389 & n3396 ) ;
  buffer buf_n3398( .i (n2533), .o (n3398) );
  assign n3399 = n3397 | n3398 ;
  buffer buf_n3400( .i (n2689), .o (n3400) );
  assign n3401 = n3399 & n3400 ;
  assign n3402 = n3381 & ~n3401 ;
  assign n3403 = ( n208 & n266 ) | ( n208 & n3402 ) | ( n266 & n3402 ) ;
  assign n3404 = ( ~n3131 & n3330 ) | ( ~n3131 & n3403 ) | ( n3330 & n3403 ) ;
  buffer buf_n3405( .i (n3404), .o (n3405) );
  buffer buf_n3406( .i (n3405), .o (n3406) );
  assign n3407 = ( n3089 & ~n3357 ) | ( n3089 & n3390 ) | ( ~n3357 & n3390 ) ;
  buffer buf_n3408( .i (n3407), .o (n3408) );
  buffer buf_n3409( .i (n3408), .o (n3409) );
  buffer buf_n3410( .i (n3409), .o (n3410) );
  assign n3411 = ( n234 & n2535 ) | ( n234 & ~n3410 ) | ( n2535 & ~n3410 ) ;
  assign n3412 = ( n234 & ~n3378 ) | ( n234 & n3410 ) | ( ~n3378 & n3410 ) ;
  assign n3413 = n3411 & ~n3412 ;
  buffer buf_n3414( .i (n3413), .o (n3414) );
  buffer buf_n3415( .i (n3414), .o (n3415) );
  buffer buf_n3416( .i (n2110), .o (n3416) );
  assign n3417 = n3414 & n3416 ;
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n3418( .i (n233), .o (n3418) );
  assign n3419 = n709 & n3418 ;
  buffer buf_n3420( .i (n3378), .o (n3420) );
  buffer buf_n3421( .i (n2535), .o (n3421) );
  assign n3422 = ( n3419 & n3420 ) | ( n3419 & n3421 ) | ( n3420 & n3421 ) ;
  buffer buf_n3423( .i (n3420), .o (n3423) );
  assign n3424 = n3422 & ~n3423 ;
  buffer buf_n3384( .i (n3383), .o (n3384) );
  buffer buf_n3385( .i (n3384), .o (n3385) );
  buffer buf_n3386( .i (n3385), .o (n3386) );
  buffer buf_n3425( .i (n24), .o (n3425) );
  assign n3426 = ( n3140 & n3210 ) | ( n3140 & n3425 ) | ( n3210 & n3425 ) ;
  buffer buf_n3427( .i (n3426), .o (n3427) );
  assign n3428 = ( n2524 & n2644 ) | ( n2524 & ~n3427 ) | ( n2644 & ~n3427 ) ;
  buffer buf_n3429( .i (n3141), .o (n3429) );
  assign n3430 = ( n2644 & n3427 ) | ( n2644 & ~n3429 ) | ( n3427 & ~n3429 ) ;
  assign n3431 = ~n3428 & n3430 ;
  buffer buf_n3432( .i (n3431), .o (n3432) );
  buffer buf_n3433( .i (n3432), .o (n3433) );
  buffer buf_n3434( .i (n3433), .o (n3434) );
  buffer buf_n3435( .i (n2526), .o (n3435) );
  buffer buf_n3436( .i (n3435), .o (n3436) );
  buffer buf_n3437( .i (n3357), .o (n3437) );
  buffer buf_n3438( .i (n3437), .o (n3438) );
  assign n3439 = ( ~n3432 & n3436 ) | ( ~n3432 & n3438 ) | ( n3436 & n3438 ) ;
  assign n3440 = n3385 & n3439 ;
  assign n3441 = ( n3386 & n3434 ) | ( n3386 & ~n3440 ) | ( n3434 & ~n3440 ) ;
  assign n3442 = n3420 | n3441 ;
  buffer buf_n3443( .i (n3368), .o (n3443) );
  buffer buf_n3444( .i (n3443), .o (n3444) );
  buffer buf_n3445( .i (n3444), .o (n3445) );
  assign n3446 = ( n3357 & n3360 ) | ( n3357 & ~n3445 ) | ( n3360 & ~n3445 ) ;
  buffer buf_n3447( .i (n3446), .o (n3447) );
  assign n3448 = ( ~n2577 & n3095 ) | ( ~n2577 & n3447 ) | ( n3095 & n3447 ) ;
  assign n3449 = ( n3095 & n3438 ) | ( n3095 & ~n3447 ) | ( n3438 & ~n3447 ) ;
  assign n3450 = n3448 & ~n3449 ;
  buffer buf_n3451( .i (n3375), .o (n3451) );
  assign n3452 = n3450 & ~n3451 ;
  assign n3453 = n3420 & ~n3452 ;
  assign n3454 = n3442 & ~n3453 ;
  assign n3455 = n3424 | n3454 ;
  assign n3456 = ( n3415 & ~n3417 ) | ( n3415 & n3455 ) | ( ~n3417 & n3455 ) ;
  assign n3457 = n121 | n3456 ;
  assign n3458 = n3378 & ~n3418 ;
  buffer buf_n3459( .i (n3377), .o (n3459) );
  buffer buf_n3460( .i (n3459), .o (n3460) );
  assign n3461 = ( n599 & n3458 ) | ( n599 & ~n3460 ) | ( n3458 & ~n3460 ) ;
  assign n3462 = n2364 & n3461 ;
  buffer buf_n3463( .i (n3201), .o (n3463) );
  assign n3464 = ( n2895 & n2987 ) | ( n2895 & ~n3463 ) | ( n2987 & ~n3463 ) ;
  buffer buf_n3465( .i (n3464), .o (n3465) );
  buffer buf_n3466( .i (n3465), .o (n3466) );
  buffer buf_n3467( .i (n3466), .o (n3467) );
  buffer buf_n3468( .i (n3467), .o (n3468) );
  buffer buf_n3469( .i (n3468), .o (n3469) );
  buffer buf_n3470( .i (n3469), .o (n3470) );
  assign n3475 = ( n3390 & ~n3445 ) | ( n3390 & n3470 ) | ( ~n3445 & n3470 ) ;
  buffer buf_n3476( .i (n3475), .o (n3476) );
  buffer buf_n3477( .i (n3476), .o (n3477) );
  buffer buf_n3478( .i (n3477), .o (n3478) );
  buffer buf_n3479( .i (n3478), .o (n3479) );
  assign n3480 = ( ~n2577 & n3260 ) | ( ~n2577 & n3476 ) | ( n3260 & n3476 ) ;
  buffer buf_n3481( .i (n3480), .o (n3481) );
  buffer buf_n3482( .i (n3481), .o (n3482) );
  buffer buf_n3471( .i (n3470), .o (n3471) );
  buffer buf_n3472( .i (n3471), .o (n3472) );
  buffer buf_n3473( .i (n3472), .o (n3473) );
  buffer buf_n3474( .i (n3473), .o (n3474) );
  assign n3483 = ~n3474 & n3481 ;
  assign n3484 = ( ~n3479 & n3482 ) | ( ~n3479 & n3483 ) | ( n3482 & n3483 ) ;
  buffer buf_n3485( .i (n2831), .o (n3485) );
  assign n3486 = n3484 | n3485 ;
  assign n3487 = ( ~n63 & n3462 ) | ( ~n63 & n3486 ) | ( n3462 & n3486 ) ;
  assign n3488 = ~n3111 & n3487 ;
  buffer buf_n3489( .i (n120), .o (n3489) );
  assign n3490 = ~n3488 & n3489 ;
  assign n3491 = n3457 & ~n3490 ;
  assign n3492 = n3405 | n3491 ;
  assign n3493 = ( ~n2713 & n3406 ) | ( ~n2713 & n3492 ) | ( n3406 & n3492 ) ;
  buffer buf_n361( .i (n360), .o (n361) );
  assign n3494 = n24 & ~n2981 ;
  buffer buf_n3495( .i (n3494), .o (n3495) );
  buffer buf_n3496( .i (n3495), .o (n3496) );
  assign n3497 = ( ~n2596 & n3444 ) | ( ~n2596 & n3496 ) | ( n3444 & n3496 ) ;
  assign n3498 = ( n3254 & ~n3443 ) | ( n3254 & n3495 ) | ( ~n3443 & n3495 ) ;
  buffer buf_n3499( .i (n2595), .o (n3499) );
  assign n3500 = ( ~n2524 & n3498 ) | ( ~n2524 & n3499 ) | ( n3498 & n3499 ) ;
  assign n3501 = n3497 | n3500 ;
  assign n3502 = ~n2821 & n3501 ;
  buffer buf_n2035( .i (n2034), .o (n2035) );
  buffer buf_n2036( .i (n2035), .o (n2036) );
  buffer buf_n2037( .i (n2036), .o (n2037) );
  buffer buf_n2038( .i (n2037), .o (n2038) );
  buffer buf_n2039( .i (n2038), .o (n2039) );
  buffer buf_n3503( .i (n3183), .o (n3503) );
  buffer buf_n3504( .i (n3503), .o (n3504) );
  assign n3505 = n2039 & ~n3504 ;
  buffer buf_n3506( .i (n3505), .o (n3506) );
  buffer buf_n3510( .i (n2508), .o (n3510) );
  buffer buf_n3511( .i (n3510), .o (n3511) );
  assign n3512 = n3506 & ~n3511 ;
  assign n3513 = n2821 & ~n3512 ;
  assign n3514 = n3502 | n3513 ;
  assign n3515 = ~n3377 & n3514 ;
  assign n3516 = ( n2854 & ~n2895 ) | ( n2854 & n3463 ) | ( ~n2895 & n3463 ) ;
  buffer buf_n3517( .i (n3516), .o (n3517) );
  buffer buf_n3518( .i (n3517), .o (n3518) );
  buffer buf_n3519( .i (n3518), .o (n3519) );
  buffer buf_n3520( .i (n3519), .o (n3520) );
  buffer buf_n3521( .i (n3520), .o (n3521) );
  buffer buf_n3522( .i (n3521), .o (n3522) );
  assign n3523 = ( n2558 & ~n3276 ) | ( n2558 & n3522 ) | ( ~n3276 & n3522 ) ;
  assign n3524 = ( ~n2558 & n3445 ) | ( ~n2558 & n3522 ) | ( n3445 & n3522 ) ;
  assign n3525 = n3523 & n3524 ;
  assign n3526 = ~n3436 & n3525 ;
  assign n3527 = n3377 & ~n3526 ;
  assign n3528 = n3515 | n3527 ;
  assign n3529 = ~n2831 & n3528 ;
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  assign n3530 = n865 & n3504 ;
  buffer buf_n3531( .i (n3530), .o (n3531) );
  buffer buf_n3532( .i (n3531), .o (n3532) );
  buffer buf_n3533( .i (n3532), .o (n3533) );
  buffer buf_n3535( .i (n3090), .o (n3535) );
  assign n3536 = ~n3533 & n3535 ;
  assign n3537 = n2121 & ~n3499 ;
  buffer buf_n3538( .i (n3537), .o (n3538) );
  assign n3539 = ~n2821 & n3538 ;
  assign n3540 = n3535 | n3539 ;
  assign n3541 = ~n3536 & n3540 ;
  assign n3542 = ~n3451 & n3541 ;
  assign n3543 = n2831 & ~n3542 ;
  assign n3544 = n3529 | n3543 ;
  buffer buf_n3545( .i (n3544), .o (n3545) );
  buffer buf_n3546( .i (n3545), .o (n3546) );
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n2321( .i (n2320), .o (n2321) );
  buffer buf_n2322( .i (n2321), .o (n2322) );
  buffer buf_n2323( .i (n2322), .o (n2323) );
  assign n3547 = n2323 | n3545 ;
  buffer buf_n3548( .i (n2762), .o (n3548) );
  assign n3549 = ( ~n21 & n3146 ) | ( ~n21 & n3548 ) | ( n3146 & n3548 ) ;
  buffer buf_n3550( .i (n3549), .o (n3550) );
  assign n3555 = ( n3268 & n3340 ) | ( n3268 & ~n3550 ) | ( n3340 & ~n3550 ) ;
  buffer buf_n3556( .i (n3555), .o (n3556) );
  buffer buf_n3557( .i (n3556), .o (n3557) );
  buffer buf_n3558( .i (n3557), .o (n3558) );
  buffer buf_n3559( .i (n3558), .o (n3559) );
  assign n3560 = ( ~n3213 & n3425 ) | ( ~n3213 & n3556 ) | ( n3425 & n3556 ) ;
  buffer buf_n3561( .i (n3560), .o (n3561) );
  buffer buf_n3562( .i (n3561), .o (n3562) );
  buffer buf_n3551( .i (n3550), .o (n3551) );
  buffer buf_n3552( .i (n3551), .o (n3552) );
  buffer buf_n3553( .i (n3552), .o (n3553) );
  buffer buf_n3554( .i (n3553), .o (n3554) );
  assign n3563 = n3554 & n3561 ;
  assign n3564 = ( ~n3559 & n3562 ) | ( ~n3559 & n3563 ) | ( n3562 & n3563 ) ;
  assign n3565 = ~n3392 & n3564 ;
  assign n3566 = n3438 | n3565 ;
  assign n3567 = ~n2314 & n3444 ;
  assign n3568 = n3360 & n3567 ;
  assign n3569 = ~n3435 & n3568 ;
  assign n3570 = n3438 & ~n3569 ;
  assign n3571 = n3566 & ~n3570 ;
  assign n3572 = n2688 | n3571 ;
  assign n3573 = ~n595 & n3437 ;
  assign n3574 = ( n596 & n612 ) | ( n596 & n3573 ) | ( n612 & n3573 ) ;
  assign n3575 = ~n3375 & n3574 ;
  assign n3576 = n2688 & ~n3575 ;
  assign n3577 = n3572 & ~n3576 ;
  assign n3578 = n3423 | n3577 ;
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  assign n3579 = ( n611 & ~n2722 ) | ( n611 & n3392 ) | ( ~n2722 & n3392 ) ;
  assign n3580 = ~n2166 & n3579 ;
  assign n3581 = n3395 & n3580 ;
  assign n3582 = ( n3070 & ~n3268 ) | ( n3070 & n3340 ) | ( ~n3268 & n3340 ) ;
  buffer buf_n3583( .i (n3582), .o (n3583) );
  buffer buf_n3584( .i (n3212), .o (n3584) );
  assign n3585 = ( ~n3311 & n3583 ) | ( ~n3311 & n3584 ) | ( n3583 & n3584 ) ;
  buffer buf_n3586( .i (n3585), .o (n3586) );
  assign n3589 = n2415 & n3586 ;
  buffer buf_n3590( .i (n3589), .o (n3590) );
  buffer buf_n3591( .i (n3590), .o (n3591) );
  buffer buf_n3587( .i (n3586), .o (n3587) );
  buffer buf_n3588( .i (n3587), .o (n3588) );
  assign n3592 = n3588 & ~n3590 ;
  assign n3593 = ( n2927 & ~n3591 ) | ( n2927 & n3592 ) | ( ~n3591 & n3592 ) ;
  assign n3594 = ( n2016 & ~n2685 ) | ( n2016 & n3593 ) | ( ~n2685 & n3593 ) ;
  assign n3595 = ( n570 & ~n3581 ) | ( n570 & n3594 ) | ( ~n3581 & n3594 ) ;
  assign n3596 = n3398 | n3595 ;
  assign n3597 = n3423 & n3596 ;
  assign n3598 = n3578 & ~n3597 ;
  assign n3599 = ( n454 & ~n2240 ) | ( n454 & n2608 ) | ( ~n2240 & n2608 ) ;
  buffer buf_n3600( .i (n3599), .o (n3600) );
  buffer buf_n3609( .i (n2782), .o (n3609) );
  assign n3610 = ~n1057 & n3609 ;
  buffer buf_n3611( .i (n3610), .o (n3611) );
  assign n3612 = ~n3600 & n3611 ;
  assign n3613 = n3119 & ~n3584 ;
  buffer buf_n3614( .i (n3613), .o (n3614) );
  assign n3616 = ( ~n1059 & n3611 ) | ( ~n1059 & n3614 ) | ( n3611 & n3614 ) ;
  buffer buf_n3617( .i (n3499), .o (n3617) );
  assign n3618 = ( n3612 & n3616 ) | ( n3612 & n3617 ) | ( n3616 & n3617 ) ;
  buffer buf_n3619( .i (n3177), .o (n3619) );
  buffer buf_n3620( .i (n3619), .o (n3620) );
  assign n3621 = n3618 | n3620 ;
  assign n3622 = n2608 & ~n3584 ;
  buffer buf_n3623( .i (n3622), .o (n3623) );
  buffer buf_n3624( .i (n3623), .o (n3624) );
  assign n3625 = n398 & n3624 ;
  assign n3626 = n3620 & ~n3625 ;
  assign n3627 = n3621 & ~n3626 ;
  buffer buf_n3628( .i (n3627), .o (n3628) );
  buffer buf_n3629( .i (n3628), .o (n3629) );
  assign n3630 = ( n654 & n2940 ) | ( n654 & n2981 ) | ( n2940 & n2981 ) ;
  buffer buf_n3631( .i (n3044), .o (n3631) );
  assign n3632 = ( n654 & ~n3269 ) | ( n654 & n3631 ) | ( ~n3269 & n3631 ) ;
  assign n3633 = ( n332 & ~n3630 ) | ( n332 & n3632 ) | ( ~n3630 & n3632 ) ;
  assign n3634 = n3214 & n3633 ;
  buffer buf_n3635( .i (n3338), .o (n3635) );
  assign n3636 = n3028 & n3635 ;
  buffer buf_n3637( .i (n3636), .o (n3637) );
  assign n3641 = n3214 | n3637 ;
  assign n3642 = ~n3634 & n3641 ;
  assign n3643 = n3619 & ~n3642 ;
  assign n3644 = n372 & n2135 ;
  assign n3645 = n3619 | n3644 ;
  assign n3646 = ~n3643 & n3645 ;
  assign n3647 = ( n1275 & n2582 ) | ( n1275 & n2888 ) | ( n2582 & n2888 ) ;
  buffer buf_n3648( .i (n3647), .o (n3648) );
  assign n3653 = ( n2853 & n2986 ) | ( n2853 & ~n3648 ) | ( n2986 & ~n3648 ) ;
  buffer buf_n3654( .i (n3653), .o (n3654) );
  buffer buf_n3655( .i (n3654), .o (n3655) );
  buffer buf_n3656( .i (n3655), .o (n3656) );
  buffer buf_n3657( .i (n3656), .o (n3657) );
  assign n3658 = ( n3337 & n3339 ) | ( n3337 & ~n3654 ) | ( n3339 & ~n3654 ) ;
  buffer buf_n3659( .i (n3658), .o (n3659) );
  buffer buf_n3660( .i (n3659), .o (n3660) );
  buffer buf_n3649( .i (n3648), .o (n3649) );
  buffer buf_n3650( .i (n3649), .o (n3650) );
  buffer buf_n3651( .i (n3650), .o (n3651) );
  buffer buf_n3652( .i (n3651), .o (n3652) );
  assign n3661 = ~n3652 & n3659 ;
  assign n3662 = ( n3657 & n3660 ) | ( n3657 & n3661 ) | ( n3660 & n3661 ) ;
  buffer buf_n3663( .i (n3662), .o (n3663) );
  buffer buf_n3664( .i (n3663), .o (n3664) );
  buffer buf_n3665( .i (n2716), .o (n3665) );
  assign n3666 = n492 & n3665 ;
  buffer buf_n3667( .i (n3666), .o (n3667) );
  buffer buf_n3668( .i (n3667), .o (n3668) );
  assign n3669 = n3663 & n3668 ;
  assign n3670 = ( n3624 & n3664 ) | ( n3624 & n3669 ) | ( n3664 & n3669 ) ;
  buffer buf_n3671( .i (n3670), .o (n3671) );
  assign n3672 = ( ~n2166 & n3646 ) | ( ~n2166 & n3671 ) | ( n3646 & n3671 ) ;
  buffer buf_n3673( .i (n3631), .o (n3673) );
  assign n3674 = n2991 & ~n3673 ;
  assign n3675 = n525 & n3368 ;
  assign n3676 = ( n2120 & n3674 ) | ( n2120 & ~n3675 ) | ( n3674 & ~n3675 ) ;
  buffer buf_n3677( .i (n2231), .o (n3677) );
  assign n3678 = ( n73 & n131 ) | ( n73 & ~n3677 ) | ( n131 & ~n3677 ) ;
  buffer buf_n3679( .i (n3678), .o (n3679) );
  assign n3687 = ( ~n2761 & n2889 ) | ( ~n2761 & n3679 ) | ( n2889 & n3679 ) ;
  buffer buf_n3688( .i (n3687), .o (n3688) );
  assign n3691 = n2987 & ~n3688 ;
  buffer buf_n3692( .i (n3691), .o (n3692) );
  buffer buf_n3693( .i (n3692), .o (n3693) );
  buffer buf_n3689( .i (n3688), .o (n3689) );
  buffer buf_n3690( .i (n3689), .o (n3690) );
  assign n3694 = n3690 | n3692 ;
  assign n3695 = ( ~n2990 & n3693 ) | ( ~n2990 & n3694 ) | ( n3693 & n3694 ) ;
  buffer buf_n3696( .i (n3695), .o (n3696) );
  buffer buf_n3697( .i (n3696), .o (n3697) );
  assign n3698 = n3215 | n3696 ;
  assign n3699 = ( n3676 & n3697 ) | ( n3676 & n3698 ) | ( n3697 & n3698 ) ;
  assign n3700 = n3390 | n3699 ;
  assign n3701 = ( ~n3311 & n3368 ) | ( ~n3311 & n3673 ) | ( n3368 & n3673 ) ;
  assign n3702 = ( n2989 & ~n3044 ) | ( n2989 & n3268 ) | ( ~n3044 & n3268 ) ;
  buffer buf_n3703( .i (n3702), .o (n3703) );
  buffer buf_n3713( .i (n2940), .o (n3713) );
  assign n3714 = ~n3703 & n3713 ;
  assign n3715 = n3701 & ~n3714 ;
  assign n3716 = ~n3499 & n3715 ;
  buffer buf_n3717( .i (n2735), .o (n3717) );
  assign n3718 = ~n3716 & n3717 ;
  assign n3719 = n3700 & ~n3718 ;
  buffer buf_n3720( .i (n3276), .o (n3720) );
  buffer buf_n3721( .i (n3720), .o (n3721) );
  assign n3722 = ( n3671 & n3719 ) | ( n3671 & n3721 ) | ( n3719 & n3721 ) ;
  assign n3723 = n3672 | n3722 ;
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  assign n3724 = n373 & n3511 ;
  assign n3725 = ( n589 & ~n1760 ) | ( n589 & n3724 ) | ( ~n1760 & n3724 ) ;
  assign n3726 = ~n590 & n3725 ;
  buffer buf_n3727( .i (n3726), .o (n3727) );
  assign n3728 = ( ~n3628 & n3723 ) | ( ~n3628 & n3727 ) | ( n3723 & n3727 ) ;
  assign n3729 = n3451 & ~n3727 ;
  assign n3730 = ( n3629 & n3728 ) | ( n3629 & ~n3729 ) | ( n3728 & ~n3729 ) ;
  assign n3731 = n3485 | n3730 ;
  buffer buf_n3732( .i (n2888), .o (n3732) );
  buffer buf_n3733( .i (n3732), .o (n3733) );
  assign n3734 = ( n2540 & ~n3201 ) | ( n2540 & n3733 ) | ( ~n3201 & n3733 ) ;
  assign n3735 = ( n2987 & ~n3548 ) | ( n2987 & n3734 ) | ( ~n3548 & n3734 ) ;
  buffer buf_n3736( .i (n3735), .o (n3736) );
  assign n3739 = n2989 & ~n3736 ;
  buffer buf_n3740( .i (n3739), .o (n3740) );
  buffer buf_n3741( .i (n3740), .o (n3741) );
  buffer buf_n3737( .i (n3736), .o (n3737) );
  buffer buf_n3738( .i (n3737), .o (n3738) );
  assign n3742 = n3738 | n3740 ;
  assign n3743 = ( ~n3317 & n3741 ) | ( ~n3317 & n3742 ) | ( n3741 & n3742 ) ;
  buffer buf_n3744( .i (n3215), .o (n3744) );
  assign n3745 = n3743 & n3744 ;
  assign n3746 = ( n2006 & ~n2718 ) | ( n2006 & n3713 ) | ( ~n2718 & n3713 ) ;
  assign n3747 = ( n2718 & n2991 ) | ( n2718 & ~n3713 ) | ( n2991 & ~n3713 ) ;
  assign n3748 = ( ~n3317 & n3746 ) | ( ~n3317 & n3747 ) | ( n3746 & n3747 ) ;
  assign n3749 = n3744 | n3748 ;
  assign n3750 = ( ~n2950 & n3745 ) | ( ~n2950 & n3749 ) | ( n3745 & n3749 ) ;
  assign n3751 = n3720 & ~n3750 ;
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n2519( .i (n2518), .o (n2519) );
  buffer buf_n3752( .i (n3269), .o (n3752) );
  assign n3753 = ( n3503 & ~n3584 ) | ( n3503 & n3752 ) | ( ~n3584 & n3752 ) ;
  assign n3754 = ~n3317 & n3753 ;
  assign n3755 = ( n1671 & n2519 ) | ( n1671 & ~n3754 ) | ( n2519 & ~n3754 ) ;
  assign n3756 = n3445 | n3755 ;
  assign n3757 = ~n3720 & n3756 ;
  assign n3758 = n3751 | n3757 ;
  assign n3759 = n2824 & ~n3758 ;
  buffer buf_n3760( .i (n3146), .o (n3760) );
  assign n3761 = ( ~n1874 & n2988 ) | ( ~n1874 & n3760 ) | ( n2988 & n3760 ) ;
  buffer buf_n3762( .i (n3761), .o (n3762) );
  buffer buf_n3763( .i (n3762), .o (n3763) );
  buffer buf_n3764( .i (n3763), .o (n3764) );
  buffer buf_n3765( .i (n3340), .o (n3765) );
  assign n3766 = ( ~n3665 & n3762 ) | ( ~n3665 & n3765 ) | ( n3762 & n3765 ) ;
  assign n3767 = n1877 | n3766 ;
  buffer buf_n3768( .i (n2990), .o (n3768) );
  buffer buf_n3769( .i (n3768), .o (n3769) );
  assign n3770 = ( n3764 & n3767 ) | ( n3764 & ~n3769 ) | ( n3767 & ~n3769 ) ;
  assign n3771 = n3275 & n3770 ;
  assign n3772 = ( ~n3262 & n3339 ) | ( ~n3262 & n3760 ) | ( n3339 & n3760 ) ;
  buffer buf_n3773( .i (n3772), .o (n3773) );
  buffer buf_n3774( .i (n3773), .o (n3774) );
  buffer buf_n3780( .i (n3262), .o (n3780) );
  buffer buf_n3781( .i (n3780), .o (n3781) );
  assign n3782 = n3773 & n3781 ;
  assign n3783 = ( ~n2629 & n3774 ) | ( ~n2629 & n3782 ) | ( n3774 & n3782 ) ;
  assign n3784 = ~n3769 & n3783 ;
  buffer buf_n3785( .i (n3137), .o (n3785) );
  assign n3786 = n3784 | n3785 ;
  assign n3787 = ~n3771 & n3786 ;
  assign n3788 = n3392 | n3787 ;
  buffer buf_n3789( .i (n2988), .o (n3789) );
  assign n3790 = ( ~n2627 & n3071 ) | ( ~n2627 & n3789 ) | ( n3071 & n3789 ) ;
  buffer buf_n3791( .i (n3790), .o (n3791) );
  buffer buf_n3792( .i (n3791), .o (n3792) );
  buffer buf_n3793( .i (n3792), .o (n3793) );
  buffer buf_n3794( .i (n3665), .o (n3794) );
  assign n3795 = ( ~n3768 & n3791 ) | ( ~n3768 & n3794 ) | ( n3791 & n3794 ) ;
  assign n3796 = ( ~n3137 & n3443 ) | ( ~n3137 & n3795 ) | ( n3443 & n3795 ) ;
  assign n3797 = n3793 & n3796 ;
  assign n3798 = ~n2950 & n3797 ;
  buffer buf_n3799( .i (n3617), .o (n3799) );
  assign n3800 = ~n3798 & n3799 ;
  assign n3801 = n3788 & ~n3800 ;
  assign n3802 = n2824 | n3801 ;
  buffer buf_n3803( .i (n2824), .o (n3803) );
  assign n3804 = ( n3759 & n3802 ) | ( n3759 & ~n3803 ) | ( n3802 & ~n3803 ) ;
  assign n3805 = ~n3398 & n3804 ;
  assign n3806 = n3485 & ~n3805 ;
  assign n3807 = n3731 & ~n3806 ;
  assign n3808 = n3598 | n3807 ;
  assign n3809 = ( ~n3546 & n3547 ) | ( ~n3546 & n3808 ) | ( n3547 & n3808 ) ;
  buffer buf_n3810( .i (n3809), .o (n3810) );
  buffer buf_n3811( .i (n3810), .o (n3811) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n3812( .i (n3789), .o (n3812) );
  assign n3813 = ~n24 & n3812 ;
  buffer buf_n3814( .i (n3813), .o (n3814) );
  buffer buf_n3815( .i (n3814), .o (n3815) );
  buffer buf_n3816( .i (n3815), .o (n3816) );
  buffer buf_n3817( .i (n3816), .o (n3817) );
  buffer buf_n3818( .i (n3817), .o (n3818) );
  buffer buf_n3819( .i (n3818), .o (n3819) );
  buffer buf_n3820( .i (n3819), .o (n3820) );
  assign n3822 = ~n2534 & n3375 ;
  assign n3823 = ( ~n964 & n3820 ) | ( ~n964 & n3822 ) | ( n3820 & n3822 ) ;
  assign n3824 = n2019 | n3823 ;
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  assign n3825 = ~n3425 & n3503 ;
  buffer buf_n3826( .i (n3825), .o (n3826) );
  buffer buf_n3827( .i (n3826), .o (n3827) );
  buffer buf_n3828( .i (n3827), .o (n3828) );
  buffer buf_n3829( .i (n3828), .o (n3829) );
  buffer buf_n3830( .i (n3829), .o (n3830) );
  assign n3831 = ( n1317 & n3819 ) | ( n1317 & ~n3830 ) | ( n3819 & ~n3830 ) ;
  assign n3832 = ~n2535 & n3831 ;
  assign n3833 = n2019 & ~n3832 ;
  assign n3834 = n3824 & ~n3833 ;
  buffer buf_n3835( .i (n3485), .o (n3835) );
  assign n3836 = n3834 | n3835 ;
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n2013( .i (n2012), .o (n2013) );
  assign n3837 = ~n2013 & n3803 ;
  assign n3838 = ( n520 & n806 ) | ( n520 & ~n3837 ) | ( n806 & ~n3837 ) ;
  buffer buf_n3839( .i (n3398), .o (n3839) );
  assign n3840 = n3838 & ~n3839 ;
  assign n3841 = n3835 & ~n3840 ;
  assign n3842 = n3836 & ~n3841 ;
  assign n3843 = n3489 | n3842 ;
  buffer buf_n2014( .i (n2013), .o (n2014) );
  buffer buf_n2015( .i (n2014), .o (n2015) );
  buffer buf_n2723( .i (n2722), .o (n2723) );
  buffer buf_n2724( .i (n2723), .o (n2724) );
  buffer buf_n2725( .i (n2724), .o (n2725) );
  buffer buf_n2726( .i (n2725), .o (n2726) );
  buffer buf_n3844( .i (n3297), .o (n3844) );
  assign n3845 = ( ~n2726 & n2793 ) | ( ~n2726 & n3844 ) | ( n2793 & n3844 ) ;
  assign n3846 = ( ~n2726 & n3460 ) | ( ~n2726 & n3844 ) | ( n3460 & n3844 ) ;
  assign n3847 = ( n2015 & n3845 ) | ( n2015 & ~n3846 ) | ( n3845 & ~n3846 ) ;
  buffer buf_n3848( .i (n2559), .o (n3848) );
  assign n3849 = n375 & ~n3848 ;
  buffer buf_n3850( .i (n3849), .o (n3850) );
  assign n3851 = n1951 & n3850 ;
  buffer buf_n3852( .i (n3851), .o (n3852) );
  buffer buf_n3853( .i (n3852), .o (n3853) );
  buffer buf_n3854( .i (n3803), .o (n3854) );
  buffer buf_n3855( .i (n3854), .o (n3855) );
  assign n3856 = n3852 | n3855 ;
  assign n3857 = ( n3847 & n3853 ) | ( n3847 & n3856 ) | ( n3853 & n3856 ) ;
  assign n3858 = ~n3111 & n3857 ;
  assign n3859 = n3489 & ~n3858 ;
  assign n3860 = n3843 & ~n3859 ;
  assign n3861 = n3810 | n3860 ;
  assign n3862 = ( n361 & n3811 ) | ( n361 & n3861 ) | ( n3811 & n3861 ) ;
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n3863( .i (n3043), .o (n3863) );
  assign n3864 = n3789 | n3863 ;
  buffer buf_n3865( .i (n3864), .o (n3865) );
  buffer buf_n3866( .i (n3865), .o (n3866) );
  buffer buf_n3867( .i (n3866), .o (n3867) );
  buffer buf_n3868( .i (n3867), .o (n3868) );
  buffer buf_n3869( .i (n3868), .o (n3869) );
  buffer buf_n3870( .i (n3869), .o (n3870) );
  buffer buf_n3871( .i (n3870), .o (n3871) );
  buffer buf_n3872( .i (n3871), .o (n3872) );
  assign n3873 = ( ~n1087 & n1436 ) | ( ~n1087 & n3872 ) | ( n1436 & n3872 ) ;
  assign n3874 = n3844 & ~n3873 ;
  assign n3875 = ~n3839 & n3874 ;
  buffer buf_n3876( .i (n3875), .o (n3876) );
  buffer buf_n3877( .i (n3876), .o (n3877) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  assign n3878 = ( n711 & n1812 ) | ( n711 & n3423 ) | ( n1812 & n3423 ) ;
  assign n3879 = ~n2640 & n3878 ;
  buffer buf_n3507( .i (n3506), .o (n3507) );
  buffer buf_n3508( .i (n3507), .o (n3508) );
  buffer buf_n3509( .i (n3508), .o (n3509) );
  assign n3880 = ~n308 & n3504 ;
  assign n3881 = ( n3255 & n3444 ) | ( n3255 & n3880 ) | ( n3444 & n3880 ) ;
  buffer buf_n3882( .i (n3443), .o (n3882) );
  buffer buf_n3883( .i (n3882), .o (n3883) );
  assign n3884 = n3881 & ~n3883 ;
  buffer buf_n3885( .i (n3884), .o (n3885) );
  buffer buf_n3886( .i (n3885), .o (n3886) );
  buffer buf_n748( .i (n747), .o (n748) );
  assign n3887 = n748 | n3885 ;
  assign n3888 = ( n3509 & n3886 ) | ( n3509 & n3887 ) | ( n3886 & n3887 ) ;
  buffer buf_n3889( .i (n3888), .o (n3889) );
  buffer buf_n3890( .i (n3889), .o (n3890) );
  buffer buf_n3891( .i (n3451), .o (n3891) );
  assign n3892 = n3889 & n3891 ;
  buffer buf_n3893( .i (n2577), .o (n3893) );
  assign n3894 = n1402 & ~n3893 ;
  assign n3895 = ~n2100 & n3894 ;
  buffer buf_n3896( .i (n3339), .o (n3896) );
  assign n3897 = ( n3465 & n3863 ) | ( n3465 & ~n3896 ) | ( n3863 & ~n3896 ) ;
  assign n3898 = ( ~n3465 & n3789 ) | ( ~n3465 & n3863 ) | ( n3789 & n3863 ) ;
  assign n3899 = n3897 & ~n3898 ;
  assign n3900 = ( n3425 & n3752 ) | ( n3425 & n3899 ) | ( n3752 & n3899 ) ;
  assign n3901 = n21 & n3463 ;
  buffer buf_n3902( .i (n3901), .o (n3902) );
  buffer buf_n3907( .i (n2988), .o (n3907) );
  assign n3908 = ( ~n2091 & n3902 ) | ( ~n2091 & n3907 ) | ( n3902 & n3907 ) ;
  assign n3909 = ~n3812 & n3908 ;
  assign n3910 = n3752 & n3909 ;
  buffer buf_n3911( .i (n20), .o (n3911) );
  buffer buf_n3912( .i (n3911), .o (n3912) );
  buffer buf_n3913( .i (n3912), .o (n3913) );
  buffer buf_n3914( .i (n3913), .o (n3914) );
  buffer buf_n3915( .i (n3914), .o (n3915) );
  buffer buf_n3916( .i (n3915), .o (n3916) );
  assign n3917 = ( n3900 & n3910 ) | ( n3900 & ~n3916 ) | ( n3910 & ~n3916 ) ;
  buffer buf_n3918( .i (n3917), .o (n3918) );
  buffer buf_n3919( .i (n3918), .o (n3919) );
  buffer buf_n3920( .i (n3919), .o (n3920) );
  buffer buf_n3921( .i (n3061), .o (n3921) );
  assign n3922 = ( n2762 & ~n3201 ) | ( n2762 & n3921 ) | ( ~n3201 & n3921 ) ;
  buffer buf_n3923( .i (n3922), .o (n3923) );
  buffer buf_n3924( .i (n3923), .o (n3924) );
  buffer buf_n3925( .i (n3924), .o (n3925) );
  buffer buf_n3926( .i (n3925), .o (n3926) );
  buffer buf_n3927( .i (n3926), .o (n3927) );
  buffer buf_n3928( .i (n3927), .o (n3928) );
  assign n3929 = ( n3215 & n3254 ) | ( n3215 & ~n3504 ) | ( n3254 & ~n3504 ) ;
  assign n3930 = n3928 & ~n3929 ;
  assign n3931 = ( ~n3511 & n3918 ) | ( ~n3511 & n3930 ) | ( n3918 & n3930 ) ;
  assign n3932 = n3620 & ~n3931 ;
  assign n3933 = ( n3535 & n3920 ) | ( n3535 & ~n3932 ) | ( n3920 & ~n3932 ) ;
  assign n3934 = n3395 | n3933 ;
  assign n3935 = ( n1739 & n2950 ) | ( n1739 & ~n3619 ) | ( n2950 & ~n3619 ) ;
  assign n3936 = n1868 & n3935 ;
  assign n3937 = ~n3436 & n3936 ;
  assign n3938 = n3395 & ~n3937 ;
  assign n3939 = n3934 & ~n3938 ;
  assign n3940 = n3895 | n3939 ;
  assign n3941 = ( n3890 & ~n3892 ) | ( n3890 & n3940 ) | ( ~n3892 & n3940 ) ;
  buffer buf_n3942( .i (n3941), .o (n3942) );
  assign n3943 = ( ~n3876 & n3879 ) | ( ~n3876 & n3942 ) | ( n3879 & n3942 ) ;
  assign n3944 = n357 & ~n3942 ;
  assign n3945 = ( n3877 & n3943 ) | ( n3877 & ~n3944 ) | ( n3943 & ~n3944 ) ;
  buffer buf_n3946( .i (n3945), .o (n3946) );
  buffer buf_n3947( .i (n3946), .o (n3947) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  assign n3948 = n123 & n3946 ;
  assign n3949 = ( n3132 & n3635 ) | ( n3132 & n3812 ) | ( n3635 & n3812 ) ;
  buffer buf_n3950( .i (n3949), .o (n3950) );
  buffer buf_n3951( .i (n3950), .o (n3951) );
  buffer buf_n3952( .i (n3951), .o (n3952) );
  buffer buf_n3957( .i (n3177), .o (n3957) );
  assign n3958 = ( n2558 & ~n3952 ) | ( n2558 & n3957 ) | ( ~n3952 & n3957 ) ;
  buffer buf_n3959( .i (n3958), .o (n3959) );
  buffer buf_n3960( .i (n3959), .o (n3960) );
  buffer buf_n3961( .i (n3960), .o (n3961) );
  buffer buf_n3962( .i (n3961), .o (n3962) );
  buffer buf_n3963( .i (n3437), .o (n3963) );
  buffer buf_n3964( .i (n3799), .o (n3964) );
  assign n3965 = ( ~n3959 & n3963 ) | ( ~n3959 & n3964 ) | ( n3963 & n3964 ) ;
  buffer buf_n3966( .i (n3965), .o (n3966) );
  buffer buf_n3967( .i (n3966), .o (n3967) );
  buffer buf_n3953( .i (n3952), .o (n3953) );
  buffer buf_n3954( .i (n3953), .o (n3954) );
  buffer buf_n3955( .i (n3954), .o (n3955) );
  buffer buf_n3956( .i (n3955), .o (n3956) );
  assign n3968 = n3956 & ~n3966 ;
  assign n3969 = ( n3962 & n3967 ) | ( n3962 & ~n3968 ) | ( n3967 & ~n3968 ) ;
  assign n3970 = ( ~n236 & n264 ) | ( ~n236 & n3969 ) | ( n264 & n3969 ) ;
  assign n3971 = ~n3535 & n3848 ;
  buffer buf_n3972( .i (n3971), .o (n3972) );
  assign n3973 = ( n1551 & n3459 ) | ( n1551 & n3972 ) | ( n3459 & n3972 ) ;
  buffer buf_n3974( .i (n3963), .o (n3974) );
  buffer buf_n3975( .i (n3974), .o (n3975) );
  buffer buf_n3976( .i (n3893), .o (n3976) );
  assign n3977 = ( n3972 & n3975 ) | ( n3972 & n3976 ) | ( n3975 & n3976 ) ;
  assign n3978 = ( n1952 & n3973 ) | ( n1952 & ~n3977 ) | ( n3973 & ~n3977 ) ;
  assign n3979 = ( n236 & n264 ) | ( n236 & ~n3978 ) | ( n264 & ~n3978 ) ;
  assign n3980 = n3970 | n3979 ;
  buffer buf_n3981( .i (n3980), .o (n3981) );
  buffer buf_n3982( .i (n3981), .o (n3982) );
  buffer buf_n3093( .i (n3092), .o (n3093) );
  assign n3983 = ( n3093 & ~n3459 ) | ( n3093 & n3976 ) | ( ~n3459 & n3976 ) ;
  assign n3984 = ( ~n3093 & n3803 ) | ( ~n3093 & n3976 ) | ( n3803 & n3976 ) ;
  assign n3985 = n3983 & ~n3984 ;
  buffer buf_n3986( .i (n3985), .o (n3986) );
  buffer buf_n3987( .i (n3986), .o (n3987) );
  assign n3988 = ( n265 & n3835 ) | ( n265 & ~n3986 ) | ( n3835 & ~n3986 ) ;
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  assign n3989 = ( ~n628 & n2793 ) | ( ~n628 & n3460 ) | ( n2793 & n3460 ) ;
  buffer buf_n3990( .i (n3976), .o (n3990) );
  assign n3991 = ( n628 & ~n3844 ) | ( n628 & n3990 ) | ( ~n3844 & n3990 ) ;
  assign n3992 = n3989 & ~n3991 ;
  assign n3993 = n265 & n3992 ;
  assign n3994 = ( n3987 & n3988 ) | ( n3987 & n3993 ) | ( n3988 & n3993 ) ;
  assign n3995 = n3981 & n3994 ;
  assign n3996 = n3609 & ~n3915 ;
  buffer buf_n3997( .i (n3996), .o (n3997) );
  buffer buf_n3998( .i (n3997), .o (n3998) );
  buffer buf_n3999( .i (n3998), .o (n3999) );
  buffer buf_n4000( .i (n3999), .o (n4000) );
  buffer buf_n4001( .i (n4000), .o (n4001) );
  buffer buf_n4002( .i (n4001), .o (n4002) );
  buffer buf_n4003( .i (n4002), .o (n4003) );
  buffer buf_n4004( .i (n4003), .o (n4004) );
  buffer buf_n4005( .i (n4004), .o (n4005) );
  buffer buf_n4006( .i (n4005), .o (n4006) );
  buffer buf_n4007( .i (n4006), .o (n4007) );
  buffer buf_n4008( .i (n4007), .o (n4008) );
  assign n4009 = ( ~n3982 & n3995 ) | ( ~n3982 & n4008 ) | ( n3995 & n4008 ) ;
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  buffer buf_n2250( .i (n2249), .o (n2250) );
  buffer buf_n4010( .i (n3429), .o (n4010) );
  assign n4011 = ( n398 & n2198 ) | ( n398 & ~n4010 ) | ( n2198 & ~n4010 ) ;
  buffer buf_n3165( .i (n3164), .o (n3165) );
  assign n4012 = n3165 & n4010 ;
  assign n4013 = ( n399 & ~n4011 ) | ( n399 & n4012 ) | ( ~n4011 & n4012 ) ;
  buffer buf_n4014( .i (n3620), .o (n4014) );
  assign n4015 = ( n3436 & n4013 ) | ( n3436 & ~n4014 ) | ( n4013 & ~n4014 ) ;
  assign n4016 = n1938 | n2899 ;
  buffer buf_n4017( .i (n4016), .o (n4017) );
  buffer buf_n4018( .i (n4017), .o (n4018) );
  buffer buf_n4019( .i (n4018), .o (n4019) );
  assign n4026 = n3916 & ~n4019 ;
  buffer buf_n4027( .i (n4026), .o (n4027) );
  assign n4034 = n2237 & n3337 ;
  buffer buf_n4035( .i (n4034), .o (n4035) );
  buffer buf_n4036( .i (n4035), .o (n4036) );
  buffer buf_n4037( .i (n4036), .o (n4037) );
  buffer buf_n4038( .i (n4037), .o (n4038) );
  buffer buf_n4039( .i (n4038), .o (n4039) );
  assign n4040 = n4027 & n4039 ;
  buffer buf_n4041( .i (n4040), .o (n4041) );
  assign n4048 = ~n4014 & n4041 ;
  buffer buf_n4049( .i (n3435), .o (n4049) );
  buffer buf_n4050( .i (n4049), .o (n4050) );
  assign n4051 = ( n4015 & n4048 ) | ( n4015 & ~n4050 ) | ( n4048 & ~n4050 ) ;
  buffer buf_n4052( .i (n4051), .o (n4052) );
  buffer buf_n4053( .i (n4052), .o (n4053) );
  buffer buf_n4054( .i (n4053), .o (n4054) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  assign n4055 = ( n758 & n1065 ) | ( n758 & n4052 ) | ( n1065 & n4052 ) ;
  assign n4056 = n2249 & ~n4055 ;
  assign n4057 = ( n2250 & n4054 ) | ( n2250 & ~n4056 ) | ( n4054 & ~n4056 ) ;
  buffer buf_n4058( .i (n4057), .o (n4058) );
  buffer buf_n4059( .i (n4058), .o (n4059) );
  assign n4060 = n358 & n4058 ;
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  assign n4061 = n715 & ~n1762 ;
  assign n4062 = n805 & n4061 ;
  buffer buf_n4063( .i (n4062), .o (n4063) );
  buffer buf_n4064( .i (n4063), .o (n4064) );
  buffer buf_n4065( .i (n4064), .o (n4065) );
  buffer buf_n4066( .i (n3503), .o (n4066) );
  assign n4067 = n2241 & ~n4066 ;
  buffer buf_n4068( .i (n4067), .o (n4068) );
  assign n4070 = ( n1154 & n4010 ) | ( n1154 & n4068 ) | ( n4010 & n4068 ) ;
  assign n4071 = ~n3437 & n4070 ;
  buffer buf_n4072( .i (n4071), .o (n4072) );
  buffer buf_n4073( .i (n4072), .o (n4073) );
  buffer buf_n4074( .i (n4073), .o (n4074) );
  buffer buf_n4075( .i (n828), .o (n4075) );
  buffer buf_n4076( .i (n4075), .o (n4076) );
  assign n4077 = ( ~n3071 & n3338 ) | ( ~n3071 & n4076 ) | ( n3338 & n4076 ) ;
  buffer buf_n4078( .i (n4077), .o (n4078) );
  assign n4083 = ( n3140 & n3673 ) | ( n3140 & ~n4078 ) | ( n3673 & ~n4078 ) ;
  buffer buf_n4084( .i (n4083), .o (n4084) );
  buffer buf_n4085( .i (n4084), .o (n4085) );
  buffer buf_n4086( .i (n4085), .o (n4086) );
  buffer buf_n4087( .i (n4086), .o (n4087) );
  buffer buf_n4088( .i (n4066), .o (n4088) );
  assign n4089 = ( n3785 & n4084 ) | ( n3785 & ~n4088 ) | ( n4084 & ~n4088 ) ;
  buffer buf_n4090( .i (n4089), .o (n4090) );
  buffer buf_n4091( .i (n4090), .o (n4091) );
  buffer buf_n4079( .i (n4078), .o (n4079) );
  buffer buf_n4080( .i (n4079), .o (n4080) );
  buffer buf_n4081( .i (n4080), .o (n4081) );
  buffer buf_n4082( .i (n4081), .o (n4082) );
  assign n4092 = n4082 | n4090 ;
  assign n4093 = ( ~n4087 & n4091 ) | ( ~n4087 & n4092 ) | ( n4091 & n4092 ) ;
  buffer buf_n4094( .i (n4014), .o (n4094) );
  assign n4095 = ( ~n4072 & n4093 ) | ( ~n4072 & n4094 ) | ( n4093 & n4094 ) ;
  buffer buf_n4096( .i (n2534), .o (n4096) );
  assign n4097 = n4095 & ~n4096 ;
  assign n4098 = ( n3421 & ~n4074 ) | ( n3421 & n4097 ) | ( ~n4074 & n4097 ) ;
  assign n4099 = ( n3839 & ~n4063 ) | ( n3839 & n4098 ) | ( ~n4063 & n4098 ) ;
  assign n4100 = n265 & n4099 ;
  assign n4101 = ( n266 & n4065 ) | ( n266 & ~n4100 ) | ( n4065 & ~n4100 ) ;
  buffer buf_n4102( .i (n4076), .o (n4102) );
  assign n4103 = ~n1943 & n4102 ;
  buffer buf_n4104( .i (n4103), .o (n4104) );
  assign n4105 = n1764 & n4104 ;
  assign n4106 = n3118 & ~n3635 ;
  buffer buf_n4107( .i (n4106), .o (n4107) );
  assign n4112 = ( ~n1945 & n4104 ) | ( ~n1945 & n4107 ) | ( n4104 & n4107 ) ;
  buffer buf_n4113( .i (n3769), .o (n4113) );
  assign n4114 = ( n4105 & n4112 ) | ( n4105 & ~n4113 ) | ( n4112 & ~n4113 ) ;
  buffer buf_n4115( .i (n4114), .o (n4115) );
  buffer buf_n4116( .i (n4115), .o (n4116) );
  assign n4117 = ( n1560 & n2460 ) | ( n1560 & ~n2782 ) | ( n2460 & ~n2782 ) ;
  buffer buf_n4118( .i (n4117), .o (n4118) );
  buffer buf_n4119( .i (n4118), .o (n4119) );
  buffer buf_n4120( .i (n4119), .o (n4120) );
  buffer buf_n4121( .i (n4120), .o (n4121) );
  assign n4126 = n4115 & n4121 ;
  assign n4127 = ( n71 & n99 ) | ( n71 & n159 ) | ( n99 & n159 ) ;
  buffer buf_n4128( .i (n4127), .o (n4128) );
  assign n4138 = ( n101 & ~n131 ) | ( n101 & n4128 ) | ( ~n131 & n4128 ) ;
  buffer buf_n4139( .i (n4138), .o (n4139) );
  assign n4142 = n2910 & ~n4139 ;
  buffer buf_n4143( .i (n4142), .o (n4143) );
  buffer buf_n4144( .i (n4143), .o (n4144) );
  buffer buf_n4140( .i (n4139), .o (n4140) );
  buffer buf_n4141( .i (n4140), .o (n4141) );
  assign n4145 = n4141 | n4143 ;
  assign n4146 = ( ~n2899 & n4144 ) | ( ~n2899 & n4145 ) | ( n4144 & n4145 ) ;
  assign n4147 = ( ~n3780 & n4076 ) | ( ~n3780 & n4146 ) | ( n4076 & n4146 ) ;
  buffer buf_n4148( .i (n4147), .o (n4148) );
  buffer buf_n4149( .i (n4148), .o (n4149) );
  buffer buf_n4150( .i (n4149), .o (n4150) );
  buffer buf_n4151( .i (n4150), .o (n4151) );
  assign n4152 = n3752 & n4148 ;
  buffer buf_n4153( .i (n4152), .o (n4153) );
  buffer buf_n4154( .i (n4153), .o (n4154) );
  assign n4155 = ( n3255 & n3429 ) | ( n3255 & ~n4153 ) | ( n3429 & ~n4153 ) ;
  assign n4156 = ( n4151 & n4154 ) | ( n4151 & ~n4155 ) | ( n4154 & ~n4155 ) ;
  assign n4157 = ( n71 & n99 ) | ( n71 & ~n129 ) | ( n99 & ~n129 ) ;
  buffer buf_n4158( .i (n4157), .o (n4158) );
  buffer buf_n4173( .i (n129), .o (n4173) );
  buffer buf_n4174( .i (n4173), .o (n4174) );
  assign n4175 = ( n3677 & n4158 ) | ( n3677 & n4174 ) | ( n4158 & n4174 ) ;
  buffer buf_n4176( .i (n4175), .o (n4176) );
  buffer buf_n4177( .i (n4176), .o (n4177) );
  buffer buf_n4178( .i (n4177), .o (n4178) );
  buffer buf_n4179( .i (n4178), .o (n4179) );
  assign n4180 = ( n2910 & n3732 ) | ( n2910 & n4176 ) | ( n3732 & n4176 ) ;
  buffer buf_n4181( .i (n4180), .o (n4181) );
  buffer buf_n4182( .i (n4181), .o (n4182) );
  buffer buf_n4159( .i (n4158), .o (n4159) );
  buffer buf_n4160( .i (n4159), .o (n4160) );
  buffer buf_n4161( .i (n4160), .o (n4161) );
  buffer buf_n4162( .i (n4161), .o (n4162) );
  assign n4183 = ~n4162 & n4181 ;
  assign n4184 = ( ~n4179 & n4182 ) | ( ~n4179 & n4183 ) | ( n4182 & n4183 ) ;
  buffer buf_n4185( .i (n3760), .o (n4185) );
  assign n4186 = ~n4184 & n4185 ;
  buffer buf_n4187( .i (n2854), .o (n4187) );
  assign n4188 = n1733 & ~n4187 ;
  assign n4189 = n4185 | n4188 ;
  assign n4190 = ~n4186 & n4189 ;
  buffer buf_n4191( .i (n4102), .o (n4191) );
  assign n4192 = n4190 | n4191 ;
  assign n4193 = ~n584 & n4035 ;
  assign n4194 = n4191 & ~n4193 ;
  assign n4195 = n4192 & ~n4194 ;
  assign n4196 = ~n3744 & n4195 ;
  assign n4197 = ( n769 & n2329 ) | ( n769 & n2888 ) | ( n2329 & n2888 ) ;
  buffer buf_n4198( .i (n4197), .o (n4198) );
  buffer buf_n4199( .i (n4198), .o (n4199) );
  buffer buf_n4200( .i (n4199), .o (n4200) );
  buffer buf_n4201( .i (n2911), .o (n4201) );
  assign n4202 = ( n3921 & ~n4198 ) | ( n3921 & n4201 ) | ( ~n4198 & n4201 ) ;
  assign n4203 = n772 | n4202 ;
  buffer buf_n4204( .i (n3733), .o (n4204) );
  buffer buf_n4205( .i (n4204), .o (n4205) );
  assign n4206 = ( ~n4200 & n4203 ) | ( ~n4200 & n4205 ) | ( n4203 & n4205 ) ;
  buffer buf_n4207( .i (n4206), .o (n4207) );
  buffer buf_n4208( .i (n4207), .o (n4208) );
  buffer buf_n4209( .i (n4187), .o (n4209) );
  buffer buf_n4210( .i (n4209), .o (n4210) );
  assign n4211 = ( ~n4102 & n4207 ) | ( ~n4102 & n4210 ) | ( n4207 & n4210 ) ;
  assign n4212 = n1687 & ~n2193 ;
  assign n4213 = ~n4102 & n4212 ;
  assign n4214 = ( ~n4208 & n4211 ) | ( ~n4208 & n4213 ) | ( n4211 & n4213 ) ;
  buffer buf_n4215( .i (n100), .o (n4215) );
  assign n4216 = n3677 & n4215 ;
  buffer buf_n4217( .i (n4216), .o (n4217) );
  buffer buf_n4218( .i (n4217), .o (n4218) );
  buffer buf_n4219( .i (n4218), .o (n4219) );
  buffer buf_n4231( .i (n4201), .o (n4231) );
  assign n4232 = ( ~n4204 & n4219 ) | ( ~n4204 & n4231 ) | ( n4219 & n4231 ) ;
  assign n4233 = ( n3921 & n4201 ) | ( n3921 & ~n4218 ) | ( n4201 & ~n4218 ) ;
  buffer buf_n4234( .i (n2853), .o (n4234) );
  assign n4235 = ( ~n4204 & n4233 ) | ( ~n4204 & n4234 ) | ( n4233 & n4234 ) ;
  assign n4236 = ~n4232 & n4235 ;
  buffer buf_n4237( .i (n4236), .o (n4237) );
  buffer buf_n4238( .i (n4237), .o (n4238) );
  buffer buf_n4239( .i (n4076), .o (n4239) );
  assign n4240 = ( n3635 & n4237 ) | ( n3635 & ~n4239 ) | ( n4237 & ~n4239 ) ;
  buffer buf_n2879( .i (n2878), .o (n2879) );
  buffer buf_n2880( .i (n2879), .o (n2880) );
  assign n4241 = ( n2190 & n2880 ) | ( n2190 & ~n4201 ) | ( n2880 & ~n4201 ) ;
  buffer buf_n4242( .i (n4241), .o (n4242) );
  buffer buf_n4243( .i (n4242), .o (n4243) );
  assign n4261 = ( n392 & n4205 ) | ( n392 & n4242 ) | ( n4205 & n4242 ) ;
  assign n4262 = ~n4243 & n4261 ;
  assign n4263 = n4239 & n4262 ;
  assign n4264 = ( n4238 & ~n4240 ) | ( n4238 & n4263 ) | ( ~n4240 & n4263 ) ;
  assign n4265 = n4214 | n4264 ;
  assign n4266 = n3744 & n4265 ;
  assign n4267 = n4196 | n4266 ;
  assign n4268 = n4156 | n4267 ;
  assign n4269 = ( n4116 & ~n4126 ) | ( n4116 & n4268 ) | ( ~n4126 & n4268 ) ;
  assign n4270 = ( n233 & ~n4050 ) | ( n233 & n4269 ) | ( ~n4050 & n4269 ) ;
  assign n4271 = ( n44 & n100 ) | ( n44 & n2231 ) | ( n100 & n2231 ) ;
  buffer buf_n4272( .i (n4271), .o (n4272) );
  assign n4285 = ( n2233 & n3187 ) | ( n2233 & ~n4272 ) | ( n3187 & ~n4272 ) ;
  buffer buf_n4286( .i (n4285), .o (n4286) );
  buffer buf_n4287( .i (n4286), .o (n4287) );
  buffer buf_n4273( .i (n4272), .o (n4273) );
  buffer buf_n4274( .i (n4273), .o (n4274) );
  buffer buf_n4288( .i (n2911), .o (n4288) );
  assign n4289 = ( n4274 & n4286 ) | ( n4274 & ~n4288 ) | ( n4286 & ~n4288 ) ;
  assign n4290 = ( ~n4234 & n4287 ) | ( ~n4234 & n4289 ) | ( n4287 & n4289 ) ;
  buffer buf_n4291( .i (n4290), .o (n4291) );
  buffer buf_n4292( .i (n4291), .o (n4292) );
  assign n4293 = ( n3780 & ~n3907 ) | ( n3780 & n4291 ) | ( ~n3907 & n4291 ) ;
  assign n4294 = n302 | n3921 ;
  assign n4295 = ( n4231 & n4234 ) | ( n4231 & ~n4294 ) | ( n4234 & ~n4294 ) ;
  assign n4296 = ~n4187 & n4295 ;
  assign n4297 = ~n3780 & n4296 ;
  assign n4298 = ( n4292 & ~n4293 ) | ( n4292 & n4297 ) | ( ~n4293 & n4297 ) ;
  buffer buf_n4299( .i (n4298), .o (n4299) );
  buffer buf_n4300( .i (n4299), .o (n4300) );
  buffer buf_n4301( .i (n4300), .o (n4301) );
  buffer buf_n4302( .i (n4191), .o (n4302) );
  assign n4303 = ( n3667 & n4299 ) | ( n3667 & ~n4302 ) | ( n4299 & ~n4302 ) ;
  assign n4304 = n2934 & ~n4303 ;
  assign n4305 = ( n2935 & n4301 ) | ( n2935 & ~n4304 ) | ( n4301 & ~n4304 ) ;
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n4306( .i (n2330), .o (n4306) );
  buffer buf_n4307( .i (n4306), .o (n4307) );
  buffer buf_n4308( .i (n4307), .o (n4308) );
  buffer buf_n4309( .i (n4308), .o (n4309) );
  assign n4310 = ( ~n3005 & n4187 ) | ( ~n3005 & n4309 ) | ( n4187 & n4309 ) ;
  buffer buf_n4311( .i (n4234), .o (n4311) );
  assign n4312 = ( ~n3005 & n3760 ) | ( ~n3005 & n4311 ) | ( n3760 & n4311 ) ;
  assign n4313 = ( n2303 & n4310 ) | ( n2303 & ~n4312 ) | ( n4310 & ~n4312 ) ;
  assign n4314 = ( n3631 & n3812 ) | ( n3631 & n4313 ) | ( n3812 & n4313 ) ;
  buffer buf_n4315( .i (n4314), .o (n4315) );
  assign n4316 = ( ~n3769 & n4302 ) | ( ~n3769 & n4315 ) | ( n4302 & n4315 ) ;
  assign n4317 = ( n3254 & n4302 ) | ( n3254 & ~n4315 ) | ( n4302 & ~n4315 ) ;
  assign n4318 = n4316 & ~n4317 ;
  buffer buf_n4319( .i (n4318), .o (n4319) );
  assign n4320 = ( ~n3799 & n4305 ) | ( ~n3799 & n4319 ) | ( n4305 & n4319 ) ;
  buffer buf_n2881( .i (n2880), .o (n2881) );
  buffer buf_n2882( .i (n2881), .o (n2882) );
  buffer buf_n2883( .i (n2882), .o (n2883) );
  buffer buf_n2884( .i (n2883), .o (n2884) );
  buffer buf_n2885( .i (n2884), .o (n2885) );
  buffer buf_n2886( .i (n2885), .o (n2886) );
  assign n4321 = ( n3609 & ~n3673 ) | ( n3609 & n3865 ) | ( ~n3673 & n3865 ) ;
  assign n4322 = ( n3609 & ~n3794 ) | ( n3609 & n3865 ) | ( ~n3794 & n3865 ) ;
  assign n4323 = ( n2886 & ~n4321 ) | ( n2886 & n4322 ) | ( ~n4321 & n4322 ) ;
  buffer buf_n4324( .i (n4075), .o (n4324) );
  buffer buf_n4325( .i (n4309), .o (n4325) );
  assign n4326 = n4324 & n4325 ;
  buffer buf_n4327( .i (n4326), .o (n4327) );
  buffer buf_n4332( .i (n3781), .o (n4332) );
  assign n4333 = ~n4327 & n4332 ;
  buffer buf_n4334( .i (n4333), .o (n4334) );
  assign n4335 = n4323 & n4334 ;
  buffer buf_n4328( .i (n4327), .o (n4328) );
  buffer buf_n4329( .i (n4328), .o (n4329) );
  buffer buf_n4129( .i (n4128), .o (n4129) );
  buffer buf_n4130( .i (n4129), .o (n4130) );
  buffer buf_n4131( .i (n4130), .o (n4131) );
  buffer buf_n4132( .i (n4131), .o (n4132) );
  buffer buf_n4133( .i (n4132), .o (n4133) );
  buffer buf_n4134( .i (n4133), .o (n4134) );
  buffer buf_n4135( .i (n4134), .o (n4135) );
  buffer buf_n4136( .i (n4135), .o (n4136) );
  buffer buf_n4137( .i (n4136), .o (n4137) );
  buffer buf_n4336( .i (n3631), .o (n4336) );
  assign n4337 = ( n3768 & n3794 ) | ( n3768 & n4336 ) | ( n3794 & n4336 ) ;
  buffer buf_n4338( .i (n3863), .o (n4338) );
  assign n4339 = ~n4210 & n4338 ;
  buffer buf_n4340( .i (n4339), .o (n4340) );
  assign n4350 = ( n4137 & ~n4337 ) | ( n4137 & n4340 ) | ( ~n4337 & n4340 ) ;
  assign n4351 = ( ~n4329 & n4334 ) | ( ~n4329 & n4350 ) | ( n4334 & n4350 ) ;
  assign n4352 = ( n4010 & n4335 ) | ( n4010 & n4351 ) | ( n4335 & n4351 ) ;
  assign n4353 = ( n3799 & n4319 ) | ( n3799 & n4352 ) | ( n4319 & n4352 ) ;
  assign n4354 = n4320 | n4353 ;
  buffer buf_n4355( .i (n232), .o (n4355) );
  assign n4356 = ( n4050 & ~n4354 ) | ( n4050 & n4355 ) | ( ~n4354 & n4355 ) ;
  assign n4357 = n4270 & ~n4356 ;
  buffer buf_n4358( .i (n4357), .o (n4358) );
  buffer buf_n4359( .i (n4358), .o (n4359) );
  buffer buf_n4360( .i (n4359), .o (n4360) );
  assign n4361 = ( n718 & n1244 ) | ( n718 & n4358 ) | ( n1244 & n4358 ) ;
  assign n4362 = n601 & ~n4361 ;
  assign n4363 = ( n602 & n4360 ) | ( n602 & ~n4362 ) | ( n4360 & ~n4362 ) ;
  assign n4364 = n4101 | n4363 ;
  assign n4365 = ( n4059 & ~n4060 ) | ( n4059 & n4364 ) | ( ~n4060 & n4364 ) ;
  assign n4366 = n4009 | n4365 ;
  assign n4367 = ( n3947 & ~n3948 ) | ( n3947 & n4366 ) | ( ~n3948 & n4366 ) ;
  buffer buf_n4244( .i (n4243), .o (n4244) );
  buffer buf_n4245( .i (n4244), .o (n4245) );
  buffer buf_n4246( .i (n4245), .o (n4246) );
  buffer buf_n4247( .i (n4246), .o (n4247) );
  buffer buf_n4248( .i (n4247), .o (n4248) );
  buffer buf_n4249( .i (n4248), .o (n4249) );
  buffer buf_n4250( .i (n4249), .o (n4250) );
  buffer buf_n4251( .i (n4250), .o (n4251) );
  buffer buf_n4252( .i (n4251), .o (n4252) );
  buffer buf_n4253( .i (n4252), .o (n4253) );
  buffer buf_n4254( .i (n4253), .o (n4254) );
  buffer buf_n4255( .i (n4254), .o (n4255) );
  buffer buf_n4256( .i (n4255), .o (n4256) );
  buffer buf_n4257( .i (n4256), .o (n4257) );
  buffer buf_n4258( .i (n4257), .o (n4258) );
  buffer buf_n4259( .i (n4258), .o (n4259) );
  buffer buf_n4260( .i (n4259), .o (n4260) );
  buffer buf_n4220( .i (n4219), .o (n4220) );
  buffer buf_n4221( .i (n4220), .o (n4221) );
  buffer buf_n4222( .i (n4221), .o (n4222) );
  buffer buf_n4223( .i (n4222), .o (n4223) );
  buffer buf_n4224( .i (n4223), .o (n4224) );
  buffer buf_n4225( .i (n4224), .o (n4225) );
  buffer buf_n4226( .i (n4225), .o (n4226) );
  buffer buf_n4227( .i (n4226), .o (n4227) );
  buffer buf_n4228( .i (n4227), .o (n4228) );
  buffer buf_n4368( .i (n4210), .o (n4368) );
  assign n4369 = n1478 & ~n4368 ;
  buffer buf_n4370( .i (n4369), .o (n4370) );
  buffer buf_n4371( .i (n4370), .o (n4371) );
  assign n4372 = ( n3429 & ~n4088 ) | ( n3429 & n4370 ) | ( ~n4088 & n4370 ) ;
  assign n4373 = ( n1481 & n4371 ) | ( n1481 & n4372 ) | ( n4371 & n4372 ) ;
  assign n4374 = n2559 & n4373 ;
  buffer buf_n2493( .i (n2492), .o (n2493) );
  buffer buf_n2494( .i (n2493), .o (n2494) );
  buffer buf_n2495( .i (n2494), .o (n2495) );
  buffer buf_n2496( .i (n2495), .o (n2496) );
  buffer buf_n2497( .i (n2496), .o (n2497) );
  assign n4375 = n3781 | n4239 ;
  buffer buf_n4376( .i (n4375), .o (n4376) );
  buffer buf_n4377( .i (n4376), .o (n4377) );
  buffer buf_n4378( .i (n4377), .o (n4378) );
  assign n4381 = ( n2497 & ~n3102 ) | ( n2497 & n4378 ) | ( ~n3102 & n4378 ) ;
  buffer buf_n4382( .i (n3255), .o (n4382) );
  buffer buf_n4383( .i (n4382), .o (n4383) );
  assign n4384 = ( n3720 & ~n4381 ) | ( n3720 & n4383 ) | ( ~n4381 & n4383 ) ;
  assign n4385 = ( ~n4228 & n4374 ) | ( ~n4228 & n4384 ) | ( n4374 & n4384 ) ;
  buffer buf_n4386( .i (n3366), .o (n4386) );
  buffer buf_n4387( .i (n4386), .o (n4387) );
  assign n4388 = ~n4385 & n4387 ;
  buffer buf_n4389( .i (n3338), .o (n4389) );
  assign n4390 = ( ~n3781 & n4338 ) | ( ~n3781 & n4389 ) | ( n4338 & n4389 ) ;
  buffer buf_n4391( .i (n4390), .o (n4391) );
  buffer buf_n4392( .i (n4391), .o (n4392) );
  buffer buf_n4393( .i (n4392), .o (n4393) );
  buffer buf_n4394( .i (n4393), .o (n4394) );
  assign n4395 = ~n4066 & n4391 ;
  buffer buf_n4396( .i (n4395), .o (n4396) );
  buffer buf_n4397( .i (n4396), .o (n4397) );
  buffer buf_n4398( .i (n3785), .o (n4398) );
  buffer buf_n4399( .i (n4332), .o (n4399) );
  buffer buf_n4400( .i (n4399), .o (n4400) );
  buffer buf_n4401( .i (n4400), .o (n4401) );
  assign n4402 = ( n4396 & ~n4398 ) | ( n4396 & n4401 ) | ( ~n4398 & n4401 ) ;
  assign n4403 = ( n4394 & n4397 ) | ( n4394 & n4402 ) | ( n4397 & n4402 ) ;
  assign n4404 = n3963 & n4403 ;
  assign n4405 = n4387 | n4404 ;
  assign n4406 = ~n4388 & n4405 ;
  assign n4407 = ( ~n2758 & n3460 ) | ( ~n2758 & n4406 ) | ( n3460 & n4406 ) ;
  assign n4408 = ~n456 & n3785 ;
  buffer buf_n4409( .i (n4336), .o (n4409) );
  assign n4410 = ( ~n455 & n3214 ) | ( ~n455 & n4409 ) | ( n3214 & n4409 ) ;
  buffer buf_n4411( .i (n4368), .o (n4411) );
  buffer buf_n4412( .i (n4411), .o (n4412) );
  assign n4413 = ( n2197 & ~n4410 ) | ( n2197 & n4412 ) | ( ~n4410 & n4412 ) ;
  assign n4414 = ( ~n4398 & n4408 ) | ( ~n4398 & n4413 ) | ( n4408 & n4413 ) ;
  buffer buf_n4415( .i (n4302), .o (n4415) );
  buffer buf_n4416( .i (n4415), .o (n4416) );
  buffer buf_n4417( .i (n4416), .o (n4417) );
  assign n4418 = n4414 | n4417 ;
  buffer buf_n4419( .i (n3794), .o (n4419) );
  assign n4420 = ~n1757 & n4419 ;
  buffer buf_n4421( .i (n4420), .o (n4421) );
  assign n4423 = ~n4398 & n4421 ;
  assign n4424 = n4417 & ~n4423 ;
  assign n4425 = n4418 & ~n4424 ;
  assign n4426 = n3893 & n4425 ;
  assign n4427 = ( n4191 & n4336 ) | ( n4191 & ~n4368 ) | ( n4336 & ~n4368 ) ;
  buffer buf_n4428( .i (n4427), .o (n4428) );
  buffer buf_n4429( .i (n4419), .o (n4429) );
  assign n4430 = ( n4412 & n4428 ) | ( n4412 & n4429 ) | ( n4428 & n4429 ) ;
  assign n4431 = n4412 & n4428 ;
  assign n4432 = n4428 | n4429 ;
  assign n4433 = ( ~n4430 & n4431 ) | ( ~n4430 & n4432 ) | ( n4431 & n4432 ) ;
  buffer buf_n4434( .i (n4401), .o (n4434) );
  assign n4435 = ~n4433 & n4434 ;
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n2153( .i (n2152), .o (n2153) );
  assign n4436 = ( n442 & n634 ) | ( n442 & ~n2153 ) | ( n634 & ~n2153 ) ;
  buffer buf_n4437( .i (n4436), .o (n4437) );
  assign n4440 = n4382 & n4437 ;
  assign n4441 = n4434 | n4440 ;
  assign n4442 = ~n4435 & n4441 ;
  assign n4443 = n3893 | n4442 ;
  buffer buf_n4444( .i (n3964), .o (n4444) );
  buffer buf_n4445( .i (n4444), .o (n4445) );
  assign n4446 = ( n4426 & n4443 ) | ( n4426 & ~n4445 ) | ( n4443 & ~n4445 ) ;
  buffer buf_n4447( .i (n3459), .o (n4447) );
  assign n4448 = ( n2758 & n4446 ) | ( n2758 & n4447 ) | ( n4446 & n4447 ) ;
  assign n4449 = n4407 & n4448 ;
  buffer buf_n4450( .i (n4449), .o (n4450) );
  buffer buf_n4451( .i (n4450), .o (n4451) );
  assign n4452 = n3111 & n4450 ;
  buffer buf_n4020( .i (n4019), .o (n4020) );
  buffer buf_n4021( .i (n4020), .o (n4021) );
  buffer buf_n4022( .i (n4021), .o (n4022) );
  assign n4453 = n3538 & ~n4022 ;
  buffer buf_n4454( .i (n4453), .o (n4454) );
  buffer buf_n4455( .i (n4454), .o (n4455) );
  buffer buf_n4456( .i (n4398), .o (n4456) );
  assign n4457 = ( n2097 & n3103 ) | ( n2097 & n4456 ) | ( n3103 & n4456 ) ;
  assign n4458 = ~n2098 & n4457 ;
  assign n4459 = n4454 | n4458 ;
  buffer buf_n4460( .i (n4050), .o (n4460) );
  assign n4461 = ( n4455 & n4459 ) | ( n4455 & ~n4460 ) | ( n4459 & ~n4460 ) ;
  buffer buf_n4462( .i (n4461), .o (n4462) );
  buffer buf_n4463( .i (n4462), .o (n4463) );
  buffer buf_n4464( .i (n4447), .o (n4464) );
  assign n4465 = ( n2321 & n4462 ) | ( n2321 & n4464 ) | ( n4462 & n4464 ) ;
  assign n4466 = ( n440 & ~n1362 ) | ( n440 & n2516 ) | ( ~n1362 & n2516 ) ;
  buffer buf_n4467( .i (n4466), .o (n4467) );
  buffer buf_n4468( .i (n3713), .o (n4468) );
  assign n4469 = n4467 & n4468 ;
  buffer buf_n4470( .i (n4469), .o (n4470) );
  buffer buf_n4471( .i (n4470), .o (n4471) );
  assign n4472 = n2910 & n4306 ;
  buffer buf_n4473( .i (n4472), .o (n4473) );
  assign n4482 = ( n3463 & ~n4231 ) | ( n3463 & n4473 ) | ( ~n4231 & n4473 ) ;
  buffer buf_n4483( .i (n4482), .o (n4483) );
  buffer buf_n4484( .i (n4483), .o (n4484) );
  buffer buf_n4485( .i (n4484), .o (n4485) );
  assign n4486 = ( n4185 & ~n4209 ) | ( n4185 & n4483 ) | ( ~n4209 & n4483 ) ;
  buffer buf_n4487( .i (n4325), .o (n4487) );
  assign n4488 = ( n4389 & ~n4486 ) | ( n4389 & n4487 ) | ( ~n4486 & n4487 ) ;
  assign n4489 = ~n4485 & n4488 ;
  assign n4490 = n4468 | n4489 ;
  buffer buf_n4491( .i (n4231), .o (n4491) );
  assign n4492 = n1045 & n4491 ;
  buffer buf_n4493( .i (n4492), .o (n4493) );
  assign n4502 = n3005 | n4491 ;
  buffer buf_n4503( .i (n4502), .o (n4503) );
  assign n4512 = ~n4493 & n4503 ;
  assign n4513 = n4368 & ~n4512 ;
  assign n4514 = n4468 & ~n4513 ;
  assign n4515 = n4490 & ~n4514 ;
  buffer buf_n4516( .i (n4210), .o (n4516) );
  assign n4517 = n1015 & ~n4516 ;
  assign n4518 = n3916 & n4517 ;
  buffer buf_n4519( .i (n4518), .o (n4519) );
  assign n4520 = ( ~n4470 & n4515 ) | ( ~n4470 & n4519 ) | ( n4515 & n4519 ) ;
  assign n4521 = n3511 & ~n4519 ;
  assign n4522 = ( n4471 & n4520 ) | ( n4471 & ~n4521 ) | ( n4520 & ~n4521 ) ;
  assign n4523 = n3848 & ~n4522 ;
  buffer buf_n3007( .i (n3006), .o (n3007) );
  buffer buf_n3008( .i (n3007), .o (n3008) );
  buffer buf_n3009( .i (n3008), .o (n3009) );
  buffer buf_n4524( .i (n3004), .o (n4524) );
  assign n4525 = ( ~n2764 & n4311 ) | ( ~n2764 & n4524 ) | ( n4311 & n4524 ) ;
  buffer buf_n4526( .i (n4525), .o (n4526) );
  buffer buf_n4527( .i (n4526), .o (n4527) );
  buffer buf_n4528( .i (n4527), .o (n4528) );
  buffer buf_n4529( .i (n4209), .o (n4529) );
  assign n4530 = ( n3765 & n4526 ) | ( n3765 & ~n4529 ) | ( n4526 & ~n4529 ) ;
  buffer buf_n4531( .i (n4389), .o (n4531) );
  assign n4532 = ( n3008 & n4530 ) | ( n3008 & ~n4531 ) | ( n4530 & ~n4531 ) ;
  assign n4533 = ( ~n3009 & n4528 ) | ( ~n3009 & n4532 ) | ( n4528 & n4532 ) ;
  assign n4534 = n4429 & n4533 ;
  buffer buf_n4535( .i (n3548), .o (n4535) );
  assign n4536 = ( n4309 & n4311 ) | ( n4309 & n4535 ) | ( n4311 & n4535 ) ;
  buffer buf_n4537( .i (n4536), .o (n4537) );
  buffer buf_n4538( .i (n4537), .o (n4538) );
  assign n4541 = ~n4529 & n4537 ;
  assign n4542 = ( ~n607 & n4538 ) | ( ~n607 & n4541 ) | ( n4538 & n4541 ) ;
  assign n4543 = n4066 & n4542 ;
  assign n4544 = n4429 | n4543 ;
  assign n4545 = ~n4534 & n4544 ;
  assign n4546 = ~n3435 & n4545 ;
  assign n4547 = n3848 | n4546 ;
  assign n4548 = ~n4523 & n4547 ;
  assign n4549 = n3975 | n4548 ;
  buffer buf_n4550( .i (n4174), .o (n4550) );
  assign n4551 = ( n1275 & n3187 ) | ( n1275 & ~n4550 ) | ( n3187 & ~n4550 ) ;
  buffer buf_n4552( .i (n4551), .o (n4552) );
  buffer buf_n4553( .i (n4552), .o (n4553) );
  buffer buf_n4558( .i (n2853), .o (n4558) );
  buffer buf_n4559( .i (n3061), .o (n4559) );
  buffer buf_n4560( .i (n4559), .o (n4560) );
  assign n4561 = ( n4553 & n4558 ) | ( n4553 & ~n4560 ) | ( n4558 & ~n4560 ) ;
  buffer buf_n4562( .i (n4561), .o (n4562) );
  assign n4565 = n4209 & ~n4562 ;
  buffer buf_n4566( .i (n4565), .o (n4566) );
  buffer buf_n4567( .i (n4566), .o (n4567) );
  buffer buf_n4563( .i (n4562), .o (n4563) );
  buffer buf_n4564( .i (n4563), .o (n4564) );
  assign n4568 = n4564 | n4566 ;
  assign n4569 = ( ~n4411 & n4567 ) | ( ~n4411 & n4568 ) | ( n4567 & n4568 ) ;
  assign n4570 = n4400 & n4569 ;
  buffer buf_n4571( .i (n3337), .o (n4571) );
  buffer buf_n4572( .i (n3043), .o (n4572) );
  assign n4573 = ( ~n3896 & n4571 ) | ( ~n3896 & n4572 ) | ( n4571 & n4572 ) ;
  buffer buf_n4574( .i (n4573), .o (n4574) );
  buffer buf_n4575( .i (n4574), .o (n4575) );
  assign n4576 = n4531 & ~n4574 ;
  assign n4577 = ( n2039 & n4575 ) | ( n2039 & ~n4576 ) | ( n4575 & ~n4576 ) ;
  assign n4578 = ~n4400 & n4577 ;
  assign n4579 = ( n4401 & ~n4570 ) | ( n4401 & n4578 ) | ( ~n4570 & n4578 ) ;
  assign n4580 = n3366 & ~n4579 ;
  buffer buf_n4581( .i (n4311), .o (n4581) );
  assign n4582 = n3896 | n4581 ;
  buffer buf_n4583( .i (n4582), .o (n4583) );
  assign n4589 = n4336 & n4583 ;
  assign n4590 = ( n608 & n2609 ) | ( n608 & ~n4589 ) | ( n2609 & ~n4589 ) ;
  assign n4591 = ~n4088 & n4590 ;
  assign n4592 = ( n274 & n1756 ) | ( n274 & ~n2119 ) | ( n1756 & ~n2119 ) ;
  buffer buf_n4593( .i (n4592), .o (n4593) );
  assign n4606 = ( n4088 & n4412 ) | ( n4088 & n4593 ) | ( n4412 & n4593 ) ;
  assign n4607 = ( n689 & n4591 ) | ( n689 & ~n4606 ) | ( n4591 & ~n4606 ) ;
  assign n4608 = n3366 | n4607 ;
  assign n4609 = ( ~n4386 & n4580 ) | ( ~n4386 & n4608 ) | ( n4580 & n4608 ) ;
  buffer buf_n4610( .i (n4049), .o (n4610) );
  assign n4611 = n4609 & ~n4610 ;
  assign n4612 = n3975 & ~n4611 ;
  assign n4613 = n4549 & ~n4612 ;
  assign n4614 = ~n4464 & n4613 ;
  assign n4615 = ( n4463 & ~n4465 ) | ( n4463 & n4614 ) | ( ~n4465 & n4614 ) ;
  buffer buf_n3680( .i (n3679), .o (n3680) );
  buffer buf_n3681( .i (n3680), .o (n3681) );
  buffer buf_n3682( .i (n3681), .o (n3682) );
  buffer buf_n3683( .i (n3682), .o (n3683) );
  buffer buf_n3684( .i (n3683), .o (n3684) );
  buffer buf_n3685( .i (n3684), .o (n3685) );
  buffer buf_n3686( .i (n3685), .o (n3686) );
  assign n4616 = ~n1586 & n3686 ;
  assign n4617 = ( ~n3510 & n4415 ) | ( ~n3510 & n4616 ) | ( n4415 & n4616 ) ;
  assign n4618 = n512 & n4531 ;
  assign n4619 = n1945 & n4618 ;
  assign n4620 = ~n3510 & n4619 ;
  assign n4621 = ( ~n4416 & n4617 ) | ( ~n4416 & n4620 ) | ( n4617 & n4620 ) ;
  buffer buf_n4622( .i (n4621), .o (n4622) );
  assign n4623 = ( ~n755 & n1401 ) | ( ~n755 & n4622 ) | ( n1401 & n4622 ) ;
  assign n4624 = ( n373 & n515 ) | ( n373 & ~n1806 ) | ( n515 & ~n1806 ) ;
  buffer buf_n4625( .i (n4624), .o (n4625) );
  assign n4631 = n4622 | n4625 ;
  assign n4632 = ( n756 & n4623 ) | ( n756 & n4631 ) | ( n4623 & n4631 ) ;
  assign n4633 = n262 | n4632 ;
  buffer buf_n4634( .i (n3002), .o (n4634) );
  buffer buf_n4635( .i (n4634), .o (n4635) );
  buffer buf_n4636( .i (n4635), .o (n4636) );
  buffer buf_n4637( .i (n4560), .o (n4637) );
  assign n4638 = ( n4205 & ~n4636 ) | ( n4205 & n4637 ) | ( ~n4636 & n4637 ) ;
  assign n4639 = ( n3907 & ~n4185 ) | ( n3907 & n4638 ) | ( ~n4185 & n4638 ) ;
  buffer buf_n4640( .i (n4639), .o (n4640) );
  assign n4643 = n3768 & ~n4640 ;
  buffer buf_n4644( .i (n4643), .o (n4644) );
  buffer buf_n4645( .i (n4644), .o (n4645) );
  buffer buf_n4641( .i (n4640), .o (n4641) );
  buffer buf_n4642( .i (n4641), .o (n4642) );
  assign n4646 = n4642 | n4644 ;
  assign n4647 = ( ~n3957 & n4645 ) | ( ~n3957 & n4646 ) | ( n4645 & n4646 ) ;
  assign n4648 = n4417 & n4647 ;
  assign n4649 = ( n2543 & n3907 ) | ( n2543 & ~n4571 ) | ( n3907 & ~n4571 ) ;
  buffer buf_n4650( .i (n4649), .o (n4650) );
  buffer buf_n4651( .i (n4650), .o (n4651) );
  buffer buf_n4652( .i (n4651), .o (n4652) );
  buffer buf_n4653( .i (n4652), .o (n4653) );
  buffer buf_n4654( .i (n3665), .o (n4654) );
  buffer buf_n4655( .i (n4338), .o (n4655) );
  assign n4656 = ( n4650 & n4654 ) | ( n4650 & n4655 ) | ( n4654 & n4655 ) ;
  buffer buf_n4657( .i (n4656), .o (n4657) );
  buffer buf_n4658( .i (n4657), .o (n4658) );
  assign n4659 = n2547 & ~n4657 ;
  assign n4660 = ( n4653 & ~n4658 ) | ( n4653 & n4659 ) | ( ~n4658 & n4659 ) ;
  assign n4661 = n4417 | n4660 ;
  assign n4662 = ( ~n3963 & n4648 ) | ( ~n3963 & n4661 ) | ( n4648 & n4661 ) ;
  assign n4663 = ~n4610 & n4662 ;
  assign n4664 = n262 & ~n4663 ;
  assign n4665 = n4633 & ~n4664 ;
  assign n4666 = n3400 | n4665 ;
  assign n4667 = ( n3101 & n3623 ) | ( n3101 & n4113 ) | ( n3623 & n4113 ) ;
  assign n4668 = ~n3957 & n4667 ;
  buffer buf_n4669( .i (n4668), .o (n4669) );
  buffer buf_n4670( .i (n4669), .o (n4670) );
  buffer buf_n4671( .i (n4670), .o (n4671) );
  assign n4672 = ( n4075 & n4309 ) | ( n4075 & n4636 ) | ( n4309 & n4636 ) ;
  buffer buf_n4673( .i (n4672), .o (n4673) );
  buffer buf_n4674( .i (n4673), .o (n4674) );
  buffer buf_n4675( .i (n4674), .o (n4675) );
  buffer buf_n4676( .i (n4675), .o (n4676) );
  buffer buf_n4677( .i (n4676), .o (n4677) );
  buffer buf_n4678( .i (n4677), .o (n4678) );
  assign n4679 = ( n3102 & n4382 ) | ( n3102 & n4401 ) | ( n4382 & n4401 ) ;
  assign n4680 = n4678 & ~n4679 ;
  assign n4681 = ( n4014 & n4669 ) | ( n4014 & n4680 ) | ( n4669 & n4680 ) ;
  assign n4682 = n4387 & ~n4681 ;
  assign n4683 = ( n4096 & n4671 ) | ( n4096 & ~n4682 ) | ( n4671 & ~n4682 ) ;
  assign n4684 = ~n3891 & n4683 ;
  assign n4685 = n3400 & ~n4684 ;
  assign n4686 = n4666 & ~n4685 ;
  assign n4687 = n4615 | n4686 ;
  assign n4688 = ( n4451 & ~n4452 ) | ( n4451 & n4687 ) | ( ~n4452 & n4687 ) ;
  buffer buf_n4689( .i (n4688), .o (n4689) );
  buffer buf_n4690( .i (n4689), .o (n4690) );
  assign n4691 = ( n45 & n2277 ) | ( n45 & n4215 ) | ( n2277 & n4215 ) ;
  buffer buf_n4692( .i (n4691), .o (n4692) );
  buffer buf_n4693( .i (n4692), .o (n4693) );
  buffer buf_n4694( .i (n4693), .o (n4694) );
  buffer buf_n4695( .i (n4694), .o (n4695) );
  buffer buf_n4696( .i (n4695), .o (n4696) );
  buffer buf_n4697( .i (n4696), .o (n4697) );
  buffer buf_n4698( .i (n4697), .o (n4698) );
  buffer buf_n4699( .i (n4698), .o (n4699) );
  buffer buf_n4700( .i (n4699), .o (n4700) );
  buffer buf_n4701( .i (n4700), .o (n4701) );
  buffer buf_n4702( .i (n4701), .o (n4702) );
  buffer buf_n4703( .i (n4702), .o (n4703) );
  buffer buf_n4704( .i (n4703), .o (n4704) );
  buffer buf_n4705( .i (n4704), .o (n4705) );
  assign n4706 = ( n3974 & n4355 ) | ( n3974 & n4444 ) | ( n4355 & n4444 ) ;
  assign n4707 = ( n570 & ~n4705 ) | ( n570 & n4706 ) | ( ~n4705 & n4706 ) ;
  buffer buf_n4708( .i (n4707), .o (n4708) );
  buffer buf_n4709( .i (n4708), .o (n4709) );
  assign n4710 = ( n264 & n4464 ) | ( n264 & ~n4708 ) | ( n4464 & ~n4708 ) ;
  assign n4711 = n4239 & n4529 ;
  buffer buf_n4712( .i (n4711), .o (n4712) );
  buffer buf_n4713( .i (n4712), .o (n4713) );
  buffer buf_n4714( .i (n4713), .o (n4714) );
  buffer buf_n4715( .i (n4714), .o (n4715) );
  buffer buf_n4716( .i (n4715), .o (n4716) );
  buffer buf_n4717( .i (n4716), .o (n4717) );
  buffer buf_n4718( .i (n4717), .o (n4718) );
  buffer buf_n4719( .i (n4434), .o (n4719) );
  buffer buf_n4720( .i (n4719), .o (n4720) );
  buffer buf_n4721( .i (n4720), .o (n4721) );
  assign n4722 = ( n4445 & n4718 ) | ( n4445 & n4721 ) | ( n4718 & n4721 ) ;
  assign n4723 = ~n263 & n4722 ;
  assign n4724 = n4464 & n4723 ;
  assign n4725 = ( n4709 & n4710 ) | ( n4709 & n4724 ) | ( n4710 & n4724 ) ;
  buffer buf_n4726( .i (n4725), .o (n4726) );
  buffer buf_n4727( .i (n4726), .o (n4727) );
  assign n4728 = ( n4325 & n4571 ) | ( n4325 & ~n4581 ) | ( n4571 & ~n4581 ) ;
  buffer buf_n4729( .i (n4728), .o (n4729) );
  buffer buf_n4730( .i (n4729), .o (n4730) );
  buffer buf_n4731( .i (n4730), .o (n4731) );
  buffer buf_n4732( .i (n4731), .o (n4732) );
  buffer buf_n4733( .i (n4732), .o (n4733) );
  buffer buf_n4738( .i (n3883), .o (n4738) );
  assign n4739 = ( n4456 & n4733 ) | ( n4456 & n4738 ) | ( n4733 & n4738 ) ;
  buffer buf_n4740( .i (n4739), .o (n4740) );
  buffer buf_n4741( .i (n4740), .o (n4741) );
  buffer buf_n4742( .i (n4741), .o (n4742) );
  buffer buf_n4743( .i (n4742), .o (n4743) );
  assign n4744 = ( n4444 & n4720 ) | ( n4444 & n4740 ) | ( n4720 & n4740 ) ;
  buffer buf_n4745( .i (n4744), .o (n4745) );
  buffer buf_n4746( .i (n4745), .o (n4746) );
  buffer buf_n4734( .i (n4733), .o (n4734) );
  buffer buf_n4735( .i (n4734), .o (n4735) );
  buffer buf_n4736( .i (n4735), .o (n4736) );
  buffer buf_n4737( .i (n4736), .o (n4737) );
  assign n4747 = n4737 & ~n4745 ;
  assign n4748 = ( n4743 & ~n4746 ) | ( n4743 & n4747 ) | ( ~n4746 & n4747 ) ;
  assign n4749 = ( ~n2640 & n3835 ) | ( ~n2640 & n4748 ) | ( n3835 & n4748 ) ;
  assign n4750 = ( n4308 & n4558 ) | ( n4308 & n4635 ) | ( n4558 & n4635 ) ;
  buffer buf_n4751( .i (n4750), .o (n4751) );
  buffer buf_n4752( .i (n4751), .o (n4752) );
  buffer buf_n4753( .i (n4752), .o (n4753) );
  buffer buf_n4754( .i (n4753), .o (n4754) );
  buffer buf_n4755( .i (n4754), .o (n4755) );
  buffer buf_n4756( .i (n4755), .o (n4756) );
  buffer buf_n4757( .i (n4756), .o (n4757) );
  buffer buf_n4758( .i (n3617), .o (n4758) );
  assign n4759 = ( ~n4738 & n4757 ) | ( ~n4738 & n4758 ) | ( n4757 & n4758 ) ;
  buffer buf_n4760( .i (n4759), .o (n4760) );
  assign n4763 = n4444 & ~n4760 ;
  buffer buf_n4764( .i (n4763), .o (n4764) );
  buffer buf_n4765( .i (n4764), .o (n4765) );
  buffer buf_n4761( .i (n4760), .o (n4761) );
  buffer buf_n4762( .i (n4761), .o (n4762) );
  assign n4766 = n4762 | n4764 ;
  assign n4767 = ( ~n148 & n4765 ) | ( ~n148 & n4766 ) | ( n4765 & n4766 ) ;
  buffer buf_n4768( .i (n3975), .o (n4768) );
  buffer buf_n4769( .i (n4768), .o (n4769) );
  buffer buf_n4770( .i (n4769), .o (n4770) );
  assign n4771 = ( n2640 & ~n4767 ) | ( n2640 & n4770 ) | ( ~n4767 & n4770 ) ;
  assign n4772 = n4749 & ~n4771 ;
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n4773( .i (n3721), .o (n4773) );
  assign n4774 = ( n749 & ~n4355 ) | ( n749 & n4773 ) | ( ~n4355 & n4773 ) ;
  buffer buf_n4775( .i (n4416), .o (n4775) );
  buffer buf_n4776( .i (n4775), .o (n4776) );
  assign n4777 = ( ~n748 & n3721 ) | ( ~n748 & n4776 ) | ( n3721 & n4776 ) ;
  assign n4778 = ( n4094 & ~n4355 ) | ( n4094 & n4777 ) | ( ~n4355 & n4777 ) ;
  assign n4779 = ~n4774 & n4778 ;
  buffer buf_n4780( .i (n4779), .o (n4780) );
  buffer buf_n4781( .i (n4780), .o (n4781) );
  assign n4782 = ( n3020 & n3839 ) | ( n3020 & n4780 ) | ( n3839 & n4780 ) ;
  buffer buf_n4783( .i (n4411), .o (n4783) );
  assign n4784 = n3882 & ~n4783 ;
  buffer buf_n4785( .i (n4784), .o (n4785) );
  buffer buf_n4786( .i (n4785), .o (n4786) );
  buffer buf_n4787( .i (n4786), .o (n4787) );
  buffer buf_n4788( .i (n4787), .o (n4788) );
  buffer buf_n4789( .i (n4094), .o (n4789) );
  assign n4790 = ( n709 & n4788 ) | ( n709 & n4789 ) | ( n4788 & n4789 ) ;
  assign n4791 = ~n4447 & n4790 ;
  assign n4792 = ~n3020 & n4791 ;
  assign n4793 = ( n4781 & ~n4782 ) | ( n4781 & n4792 ) | ( ~n4782 & n4792 ) ;
  buffer buf_n4794( .i (n4793), .o (n4794) );
  assign n4795 = ( ~n4726 & n4772 ) | ( ~n4726 & n4794 ) | ( n4772 & n4794 ) ;
  assign n4796 = n3025 & ~n4794 ;
  assign n4797 = ( n4727 & n4795 ) | ( n4727 & ~n4796 ) | ( n4795 & ~n4796 ) ;
  assign n4798 = n4689 | n4797 ;
  assign n4799 = ( ~n4260 & n4690 ) | ( ~n4260 & n4798 ) | ( n4690 & n4798 ) ;
  buffer buf_n1405( .i (n1404), .o (n1405) );
  assign n4800 = ( n689 & ~n801 ) | ( n689 & n2778 ) | ( ~n801 & n2778 ) ;
  assign n4801 = ( n690 & ~n4456 ) | ( n690 & n4800 ) | ( ~n4456 & n4800 ) ;
  assign n4802 = n4776 & ~n4801 ;
  assign n4803 = ~n4610 & n4802 ;
  buffer buf_n4804( .i (n4803), .o (n4804) );
  buffer buf_n4805( .i (n4804), .o (n4805) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  assign n4806 = n1569 & ~n4804 ;
  assign n4807 = ( n1405 & n4805 ) | ( n1405 & ~n4806 ) | ( n4805 & ~n4806 ) ;
  buffer buf_n4808( .i (n4807), .o (n4808) );
  buffer buf_n4809( .i (n4808), .o (n4809) );
  assign n4810 = n1404 & n2248 ;
  assign n4811 = n404 & n4810 ;
  assign n4812 = n542 | n4386 ;
  assign n4813 = ( ~n2724 & n3105 ) | ( ~n2724 & n4812 ) | ( n3105 & n4812 ) ;
  assign n4814 = ( n370 & n1429 ) | ( n370 & ~n2885 ) | ( n1429 & ~n2885 ) ;
  buffer buf_n4815( .i (n4324), .o (n4815) );
  buffer buf_n4816( .i (n4815), .o (n4816) );
  buffer buf_n4817( .i (n4816), .o (n4817) );
  buffer buf_n4818( .i (n4205), .o (n4818) );
  buffer buf_n4819( .i (n4818), .o (n4819) );
  buffer buf_n4820( .i (n4819), .o (n4820) );
  buffer buf_n4821( .i (n4820), .o (n4821) );
  assign n4822 = ( n4814 & n4817 ) | ( n4814 & ~n4821 ) | ( n4817 & ~n4821 ) ;
  buffer buf_n4823( .i (n4822), .o (n4823) );
  buffer buf_n4824( .i (n4823), .o (n4824) );
  assign n4825 = ~n4416 & n4823 ;
  buffer buf_n4826( .i (n3957), .o (n4826) );
  assign n4827 = ( n4824 & n4825 ) | ( n4824 & n4826 ) | ( n4825 & n4826 ) ;
  buffer buf_n4828( .i (n4827), .o (n4828) );
  buffer buf_n4829( .i (n4828), .o (n4829) );
  buffer buf_n4830( .i (n4383), .o (n4830) );
  buffer buf_n4831( .i (n4830), .o (n4831) );
  assign n4832 = n4828 | n4831 ;
  assign n4833 = ( n4813 & n4829 ) | ( n4813 & n4832 ) | ( n4829 & n4832 ) ;
  assign n4834 = ( n2689 & ~n3891 ) | ( n2689 & n4833 ) | ( ~n3891 & n4833 ) ;
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n2155( .i (n2154), .o (n2155) );
  buffer buf_n4835( .i (n4531), .o (n4835) );
  buffer buf_n4836( .i (n4835), .o (n4836) );
  assign n4837 = ( ~n309 & n4415 ) | ( ~n309 & n4836 ) | ( n4415 & n4836 ) ;
  buffer buf_n4838( .i (n4419), .o (n4838) );
  assign n4839 = ( ~n309 & n4836 ) | ( ~n309 & n4838 ) | ( n4836 & n4838 ) ;
  assign n4840 = ( n2155 & n4837 ) | ( n2155 & ~n4839 ) | ( n4837 & ~n4839 ) ;
  assign n4841 = ~n4383 & n4840 ;
  buffer buf_n4842( .i (n4841), .o (n4842) );
  buffer buf_n4843( .i (n4842), .o (n4843) );
  buffer buf_n4844( .i (n4415), .o (n4844) );
  buffer buf_n4845( .i (n4113), .o (n4845) );
  assign n4846 = ( n4382 & n4844 ) | ( n4382 & ~n4845 ) | ( n4844 & ~n4845 ) ;
  buffer buf_n4847( .i (n4846), .o (n4847) );
  assign n4851 = n3408 & n4847 ;
  assign n4852 = n4842 | n4851 ;
  assign n4853 = ( ~n4445 & n4843 ) | ( ~n4445 & n4852 ) | ( n4843 & n4852 ) ;
  buffer buf_n4854( .i (n2688), .o (n4854) );
  assign n4855 = ( n3891 & ~n4853 ) | ( n3891 & n4854 ) | ( ~n4853 & n4854 ) ;
  assign n4856 = n4834 & ~n4855 ;
  assign n4857 = ( ~n356 & n4811 ) | ( ~n356 & n4856 ) | ( n4811 & n4856 ) ;
  assign n4858 = ~n4808 & n4857 ;
  assign n4859 = ( ~n358 & n4809 ) | ( ~n358 & n4858 ) | ( n4809 & n4858 ) ;
  buffer buf_n4860( .i (n4859), .o (n4860) );
  buffer buf_n4861( .i (n4860), .o (n4861) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n2498( .i (n2497), .o (n2498) );
  buffer buf_n2499( .i (n2498), .o (n2499) );
  assign n4862 = ( n2499 & n3721 ) | ( n2499 & n4049 ) | ( n3721 & n4049 ) ;
  buffer buf_n4863( .i (n3510), .o (n4863) );
  buffer buf_n4864( .i (n4863), .o (n4864) );
  assign n4865 = ( ~n2498 & n4456 ) | ( ~n2498 & n4864 ) | ( n4456 & n4864 ) ;
  assign n4866 = ( n3964 & ~n4719 ) | ( n3964 & n4865 ) | ( ~n4719 & n4865 ) ;
  assign n4867 = ~n4862 & n4866 ;
  assign n4868 = n926 & ~n4783 ;
  assign n4869 = ( ~n3617 & n4863 ) | ( ~n3617 & n4868 ) | ( n4863 & n4868 ) ;
  assign n4870 = ~n4864 & n4869 ;
  buffer buf_n4871( .i (n4870), .o (n4871) );
  buffer buf_n4872( .i (n4871), .o (n4872) );
  buffer buf_n4873( .i (n232), .o (n4873) );
  assign n4874 = n4871 | n4873 ;
  assign n4875 = ( n4867 & n4872 ) | ( n4867 & n4874 ) | ( n4872 & n4874 ) ;
  assign n4876 = n4768 | n4875 ;
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  assign n4877 = n3896 & n4581 ;
  buffer buf_n4878( .i (n4877), .o (n4878) );
  buffer buf_n4879( .i (n4878), .o (n4879) );
  buffer buf_n4880( .i (n4879), .o (n4880) );
  buffer buf_n4881( .i (n4880), .o (n4881) );
  buffer buf_n4882( .i (n4881), .o (n4882) );
  buffer buf_n4883( .i (n4882), .o (n4883) );
  buffer buf_n4884( .i (n4883), .o (n4884) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n4887( .i (n4783), .o (n4887) );
  buffer buf_n4888( .i (n4887), .o (n4888) );
  buffer buf_n4889( .i (n4888), .o (n4889) );
  assign n4890 = ~n672 & n4889 ;
  assign n4891 = ( n661 & n4884 ) | ( n661 & ~n4890 ) | ( n4884 & ~n4890 ) ;
  assign n4892 = ~n4460 & n4891 ;
  assign n4893 = n4768 & ~n4892 ;
  assign n4894 = n4876 & ~n4893 ;
  buffer buf_n4895( .i (n4447), .o (n4895) );
  buffer buf_n4896( .i (n4895), .o (n4896) );
  assign n4897 = n4894 | n4896 ;
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n4898( .i (n4836), .o (n4898) );
  assign n4899 = ( n610 & n4844 ) | ( n610 & ~n4898 ) | ( n4844 & ~n4898 ) ;
  assign n4900 = ( n609 & ~n3882 ) | ( n609 & n4836 ) | ( ~n3882 & n4836 ) ;
  buffer buf_n4901( .i (n4400), .o (n4901) );
  assign n4902 = ( n4844 & ~n4900 ) | ( n4844 & n4901 ) | ( ~n4900 & n4901 ) ;
  assign n4903 = ~n4899 & n4902 ;
  buffer buf_n4904( .i (n4903), .o (n4904) );
  buffer buf_n4905( .i (n4904), .o (n4905) );
  buffer buf_n4906( .i (n4905), .o (n4906) );
  buffer buf_n4907( .i (n3964), .o (n4907) );
  assign n4908 = ( n930 & n4904 ) | ( n930 & ~n4907 ) | ( n4904 & ~n4907 ) ;
  assign n4909 = n839 & ~n4908 ;
  assign n4910 = ( n840 & n4906 ) | ( n840 & ~n4909 ) | ( n4906 & ~n4909 ) ;
  buffer buf_n4911( .i (n4460), .o (n4911) );
  buffer buf_n4912( .i (n4911), .o (n4912) );
  assign n4913 = n4910 & ~n4912 ;
  assign n4914 = n4896 & ~n4913 ;
  assign n4915 = n4897 & ~n4914 ;
  assign n4916 = n181 | n4915 ;
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  assign n4917 = ( n281 & n1370 ) | ( n281 & ~n4788 ) | ( n1370 & ~n4788 ) ;
  assign n4918 = ~n747 & n4826 ;
  buffer buf_n4919( .i (n4918), .o (n4919) );
  buffer buf_n4920( .i (n4919), .o (n4920) );
  buffer buf_n4921( .i (n4920), .o (n4921) );
  assign n4922 = n4917 & n4921 ;
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  assign n4923 = n278 & ~n4888 ;
  buffer buf_n4924( .i (n4923), .o (n4924) );
  buffer buf_n4925( .i (n4924), .o (n4925) );
  buffer buf_n4926( .i (n4925), .o (n4926) );
  assign n4927 = ( ~n751 & n4921 ) | ( ~n751 & n4926 ) | ( n4921 & n4926 ) ;
  assign n4928 = ( n4769 & n4922 ) | ( n4769 & n4927 ) | ( n4922 & n4927 ) ;
  assign n4929 = n4919 & n4924 ;
  assign n4930 = n928 & n4888 ;
  buffer buf_n4931( .i (n4930), .o (n4931) );
  assign n4937 = ( ~n749 & n4919 ) | ( ~n749 & n4931 ) | ( n4919 & n4931 ) ;
  buffer buf_n4938( .i (n3974), .o (n4938) );
  assign n4939 = ( n4929 & n4937 ) | ( n4929 & n4938 ) | ( n4937 & n4938 ) ;
  buffer buf_n4940( .i (n4939), .o (n4940) );
  buffer buf_n4941( .i (n4940), .o (n4941) );
  assign n4942 = n148 & ~n4940 ;
  assign n4943 = ( n4928 & n4941 ) | ( n4928 & ~n4942 ) | ( n4941 & ~n4942 ) ;
  buffer buf_n4944( .i (n3416), .o (n4944) );
  assign n4945 = n4943 & ~n4944 ;
  assign n4946 = n181 & ~n4945 ;
  assign n4947 = n4916 & ~n4946 ;
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  assign n4948 = ~n341 & n1812 ;
  buffer buf_n4949( .i (n2761), .o (n4949) );
  assign n4950 = ( n2584 & n4634 ) | ( n2584 & ~n4949 ) | ( n4634 & ~n4949 ) ;
  buffer buf_n4951( .i (n4950), .o (n4951) );
  assign n4954 = n4636 & ~n4951 ;
  buffer buf_n4955( .i (n4954), .o (n4955) );
  buffer buf_n4956( .i (n4955), .o (n4956) );
  buffer buf_n4952( .i (n4951), .o (n4952) );
  buffer buf_n4953( .i (n4952), .o (n4953) );
  assign n4957 = n4953 | n4955 ;
  buffer buf_n4958( .i (n4389), .o (n4958) );
  assign n4959 = ( n4956 & n4957 ) | ( n4956 & ~n4958 ) | ( n4957 & ~n4958 ) ;
  assign n4960 = ~n4817 & n4959 ;
  assign n4961 = n4468 & ~n4817 ;
  buffer buf_n4962( .i (n4204), .o (n4962) );
  buffer buf_n4963( .i (n4308), .o (n4963) );
  assign n4964 = ( n4636 & ~n4962 ) | ( n4636 & n4963 ) | ( ~n4962 & n4963 ) ;
  buffer buf_n4965( .i (n4964), .o (n4965) );
  buffer buf_n4966( .i (n4965), .o (n4966) );
  assign n4967 = n4819 & n4965 ;
  assign n4968 = ( ~n1048 & n4966 ) | ( ~n1048 & n4967 ) | ( n4966 & n4967 ) ;
  buffer buf_n4969( .i (n3765), .o (n4969) );
  buffer buf_n4970( .i (n4969), .o (n4970) );
  assign n4971 = ( ~n4817 & n4968 ) | ( ~n4817 & n4970 ) | ( n4968 & n4970 ) ;
  assign n4972 = ( n4960 & ~n4961 ) | ( n4960 & n4971 ) | ( ~n4961 & n4971 ) ;
  assign n4973 = n4887 & n4972 ;
  buffer buf_n4974( .i (n2277), .o (n4974) );
  assign n4975 = ( n46 & ~n4550 ) | ( n46 & n4974 ) | ( ~n4550 & n4974 ) ;
  buffer buf_n4976( .i (n4975), .o (n4976) );
  assign n4981 = ( ~n4307 & n4634 ) | ( ~n4307 & n4976 ) | ( n4634 & n4976 ) ;
  buffer buf_n4982( .i (n4981), .o (n4982) );
  buffer buf_n4983( .i (n4982), .o (n4983) );
  buffer buf_n4984( .i (n4983), .o (n4984) );
  buffer buf_n4985( .i (n4984), .o (n4985) );
  assign n4986 = ( n4075 & n4535 ) | ( n4075 & n4982 ) | ( n4535 & n4982 ) ;
  buffer buf_n4987( .i (n4986), .o (n4987) );
  buffer buf_n4988( .i (n4987), .o (n4988) );
  buffer buf_n4977( .i (n4976), .o (n4977) );
  buffer buf_n4978( .i (n4977), .o (n4978) );
  buffer buf_n4979( .i (n4978), .o (n4979) );
  buffer buf_n4980( .i (n4979), .o (n4980) );
  assign n4989 = n4980 & ~n4987 ;
  assign n4990 = ( n4985 & ~n4988 ) | ( n4985 & n4989 ) | ( ~n4988 & n4989 ) ;
  assign n4991 = n4821 & ~n4990 ;
  assign n4992 = n924 & n4816 ;
  assign n4993 = n4821 | n4992 ;
  assign n4994 = ~n4991 & n4993 ;
  assign n4995 = n4887 | n4994 ;
  assign n4996 = ( ~n4888 & n4973 ) | ( ~n4888 & n4995 ) | ( n4973 & n4995 ) ;
  assign n4997 = n4830 & n4996 ;
  buffer buf_n4554( .i (n4553), .o (n4554) );
  buffer buf_n4555( .i (n4554), .o (n4555) );
  buffer buf_n4556( .i (n4555), .o (n4556) );
  buffer buf_n4557( .i (n4556), .o (n4557) );
  assign n4998 = n4557 & n4820 ;
  assign n4999 = n4529 | n4556 ;
  assign n5000 = ( n4820 & ~n4958 ) | ( n4820 & n4999 ) | ( ~n4958 & n4999 ) ;
  assign n5001 = ~n4998 & n5000 ;
  buffer buf_n5002( .i (n4816), .o (n5002) );
  buffer buf_n5003( .i (n5002), .o (n5003) );
  buffer buf_n5004( .i (n4399), .o (n5004) );
  assign n5005 = ( n5001 & n5003 ) | ( n5001 & ~n5004 ) | ( n5003 & ~n5004 ) ;
  assign n5006 = n425 & ~n4969 ;
  buffer buf_n5007( .i (n4581), .o (n5007) );
  buffer buf_n5008( .i (n4571), .o (n5008) );
  assign n5009 = ( ~n424 & n5007 ) | ( ~n424 & n5008 ) | ( n5007 & n5008 ) ;
  assign n5010 = ( n1057 & n4969 ) | ( n1057 & ~n5009 ) | ( n4969 & ~n5009 ) ;
  assign n5011 = ( n4970 & n5006 ) | ( n4970 & ~n5010 ) | ( n5006 & ~n5010 ) ;
  assign n5012 = ( n5003 & n5004 ) | ( n5003 & ~n5011 ) | ( n5004 & ~n5011 ) ;
  assign n5013 = n5005 & ~n5012 ;
  buffer buf_n2860( .i (n2859), .o (n2860) );
  buffer buf_n2861( .i (n2860), .o (n2861) );
  buffer buf_n2862( .i (n2861), .o (n2862) );
  buffer buf_n2863( .i (n2862), .o (n2863) );
  buffer buf_n2864( .i (n2863), .o (n2864) );
  buffer buf_n2865( .i (n2864), .o (n2865) );
  assign n5014 = ( ~n926 & n2865 ) | ( ~n926 & n5003 ) | ( n2865 & n5003 ) ;
  assign n5015 = n927 & n5014 ;
  assign n5016 = n5013 | n5015 ;
  assign n5017 = ~n4830 & n5016 ;
  assign n5018 = n4997 | n5017 ;
  assign n5019 = ~n4460 & n5018 ;
  buffer buf_n5020( .i (n5019), .o (n5020) );
  buffer buf_n5021( .i (n5020), .o (n5021) );
  assign n5022 = n718 | n5020 ;
  assign n5023 = ( n4948 & n5021 ) | ( n4948 & n5022 ) | ( n5021 & n5022 ) ;
  assign n5024 = n180 & ~n5023 ;
  assign n5025 = ( ~n4535 & n4962 ) | ( ~n4535 & n4963 ) | ( n4962 & n4963 ) ;
  buffer buf_n5026( .i (n5025), .o (n5026) );
  buffer buf_n5027( .i (n5026), .o (n5027) );
  buffer buf_n5028( .i (n5027), .o (n5028) );
  buffer buf_n5029( .i (n5028), .o (n5029) );
  buffer buf_n5030( .i (n5029), .o (n5030) );
  assign n5031 = ( ~n4845 & n4898 ) | ( ~n4845 & n5030 ) | ( n4898 & n5030 ) ;
  assign n5032 = ( n4898 & n4901 ) | ( n4898 & ~n5030 ) | ( n4901 & ~n5030 ) ;
  assign n5033 = n5031 & ~n5032 ;
  buffer buf_n5034( .i (n5033), .o (n5034) );
  buffer buf_n5035( .i (n5034), .o (n5035) );
  assign n5036 = ( n3974 & n4831 ) | ( n3974 & ~n5034 ) | ( n4831 & ~n5034 ) ;
  assign n5037 = n541 & n4758 ;
  assign n5038 = n612 & n5037 ;
  assign n5039 = n4831 & n5038 ;
  assign n5040 = ( n5035 & n5036 ) | ( n5035 & n5039 ) | ( n5036 & n5039 ) ;
  buffer buf_n5041( .i (n4758), .o (n5041) );
  assign n5042 = ( n4776 & n4830 ) | ( n4776 & n5041 ) | ( n4830 & n5041 ) ;
  buffer buf_n5043( .i (n4535), .o (n5043) );
  assign n5044 = ( n4325 & n4818 ) | ( n4325 & n5043 ) | ( n4818 & n5043 ) ;
  assign n5045 = ( n4487 & ~n5007 ) | ( n4487 & n5044 ) | ( ~n5007 & n5044 ) ;
  buffer buf_n5046( .i (n5045), .o (n5046) );
  assign n5049 = n4399 & ~n5046 ;
  buffer buf_n5050( .i (n5049), .o (n5050) );
  buffer buf_n5051( .i (n5050), .o (n5051) );
  buffer buf_n5047( .i (n5046), .o (n5047) );
  buffer buf_n5048( .i (n5047), .o (n5048) );
  assign n5052 = n5048 | n5050 ;
  assign n5053 = ( ~n4434 & n5051 ) | ( ~n4434 & n5052 ) | ( n5051 & n5052 ) ;
  assign n5054 = n4844 | n4898 ;
  buffer buf_n5055( .i (n5054), .o (n5055) );
  buffer buf_n5057( .i (n4383), .o (n5057) );
  assign n5058 = ( n5053 & n5055 ) | ( n5053 & n5057 ) | ( n5055 & n5057 ) ;
  assign n5059 = ~n5042 & n5058 ;
  buffer buf_n5060( .i (n5059), .o (n5060) );
  assign n5061 = ( ~n4854 & n5040 ) | ( ~n4854 & n5060 ) | ( n5040 & n5060 ) ;
  assign n5062 = n3765 & ~n4819 ;
  buffer buf_n5063( .i (n5062), .o (n5063) );
  buffer buf_n5064( .i (n5063), .o (n5064) );
  buffer buf_n5070( .i (n4409), .o (n5070) );
  assign n5071 = ( n4113 & n5064 ) | ( n4113 & n5070 ) | ( n5064 & n5070 ) ;
  assign n5072 = ( n5003 & n5064 ) | ( n5003 & n5070 ) | ( n5064 & n5070 ) ;
  assign n5073 = ( n1947 & n5071 ) | ( n1947 & ~n5072 ) | ( n5071 & ~n5072 ) ;
  buffer buf_n5074( .i (n4901), .o (n5074) );
  assign n5075 = ~n5073 & n5074 ;
  assign n5076 = n4655 & ~n4816 ;
  buffer buf_n5077( .i (n5076), .o (n5077) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  assign n5081 = n2260 & n5002 ;
  buffer buf_n5082( .i (n5002), .o (n5082) );
  assign n5083 = ( n5077 & ~n5081 ) | ( n5077 & n5082 ) | ( ~n5081 & n5082 ) ;
  assign n5084 = n4845 & ~n5083 ;
  assign n5085 = n5074 | n5084 ;
  assign n5086 = ~n5075 & n5085 ;
  assign n5087 = n4907 & ~n5086 ;
  assign n5088 = ( n664 & ~n4332 ) | ( n664 & n4655 ) | ( ~n4332 & n4655 ) ;
  buffer buf_n5089( .i (n5088), .o (n5089) );
  buffer buf_n5090( .i (n5089), .o (n5090) );
  buffer buf_n5091( .i (n5090), .o (n5091) );
  assign n5092 = ( n5004 & ~n5082 ) | ( n5004 & n5089 ) | ( ~n5082 & n5089 ) ;
  buffer buf_n5093( .i (n5070), .o (n5093) );
  assign n5094 = ( n3883 & ~n5092 ) | ( n3883 & n5093 ) | ( ~n5092 & n5093 ) ;
  assign n5095 = ~n5091 & n5094 ;
  buffer buf_n5096( .i (n4826), .o (n5096) );
  assign n5097 = n5095 & n5096 ;
  assign n5098 = n4907 | n5097 ;
  assign n5099 = ~n5087 & n5098 ;
  assign n5100 = ( n4854 & n5060 ) | ( n4854 & n5099 ) | ( n5060 & n5099 ) ;
  assign n5101 = n5061 | n5100 ;
  assign n5102 = ~n3416 & n5101 ;
  assign n5103 = n180 | n5102 ;
  assign n5104 = ~n5024 & n5103 ;
  assign n5105 = n432 & n805 ;
  assign n5106 = ( n2127 & n4768 ) | ( n2127 & n5105 ) | ( n4768 & n5105 ) ;
  assign n5107 = ~n4769 & n5106 ;
  buffer buf_n5108( .i (n5107), .o (n5108) );
  buffer buf_n5109( .i (n5108), .o (n5109) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n5110( .i (n4831), .o (n5110) );
  assign n5111 = ( n662 & n4789 ) | ( n662 & n5110 ) | ( n4789 & n5110 ) ;
  buffer buf_n5112( .i (n4789), .o (n5112) );
  assign n5113 = n5111 & ~n5112 ;
  assign n5114 = ( ~n3400 & n4769 ) | ( ~n3400 & n5113 ) | ( n4769 & n5113 ) ;
  buffer buf_n5115( .i (n4491), .o (n5115) );
  buffer buf_n5116( .i (n5115), .o (n5116) );
  assign n5117 = ( n4815 & n5008 ) | ( n4815 & ~n5116 ) | ( n5008 & ~n5116 ) ;
  buffer buf_n5118( .i (n4815), .o (n5118) );
  assign n5119 = ( ~n4969 & n5117 ) | ( ~n4969 & n5118 ) | ( n5117 & n5118 ) ;
  buffer buf_n5120( .i (n5119), .o (n5120) );
  assign n5123 = n5082 & ~n5120 ;
  buffer buf_n5124( .i (n5123), .o (n5124) );
  buffer buf_n5125( .i (n5124), .o (n5125) );
  buffer buf_n5121( .i (n5120), .o (n5121) );
  buffer buf_n5122( .i (n5121), .o (n5122) );
  assign n5126 = n5122 | n5124 ;
  assign n5127 = ( ~n4776 & n5125 ) | ( ~n4776 & n5126 ) | ( n5125 & n5126 ) ;
  buffer buf_n5128( .i (n5127), .o (n5128) );
  buffer buf_n5129( .i (n5128), .o (n5129) );
  assign n5130 = ( ~n4789 & n5110 ) | ( ~n4789 & n5128 ) | ( n5110 & n5128 ) ;
  assign n5131 = ( n4288 & ~n4634 ) | ( n4288 & n4949 ) | ( ~n4634 & n4949 ) ;
  buffer buf_n5132( .i (n5131), .o (n5132) );
  buffer buf_n5133( .i (n5132), .o (n5133) );
  assign n5134 = ~n4491 & n5132 ;
  buffer buf_n5135( .i (n4635), .o (n5135) );
  buffer buf_n5136( .i (n5135), .o (n5136) );
  assign n5137 = ( n5133 & n5134 ) | ( n5133 & n5136 ) | ( n5134 & n5136 ) ;
  buffer buf_n5138( .i (n5137), .o (n5138) );
  buffer buf_n5139( .i (n5138), .o (n5139) );
  buffer buf_n5140( .i (n5139), .o (n5140) );
  buffer buf_n5141( .i (n5140), .o (n5141) );
  buffer buf_n5142( .i (n5141), .o (n5142) );
  buffer buf_n5143( .i (n5142), .o (n5143) );
  buffer buf_n5145( .i (n4775), .o (n5145) );
  assign n5146 = n5143 & ~n5145 ;
  assign n5147 = ~n4094 & n5146 ;
  assign n5148 = ~n5110 & n5147 ;
  assign n5149 = ( n5129 & ~n5130 ) | ( n5129 & n5148 ) | ( ~n5130 & n5148 ) ;
  buffer buf_n5150( .i (n4854), .o (n5150) );
  assign n5151 = n5149 & ~n5150 ;
  assign n5152 = ( ~n4770 & n5114 ) | ( ~n4770 & n5151 ) | ( n5114 & n5151 ) ;
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n5153( .i (n716), .o (n5153) );
  assign n5154 = n2046 & n5153 ;
  assign n5155 = n379 & n5154 ;
  buffer buf_n5156( .i (n5155), .o (n5156) );
  assign n5157 = ( ~n5108 & n5152 ) | ( ~n5108 & n5156 ) | ( n5152 & n5156 ) ;
  assign n5158 = n4944 & ~n5156 ;
  assign n5159 = ( n5109 & n5157 ) | ( n5109 & ~n5158 ) | ( n5157 & ~n5158 ) ;
  assign n5160 = n5104 | n5159 ;
  assign n5161 = ( ~n4860 & n4947 ) | ( ~n4860 & n5160 ) | ( n4947 & n5160 ) ;
  assign n5162 = n4861 | n5161 ;
  buffer buf_n5163( .i (n47), .o (n5163) );
  buffer buf_n5164( .i (n5163), .o (n5164) );
  buffer buf_n5165( .i (n4288), .o (n5165) );
  assign n5166 = n5164 & ~n5165 ;
  buffer buf_n5167( .i (n5166), .o (n5167) );
  buffer buf_n5168( .i (n5167), .o (n5168) );
  buffer buf_n5169( .i (n5168), .o (n5169) );
  buffer buf_n5170( .i (n5169), .o (n5170) );
  buffer buf_n5171( .i (n5170), .o (n5171) );
  buffer buf_n5172( .i (n5171), .o (n5172) );
  buffer buf_n5173( .i (n5172), .o (n5173) );
  buffer buf_n5174( .i (n5173), .o (n5174) );
  buffer buf_n5175( .i (n5174), .o (n5175) );
  buffer buf_n5176( .i (n5175), .o (n5176) );
  buffer buf_n5177( .i (n5176), .o (n5177) );
  buffer buf_n5178( .i (n4773), .o (n5178) );
  buffer buf_n5179( .i (n5178), .o (n5179) );
  assign n5180 = ( ~n4911 & n5177 ) | ( ~n4911 & n5179 ) | ( n5177 & n5179 ) ;
  buffer buf_n5181( .i (n4938), .o (n5181) );
  assign n5182 = ( ~n5177 & n5179 ) | ( ~n5177 & n5181 ) | ( n5179 & n5181 ) ;
  assign n5183 = ( n178 & n5180 ) | ( n178 & ~n5182 ) | ( n5180 & ~n5182 ) ;
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n5184( .i (n5145), .o (n5184) );
  assign n5185 = ( n827 & ~n4873 ) | ( n827 & n5184 ) | ( ~n4873 & n5184 ) ;
  assign n5186 = ~n4938 & n5185 ;
  buffer buf_n5187( .i (n5186), .o (n5187) );
  buffer buf_n5188( .i (n5187), .o (n5188) );
  assign n5189 = n236 | n5187 ;
  assign n5190 = ( n5183 & n5188 ) | ( n5183 & n5189 ) | ( n5188 & n5189 ) ;
  assign n5191 = n92 | n5190 ;
  buffer buf_n4885( .i (n4884), .o (n4885) );
  buffer buf_n4886( .i (n4885), .o (n4886) );
  assign n5192 = ( n3421 & n4886 ) | ( n3421 & ~n5181 ) | ( n4886 & ~n5181 ) ;
  assign n5193 = ( n4885 & n4938 ) | ( n4885 & ~n5178 ) | ( n4938 & ~n5178 ) ;
  buffer buf_n5194( .i (n3418), .o (n5194) );
  assign n5195 = ( n3421 & ~n5193 ) | ( n3421 & n5194 ) | ( ~n5193 & n5194 ) ;
  assign n5196 = ~n5192 & n5195 ;
  assign n5197 = ~n3416 & n5196 ;
  assign n5198 = n92 & ~n5197 ;
  assign n5199 = n5191 & ~n5198 ;
  buffer buf_n5200( .i (n5199), .o (n5200) );
  buffer buf_n5201( .i (n5200), .o (n5201) );
  assign n5202 = ( n670 & ~n1806 ) | ( n670 & n2611 ) | ( ~n1806 & n2611 ) ;
  buffer buf_n5203( .i (n5202), .o (n5203) );
  buffer buf_n5204( .i (n5203), .o (n5204) );
  buffer buf_n5205( .i (n5204), .o (n5205) );
  buffer buf_n5206( .i (n5205), .o (n5206) );
  buffer buf_n5207( .i (n5206), .o (n5207) );
  buffer buf_n5208( .i (n5207), .o (n5208) );
  buffer buf_n5209( .i (n5208), .o (n5209) );
  buffer buf_n5210( .i (n5209), .o (n5210) );
  buffer buf_n5211( .i (n5210), .o (n5211) );
  buffer buf_n5212( .i (n5211), .o (n5212) );
  assign n5213 = n5200 & ~n5212 ;
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n3190( .i (n3189), .o (n3190) );
  buffer buf_n3191( .i (n3190), .o (n3191) );
  buffer buf_n3192( .i (n3191), .o (n3192) );
  buffer buf_n3193( .i (n3192), .o (n3193) );
  buffer buf_n3194( .i (n3193), .o (n3194) );
  buffer buf_n3195( .i (n3194), .o (n3195) );
  buffer buf_n3196( .i (n3195), .o (n3196) );
  buffer buf_n3197( .i (n3196), .o (n3197) );
  buffer buf_n3198( .i (n3197), .o (n3198) );
  buffer buf_n3199( .i (n3198), .o (n3199) );
  buffer buf_n3200( .i (n3199), .o (n3200) );
  assign n5214 = ( ~n3548 & n4558 ) | ( ~n3548 & n5164 ) | ( n4558 & n5164 ) ;
  buffer buf_n5215( .i (n5214), .o (n5215) );
  buffer buf_n5216( .i (n5215), .o (n5216) );
  buffer buf_n5217( .i (n5216), .o (n5217) );
  buffer buf_n5218( .i (n5217), .o (n5218) );
  buffer buf_n5219( .i (n5218), .o (n5219) );
  buffer buf_n5220( .i (n5219), .o (n5220) );
  buffer buf_n5221( .i (n5220), .o (n5221) );
  buffer buf_n5222( .i (n5221), .o (n5222) );
  buffer buf_n5223( .i (n5222), .o (n5223) );
  assign n5224 = n3200 & ~n5223 ;
  buffer buf_n5225( .i (n4610), .o (n5225) );
  assign n5226 = n5224 | n5225 ;
  buffer buf_n4584( .i (n4583), .o (n4584) );
  buffer buf_n4585( .i (n4584), .o (n4585) );
  buffer buf_n4586( .i (n4585), .o (n4586) );
  buffer buf_n4587( .i (n4586), .o (n4587) );
  buffer buf_n4588( .i (n4587), .o (n4588) );
  assign n5227 = n4588 | n5041 ;
  assign n5228 = n5184 | n5227 ;
  assign n5229 = n5225 & n5228 ;
  assign n5230 = n5226 & ~n5229 ;
  buffer buf_n5231( .i (n5230), .o (n5231) );
  buffer buf_n5232( .i (n5231), .o (n5232) );
  buffer buf_n3601( .i (n3600), .o (n3601) );
  buffer buf_n3602( .i (n3601), .o (n3602) );
  buffer buf_n3603( .i (n3602), .o (n3603) );
  buffer buf_n3604( .i (n3603), .o (n3604) );
  buffer buf_n3605( .i (n3604), .o (n3605) );
  buffer buf_n3606( .i (n3605), .o (n3606) );
  buffer buf_n3607( .i (n3606), .o (n3607) );
  buffer buf_n3608( .i (n3607), .o (n3608) );
  assign n5233 = n3608 & n5231 ;
  assign n5234 = n519 & n709 ;
  assign n5235 = ( n403 & ~n932 ) | ( n403 & n5234 ) | ( ~n932 & n5234 ) ;
  assign n5236 = n933 & n5235 ;
  buffer buf_n5237( .i (n4558), .o (n5237) );
  buffer buf_n5238( .i (n4949), .o (n5238) );
  buffer buf_n5239( .i (n5238), .o (n5239) );
  assign n5240 = ( n4963 & ~n5237 ) | ( n4963 & n5239 ) | ( ~n5237 & n5239 ) ;
  buffer buf_n5241( .i (n5240), .o (n5241) );
  buffer buf_n5242( .i (n5241), .o (n5242) );
  buffer buf_n5243( .i (n5242), .o (n5243) );
  buffer buf_n5244( .i (n5243), .o (n5244) );
  assign n5246 = ( n4783 & ~n5004 ) | ( n4783 & n5244 ) | ( ~n5004 & n5244 ) ;
  assign n5247 = ~n4409 & n5243 ;
  assign n5248 = ( ~n3882 & n5244 ) | ( ~n3882 & n5247 ) | ( n5244 & n5247 ) ;
  assign n5249 = n5246 | n5248 ;
  assign n5250 = n4775 & n5249 ;
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  assign n5251 = n553 | n4887 ;
  assign n5252 = ~n4775 & n5251 ;
  assign n5253 = n5250 | n5252 ;
  assign n5254 = n4907 & ~n5253 ;
  assign n5255 = ~n44 & n246 ;
  buffer buf_n5256( .i (n5255), .o (n5256) );
  buffer buf_n5257( .i (n5256), .o (n5257) );
  buffer buf_n5258( .i (n5257), .o (n5258) );
  buffer buf_n5259( .i (n5258), .o (n5259) );
  buffer buf_n5260( .i (n5259), .o (n5260) );
  buffer buf_n5261( .i (n5260), .o (n5261) );
  buffer buf_n5262( .i (n5261), .o (n5262) );
  buffer buf_n5263( .i (n5262), .o (n5263) );
  buffer buf_n5264( .i (n5263), .o (n5264) );
  buffer buf_n5265( .i (n5264), .o (n5265) );
  buffer buf_n5266( .i (n5265), .o (n5266) );
  buffer buf_n5267( .i (n5266), .o (n5267) );
  assign n5268 = ( n1363 & n4655 ) | ( n1363 & n5263 ) | ( n4655 & n5263 ) ;
  buffer buf_n5269( .i (n5268), .o (n5269) );
  buffer buf_n5270( .i (n5269), .o (n5270) );
  buffer buf_n5271( .i (n5270), .o (n5271) );
  buffer buf_n5272( .i (n4411), .o (n5272) );
  assign n5273 = ( ~n5070 & n5269 ) | ( ~n5070 & n5272 ) | ( n5269 & n5272 ) ;
  assign n5274 = ( ~n4901 & n5266 ) | ( ~n4901 & n5273 ) | ( n5266 & n5273 ) ;
  assign n5275 = ( ~n5267 & n5271 ) | ( ~n5267 & n5274 ) | ( n5271 & n5274 ) ;
  assign n5276 = ~n552 & n834 ;
  buffer buf_n5277( .i (n5276), .o (n5277) );
  buffer buf_n5278( .i (n5277), .o (n5278) );
  assign n5279 = n4738 | n5277 ;
  assign n5280 = ( n5275 & n5278 ) | ( n5275 & n5279 ) | ( n5278 & n5279 ) ;
  buffer buf_n5281( .i (n5041), .o (n5281) );
  assign n5282 = n5280 | n5281 ;
  assign n5283 = ( ~n4445 & n5254 ) | ( ~n4445 & n5282 ) | ( n5254 & n5282 ) ;
  buffer buf_n5284( .i (n4096), .o (n5284) );
  assign n5285 = ( ~n4911 & n5283 ) | ( ~n4911 & n5284 ) | ( n5283 & n5284 ) ;
  buffer buf_n5286( .i (n5043), .o (n5286) );
  buffer buf_n5287( .i (n5286), .o (n5287) );
  assign n5288 = ~n3011 & n5287 ;
  assign n5289 = ~n4409 & n5288 ;
  buffer buf_n5290( .i (n5289), .o (n5290) );
  buffer buf_n5291( .i (n5290), .o (n5291) );
  buffer buf_n5292( .i (n5272), .o (n5292) );
  assign n5293 = n5290 & ~n5292 ;
  buffer buf_n5294( .i (n4338), .o (n5294) );
  buffer buf_n5295( .i (n5294), .o (n5295) );
  assign n5296 = n396 & n5295 ;
  assign n5297 = ~n334 & n5296 ;
  buffer buf_n5298( .i (n3187), .o (n5298) );
  buffer buf_n5299( .i (n5298), .o (n5299) );
  buffer buf_n5300( .i (n3002), .o (n5300) );
  assign n5301 = ( n4307 & n5299 ) | ( n4307 & ~n5300 ) | ( n5299 & ~n5300 ) ;
  buffer buf_n5302( .i (n5301), .o (n5302) );
  assign n5307 = ( ~n5237 & n5239 ) | ( ~n5237 & n5302 ) | ( n5239 & n5302 ) ;
  buffer buf_n5308( .i (n5307), .o (n5308) );
  buffer buf_n5309( .i (n5308), .o (n5309) );
  buffer buf_n5310( .i (n5309), .o (n5310) );
  buffer buf_n5311( .i (n5310), .o (n5311) );
  assign n5312 = ( n4487 & ~n5008 ) | ( n4487 & n5308 ) | ( ~n5008 & n5308 ) ;
  buffer buf_n5313( .i (n5312), .o (n5313) );
  buffer buf_n5314( .i (n5313), .o (n5314) );
  buffer buf_n5303( .i (n5302), .o (n5303) );
  buffer buf_n5304( .i (n5303), .o (n5304) );
  buffer buf_n5305( .i (n5304), .o (n5305) );
  buffer buf_n5306( .i (n5305), .o (n5306) );
  assign n5315 = ~n5306 & n5313 ;
  assign n5316 = ( ~n5311 & n5314 ) | ( ~n5311 & n5315 ) | ( n5314 & n5315 ) ;
  assign n5317 = n5297 | n5316 ;
  assign n5318 = ( n5291 & ~n5293 ) | ( n5291 & n5317 ) | ( ~n5293 & n5317 ) ;
  assign n5319 = n5145 | n5318 ;
  buffer buf_n5320( .i (n4399), .o (n5320) );
  assign n5321 = n5272 & ~n5320 ;
  buffer buf_n5322( .i (n4516), .o (n5322) );
  assign n5323 = ( n1479 & ~n4970 ) | ( n1479 & n5322 ) | ( ~n4970 & n5322 ) ;
  assign n5324 = n1480 | n5323 ;
  assign n5325 = ~n5321 & n5324 ;
  buffer buf_n5326( .i (n5093), .o (n5326) );
  assign n5327 = n5325 & ~n5326 ;
  assign n5328 = n5145 & ~n5327 ;
  assign n5329 = n5319 & ~n5328 ;
  assign n5330 = ( n3583 & ~n4332 ) | ( n3583 & n5294 ) | ( ~n4332 & n5294 ) ;
  buffer buf_n5331( .i (n5330), .o (n5331) );
  assign n5334 = n5320 & n5331 ;
  buffer buf_n5335( .i (n5334), .o (n5335) );
  buffer buf_n5336( .i (n5335), .o (n5336) );
  buffer buf_n5332( .i (n5331), .o (n5332) );
  buffer buf_n5333( .i (n5332), .o (n5333) );
  assign n5337 = n5333 & ~n5335 ;
  assign n5338 = ( n4719 & ~n5336 ) | ( n4719 & n5337 ) | ( ~n5336 & n5337 ) ;
  assign n5339 = ( n4773 & ~n5281 ) | ( n4773 & n5338 ) | ( ~n5281 & n5338 ) ;
  assign n5340 = ( n402 & ~n5329 ) | ( n402 & n5339 ) | ( ~n5329 & n5339 ) ;
  assign n5341 = ( n4911 & n5284 ) | ( n4911 & n5340 ) | ( n5284 & n5340 ) ;
  assign n5342 = n5285 & ~n5341 ;
  assign n5343 = n5236 | n5342 ;
  assign n5344 = ( n5232 & ~n5233 ) | ( n5232 & n5343 ) | ( ~n5233 & n5343 ) ;
  assign n5345 = n93 | n5344 ;
  buffer buf_n4341( .i (n4340), .o (n4341) );
  buffer buf_n4342( .i (n4341), .o (n4342) );
  buffer buf_n4343( .i (n4342), .o (n4343) );
  buffer buf_n4344( .i (n4343), .o (n4344) );
  buffer buf_n4345( .i (n4344), .o (n4345) );
  buffer buf_n4346( .i (n4345), .o (n4346) );
  buffer buf_n4347( .i (n4346), .o (n4347) );
  buffer buf_n4348( .i (n4347), .o (n4348) );
  buffer buf_n4349( .i (n4348), .o (n4349) );
  buffer buf_n5346( .i (n5237), .o (n5346) );
  buffer buf_n5347( .i (n4963), .o (n5347) );
  assign n5348 = ( n1161 & ~n5346 ) | ( n1161 & n5347 ) | ( ~n5346 & n5347 ) ;
  buffer buf_n5349( .i (n5348), .o (n5349) );
  buffer buf_n5350( .i (n5349), .o (n5350) );
  buffer buf_n5351( .i (n5350), .o (n5351) );
  buffer buf_n5352( .i (n5351), .o (n5352) );
  assign n5353 = ( n4654 & n5287 ) | ( n4654 & n5349 ) | ( n5287 & n5349 ) ;
  buffer buf_n5354( .i (n5353), .o (n5354) );
  buffer buf_n5355( .i (n5354), .o (n5355) );
  assign n5356 = ~n1165 & n5354 ;
  assign n5357 = ( ~n5352 & n5355 ) | ( ~n5352 & n5356 ) | ( n5355 & n5356 ) ;
  buffer buf_n5358( .i (n5082), .o (n5358) );
  buffer buf_n5359( .i (n5358), .o (n5359) );
  assign n5360 = n5357 | n5359 ;
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  assign n5361 = n895 | n5292 ;
  assign n5362 = n5359 & n5361 ;
  assign n5363 = n5360 & ~n5362 ;
  assign n5364 = n5281 & n5363 ;
  buffer buf_n5365( .i (n4215), .o (n5365) );
  assign n5366 = ( n2188 & n4974 ) | ( n2188 & ~n5365 ) | ( n4974 & ~n5365 ) ;
  buffer buf_n5367( .i (n5366), .o (n5367) );
  assign n5373 = ( n4288 & n5163 ) | ( n4288 & ~n5367 ) | ( n5163 & ~n5367 ) ;
  buffer buf_n5374( .i (n5373), .o (n5374) );
  buffer buf_n5375( .i (n5374), .o (n5375) );
  buffer buf_n5376( .i (n5375), .o (n5376) );
  buffer buf_n5377( .i (n5376), .o (n5377) );
  buffer buf_n5378( .i (n5377), .o (n5378) );
  buffer buf_n5368( .i (n5367), .o (n5368) );
  buffer buf_n5369( .i (n5368), .o (n5369) );
  buffer buf_n5370( .i (n5369), .o (n5370) );
  buffer buf_n5379( .i (n5165), .o (n5379) );
  assign n5380 = ( n5239 & n5374 ) | ( n5239 & ~n5379 ) | ( n5374 & ~n5379 ) ;
  assign n5381 = n5370 & n5380 ;
  buffer buf_n5382( .i (n5381), .o (n5382) );
  buffer buf_n5383( .i (n5382), .o (n5383) );
  assign n5384 = n5118 & ~n5382 ;
  assign n5385 = ( n5378 & n5383 ) | ( n5378 & ~n5384 ) | ( n5383 & ~n5384 ) ;
  assign n5386 = n5320 & n5385 ;
  buffer buf_n5387( .i (n5386), .o (n5387) );
  buffer buf_n5388( .i (n5387), .o (n5388) );
  buffer buf_n5389( .i (n5164), .o (n5389) );
  assign n5390 = ( ~n5237 & n5239 ) | ( ~n5237 & n5389 ) | ( n5239 & n5389 ) ;
  buffer buf_n5391( .i (n5299), .o (n5391) );
  buffer buf_n5392( .i (n5391), .o (n5392) );
  buffer buf_n5393( .i (n4308), .o (n5393) );
  assign n5394 = ( ~n5389 & n5392 ) | ( ~n5389 & n5393 ) | ( n5392 & n5393 ) ;
  assign n5395 = n5390 | n5394 ;
  buffer buf_n5396( .i (n5395), .o (n5396) );
  buffer buf_n5397( .i (n5396), .o (n5397) );
  buffer buf_n5398( .i (n5397), .o (n5398) );
  buffer buf_n5399( .i (n5398), .o (n5399) );
  buffer buf_n5400( .i (n5399), .o (n5400) );
  assign n5401 = ~n5387 & n5400 ;
  assign n5402 = ( n4386 & n5388 ) | ( n4386 & ~n5401 ) | ( n5388 & ~n5401 ) ;
  assign n5403 = n5281 | n5402 ;
  buffer buf_n5404( .i (n5041), .o (n5404) );
  buffer buf_n5405( .i (n5404), .o (n5405) );
  assign n5406 = ( n5364 & n5403 ) | ( n5364 & ~n5405 ) | ( n5403 & ~n5405 ) ;
  assign n5407 = n3854 & ~n5406 ;
  assign n5408 = n4324 & n5115 ;
  buffer buf_n5409( .i (n5408), .o (n5409) );
  buffer buf_n5410( .i (n5409), .o (n5410) );
  buffer buf_n5411( .i (n5410), .o (n5411) );
  buffer buf_n5412( .i (n5411), .o (n5412) );
  buffer buf_n5413( .i (n5412), .o (n5413) );
  assign n5414 = n4838 & n5272 ;
  assign n5415 = ( ~n3883 & n5358 ) | ( ~n3883 & n5414 ) | ( n5358 & n5414 ) ;
  assign n5416 = ( n2633 & ~n5413 ) | ( n2633 & n5415 ) | ( ~n5413 & n5415 ) ;
  buffer buf_n5417( .i (n4758), .o (n5417) );
  assign n5418 = n5416 & n5417 ;
  buffer buf_n4438( .i (n4437), .o (n4438) );
  buffer buf_n4439( .i (n4438), .o (n4439) );
  buffer buf_n5419( .i (n4738), .o (n5419) );
  assign n5420 = ( n4439 & n5417 ) | ( n4439 & ~n5419 ) | ( n5417 & ~n5419 ) ;
  assign n5421 = ( ~n661 & n5418 ) | ( ~n661 & n5420 ) | ( n5418 & n5420 ) ;
  assign n5422 = n4721 & n5421 ;
  assign n5423 = n3854 | n5422 ;
  assign n5424 = ~n5407 & n5423 ;
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n5425( .i (n5359), .o (n5425) );
  assign n5426 = ( n1615 & n4719 ) | ( n1615 & ~n5425 ) | ( n4719 & ~n5425 ) ;
  buffer buf_n5427( .i (n4970), .o (n5427) );
  buffer buf_n5428( .i (n5427), .o (n5428) );
  buffer buf_n5429( .i (n5428), .o (n5429) );
  assign n5430 = ( ~n1614 & n5074 ) | ( ~n1614 & n5429 ) | ( n5074 & n5429 ) ;
  assign n5431 = ( n5417 & ~n5425 ) | ( n5417 & n5430 ) | ( ~n5425 & n5430 ) ;
  assign n5432 = ~n5426 & n5431 ;
  assign n5433 = n4096 & ~n5432 ;
  buffer buf_n5056( .i (n5055), .o (n5056) );
  assign n5434 = n280 & ~n5056 ;
  buffer buf_n5435( .i (n4387), .o (n5435) );
  assign n5436 = n5434 | n5435 ;
  assign n5437 = ~n5433 & n5436 ;
  assign n5438 = ( n3855 & ~n5150 ) | ( n3855 & n5437 ) | ( ~n5150 & n5437 ) ;
  assign n5439 = ( ~n4349 & n5424 ) | ( ~n4349 & n5438 ) | ( n5424 & n5438 ) ;
  assign n5440 = ~n4944 & n5439 ;
  assign n5441 = n93 & ~n5440 ;
  assign n5442 = n5345 & ~n5441 ;
  assign n5443 = ( n5043 & n5136 ) | ( n5043 & ~n5346 ) | ( n5136 & ~n5346 ) ;
  buffer buf_n5444( .i (n5443), .o (n5444) );
  buffer buf_n5445( .i (n5444), .o (n5445) );
  assign n5452 = ( n5002 & n5322 ) | ( n5002 & n5445 ) | ( n5322 & n5445 ) ;
  buffer buf_n5453( .i (n5452), .o (n5453) );
  buffer buf_n5454( .i (n5453), .o (n5454) );
  buffer buf_n5455( .i (n5454), .o (n5455) );
  buffer buf_n5446( .i (n5445), .o (n5446) );
  buffer buf_n5447( .i (n5446), .o (n5447) );
  buffer buf_n5448( .i (n5447), .o (n5448) );
  assign n5456 = ( n5292 & n5428 ) | ( n5292 & ~n5453 ) | ( n5428 & ~n5453 ) ;
  assign n5457 = n5448 & n5456 ;
  assign n5458 = ( n5425 & ~n5455 ) | ( n5425 & n5457 ) | ( ~n5455 & n5457 ) ;
  buffer buf_n5459( .i (n5096), .o (n5459) );
  assign n5460 = ~n5458 & n5459 ;
  assign n5461 = ~n1472 & n5292 ;
  buffer buf_n5462( .i (n4835), .o (n5462) );
  buffer buf_n5463( .i (n5462), .o (n5463) );
  buffer buf_n5464( .i (n5463), .o (n5464) );
  assign n5465 = ( ~n1473 & n5461 ) | ( ~n1473 & n5464 ) | ( n5461 & n5464 ) ;
  assign n5466 = n5425 & n5465 ;
  assign n5467 = n5459 | n5466 ;
  assign n5468 = ~n5460 & n5467 ;
  assign n5469 = n3854 & ~n5468 ;
  buffer buf_n5470( .i (n5118), .o (n5470) );
  assign n5471 = ( ~n3950 & n5322 ) | ( ~n3950 & n5470 ) | ( n5322 & n5470 ) ;
  buffer buf_n5472( .i (n5471), .o (n5472) );
  buffer buf_n5473( .i (n5472), .o (n5473) );
  buffer buf_n5474( .i (n5473), .o (n5474) );
  buffer buf_n5475( .i (n5474), .o (n5475) );
  assign n5476 = ( n4845 & n5463 ) | ( n4845 & ~n5472 ) | ( n5463 & ~n5472 ) ;
  buffer buf_n5477( .i (n5476), .o (n5477) );
  buffer buf_n5478( .i (n5477), .o (n5478) );
  assign n5479 = ~n3954 & n5477 ;
  assign n5480 = ( n5475 & n5478 ) | ( n5475 & n5479 ) | ( n5478 & n5479 ) ;
  assign n5481 = ~n3418 & n5480 ;
  buffer buf_n5482( .i (n5110), .o (n5482) );
  assign n5483 = n5481 | n5482 ;
  assign n5484 = ~n5469 & n5483 ;
  buffer buf_n5485( .i (n4912), .o (n5485) );
  assign n5486 = n5484 | n5485 ;
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n5487( .i (n402), .o (n5487) );
  assign n5488 = ~n2101 & n5487 ;
  assign n5489 = ~n316 & n5488 ;
  assign n5490 = n5485 & ~n5489 ;
  assign n5491 = n5486 & ~n5490 ;
  assign n5492 = n181 & n5491 ;
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n5493( .i (n4821), .o (n5493) );
  buffer buf_n5494( .i (n5493), .o (n5494) );
  buffer buf_n5495( .i (n5322), .o (n5495) );
  buffer buf_n5496( .i (n5495), .o (n5496) );
  assign n5497 = ( n5093 & n5494 ) | ( n5093 & ~n5496 ) | ( n5494 & ~n5496 ) ;
  buffer buf_n5498( .i (n5497), .o (n5498) );
  buffer buf_n5499( .i (n5498), .o (n5499) );
  buffer buf_n5500( .i (n5499), .o (n5500) );
  buffer buf_n5501( .i (n5500), .o (n5501) );
  assign n5502 = n5057 & ~n5498 ;
  buffer buf_n5503( .i (n5502), .o (n5503) );
  buffer buf_n5504( .i (n5503), .o (n5504) );
  buffer buf_n5505( .i (n5184), .o (n5505) );
  buffer buf_n5506( .i (n5459), .o (n5506) );
  assign n5507 = ( n5503 & n5505 ) | ( n5503 & n5506 ) | ( n5505 & n5506 ) ;
  assign n5508 = ( ~n5501 & n5504 ) | ( ~n5501 & n5507 ) | ( n5504 & n5507 ) ;
  assign n5509 = ( ~n1201 & n4912 ) | ( ~n1201 & n5508 ) | ( n4912 & n5508 ) ;
  buffer buf_n5510( .i (n708), .o (n5510) );
  assign n5511 = ( n4346 & n5506 ) | ( n4346 & n5510 ) | ( n5506 & n5510 ) ;
  assign n5512 = ~n5112 & n5511 ;
  assign n5513 = ~n1201 & n5512 ;
  assign n5514 = ( ~n5485 & n5509 ) | ( ~n5485 & n5513 ) | ( n5509 & n5513 ) ;
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n5515( .i (n4572), .o (n5515) );
  assign n5516 = n394 & ~n5515 ;
  buffer buf_n5517( .i (n5516), .o (n5517) );
  buffer buf_n5518( .i (n5517), .o (n5518) );
  buffer buf_n5519( .i (n5518), .o (n5519) );
  buffer buf_n5520( .i (n5519), .o (n5520) );
  buffer buf_n5521( .i (n5520), .o (n5521) );
  buffer buf_n5522( .i (n5521), .o (n5522) );
  buffer buf_n5523( .i (n5522), .o (n5523) );
  buffer buf_n5524( .i (n5523), .o (n5524) );
  buffer buf_n5525( .i (n5524), .o (n5525) );
  assign n5526 = n1405 & ~n5525 ;
  buffer buf_n4229( .i (n4228), .o (n4229) );
  buffer buf_n4230( .i (n4229), .o (n4230) );
  assign n5527 = ( n757 & n4230 ) | ( n757 & n5405 ) | ( n4230 & n5405 ) ;
  assign n5528 = ~n3990 & n5527 ;
  buffer buf_n5529( .i (n5287), .o (n5529) );
  assign n5530 = ( ~n4224 & n5470 ) | ( ~n4224 & n5529 ) | ( n5470 & n5529 ) ;
  buffer buf_n5531( .i (n5530), .o (n5531) );
  buffer buf_n5532( .i (n5531), .o (n5532) );
  buffer buf_n5533( .i (n5532), .o (n5533) );
  assign n5534 = ( ~n5358 & n5496 ) | ( ~n5358 & n5531 ) | ( n5496 & n5531 ) ;
  assign n5535 = ( n5326 & ~n5429 ) | ( n5326 & n5534 ) | ( ~n5429 & n5534 ) ;
  assign n5536 = n5533 & n5535 ;
  assign n5537 = n3531 & ~n5358 ;
  buffer buf_n5538( .i (n5537), .o (n5538) );
  buffer buf_n5539( .i (n5538), .o (n5539) );
  assign n5540 = n5417 & ~n5538 ;
  assign n5541 = ( n5536 & n5539 ) | ( n5536 & ~n5540 ) | ( n5539 & ~n5540 ) ;
  assign n5542 = ( ~n5225 & n5506 ) | ( ~n5225 & n5541 ) | ( n5506 & n5541 ) ;
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n5543( .i (n5470), .o (n5543) );
  buffer buf_n5544( .i (n5543), .o (n5544) );
  assign n5545 = ( ~n4586 & n5428 ) | ( ~n4586 & n5544 ) | ( n5428 & n5544 ) ;
  assign n5546 = ( ~n4586 & n5093 ) | ( ~n4586 & n5544 ) | ( n5093 & n5544 ) ;
  assign n5547 = ( n2263 & n5545 ) | ( n2263 & ~n5546 ) | ( n5545 & ~n5546 ) ;
  buffer buf_n5548( .i (n5464), .o (n5548) );
  assign n5549 = n5547 | n5548 ;
  assign n5550 = n836 & n2042 ;
  assign n5551 = n5548 & ~n5550 ;
  assign n5552 = n5549 & ~n5551 ;
  assign n5553 = ( n5225 & n5506 ) | ( n5225 & ~n5552 ) | ( n5506 & ~n5552 ) ;
  assign n5554 = n5542 & ~n5553 ;
  assign n5555 = n5528 | n5554 ;
  assign n5556 = ( n1406 & ~n5526 ) | ( n1406 & n5555 ) | ( ~n5526 & n5555 ) ;
  assign n5557 = n5514 | n5556 ;
  assign n5558 = ~n181 & n5557 ;
  assign n5559 = n5492 | n5558 ;
  assign n5560 = n5442 | n5559 ;
  assign n5561 = ( n5201 & ~n5213 ) | ( n5201 & n5560 ) | ( ~n5213 & n5560 ) ;
  buffer buf_n5562( .i (n5295), .o (n5562) );
  buffer buf_n5563( .i (n5562), .o (n5563) );
  assign n5564 = ( ~n3717 & n5496 ) | ( ~n3717 & n5563 ) | ( n5496 & n5563 ) ;
  buffer buf_n5565( .i (n5564), .o (n5565) );
  assign n5566 = ( ~n5057 & n5548 ) | ( ~n5057 & n5565 ) | ( n5548 & n5565 ) ;
  assign n5567 = ( n4889 & n5548 ) | ( n4889 & ~n5565 ) | ( n5548 & ~n5565 ) ;
  assign n5568 = n5566 & ~n5567 ;
  buffer buf_n5569( .i (n5568), .o (n5569) );
  buffer buf_n5570( .i (n5569), .o (n5570) );
  buffer buf_n5571( .i (n4049), .o (n5571) );
  buffer buf_n5572( .i (n5571), .o (n5572) );
  buffer buf_n5573( .i (n5572), .o (n5573) );
  assign n5574 = ( ~n5181 & n5569 ) | ( ~n5181 & n5573 ) | ( n5569 & n5573 ) ;
  buffer buf_n4023( .i (n4022), .o (n4023) );
  buffer buf_n4024( .i (n4023), .o (n4024) );
  buffer buf_n4025( .i (n4024), .o (n4025) );
  assign n5575 = n3850 & ~n4025 ;
  assign n5576 = ~n5573 & n5575 ;
  assign n5577 = ( n5570 & ~n5574 ) | ( n5570 & n5576 ) | ( ~n5574 & n5576 ) ;
  buffer buf_n5578( .i (n5577), .o (n5578) );
  buffer buf_n5579( .i (n5578), .o (n5579) );
  buffer buf_n4042( .i (n4041), .o (n4042) );
  buffer buf_n4043( .i (n4042), .o (n4043) );
  buffer buf_n4044( .i (n4043), .o (n4044) );
  buffer buf_n4045( .i (n4044), .o (n4045) );
  buffer buf_n4046( .i (n4045), .o (n4046) );
  buffer buf_n4047( .i (n4046), .o (n4047) );
  assign n5580 = ( n4516 & n4654 ) | ( n4516 & n5294 ) | ( n4654 & n5294 ) ;
  assign n5581 = ( ~n4835 & n5295 ) | ( ~n4835 & n5580 ) | ( n5295 & n5580 ) ;
  buffer buf_n5582( .i (n5581), .o (n5582) );
  assign n5585 = n5563 & ~n5582 ;
  buffer buf_n5586( .i (n5585), .o (n5586) );
  buffer buf_n5587( .i (n5586), .o (n5587) );
  buffer buf_n5583( .i (n5582), .o (n5583) );
  buffer buf_n5584( .i (n5583), .o (n5584) );
  assign n5588 = n5584 | n5586 ;
  buffer buf_n5589( .i (n5057), .o (n5589) );
  assign n5590 = ( n5587 & n5588 ) | ( n5587 & ~n5589 ) | ( n5588 & ~n5589 ) ;
  buffer buf_n5591( .i (n5590), .o (n5591) );
  buffer buf_n5592( .i (n5591), .o (n5592) );
  buffer buf_n3821( .i (n3820), .o (n3821) );
  assign n5593 = ( n3821 & n5181 ) | ( n3821 & ~n5591 ) | ( n5181 & ~n5591 ) ;
  assign n5594 = n5592 & n5593 ;
  buffer buf_n5595( .i (n5594), .o (n5595) );
  assign n5596 = ( n4047 & ~n5578 ) | ( n4047 & n5595 ) | ( ~n5578 & n5595 ) ;
  buffer buf_n5597( .i (n4896), .o (n5597) );
  assign n5598 = ~n5595 & n5597 ;
  assign n5599 = ( n5579 & n5596 ) | ( n5579 & ~n5598 ) | ( n5596 & ~n5598 ) ;
  buffer buf_n5600( .i (n5599), .o (n5600) );
  buffer buf_n5601( .i (n5600), .o (n5601) );
  buffer buf_n5602( .i (n359), .o (n5602) );
  assign n5603 = n5600 & ~n5602 ;
  buffer buf_n5604( .i (n4487), .o (n5604) );
  buffer buf_n5605( .i (n5604), .o (n5605) );
  assign n5606 = ( ~n1572 & n4419 ) | ( ~n1572 & n5605 ) | ( n4419 & n5605 ) ;
  assign n5607 = ( n1571 & ~n3915 ) | ( n1571 & n4654 ) | ( ~n3915 & n4654 ) ;
  buffer buf_n5608( .i (n4820), .o (n5608) );
  assign n5609 = ( n5605 & n5607 ) | ( n5605 & ~n5608 ) | ( n5607 & ~n5608 ) ;
  assign n5610 = n5606 & ~n5609 ;
  assign n5611 = ~n5428 & n5610 ;
  buffer buf_n5612( .i (n5611), .o (n5612) );
  buffer buf_n5613( .i (n5612), .o (n5613) );
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n2211( .i (n2210), .o (n2211) );
  buffer buf_n2212( .i (n2211), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  buffer buf_n5065( .i (n5064), .o (n5065) );
  buffer buf_n5066( .i (n5065), .o (n5066) );
  buffer buf_n5614( .i (n3717), .o (n5614) );
  assign n5615 = ( n2213 & n5066 ) | ( n2213 & ~n5614 ) | ( n5066 & ~n5614 ) ;
  assign n5616 = n5612 | n5615 ;
  assign n5617 = ( n5571 & n5613 ) | ( n5571 & n5616 ) | ( n5613 & n5616 ) ;
  assign n5618 = n5405 & ~n5617 ;
  buffer buf_n3775( .i (n3774), .o (n3775) );
  buffer buf_n3776( .i (n3775), .o (n3776) );
  buffer buf_n3777( .i (n3776), .o (n3777) );
  buffer buf_n3778( .i (n3777), .o (n3778) );
  buffer buf_n3779( .i (n3778), .o (n3779) );
  assign n5619 = n3776 & ~n5427 ;
  buffer buf_n5620( .i (n5619), .o (n5620) );
  buffer buf_n5621( .i (n5620), .o (n5621) );
  assign n5622 = ( n4826 & n5614 ) | ( n4826 & ~n5620 ) | ( n5614 & ~n5620 ) ;
  assign n5623 = ( n3779 & n5621 ) | ( n3779 & ~n5622 ) | ( n5621 & ~n5622 ) ;
  assign n5624 = ~n5571 & n5623 ;
  assign n5625 = n5405 | n5624 ;
  assign n5626 = ~n5618 & n5625 ;
  buffer buf_n5627( .i (n5626), .o (n5627) );
  buffer buf_n5628( .i (n5627), .o (n5628) );
  assign n5629 = n4770 & n5627 ;
  buffer buf_n1007( .i (n1006), .o (n1007) );
  assign n5630 = ( n929 & n1007 ) | ( n929 & n2738 ) | ( n1007 & n2738 ) ;
  buffer buf_n5631( .i (n929), .o (n5631) );
  assign n5632 = ( ~n4720 & n5630 ) | ( ~n4720 & n5631 ) | ( n5630 & n5631 ) ;
  buffer buf_n5633( .i (n5632), .o (n5633) );
  buffer buf_n5634( .i (n5633), .o (n5634) );
  assign n5635 = ( ~n734 & n3990 ) | ( ~n734 & n5633 ) | ( n3990 & n5633 ) ;
  assign n5636 = n5634 & ~n5635 ;
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n2846( .i (n2845), .o (n2846) );
  buffer buf_n2847( .i (n2846), .o (n2847) );
  buffer buf_n2848( .i (n2847), .o (n2848) );
  assign n5637 = ( n2848 & n3013 ) | ( n2848 & n5543 ) | ( n3013 & n5543 ) ;
  assign n5638 = ~n3014 & n5637 ;
  buffer buf_n5639( .i (n5638), .o (n5639) );
  buffer buf_n5640( .i (n5639), .o (n5640) );
  buffer buf_n5641( .i (n5640), .o (n5641) );
  buffer buf_n2520( .i (n2519), .o (n2520) );
  buffer buf_n2521( .i (n2520), .o (n2521) );
  buffer buf_n2522( .i (n2521), .o (n2522) );
  buffer buf_n5642( .i (n5464), .o (n5642) );
  assign n5643 = ( n2522 & n5639 ) | ( n2522 & ~n5642 ) | ( n5639 & ~n5642 ) ;
  assign n5644 = n543 & ~n5643 ;
  assign n5645 = ( n544 & n5641 ) | ( n544 & ~n5644 ) | ( n5641 & ~n5644 ) ;
  assign n5646 = n5573 | n5645 ;
  buffer buf_n4504( .i (n4503), .o (n4504) );
  buffer buf_n4505( .i (n4504), .o (n4505) );
  buffer buf_n4506( .i (n4505), .o (n4506) );
  buffer buf_n4507( .i (n4506), .o (n4507) );
  buffer buf_n4508( .i (n4507), .o (n4508) );
  buffer buf_n4509( .i (n4508), .o (n4509) );
  buffer buf_n4510( .i (n4509), .o (n4510) );
  buffer buf_n4511( .i (n4510), .o (n4511) );
  assign n5647 = n314 | n4511 ;
  assign n5648 = n5573 & n5647 ;
  assign n5649 = n5646 & ~n5648 ;
  assign n5650 = n5636 | n5649 ;
  assign n5651 = ( n5628 & ~n5629 ) | ( n5628 & n5650 ) | ( ~n5629 & n5650 ) ;
  assign n5652 = n3489 | n5651 ;
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n5653( .i (n5614), .o (n5653) );
  assign n5654 = ( n962 & ~n5419 ) | ( n962 & n5653 ) | ( ~n5419 & n5653 ) ;
  buffer buf_n5655( .i (n5074), .o (n5655) );
  assign n5656 = ( ~n962 & n5419 ) | ( ~n962 & n5655 ) | ( n5419 & n5655 ) ;
  assign n5657 = ( ~n460 & n5654 ) | ( ~n460 & n5656 ) | ( n5654 & n5656 ) ;
  buffer buf_n5658( .i (n5404), .o (n5658) );
  assign n5659 = ~n5657 & n5658 ;
  buffer buf_n613( .i (n612), .o (n613) );
  assign n5660 = n613 & n5459 ;
  assign n5661 = n5658 | n5660 ;
  assign n5662 = ~n5659 & n5661 ;
  buffer buf_n5663( .i (n5505), .o (n5663) );
  buffer buf_n5664( .i (n5663), .o (n5664) );
  assign n5665 = n5662 & n5664 ;
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  assign n5666 = ( n1384 & n4838 ) | ( n1384 & ~n5064 ) | ( n4838 & ~n5064 ) ;
  buffer buf_n5667( .i (n5666), .o (n5667) );
  buffer buf_n5668( .i (n5667), .o (n5668) );
  buffer buf_n5669( .i (n5668), .o (n5669) );
  assign n5670 = ( n5429 & ~n5614 ) | ( n5429 & n5667 ) | ( ~n5614 & n5667 ) ;
  assign n5671 = ( n1387 & ~n5096 ) | ( n1387 & n5670 ) | ( ~n5096 & n5670 ) ;
  assign n5672 = ( ~n1388 & n5669 ) | ( ~n1388 & n5671 ) | ( n5669 & n5671 ) ;
  assign n5673 = ~n5658 & n5672 ;
  buffer buf_n5674( .i (n5096), .o (n5674) );
  assign n5675 = n1215 & ~n5674 ;
  assign n5676 = n5658 & ~n5675 ;
  assign n5677 = n5673 | n5676 ;
  assign n5678 = ~n5664 & n5677 ;
  assign n5679 = ( n4770 & ~n5665 ) | ( n4770 & n5678 ) | ( ~n5665 & n5678 ) ;
  assign n5680 = n4944 | n5679 ;
  buffer buf_n5681( .i (n120), .o (n5681) );
  assign n5682 = n5680 & n5681 ;
  assign n5683 = n5652 & ~n5682 ;
  assign n5684 = ( n3135 & n5493 ) | ( n3135 & ~n5495 ) | ( n5493 & ~n5495 ) ;
  buffer buf_n5685( .i (n5684), .o (n5685) );
  buffer buf_n5686( .i (n5494), .o (n5686) );
  assign n5687 = n5685 | n5686 ;
  assign n5688 = n5685 & n5686 ;
  assign n5689 = n5687 & ~n5688 ;
  buffer buf_n5690( .i (n5689), .o (n5690) );
  buffer buf_n5691( .i (n5690), .o (n5691) );
  buffer buf_n5692( .i (n4873), .o (n5692) );
  assign n5693 = ( n5572 & n5690 ) | ( n5572 & ~n5692 ) | ( n5690 & ~n5692 ) ;
  buffer buf_n3534( .i (n3533), .o (n3534) );
  assign n5694 = ~n313 & n3534 ;
  assign n5695 = ~n5572 & n5694 ;
  assign n5696 = ( n5691 & ~n5693 ) | ( n5691 & n5695 ) | ( ~n5693 & n5695 ) ;
  buffer buf_n5697( .i (n5696), .o (n5697) );
  buffer buf_n5698( .i (n5697), .o (n5698) );
  assign n5699 = ( n1404 & n2775 ) | ( n1404 & n5179 ) | ( n2775 & n5179 ) ;
  assign n5700 = ~n5150 & n5699 ;
  buffer buf_n2837( .i (n2836), .o (n2837) );
  buffer buf_n2838( .i (n2837), .o (n2838) );
  assign n5701 = n918 & ~n2838 ;
  assign n5702 = ( n3517 & n5043 ) | ( n3517 & n5115 ) | ( n5043 & n5115 ) ;
  buffer buf_n5703( .i (n5702), .o (n5703) );
  buffer buf_n5704( .i (n5703), .o (n5704) );
  buffer buf_n5705( .i (n5704), .o (n5705) );
  assign n5706 = ( n4958 & n5287 ) | ( n4958 & ~n5703 ) | ( n5287 & ~n5703 ) ;
  assign n5707 = n3520 | n5706 ;
  assign n5708 = ( n4838 & ~n5705 ) | ( n4838 & n5707 ) | ( ~n5705 & n5707 ) ;
  assign n5709 = n5563 & ~n5708 ;
  assign n5710 = ~n5686 & n5709 ;
  buffer buf_n4163( .i (n4162), .o (n4163) );
  buffer buf_n4164( .i (n4163), .o (n4164) );
  buffer buf_n5711( .i (n5238), .o (n5711) );
  buffer buf_n5712( .i (n5711), .o (n5712) );
  assign n5713 = ( n4164 & n4818 ) | ( n4164 & ~n5712 ) | ( n4818 & ~n5712 ) ;
  buffer buf_n5714( .i (n5713), .o (n5714) );
  buffer buf_n5717( .i (n4819), .o (n5717) );
  assign n5718 = ~n5714 & n5717 ;
  buffer buf_n5719( .i (n5718), .o (n5719) );
  buffer buf_n5720( .i (n5719), .o (n5720) );
  buffer buf_n5715( .i (n5714), .o (n5715) );
  buffer buf_n5716( .i (n5715), .o (n5716) );
  assign n5721 = n5716 | n5719 ;
  assign n5722 = ( ~n5494 & n5720 ) | ( ~n5494 & n5721 ) | ( n5720 & n5721 ) ;
  assign n5723 = n5517 & ~n5608 ;
  buffer buf_n5724( .i (n5723), .o (n5724) );
  buffer buf_n5725( .i (n5724), .o (n5725) );
  assign n5726 = n5563 | n5724 ;
  assign n5727 = ( n5722 & n5725 ) | ( n5722 & n5726 ) | ( n5725 & n5726 ) ;
  assign n5728 = n5710 | n5727 ;
  assign n5729 = ( n919 & ~n5701 ) | ( n919 & n5728 ) | ( ~n5701 & n5728 ) ;
  assign n5730 = ( n5505 & ~n5572 ) | ( n5505 & n5729 ) | ( ~n5572 & n5729 ) ;
  assign n5731 = ( n4572 & ~n5346 ) | ( n4572 & n5712 ) | ( ~n5346 & n5712 ) ;
  buffer buf_n5732( .i (n5731), .o (n5732) );
  buffer buf_n5733( .i (n5732), .o (n5733) );
  buffer buf_n5734( .i (n5733), .o (n5734) );
  buffer buf_n5735( .i (n5286), .o (n5735) );
  assign n5736 = n5732 & n5735 ;
  buffer buf_n5737( .i (n4516), .o (n5737) );
  assign n5738 = ( n4835 & n5736 ) | ( n4835 & ~n5737 ) | ( n5736 & ~n5737 ) ;
  assign n5739 = ( n1431 & n5734 ) | ( n1431 & ~n5738 ) | ( n5734 & ~n5738 ) ;
  assign n5740 = n3717 | n5739 ;
  assign n5741 = n565 & ~n2095 ;
  buffer buf_n5742( .i (n5116), .o (n5742) );
  buffer buf_n5743( .i (n5742), .o (n5743) );
  buffer buf_n5744( .i (n5743), .o (n5744) );
  buffer buf_n5745( .i (n5744), .o (n5745) );
  assign n5746 = ~n5741 & n5745 ;
  assign n5747 = n5740 & ~n5746 ;
  buffer buf_n5748( .i (n5686), .o (n5748) );
  assign n5749 = n5747 | n5748 ;
  buffer buf_n2058( .i (n2057), .o (n2058) );
  assign n5750 = n399 & n2058 ;
  assign n5751 = n5748 & ~n5750 ;
  assign n5752 = n5749 & ~n5751 ;
  buffer buf_n5753( .i (n5571), .o (n5753) );
  assign n5754 = ( n5505 & ~n5752 ) | ( n5505 & n5753 ) | ( ~n5752 & n5753 ) ;
  assign n5755 = n5730 & ~n5754 ;
  buffer buf_n5756( .i (n5755), .o (n5756) );
  assign n5757 = ( ~n5697 & n5700 ) | ( ~n5697 & n5756 ) | ( n5700 & n5756 ) ;
  assign n5758 = n4255 & ~n5756 ;
  assign n5759 = ( n5698 & n5757 ) | ( n5698 & ~n5758 ) | ( n5757 & ~n5758 ) ;
  assign n5760 = n267 & ~n5759 ;
  buffer buf_n2803( .i (n2802), .o (n2803) );
  buffer buf_n2804( .i (n2803), .o (n2804) );
  buffer buf_n2805( .i (n2804), .o (n2805) );
  buffer buf_n2806( .i (n2805), .o (n2806) );
  buffer buf_n2807( .i (n2806), .o (n2807) );
  buffer buf_n5761( .i (n5496), .o (n5761) );
  assign n5762 = n2807 | n5761 ;
  buffer buf_n2812( .i (n2811), .o (n2812) );
  assign n5763 = n2812 & n5761 ;
  assign n5764 = n5762 & ~n5763 ;
  assign n5765 = n5404 & ~n5764 ;
  assign n5766 = n1007 & n4889 ;
  assign n5767 = n5404 | n5766 ;
  assign n5768 = ~n5765 & n5767 ;
  buffer buf_n5769( .i (n5745), .o (n5769) );
  assign n5770 = n917 & ~n5769 ;
  assign n5771 = n2124 & n5770 ;
  buffer buf_n5772( .i (n5771), .o (n5772) );
  buffer buf_n5773( .i (n5772), .o (n5773) );
  buffer buf_n5774( .i (n5589), .o (n5774) );
  assign n5775 = ~n5772 & n5774 ;
  assign n5776 = ( n5768 & n5773 ) | ( n5768 & ~n5775 ) | ( n5773 & ~n5775 ) ;
  assign n5777 = ( n5135 & ~n5379 ) | ( n5135 & n5392 ) | ( ~n5379 & n5392 ) ;
  assign n5778 = ( n5346 & ~n5712 ) | ( n5346 & n5777 ) | ( ~n5712 & n5777 ) ;
  buffer buf_n5779( .i (n5778), .o (n5779) );
  buffer buf_n5782( .i (n5007), .o (n5782) );
  assign n5783 = ~n5779 & n5782 ;
  buffer buf_n5784( .i (n5783), .o (n5784) );
  buffer buf_n5785( .i (n5784), .o (n5785) );
  buffer buf_n5780( .i (n5779), .o (n5780) );
  buffer buf_n5781( .i (n5780), .o (n5781) );
  assign n5786 = n5781 | n5784 ;
  buffer buf_n5787( .i (n5495), .o (n5787) );
  assign n5788 = ( n5785 & n5786 ) | ( n5785 & ~n5787 ) | ( n5786 & ~n5787 ) ;
  buffer buf_n5789( .i (n5494), .o (n5789) );
  assign n5790 = ( n5326 & n5788 ) | ( n5326 & n5789 ) | ( n5788 & n5789 ) ;
  buffer buf_n5791( .i (n5790), .o (n5791) );
  assign n5792 = ( n5184 & ~n5589 ) | ( n5184 & n5791 ) | ( ~n5589 & n5791 ) ;
  buffer buf_n5793( .i (n5359), .o (n5793) );
  buffer buf_n5794( .i (n5793), .o (n5794) );
  assign n5795 = ( n5674 & ~n5791 ) | ( n5674 & n5794 ) | ( ~n5791 & n5794 ) ;
  assign n5796 = n5792 & ~n5795 ;
  buffer buf_n5797( .i (n5796), .o (n5797) );
  assign n5798 = ( ~n5664 & n5776 ) | ( ~n5664 & n5797 ) | ( n5776 & n5797 ) ;
  assign n5799 = ~n4637 & n5392 ;
  buffer buf_n5800( .i (n5799), .o (n5800) );
  buffer buf_n5801( .i (n5800), .o (n5801) );
  buffer buf_n5802( .i (n5801), .o (n5802) );
  buffer buf_n5803( .i (n5802), .o (n5803) );
  assign n5807 = ( n5427 & ~n5462 ) | ( n5427 & n5803 ) | ( ~n5462 & n5803 ) ;
  assign n5808 = ( n5295 & ~n5529 ) | ( n5295 & n5802 ) | ( ~n5529 & n5802 ) ;
  assign n5809 = ( n5462 & ~n5495 ) | ( n5462 & n5808 ) | ( ~n5495 & n5808 ) ;
  assign n5810 = n5807 | n5809 ;
  buffer buf_n5811( .i (n5810), .o (n5811) );
  buffer buf_n5812( .i (n5811), .o (n5812) );
  assign n5813 = n5748 | n5811 ;
  buffer buf_n1693( .i (n1692), .o (n1693) );
  assign n5814 = n1693 & n2042 ;
  assign n5815 = ( ~n4637 & n4962 ) | ( ~n4637 & n5392 ) | ( n4962 & n5392 ) ;
  buffer buf_n5816( .i (n5815), .o (n5816) );
  buffer buf_n5824( .i (n4818), .o (n5824) );
  assign n5825 = ( ~n5286 & n5816 ) | ( ~n5286 & n5824 ) | ( n5816 & n5824 ) ;
  buffer buf_n5826( .i (n5825), .o (n5826) );
  assign n5829 = n5608 & ~n5826 ;
  buffer buf_n5830( .i (n5829), .o (n5830) );
  buffer buf_n5831( .i (n5830), .o (n5831) );
  buffer buf_n5827( .i (n5826), .o (n5827) );
  buffer buf_n5828( .i (n5827), .o (n5828) );
  assign n5832 = n5828 | n5830 ;
  assign n5833 = ( ~n5789 & n5831 ) | ( ~n5789 & n5832 ) | ( n5831 & n5832 ) ;
  assign n5834 = n5814 | n5833 ;
  assign n5835 = ( ~n5812 & n5813 ) | ( ~n5812 & n5834 ) | ( n5813 & n5834 ) ;
  assign n5836 = n5435 & ~n5835 ;
  assign n5837 = ( n527 & n5427 ) | ( n527 & ~n5446 ) | ( n5427 & ~n5446 ) ;
  buffer buf_n5838( .i (n5837), .o (n5838) );
  buffer buf_n5839( .i (n5838), .o (n5839) );
  assign n5840 = ( n5448 & ~n5789 ) | ( n5448 & n5838 ) | ( ~n5789 & n5838 ) ;
  assign n5841 = ( ~n5419 & n5839 ) | ( ~n5419 & n5840 ) | ( n5839 & n5840 ) ;
  assign n5842 = n5589 | n5841 ;
  assign n5843 = ~n5435 & n5842 ;
  assign n5844 = n5836 | n5843 ;
  assign n5845 = ( n5664 & n5797 ) | ( n5664 & ~n5844 ) | ( n5797 & ~n5844 ) ;
  assign n5846 = n5798 | n5845 ;
  buffer buf_n5847( .i (n5485), .o (n5847) );
  assign n5848 = n5846 & ~n5847 ;
  assign n5849 = n267 | n5848 ;
  assign n5850 = ~n5760 & n5849 ;
  assign n5851 = n5683 | n5850 ;
  assign n5852 = ( n5601 & ~n5603 ) | ( n5601 & n5851 ) | ( ~n5603 & n5851 ) ;
  assign n5853 = n3916 & n5737 ;
  buffer buf_n5854( .i (n5853), .o (n5854) );
  buffer buf_n5855( .i (n5854), .o (n5855) );
  assign n5856 = ( ~n5464 & n5769 ) | ( ~n5464 & n5855 ) | ( n5769 & n5855 ) ;
  assign n5857 = ( n5745 & n5787 ) | ( n5745 & ~n5854 ) | ( n5787 & ~n5854 ) ;
  buffer buf_n5858( .i (n5463), .o (n5858) );
  assign n5859 = ( n4864 & n5857 ) | ( n4864 & ~n5858 ) | ( n5857 & ~n5858 ) ;
  assign n5860 = ~n5856 & n5859 ;
  buffer buf_n5861( .i (n5860), .o (n5861) );
  buffer buf_n5862( .i (n5861), .o (n5862) );
  buffer buf_n5863( .i (n5794), .o (n5863) );
  buffer buf_n5864( .i (n5674), .o (n5864) );
  assign n5865 = ( n5861 & n5863 ) | ( n5861 & n5864 ) | ( n5863 & n5864 ) ;
  buffer buf_n2463( .i (n2462), .o (n2463) );
  buffer buf_n2464( .i (n2463), .o (n2464) );
  buffer buf_n2465( .i (n2464), .o (n2465) );
  buffer buf_n2466( .i (n2465), .o (n2466) );
  assign n5866 = ( n731 & n2466 ) | ( n731 & n5642 ) | ( n2466 & n5642 ) ;
  buffer buf_n5867( .i (n5642), .o (n5867) );
  assign n5868 = n5866 & ~n5867 ;
  assign n5869 = ~n5864 & n5868 ;
  assign n5870 = ( n5862 & ~n5865 ) | ( n5862 & n5869 ) | ( ~n5865 & n5869 ) ;
  buffer buf_n5871( .i (n5870), .o (n5871) );
  buffer buf_n5872( .i (n5871), .o (n5872) );
  buffer buf_n5873( .i (n5872), .o (n5873) );
  assign n5874 = ( ~n119 & n601 ) | ( ~n119 & n5871 ) | ( n601 & n5871 ) ;
  assign n5875 = n761 & ~n5874 ;
  assign n5876 = ( n762 & n5873 ) | ( n762 & ~n5875 ) | ( n5873 & ~n5875 ) ;
  buffer buf_n5877( .i (n5876), .o (n5877) );
  buffer buf_n5878( .i (n5877), .o (n5878) );
  assign n5879 = n2712 & n5877 ;
  buffer buf_n523( .i (n522), .o (n523) );
  assign n5880 = ( ~n2145 & n2298 ) | ( ~n2145 & n5256 ) | ( n2298 & n5256 ) ;
  buffer buf_n5881( .i (n4974), .o (n5881) );
  assign n5882 = ( n5298 & n5880 ) | ( n5298 & ~n5881 ) | ( n5880 & ~n5881 ) ;
  buffer buf_n5883( .i (n5882), .o (n5883) );
  buffer buf_n5884( .i (n5883), .o (n5884) );
  assign n5885 = ~n5391 & n5883 ;
  assign n5886 = ( n5711 & n5884 ) | ( n5711 & n5885 ) | ( n5884 & n5885 ) ;
  buffer buf_n5887( .i (n5886), .o (n5887) );
  buffer buf_n5888( .i (n5887), .o (n5888) );
  assign n5889 = n4017 & ~n5887 ;
  assign n5890 = ( n1303 & n5888 ) | ( n1303 & ~n5889 ) | ( n5888 & ~n5889 ) ;
  buffer buf_n5891( .i (n5294), .o (n5891) );
  assign n5892 = ~n5890 & n5891 ;
  assign n5893 = ~n5396 & n5742 ;
  assign n5894 = n5891 | n5893 ;
  assign n5895 = ~n5892 & n5894 ;
  buffer buf_n5896( .i (n5493), .o (n5896) );
  assign n5897 = n5895 & ~n5896 ;
  buffer buf_n5898( .i (n2230), .o (n5898) );
  buffer buf_n5899( .i (n5898), .o (n5899) );
  assign n5900 = ( ~n2329 & n2330 ) | ( ~n2329 & n5899 ) | ( n2330 & n5899 ) ;
  buffer buf_n5901( .i (n5900), .o (n5901) );
  buffer buf_n5902( .i (n5901), .o (n5902) );
  buffer buf_n5903( .i (n5902), .o (n5903) );
  buffer buf_n5904( .i (n5903), .o (n5904) );
  assign n5906 = ( n5347 & n5712 ) | ( n5347 & ~n5904 ) | ( n5712 & ~n5904 ) ;
  buffer buf_n5907( .i (n5711), .o (n5907) );
  assign n5908 = ( ~n5115 & n5904 ) | ( ~n5115 & n5907 ) | ( n5904 & n5907 ) ;
  assign n5909 = n5906 & ~n5908 ;
  assign n5910 = ( ~n5118 & n5782 ) | ( ~n5118 & n5909 ) | ( n5782 & n5909 ) ;
  buffer buf_n5911( .i (n5379), .o (n5911) );
  assign n5912 = n344 & n5911 ;
  assign n5913 = ~n5515 & n5912 ;
  buffer buf_n5914( .i (n4815), .o (n5914) );
  assign n5915 = ( n5782 & n5913 ) | ( n5782 & n5914 ) | ( n5913 & n5914 ) ;
  assign n5916 = n5910 & n5915 ;
  assign n5917 = n3029 & ~n5914 ;
  assign n5918 = n442 & n5917 ;
  assign n5919 = n5916 | n5918 ;
  assign n5920 = n5896 & n5919 ;
  assign n5921 = n5897 | n5920 ;
  buffer buf_n5922( .i (n5921), .o (n5922) );
  buffer buf_n5923( .i (n5922), .o (n5923) );
  buffer buf_n5924( .i (n3733), .o (n5924) );
  assign n5925 = ( n2913 & ~n4560 ) | ( n2913 & n5924 ) | ( ~n4560 & n5924 ) ;
  buffer buf_n5926( .i (n5925), .o (n5926) );
  buffer buf_n5929( .i (n4962), .o (n5929) );
  assign n5930 = ~n5926 & n5929 ;
  buffer buf_n5931( .i (n5930), .o (n5931) );
  buffer buf_n5932( .i (n5931), .o (n5932) );
  buffer buf_n5927( .i (n5926), .o (n5927) );
  buffer buf_n5928( .i (n5927), .o (n5928) );
  assign n5933 = n5928 | n5931 ;
  assign n5934 = ( ~n5608 & n5932 ) | ( ~n5608 & n5933 ) | ( n5932 & n5933 ) ;
  buffer buf_n5935( .i (n5934), .o (n5935) );
  buffer buf_n5936( .i (n5935), .o (n5936) );
  assign n5937 = ( n349 & n5544 ) | ( n349 & n5935 ) | ( n5544 & n5935 ) ;
  assign n5938 = n744 & ~n5737 ;
  assign n5939 = n2242 & n5938 ;
  assign n5940 = ~n349 & n5939 ;
  assign n5941 = ( n5936 & ~n5937 ) | ( n5936 & n5940 ) | ( ~n5937 & n5940 ) ;
  assign n5942 = n536 & ~n5116 ;
  assign n5943 = ~n330 & n4572 ;
  buffer buf_n5944( .i (n5943), .o (n5944) );
  assign n5955 = n5942 & n5944 ;
  buffer buf_n5956( .i (n5955), .o (n5956) );
  buffer buf_n5957( .i (n5956), .o (n5957) );
  buffer buf_n5958( .i (n5957), .o (n5958) );
  assign n5959 = ( ~n5493 & n5543 ) | ( ~n5493 & n5956 ) | ( n5543 & n5956 ) ;
  assign n5960 = n3032 & ~n5959 ;
  assign n5961 = ( n3033 & n5958 ) | ( n3033 & ~n5960 ) | ( n5958 & ~n5960 ) ;
  buffer buf_n5962( .i (n4864), .o (n5962) );
  assign n5963 = ( n5941 & n5961 ) | ( n5941 & ~n5962 ) | ( n5961 & ~n5962 ) ;
  assign n5964 = ~n5922 & n5963 ;
  assign n5965 = ( ~n5753 & n5923 ) | ( ~n5753 & n5964 ) | ( n5923 & n5964 ) ;
  buffer buf_n5966( .i (n5965), .o (n5966) );
  buffer buf_n5967( .i (n5966), .o (n5967) );
  buffer buf_n5968( .i (n5967), .o (n5968) );
  assign n5969 = ( n718 & n933 ) | ( n718 & n5966 ) | ( n933 & n5966 ) ;
  assign n5970 = n522 & ~n5969 ;
  assign n5971 = ( n523 & n5968 ) | ( n523 & ~n5970 ) | ( n5968 & ~n5970 ) ;
  buffer buf_n2102( .i (n2101), .o (n2102) );
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n5972( .i (n5899), .o (n5972) );
  assign n5973 = ( n969 & ~n5881 ) | ( n969 & n5972 ) | ( ~n5881 & n5972 ) ;
  buffer buf_n5974( .i (n5973), .o (n5974) );
  assign n5977 = n5238 & n5974 ;
  buffer buf_n5978( .i (n5977), .o (n5978) );
  buffer buf_n5979( .i (n5978), .o (n5979) );
  buffer buf_n5975( .i (n5974), .o (n5975) );
  buffer buf_n5976( .i (n5975), .o (n5976) );
  assign n5980 = n5976 & ~n5978 ;
  assign n5981 = ( n5286 & ~n5979 ) | ( n5286 & n5980 ) | ( ~n5979 & n5980 ) ;
  assign n5982 = n4958 & ~n5981 ;
  buffer buf_n5983( .i (n5717), .o (n5983) );
  assign n5984 = n5982 & n5983 ;
  buffer buf_n5985( .i (n5984), .o (n5985) );
  buffer buf_n5986( .i (n5985), .o (n5986) );
  assign n5987 = n2836 | n5985 ;
  assign n5988 = ( ~n2358 & n5986 ) | ( ~n2358 & n5987 ) | ( n5986 & n5987 ) ;
  assign n5989 = ( n5793 & ~n5962 ) | ( n5793 & n5988 ) | ( ~n5962 & n5988 ) ;
  assign n5990 = ( ~n3923 & n5379 ) | ( ~n3923 & n5711 ) | ( n5379 & n5711 ) ;
  buffer buf_n5991( .i (n5990), .o (n5991) );
  buffer buf_n5992( .i (n5991), .o (n5992) );
  buffer buf_n5993( .i (n5992), .o (n5993) );
  buffer buf_n5994( .i (n5993), .o (n5994) );
  assign n5995 = ( n5008 & ~n5515 ) | ( n5008 & n5991 ) | ( ~n5515 & n5991 ) ;
  buffer buf_n5996( .i (n5995), .o (n5996) );
  buffer buf_n5997( .i (n5996), .o (n5997) );
  assign n5998 = n3927 | n5996 ;
  assign n5999 = ( ~n5994 & n5997 ) | ( ~n5994 & n5998 ) | ( n5997 & n5998 ) ;
  assign n6000 = n5787 | n5999 ;
  assign n6001 = n5789 | n6000 ;
  assign n6002 = ( n5793 & n5962 ) | ( n5793 & n6001 ) | ( n5962 & n6001 ) ;
  assign n6003 = n5989 & ~n6002 ;
  buffer buf_n6004( .i (n6003), .o (n6004) );
  buffer buf_n6005( .i (n6004), .o (n6005) );
  buffer buf_n6006( .i (n6005), .o (n6006) );
  assign n6007 = ( n378 & n5153 ) | ( n378 & n6004 ) | ( n5153 & n6004 ) ;
  assign n6008 = n2102 | n6007 ;
  assign n6009 = ( ~n2103 & n6006 ) | ( ~n2103 & n6008 ) | ( n6006 & n6008 ) ;
  buffer buf_n6010( .i (n6009), .o (n6010) );
  assign n6011 = ( n151 & n5971 ) | ( n151 & n6010 ) | ( n5971 & n6010 ) ;
  buffer buf_n6012( .i (n5515), .o (n6012) );
  assign n6013 = ( n5242 & ~n5604 ) | ( n5242 & n6012 ) | ( ~n5604 & n6012 ) ;
  buffer buf_n6014( .i (n6013), .o (n6014) );
  buffer buf_n6015( .i (n6014), .o (n6015) );
  buffer buf_n6016( .i (n6015), .o (n6016) );
  buffer buf_n5245( .i (n5244), .o (n5245) );
  buffer buf_n6017( .i (n5529), .o (n6017) );
  assign n6018 = ( n5320 & n6014 ) | ( n5320 & ~n6017 ) | ( n6014 & ~n6017 ) ;
  assign n6019 = ~n5245 & n6018 ;
  assign n6020 = ( ~n5326 & n6016 ) | ( ~n5326 & n6019 ) | ( n6016 & n6019 ) ;
  assign n6021 = n5793 | n6020 ;
  assign n6022 = n1239 & ~n5761 ;
  buffer buf_n6023( .i (n5544), .o (n6023) );
  buffer buf_n6024( .i (n6023), .o (n6024) );
  assign n6025 = ~n6022 & n6024 ;
  assign n6026 = n6021 & ~n6025 ;
  assign n6027 = ( n842 & n5529 ) | ( n842 & n5605 ) | ( n5529 & n5605 ) ;
  buffer buf_n6028( .i (n6027), .o (n6028) );
  buffer buf_n6029( .i (n5562), .o (n6029) );
  buffer buf_n6030( .i (n6017), .o (n6030) );
  assign n6031 = ( n6028 & n6029 ) | ( n6028 & ~n6030 ) | ( n6029 & ~n6030 ) ;
  buffer buf_n6032( .i (n5605), .o (n6032) );
  buffer buf_n6033( .i (n6032), .o (n6033) );
  assign n6034 = ( ~n6028 & n6029 ) | ( ~n6028 & n6033 ) | ( n6029 & n6033 ) ;
  assign n6035 = n6031 & ~n6034 ;
  buffer buf_n6036( .i (n6035), .o (n6036) );
  buffer buf_n6037( .i (n6036), .o (n6037) );
  buffer buf_n6038( .i (n5962), .o (n6038) );
  assign n6039 = ~n6036 & n6038 ;
  assign n6040 = ( n6026 & n6037 ) | ( n6026 & ~n6039 ) | ( n6037 & ~n6039 ) ;
  assign n6041 = n5112 | n6040 ;
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  assign n6042 = ~n638 & n2181 ;
  buffer buf_n6043( .i (n5347), .o (n6043) );
  assign n6044 = n5007 | n6043 ;
  buffer buf_n6045( .i (n6044), .o (n6045) );
  buffer buf_n6046( .i (n6045), .o (n6046) );
  buffer buf_n6047( .i (n6046), .o (n6047) );
  buffer buf_n6048( .i (n5737), .o (n6048) );
  assign n6049 = ( n4341 & ~n5543 ) | ( n4341 & n6048 ) | ( ~n5543 & n6048 ) ;
  buffer buf_n6050( .i (n5470), .o (n6050) );
  assign n6051 = ( ~n4341 & n6032 ) | ( ~n4341 & n6050 ) | ( n6032 & n6050 ) ;
  assign n6052 = ( ~n6047 & n6049 ) | ( ~n6047 & n6051 ) | ( n6049 & n6051 ) ;
  assign n6053 = ~n5429 & n6052 ;
  buffer buf_n6054( .i (n4637), .o (n6054) );
  buffer buf_n6055( .i (n6054), .o (n6055) );
  assign n6056 = ( n2092 & n2258 ) | ( n2092 & ~n6055 ) | ( n2258 & ~n6055 ) ;
  buffer buf_n6057( .i (n6056), .o (n6057) );
  buffer buf_n6068( .i (n5782), .o (n6068) );
  buffer buf_n6069( .i (n5604), .o (n6069) );
  assign n6070 = ( ~n6057 & n6068 ) | ( ~n6057 & n6069 ) | ( n6068 & n6069 ) ;
  buffer buf_n6071( .i (n6070), .o (n6071) );
  buffer buf_n6072( .i (n6050), .o (n6072) );
  assign n6073 = ( ~n5787 & n6071 ) | ( ~n5787 & n6072 ) | ( n6071 & n6072 ) ;
  assign n6074 = ( n6033 & ~n6071 ) | ( n6033 & n6072 ) | ( ~n6071 & n6072 ) ;
  assign n6075 = n6073 & ~n6074 ;
  assign n6076 = n6053 | n6075 ;
  assign n6077 = ( n2182 & ~n6042 ) | ( n2182 & n6076 ) | ( ~n6042 & n6076 ) ;
  assign n6078 = ~n5753 & n6077 ;
  assign n6079 = n5112 & ~n6078 ;
  assign n6080 = n6041 & ~n6079 ;
  assign n6081 = n179 | n6080 ;
  assign n6082 = ( n2038 & n4878 ) | ( n2038 & n5604 ) | ( n4878 & n5604 ) ;
  buffer buf_n6083( .i (n6082), .o (n6083) );
  buffer buf_n6084( .i (n6083), .o (n6084) );
  buffer buf_n6085( .i (n6084), .o (n6085) );
  assign n6086 = ( n6032 & n6048 ) | ( n6032 & ~n6083 ) | ( n6048 & ~n6083 ) ;
  assign n6087 = ( ~n2041 & n6030 ) | ( ~n2041 & n6086 ) | ( n6030 & n6086 ) ;
  assign n6088 = ( n2042 & ~n6085 ) | ( n2042 & n6087 ) | ( ~n6085 & n6087 ) ;
  assign n6089 = n6024 & ~n6088 ;
  assign n6090 = n946 & n6030 ;
  assign n6091 = n945 | n5562 ;
  assign n6092 = ( n6030 & n6033 ) | ( n6030 & n6091 ) | ( n6033 & n6091 ) ;
  assign n6093 = ~n6090 & n6092 ;
  assign n6094 = n6024 | n6093 ;
  assign n6095 = ( ~n5794 & n6089 ) | ( ~n5794 & n6094 ) | ( n6089 & n6094 ) ;
  assign n6096 = n5864 & ~n6095 ;
  buffer buf_n6097( .i (n6029), .o (n6097) );
  assign n6098 = ~n350 & n6097 ;
  assign n6099 = ( ~n351 & n4889 ) | ( ~n351 & n6098 ) | ( n4889 & n6098 ) ;
  assign n6100 = ~n5794 & n6099 ;
  assign n6101 = n5864 | n6100 ;
  assign n6102 = ~n6096 & n6101 ;
  assign n6103 = ~n4912 & n6102 ;
  assign n6104 = n179 & ~n6103 ;
  assign n6105 = n6081 & ~n6104 ;
  assign n6106 = ( ~n151 & n6010 ) | ( ~n151 & n6105 ) | ( n6010 & n6105 ) ;
  assign n6107 = n6011 | n6106 ;
  assign n6108 = n5824 & n6055 ;
  buffer buf_n6109( .i (n6108), .o (n6109) );
  buffer buf_n6113( .i (n5136), .o (n6113) );
  buffer buf_n6114( .i (n6113), .o (n6114) );
  buffer buf_n6115( .i (n6114), .o (n6115) );
  assign n6116 = ( n6069 & n6109 ) | ( n6069 & n6115 ) | ( n6109 & n6115 ) ;
  buffer buf_n6117( .i (n6116), .o (n6117) );
  assign n6118 = n5463 | n6117 ;
  buffer buf_n6119( .i (n5462), .o (n6119) );
  assign n6120 = n6117 & n6119 ;
  assign n6121 = n6118 & ~n6120 ;
  assign n6122 = n5653 | n6121 ;
  assign n6123 = n1829 & n6032 ;
  assign n6124 = ( n2497 & n6033 ) | ( n2497 & ~n6123 ) | ( n6033 & ~n6123 ) ;
  buffer buf_n6125( .i (n5896), .o (n6125) );
  assign n6126 = n6124 | n6125 ;
  assign n6127 = n5653 & n6126 ;
  assign n6128 = n6122 & ~n6127 ;
  assign n6129 = n5863 & ~n6128 ;
  assign n6130 = ( ~n2244 & n5858 ) | ( ~n2244 & n6125 ) | ( n5858 & n6125 ) ;
  assign n6131 = ( n2243 & n5896 ) | ( n2243 & ~n6029 ) | ( n5896 & ~n6029 ) ;
  assign n6132 = ( ~n5769 & n5858 ) | ( ~n5769 & n6131 ) | ( n5858 & n6131 ) ;
  assign n6133 = n6130 & ~n6132 ;
  assign n6134 = ~n4720 & n6133 ;
  assign n6135 = n5863 | n6134 ;
  assign n6136 = ~n6129 & n6135 ;
  assign n6137 = n5150 & n6136 ;
  assign n6138 = ( n5136 & n5347 ) | ( n5136 & n5911 ) | ( n5347 & n5911 ) ;
  assign n6139 = ( n6043 & ~n6055 ) | ( n6043 & n6138 ) | ( ~n6055 & n6138 ) ;
  buffer buf_n6140( .i (n6139), .o (n6140) );
  assign n6143 = n6069 & ~n6140 ;
  buffer buf_n6144( .i (n6143), .o (n6144) );
  buffer buf_n6145( .i (n6144), .o (n6145) );
  buffer buf_n6141( .i (n6140), .o (n6141) );
  buffer buf_n6142( .i (n6141), .o (n6142) );
  assign n6146 = n6142 | n6144 ;
  buffer buf_n6147( .i (n6069), .o (n6147) );
  buffer buf_n6148( .i (n6147), .o (n6148) );
  buffer buf_n6149( .i (n6148), .o (n6149) );
  assign n6150 = ( n6145 & n6146 ) | ( n6145 & ~n6149 ) | ( n6146 & ~n6149 ) ;
  assign n6151 = n6024 & ~n6150 ;
  assign n6152 = n2521 & ~n5858 ;
  buffer buf_n6153( .i (n6023), .o (n6153) );
  assign n6154 = n6152 | n6153 ;
  assign n6155 = ~n6151 & n6154 ;
  buffer buf_n6156( .i (n5562), .o (n6156) );
  assign n6157 = n2520 & ~n6156 ;
  assign n6158 = n2009 & n6072 ;
  assign n6159 = n6157 & n6158 ;
  buffer buf_n6160( .i (n6159), .o (n6160) );
  buffer buf_n6161( .i (n6160), .o (n6161) );
  assign n6162 = n5674 & ~n6160 ;
  assign n6163 = ( n6155 & n6161 ) | ( n6155 & ~n6162 ) | ( n6161 & ~n6162 ) ;
  buffer buf_n6164( .i (n5983), .o (n6164) );
  buffer buf_n6165( .i (n6115), .o (n6165) );
  assign n6166 = ( ~n6147 & n6164 ) | ( ~n6147 & n6165 ) | ( n6164 & n6165 ) ;
  buffer buf_n6167( .i (n6166), .o (n6167) );
  buffer buf_n6168( .i (n6119), .o (n6168) );
  assign n6169 = ( n6097 & n6167 ) | ( n6097 & ~n6168 ) | ( n6167 & ~n6168 ) ;
  assign n6170 = ( n6097 & n6125 ) | ( n6097 & ~n6167 ) | ( n6125 & ~n6167 ) ;
  assign n6171 = n6169 & ~n6170 ;
  buffer buf_n6172( .i (n6153), .o (n6172) );
  assign n6173 = n6171 | n6172 ;
  buffer buf_n4108( .i (n4107), .o (n4108) );
  buffer buf_n4109( .i (n4108), .o (n4109) );
  buffer buf_n4110( .i (n4109), .o (n4110) );
  buffer buf_n4111( .i (n4110), .o (n4111) );
  assign n6174 = n4111 & n5748 ;
  assign n6175 = n6172 & ~n6174 ;
  assign n6176 = n6173 & ~n6175 ;
  assign n6177 = n6163 | n6176 ;
  buffer buf_n6178( .i (n5179), .o (n6178) );
  assign n6179 = n6177 & ~n6178 ;
  assign n6180 = n6137 | n6179 ;
  buffer buf_n6181( .i (n6180), .o (n6181) );
  buffer buf_n6182( .i (n6181), .o (n6182) );
  assign n6183 = n3025 & n6181 ;
  buffer buf_n6184( .i (n4721), .o (n6184) );
  assign n6185 = ( n1266 & n5482 ) | ( n1266 & n6184 ) | ( n5482 & n6184 ) ;
  buffer buf_n6186( .i (n6185), .o (n6186) );
  assign n6187 = ( n179 & ~n207 ) | ( n179 & n6186 ) | ( ~n207 & n6186 ) ;
  buffer buf_n6188( .i (n5284), .o (n6188) );
  buffer buf_n6189( .i (n6188), .o (n6189) );
  buffer buf_n6190( .i (n6184), .o (n6190) );
  buffer buf_n6191( .i (n6190), .o (n6191) );
  assign n6192 = ( ~n6186 & n6189 ) | ( ~n6186 & n6191 ) | ( n6189 & n6191 ) ;
  assign n6193 = n6187 & ~n6192 ;
  buffer buf_n2251( .i (n2250), .o (n2251) );
  assign n6194 = ( n5745 & ~n6072 ) | ( n5745 & n6119 ) | ( ~n6072 & n6119 ) ;
  buffer buf_n6195( .i (n6050), .o (n6195) );
  buffer buf_n6196( .i (n5744), .o (n6196) );
  assign n6197 = ( n6156 & ~n6195 ) | ( n6156 & n6196 ) | ( ~n6195 & n6196 ) ;
  assign n6198 = n6194 & ~n6197 ;
  buffer buf_n6199( .i (n5761), .o (n6199) );
  assign n6200 = n6198 & n6199 ;
  buffer buf_n6201( .i (n6125), .o (n6201) );
  buffer buf_n6202( .i (n6201), .o (n6202) );
  assign n6203 = ( n6038 & n6200 ) | ( n6038 & n6202 ) | ( n6200 & n6202 ) ;
  assign n6204 = ~n5753 & n6203 ;
  buffer buf_n6205( .i (n6204), .o (n6205) );
  buffer buf_n6206( .i (n6205), .o (n6206) );
  buffer buf_n6207( .i (n6206), .o (n6207) );
  assign n6208 = ( ~n695 & n1405 ) | ( ~n695 & n6205 ) | ( n1405 & n6205 ) ;
  assign n6209 = n2250 & ~n6208 ;
  assign n6210 = ( n2251 & n6207 ) | ( n2251 & ~n6209 ) | ( n6207 & ~n6209 ) ;
  assign n6211 = n6193 | n6210 ;
  assign n6212 = ( n6182 & ~n6183 ) | ( n6182 & n6211 ) | ( ~n6183 & n6211 ) ;
  assign n6213 = n6107 | n6212 ;
  assign n6214 = ( n5878 & ~n5879 ) | ( n5878 & n6213 ) | ( ~n5879 & n6213 ) ;
  buffer buf_n735( .i (n734), .o (n735) );
  assign n6215 = ( n5642 & n5653 ) | ( n5642 & n6199 ) | ( n5653 & n6199 ) ;
  buffer buf_n6216( .i (n6215), .o (n6216) );
  buffer buf_n6217( .i (n6216), .o (n6217) );
  assign n6218 = ~n5435 & n6216 ;
  assign n6219 = ( ~n3990 & n6217 ) | ( ~n3990 & n6218 ) | ( n6217 & n6218 ) ;
  assign n6220 = n735 & n6219 ;
  buffer buf_n6221( .i (n6220), .o (n6221) );
  buffer buf_n6222( .i (n6221), .o (n6222) );
  buffer buf_n6223( .i (n5972), .o (n6223) );
  assign n6224 = ( n5163 & n5299 ) | ( n5163 & ~n6223 ) | ( n5299 & ~n6223 ) ;
  buffer buf_n6225( .i (n6224), .o (n6225) );
  buffer buf_n6226( .i (n6225), .o (n6226) );
  buffer buf_n6227( .i (n6226), .o (n6227) );
  buffer buf_n6228( .i (n6227), .o (n6228) );
  buffer buf_n6229( .i (n6228), .o (n6229) );
  buffer buf_n6230( .i (n6229), .o (n6230) );
  buffer buf_n6231( .i (n6230), .o (n6231) );
  buffer buf_n6232( .i (n6231), .o (n6232) );
  buffer buf_n6233( .i (n6232), .o (n6233) );
  buffer buf_n6234( .i (n6233), .o (n6234) );
  assign n6238 = ( n6038 & ~n6172 ) | ( n6038 & n6234 ) | ( ~n6172 & n6234 ) ;
  buffer buf_n6239( .i (n6238), .o (n6239) );
  buffer buf_n6240( .i (n6239), .o (n6240) );
  buffer buf_n6241( .i (n6240), .o (n6241) );
  buffer buf_n6235( .i (n6234), .o (n6235) );
  buffer buf_n6236( .i (n6235), .o (n6236) );
  buffer buf_n6237( .i (n6236), .o (n6237) );
  buffer buf_n6242( .i (n5178), .o (n6242) );
  assign n6243 = ( n5663 & n6239 ) | ( n5663 & ~n6242 ) | ( n6239 & ~n6242 ) ;
  assign n6244 = ~n6237 & n6243 ;
  buffer buf_n6245( .i (n6038), .o (n6245) );
  buffer buf_n6246( .i (n6245), .o (n6246) );
  buffer buf_n6247( .i (n6246), .o (n6247) );
  buffer buf_n6248( .i (n6247), .o (n6248) );
  assign n6249 = ( n6241 & n6244 ) | ( n6241 & ~n6248 ) | ( n6244 & ~n6248 ) ;
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n3166( .i (n3165), .o (n3166) );
  buffer buf_n3167( .i (n3166), .o (n3167) );
  buffer buf_n3168( .i (n3167), .o (n3168) );
  buffer buf_n3169( .i (n3168), .o (n3169) );
  buffer buf_n3170( .i (n3169), .o (n3170) );
  assign n6250 = n3170 & ~n6246 ;
  assign n6251 = n546 & n6250 ;
  buffer buf_n6252( .i (n6251), .o (n6252) );
  assign n6253 = ( ~n6221 & n6249 ) | ( ~n6221 & n6252 ) | ( n6249 & n6252 ) ;
  assign n6254 = n5597 & ~n6252 ;
  assign n6255 = ( n6222 & n6253 ) | ( n6222 & ~n6254 ) | ( n6253 & ~n6254 ) ;
  buffer buf_n6256( .i (n6255), .o (n6256) );
  buffer buf_n6257( .i (n6256), .o (n6257) );
  buffer buf_n4594( .i (n4593), .o (n4594) );
  buffer buf_n4595( .i (n4594), .o (n4595) );
  buffer buf_n4596( .i (n4595), .o (n4596) );
  buffer buf_n4597( .i (n4596), .o (n4597) );
  buffer buf_n4598( .i (n4597), .o (n4598) );
  buffer buf_n4599( .i (n4598), .o (n4599) );
  buffer buf_n4600( .i (n4599), .o (n4600) );
  buffer buf_n4601( .i (n4600), .o (n4601) );
  buffer buf_n4602( .i (n4601), .o (n4602) );
  buffer buf_n4603( .i (n4602), .o (n4603) );
  buffer buf_n4604( .i (n4603), .o (n4604) );
  buffer buf_n4605( .i (n4604), .o (n4605) );
  assign n6258 = n4605 & n6256 ;
  buffer buf_n6259( .i (n5907), .o (n6259) );
  assign n6260 = n742 & ~n6259 ;
  assign n6261 = ( n6012 & n6114 ) | ( n6012 & n6260 ) | ( n6114 & n6260 ) ;
  assign n6262 = ~n6115 & n6261 ;
  buffer buf_n6263( .i (n6262), .o (n6263) );
  buffer buf_n6264( .i (n6263), .o (n6264) );
  buffer buf_n6265( .i (n6264), .o (n6265) );
  assign n6266 = ( ~n310 & n2041 ) | ( ~n310 & n6263 ) | ( n2041 & n6263 ) ;
  assign n6267 = n6168 & ~n6266 ;
  buffer buf_n6268( .i (n6168), .o (n6268) );
  assign n6269 = ( n6265 & ~n6267 ) | ( n6265 & n6268 ) | ( ~n6267 & n6268 ) ;
  assign n6270 = n4773 & ~n6269 ;
  buffer buf_n3136( .i (n3135), .o (n3136) );
  buffer buf_n6271( .i (n6017), .o (n6271) );
  assign n6272 = ( n3136 & n6119 ) | ( n3136 & ~n6271 ) | ( n6119 & ~n6271 ) ;
  buffer buf_n6273( .i (n6164), .o (n6273) );
  assign n6274 = ( n3136 & ~n6271 ) | ( n3136 & n6273 ) | ( ~n6271 & n6273 ) ;
  assign n6275 = ( n2010 & n6272 ) | ( n2010 & ~n6274 ) | ( n6272 & ~n6274 ) ;
  buffer buf_n6276( .i (n6097), .o (n6276) );
  assign n6277 = n6275 & n6276 ;
  buffer buf_n6278( .i (n6199), .o (n6278) );
  assign n6279 = n6277 | n6278 ;
  assign n6280 = ~n6270 & n6279 ;
  buffer buf_n6281( .i (n6280), .o (n6281) );
  buffer buf_n6282( .i (n6281), .o (n6282) );
  assign n6283 = n6190 & n6281 ;
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  assign n6284 = ~n591 & n613 ;
  assign n6285 = ( ~n1725 & n5863 ) | ( ~n1725 & n6284 ) | ( n5863 & n6284 ) ;
  assign n6286 = ~n5663 & n6285 ;
  buffer buf_n5371( .i (n5370), .o (n5371) );
  buffer buf_n5372( .i (n5371), .o (n5372) );
  assign n6287 = ( n440 & n6055 ) | ( n440 & n6259 ) | ( n6055 & n6259 ) ;
  assign n6288 = n5372 & ~n6287 ;
  buffer buf_n6289( .i (n5914), .o (n6289) );
  assign n6290 = n6288 & n6289 ;
  buffer buf_n6291( .i (n6054), .o (n6291) );
  assign n6292 = ( ~n5116 & n5800 ) | ( ~n5116 & n6291 ) | ( n5800 & n6291 ) ;
  buffer buf_n6293( .i (n5911), .o (n6293) );
  assign n6294 = ( n5800 & n6259 ) | ( n5800 & ~n6293 ) | ( n6259 & ~n6293 ) ;
  assign n6295 = ( n2038 & n6292 ) | ( n2038 & ~n6294 ) | ( n6292 & ~n6294 ) ;
  assign n6296 = n6289 | n6295 ;
  assign n6297 = ( ~n6050 & n6290 ) | ( ~n6050 & n6296 ) | ( n6290 & n6296 ) ;
  assign n6298 = n6148 & ~n6297 ;
  buffer buf_n6299( .i (n5391), .o (n6299) );
  buffer buf_n6300( .i (n6299), .o (n6300) );
  assign n6301 = ( n2117 & n5215 ) | ( n2117 & ~n6300 ) | ( n5215 & ~n6300 ) ;
  buffer buf_n6302( .i (n6301), .o (n6302) );
  buffer buf_n6303( .i (n6302), .o (n6303) );
  assign n6304 = ( n5217 & n6012 ) | ( n5217 & ~n6302 ) | ( n6012 & ~n6302 ) ;
  assign n6305 = ( n6068 & n6303 ) | ( n6068 & ~n6304 ) | ( n6303 & ~n6304 ) ;
  assign n6306 = n5744 & n6305 ;
  assign n6307 = n6148 | n6306 ;
  assign n6308 = ~n6298 & n6307 ;
  assign n6309 = n6201 & n6308 ;
  assign n6310 = ( n2174 & n5167 ) | ( n2174 & n6300 ) | ( n5167 & n6300 ) ;
  buffer buf_n6311( .i (n6300), .o (n6311) );
  assign n6312 = n6310 & ~n6311 ;
  buffer buf_n6313( .i (n6312), .o (n6313) );
  buffer buf_n6314( .i (n6313), .o (n6314) );
  buffer buf_n6315( .i (n6314), .o (n6315) );
  assign n6316 = ( n3063 & n5164 ) | ( n3063 & n5238 ) | ( n5164 & n5238 ) ;
  buffer buf_n6317( .i (n6316), .o (n6317) );
  buffer buf_n6318( .i (n6317), .o (n6318) );
  buffer buf_n6319( .i (n6318), .o (n6319) );
  assign n6320 = ( n5907 & n6054 ) | ( n5907 & ~n6317 ) | ( n6054 & ~n6317 ) ;
  assign n6321 = n6293 & n6320 ;
  assign n6322 = ( n5914 & ~n6319 ) | ( n5914 & n6321 ) | ( ~n6319 & n6321 ) ;
  assign n6323 = ( n6068 & n6313 ) | ( n6068 & n6322 ) | ( n6313 & n6322 ) ;
  assign n6324 = n6147 & ~n6323 ;
  assign n6325 = ( n6148 & n6315 ) | ( n6148 & ~n6324 ) | ( n6315 & ~n6324 ) ;
  buffer buf_n6326( .i (n5163), .o (n6326) );
  buffer buf_n6327( .i (n4307), .o (n6327) );
  assign n6328 = ( ~n5391 & n6326 ) | ( ~n5391 & n6327 ) | ( n6326 & n6327 ) ;
  buffer buf_n6329( .i (n4949), .o (n6329) );
  buffer buf_n6330( .i (n6329), .o (n6330) );
  assign n6331 = ( n5389 & n6328 ) | ( n5389 & ~n6330 ) | ( n6328 & ~n6330 ) ;
  buffer buf_n6332( .i (n6331), .o (n6332) );
  buffer buf_n6335( .i (n4324), .o (n6335) );
  assign n6336 = ~n6332 & n6335 ;
  buffer buf_n6337( .i (n6336), .o (n6337) );
  buffer buf_n6338( .i (n6337), .o (n6338) );
  buffer buf_n6333( .i (n6332), .o (n6333) );
  buffer buf_n6334( .i (n6333), .o (n6334) );
  assign n6339 = n6334 | n6337 ;
  buffer buf_n6340( .i (n6289), .o (n6340) );
  assign n6341 = ( n6338 & n6339 ) | ( n6338 & ~n6340 ) | ( n6339 & ~n6340 ) ;
  assign n6342 = ( n6156 & n6196 ) | ( n6156 & n6341 ) | ( n6196 & n6341 ) ;
  assign n6343 = ( ~n2244 & n6325 ) | ( ~n2244 & n6342 ) | ( n6325 & n6342 ) ;
  assign n6344 = n6201 | n6343 ;
  assign n6345 = ( ~n6202 & n6309 ) | ( ~n6202 & n6344 ) | ( n6309 & n6344 ) ;
  buffer buf_n6346( .i (n5867), .o (n6346) );
  assign n6347 = n6345 & n6346 ;
  buffer buf_n6348( .i (n5924), .o (n6348) );
  buffer buf_n6349( .i (n5165), .o (n6349) );
  assign n6350 = ( n6225 & n6348 ) | ( n6225 & ~n6349 ) | ( n6348 & ~n6349 ) ;
  buffer buf_n6351( .i (n6350), .o (n6351) );
  assign n6354 = n6293 & n6351 ;
  buffer buf_n6355( .i (n6354), .o (n6355) );
  buffer buf_n6356( .i (n6355), .o (n6356) );
  buffer buf_n6352( .i (n6351), .o (n6352) );
  buffer buf_n6353( .i (n6352), .o (n6353) );
  assign n6357 = n6353 & ~n6355 ;
  assign n6358 = ( n5744 & ~n6356 ) | ( n5744 & n6357 ) | ( ~n6356 & n6357 ) ;
  buffer buf_n6359( .i (n6358), .o (n6359) );
  buffer buf_n6360( .i (n6359), .o (n6360) );
  assign n6361 = n2180 & ~n6359 ;
  assign n6362 = ( n2138 & ~n6360 ) | ( n2138 & n6361 ) | ( ~n6360 & n6361 ) ;
  buffer buf_n6363( .i (n47), .o (n6363) );
  buffer buf_n6364( .i (n4306), .o (n6364) );
  assign n6365 = ( ~n5901 & n6363 ) | ( ~n5901 & n6364 ) | ( n6363 & n6364 ) ;
  buffer buf_n6366( .i (n6365), .o (n6366) );
  buffer buf_n6367( .i (n6366), .o (n6367) );
  buffer buf_n6368( .i (n6367), .o (n6368) );
  buffer buf_n6369( .i (n6368), .o (n6369) );
  buffer buf_n6370( .i (n4560), .o (n6370) );
  assign n6371 = ( ~n6349 & n6366 ) | ( ~n6349 & n6370 ) | ( n6366 & n6370 ) ;
  buffer buf_n6372( .i (n6371), .o (n6372) );
  buffer buf_n6373( .i (n6372), .o (n6373) );
  buffer buf_n5905( .i (n5904), .o (n5905) );
  assign n6374 = n5905 & n6372 ;
  assign n6375 = ( ~n6369 & n6373 ) | ( ~n6369 & n6374 ) | ( n6373 & n6374 ) ;
  assign n6376 = n2173 & ~n5389 ;
  assign n6377 = ~n5911 & n6376 ;
  buffer buf_n6378( .i (n6377), .o (n6378) );
  buffer buf_n6379( .i (n6378), .o (n6379) );
  assign n6380 = n5735 & ~n6378 ;
  assign n6381 = ( n6375 & n6379 ) | ( n6375 & ~n6380 ) | ( n6379 & ~n6380 ) ;
  assign n6382 = n6048 & ~n6381 ;
  assign n6383 = n2060 & n6289 ;
  assign n6384 = n6048 | n6383 ;
  assign n6385 = ~n6382 & n6384 ;
  buffer buf_n6386( .i (n6273), .o (n6386) );
  assign n6387 = n6385 & ~n6386 ;
  buffer buf_n6388( .i (n6043), .o (n6388) );
  buffer buf_n6389( .i (n6388), .o (n6389) );
  assign n6390 = ( n634 & ~n2834 ) | ( n634 & n6389 ) | ( ~n2834 & n6389 ) ;
  assign n6391 = ( n1103 & n5907 ) | ( n1103 & ~n6054 ) | ( n5907 & ~n6054 ) ;
  buffer buf_n6392( .i (n6370), .o (n6392) );
  assign n6393 = ( n1103 & ~n6300 ) | ( n1103 & n6392 ) | ( ~n6300 & n6392 ) ;
  assign n6394 = n6391 | n6393 ;
  buffer buf_n6395( .i (n6335), .o (n6395) );
  assign n6396 = ~n6394 & n6395 ;
  assign n6397 = n6389 & n6396 ;
  assign n6398 = ( n2835 & n6390 ) | ( n2835 & n6397 ) | ( n6390 & n6397 ) ;
  buffer buf_n6399( .i (n6395), .o (n6399) );
  assign n6400 = n2177 & n6399 ;
  assign n6401 = n443 & n6400 ;
  assign n6402 = n6398 | n6401 ;
  assign n6403 = n6386 & n6402 ;
  assign n6404 = n6387 | n6403 ;
  assign n6405 = n6362 | n6404 ;
  assign n6406 = ~n6346 & n6405 ;
  assign n6407 = n6347 | n6406 ;
  assign n6408 = n6286 | n6407 ;
  assign n6409 = ( n6282 & ~n6283 ) | ( n6282 & n6408 ) | ( ~n6283 & n6408 ) ;
  buffer buf_n6410( .i (n6409), .o (n6410) );
  buffer buf_n6411( .i (n6410), .o (n6411) );
  assign n6412 = n3025 & n6410 ;
  assign n6413 = n4729 & ~n5444 ;
  assign n6414 = n3814 & n6413 ;
  buffer buf_n6415( .i (n6414), .o (n6415) );
  buffer buf_n6416( .i (n6415), .o (n6416) );
  buffer buf_n6417( .i (n6416), .o (n6417) );
  buffer buf_n3903( .i (n3902), .o (n3903) );
  buffer buf_n3904( .i (n3903), .o (n3904) );
  buffer buf_n3905( .i (n3904), .o (n3905) );
  buffer buf_n3906( .i (n3905), .o (n3906) );
  assign n6418 = n586 & n6115 ;
  assign n6419 = ( n3906 & n3997 ) | ( n3906 & ~n6418 ) | ( n3997 & ~n6418 ) ;
  buffer buf_n6420( .i (n6147), .o (n6420) );
  assign n6421 = ( n6415 & n6419 ) | ( n6415 & ~n6420 ) | ( n6419 & ~n6420 ) ;
  buffer buf_n6422( .i (n6271), .o (n6422) );
  assign n6423 = ~n6421 & n6422 ;
  buffer buf_n6424( .i (n6422), .o (n6424) );
  assign n6425 = ( n6417 & ~n6423 ) | ( n6417 & n6424 ) | ( ~n6423 & n6424 ) ;
  buffer buf_n6426( .i (n5769), .o (n6426) );
  buffer buf_n6427( .i (n6426), .o (n6427) );
  assign n6428 = n6425 & n6427 ;
  buffer buf_n6429( .i (n6428), .o (n6429) );
  buffer buf_n6430( .i (n6429), .o (n6430) );
  buffer buf_n2467( .i (n2466), .o (n2467) );
  assign n6431 = ( n2467 & n5631 ) | ( n2467 & n5867 ) | ( n5631 & n5867 ) ;
  assign n6432 = ~n6346 & n6431 ;
  assign n6433 = n6429 | n6432 ;
  assign n6434 = ( ~n6247 & n6430 ) | ( ~n6247 & n6433 ) | ( n6430 & n6433 ) ;
  buffer buf_n6435( .i (n5663), .o (n6435) );
  buffer buf_n6436( .i (n6435), .o (n6436) );
  assign n6437 = n6434 | n6436 ;
  assign n6438 = ( n1368 & n6199 ) | ( n1368 & n6268 ) | ( n6199 & n6268 ) ;
  assign n6439 = ( n1368 & ~n6201 ) | ( n1368 & n6268 ) | ( ~n6201 & n6268 ) ;
  buffer buf_n6440( .i (n590), .o (n6440) );
  assign n6441 = ( ~n6438 & n6439 ) | ( ~n6438 & n6440 ) | ( n6439 & n6440 ) ;
  buffer buf_n2936( .i (n2935), .o (n2936) );
  buffer buf_n6442( .i (n6389), .o (n6442) );
  assign n6443 = n372 & ~n6442 ;
  buffer buf_n6444( .i (n6443), .o (n6444) );
  assign n6448 = n2936 & n6444 ;
  buffer buf_n6449( .i (n6448), .o (n6449) );
  buffer buf_n6450( .i (n6449), .o (n6450) );
  assign n6451 = n6427 & ~n6449 ;
  assign n6452 = ( n6441 & ~n6450 ) | ( n6441 & n6451 ) | ( ~n6450 & n6451 ) ;
  assign n6453 = n407 & n1308 ;
  buffer buf_n6454( .i (n6453), .o (n6454) );
  buffer buf_n6455( .i (n6454), .o (n6455) );
  assign n6456 = n5692 | n6454 ;
  assign n6457 = ( ~n6452 & n6455 ) | ( ~n6452 & n6456 ) | ( n6455 & n6456 ) ;
  assign n6458 = ~n6247 & n6457 ;
  assign n6459 = n6436 & ~n6458 ;
  assign n6460 = n6437 & ~n6459 ;
  assign n6461 = n3041 | n6460 ;
  assign n6462 = ( n6411 & ~n6412 ) | ( n6411 & n6461 ) | ( ~n6412 & n6461 ) ;
  buffer buf_n6445( .i (n6444), .o (n6445) );
  buffer buf_n6446( .i (n6445), .o (n6446) );
  buffer buf_n6447( .i (n6446), .o (n6447) );
  assign n6463 = ( ~n5178 & n6245 ) | ( ~n5178 & n6447 ) | ( n6245 & n6447 ) ;
  buffer buf_n2373( .i (n2372), .o (n2373) );
  buffer buf_n6464( .i (n6114), .o (n6464) );
  assign n6465 = ( n2373 & ~n6389 ) | ( n2373 & n6464 ) | ( ~n6389 & n6464 ) ;
  buffer buf_n6466( .i (n6465), .o (n6466) );
  buffer buf_n6469( .i (n6165), .o (n6469) );
  assign n6470 = ~n6466 & n6469 ;
  buffer buf_n6471( .i (n6470), .o (n6471) );
  buffer buf_n6472( .i (n6471), .o (n6472) );
  buffer buf_n6467( .i (n6466), .o (n6467) );
  buffer buf_n6468( .i (n6467), .o (n6468) );
  assign n6473 = n6468 | n6471 ;
  assign n6474 = ( ~n5867 & n6472 ) | ( ~n5867 & n6473 ) | ( n6472 & n6473 ) ;
  buffer buf_n6475( .i (n6278), .o (n6475) );
  assign n6476 = ( n6245 & ~n6474 ) | ( n6245 & n6475 ) | ( ~n6474 & n6475 ) ;
  assign n6477 = n6463 & ~n6476 ;
  buffer buf_n6478( .i (n6477), .o (n6478) );
  buffer buf_n6479( .i (n6478), .o (n6479) );
  buffer buf_n6480( .i (n6427), .o (n6480) );
  assign n6481 = n2615 & n6480 ;
  assign n6482 = ( n1065 & n6246 ) | ( n1065 & n6481 ) | ( n6246 & n6481 ) ;
  assign n6483 = ~n6247 & n6482 ;
  buffer buf_n6484( .i (n6196), .o (n6484) );
  assign n6485 = n4508 & ~n6484 ;
  assign n6486 = ( n4509 & ~n5203 ) | ( n4509 & n6485 ) | ( ~n5203 & n6485 ) ;
  buffer buf_n6487( .i (n6486), .o (n6487) );
  buffer buf_n6488( .i (n6487), .o (n6488) );
  buffer buf_n6489( .i (n6172), .o (n6489) );
  assign n6490 = ( n4002 & n6487 ) | ( n4002 & n6489 ) | ( n6487 & n6489 ) ;
  assign n6491 = ~n6488 & n6490 ;
  buffer buf_n6492( .i (n6491), .o (n6492) );
  assign n6493 = ( ~n6478 & n6483 ) | ( ~n6478 & n6492 ) | ( n6483 & n6492 ) ;
  assign n6494 = n6436 & ~n6492 ;
  assign n6495 = ( n6479 & n6493 ) | ( n6479 & ~n6494 ) | ( n6493 & ~n6494 ) ;
  assign n6496 = n93 | n6495 ;
  buffer buf_n3280( .i (n3279), .o (n3280) );
  buffer buf_n3281( .i (n3280), .o (n3281) );
  buffer buf_n3282( .i (n3281), .o (n3282) );
  buffer buf_n3283( .i (n3282), .o (n3283) );
  buffer buf_n3284( .i (n3283), .o (n3284) );
  buffer buf_n3285( .i (n3284), .o (n3285) );
  buffer buf_n3286( .i (n3285), .o (n3286) );
  buffer buf_n3287( .i (n3286), .o (n3287) );
  buffer buf_n3288( .i (n3287), .o (n3288) );
  buffer buf_n6497( .i (n6388), .o (n6497) );
  assign n6498 = ( n5743 & n6068 ) | ( n5743 & ~n6497 ) | ( n6068 & ~n6497 ) ;
  buffer buf_n6499( .i (n6498), .o (n6499) );
  buffer buf_n6504( .i (n6311), .o (n6504) );
  buffer buf_n6505( .i (n6504), .o (n6505) );
  buffer buf_n6506( .i (n6505), .o (n6506) );
  buffer buf_n6507( .i (n6506), .o (n6507) );
  assign n6508 = ( n6156 & n6499 ) | ( n6156 & ~n6507 ) | ( n6499 & ~n6507 ) ;
  buffer buf_n6509( .i (n5891), .o (n6509) );
  buffer buf_n6510( .i (n6509), .o (n6510) );
  assign n6511 = ( n6196 & ~n6499 ) | ( n6196 & n6510 ) | ( ~n6499 & n6510 ) ;
  assign n6512 = n6508 & ~n6511 ;
  assign n6513 = ( n6153 & ~n6268 ) | ( n6153 & n6512 ) | ( ~n6268 & n6512 ) ;
  assign n6514 = ( n5743 & n6497 ) | ( n5743 & n6505 ) | ( n6497 & n6505 ) ;
  buffer buf_n6515( .i (n6514), .o (n6515) );
  assign n6516 = ( n6507 & n6510 ) | ( n6507 & ~n6515 ) | ( n6510 & ~n6515 ) ;
  buffer buf_n6517( .i (n5743), .o (n6517) );
  buffer buf_n6518( .i (n6517), .o (n6518) );
  assign n6519 = ( n6510 & n6515 ) | ( n6510 & ~n6518 ) | ( n6515 & ~n6518 ) ;
  assign n6520 = ~n6516 & n6519 ;
  buffer buf_n6521( .i (n6168), .o (n6521) );
  assign n6522 = ( n6153 & ~n6520 ) | ( n6153 & n6521 ) | ( ~n6520 & n6521 ) ;
  assign n6523 = n6513 & ~n6522 ;
  buffer buf_n6524( .i (n6523), .o (n6524) );
  buffer buf_n6525( .i (n6524), .o (n6525) );
  buffer buf_n6526( .i (n6525), .o (n6526) );
  buffer buf_n6527( .i (n6489), .o (n6527) );
  assign n6528 = ( n5487 & n6524 ) | ( n5487 & ~n6527 ) | ( n6524 & ~n6527 ) ;
  assign n6529 = n3287 | n6528 ;
  assign n6530 = ( ~n3288 & n6526 ) | ( ~n3288 & n6529 ) | ( n6526 & n6529 ) ;
  assign n6531 = ~n5847 & n6530 ;
  assign n6532 = n93 & ~n6531 ;
  assign n6533 = n6496 & ~n6532 ;
  assign n6534 = n6462 | n6533 ;
  assign n6535 = ( n6257 & ~n6258 ) | ( n6257 & n6534 ) | ( ~n6258 & n6534 ) ;
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  assign n6536 = ( n4673 & ~n6043 ) | ( n4673 & n6293 ) | ( ~n6043 & n6293 ) ;
  buffer buf_n6537( .i (n6536), .o (n6537) );
  buffer buf_n6538( .i (n6537), .o (n6538) );
  buffer buf_n6539( .i (n6538), .o (n6539) );
  buffer buf_n6540( .i (n6539), .o (n6540) );
  assign n6541 = ( n6399 & n6464 ) | ( n6399 & n6537 ) | ( n6464 & n6537 ) ;
  buffer buf_n6542( .i (n6541), .o (n6542) );
  buffer buf_n6543( .i (n6542), .o (n6543) );
  assign n6544 = ~n4677 & n6542 ;
  assign n6545 = ( ~n6540 & n6543 ) | ( ~n6540 & n6544 ) | ( n6543 & n6544 ) ;
  buffer buf_n6546( .i (n6507), .o (n6546) );
  buffer buf_n6547( .i (n6546), .o (n6547) );
  assign n6548 = ~n6545 & n6547 ;
  buffer buf_n4494( .i (n4493), .o (n4494) );
  buffer buf_n4495( .i (n4494), .o (n4495) );
  buffer buf_n4496( .i (n4495), .o (n4496) );
  buffer buf_n4497( .i (n4496), .o (n4497) );
  buffer buf_n4498( .i (n4497), .o (n4498) );
  assign n6549 = n4498 & ~n6023 ;
  assign n6550 = n6547 | n6549 ;
  assign n6551 = ~n6548 & n6550 ;
  buffer buf_n6552( .i (n6202), .o (n6552) );
  assign n6553 = ( ~n6245 & n6551 ) | ( ~n6245 & n6552 ) | ( n6551 & n6552 ) ;
  assign n6554 = ~n4712 & n6505 ;
  buffer buf_n6555( .i (n6554), .o (n6555) );
  assign n6556 = ~n6518 & n6555 ;
  assign n6557 = ( ~n4714 & n6420 ) | ( ~n4714 & n6555 ) | ( n6420 & n6555 ) ;
  assign n6558 = ( n6023 & n6556 ) | ( n6023 & n6557 ) | ( n6556 & n6557 ) ;
  assign n6559 = n6521 | n6558 ;
  assign n6560 = n4118 | n6497 ;
  buffer buf_n6561( .i (n6560), .o (n6561) );
  buffer buf_n6562( .i (n6561), .o (n6562) );
  buffer buf_n6563( .i (n6195), .o (n6563) );
  assign n6564 = ~n6562 & n6563 ;
  assign n6565 = n6521 & ~n6564 ;
  assign n6566 = n6559 & ~n6565 ;
  buffer buf_n6567( .i (n4863), .o (n6567) );
  buffer buf_n6568( .i (n6567), .o (n6568) );
  buffer buf_n6569( .i (n6568), .o (n6569) );
  buffer buf_n6570( .i (n6569), .o (n6570) );
  assign n6571 = ( n6552 & ~n6566 ) | ( n6552 & n6570 ) | ( ~n6566 & n6570 ) ;
  assign n6572 = n6553 & ~n6571 ;
  assign n6573 = ( ~n1403 & n1789 ) | ( ~n1403 & n6480 ) | ( n1789 & n6480 ) ;
  buffer buf_n6574( .i (n1403), .o (n6574) );
  assign n6575 = n6573 & n6574 ;
  assign n6576 = n6572 | n6575 ;
  buffer buf_n6577( .i (n6576), .o (n6577) );
  buffer buf_n6578( .i (n6577), .o (n6578) );
  assign n6579 = ( ~n208 & n238 ) | ( ~n208 & n6577 ) | ( n238 & n6577 ) ;
  assign n6580 = ( n2050 & n6578 ) | ( n2050 & ~n6579 ) | ( n6578 & ~n6579 ) ;
  buffer buf_n6581( .i (n6580), .o (n6581) );
  buffer buf_n6582( .i (n6581), .o (n6582) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n6583( .i (n5393), .o (n6583) );
  buffer buf_n6584( .i (n6583), .o (n6584) );
  assign n6585 = ( n1119 & ~n6291 ) | ( n1119 & n6584 ) | ( ~n6291 & n6584 ) ;
  buffer buf_n6586( .i (n6585), .o (n6586) );
  assign n6589 = n6497 & ~n6586 ;
  buffer buf_n6590( .i (n6589), .o (n6590) );
  buffer buf_n6591( .i (n6590), .o (n6591) );
  buffer buf_n6587( .i (n6586), .o (n6587) );
  buffer buf_n6588( .i (n6587), .o (n6588) );
  assign n6592 = n6588 | n6590 ;
  assign n6593 = ( ~n6149 & n6591 ) | ( ~n6149 & n6592 ) | ( n6591 & n6592 ) ;
  assign n6594 = n6521 & n6593 ;
  buffer buf_n6595( .i (n6563), .o (n6595) );
  buffer buf_n6596( .i (n6595), .o (n6596) );
  assign n6597 = ~n6594 & n6596 ;
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  assign n6598 = ~n555 & n568 ;
  assign n6599 = n6596 | n6598 ;
  assign n6600 = ~n6597 & n6599 ;
  buffer buf_n6601( .i (n6552), .o (n6601) );
  assign n6602 = ( ~n6246 & n6600 ) | ( ~n6246 & n6601 ) | ( n6600 & n6601 ) ;
  buffer buf_n6603( .i (n6330), .o (n6603) );
  assign n6604 = ( n3308 & n6392 ) | ( n3308 & ~n6603 ) | ( n6392 & ~n6603 ) ;
  buffer buf_n6605( .i (n6604), .o (n6605) );
  assign n6608 = n6012 & ~n6605 ;
  buffer buf_n6609( .i (n6608), .o (n6609) );
  buffer buf_n6610( .i (n6609), .o (n6610) );
  buffer buf_n6606( .i (n6605), .o (n6606) );
  buffer buf_n6607( .i (n6606), .o (n6607) );
  assign n6611 = n6607 | n6609 ;
  assign n6612 = ( ~n6510 & n6610 ) | ( ~n6510 & n6611 ) | ( n6610 & n6611 ) ;
  assign n6613 = n6563 | n6612 ;
  buffer buf_n3638( .i (n3637), .o (n3638) );
  buffer buf_n3639( .i (n3638), .o (n3639) );
  buffer buf_n3640( .i (n3639), .o (n3640) );
  assign n6614 = ~n3640 & n6563 ;
  assign n6615 = n6613 & ~n6614 ;
  assign n6616 = n6278 | n6615 ;
  assign n6617 = ( n4393 & n6271 ) | ( n4393 & ~n6469 ) | ( n6271 & ~n6469 ) ;
  buffer buf_n6618( .i (n6017), .o (n6618) );
  assign n6619 = ( n4393 & n6420 ) | ( n4393 & ~n6618 ) | ( n6420 & ~n6618 ) ;
  assign n6620 = n6617 & n6619 ;
  assign n6621 = n6595 & n6620 ;
  assign n6622 = n6278 & ~n6621 ;
  assign n6623 = n6616 & ~n6622 ;
  buffer buf_n6624( .i (n6570), .o (n6624) );
  assign n6625 = ( n6601 & ~n6623 ) | ( n6601 & n6624 ) | ( ~n6623 & n6624 ) ;
  assign n6626 = n6602 & ~n6625 ;
  buffer buf_n6627( .i (n6626), .o (n6627) );
  buffer buf_n6628( .i (n6627), .o (n6628) );
  buffer buf_n6629( .i (n6628), .o (n6629) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n720( .i (n719), .o (n720) );
  assign n6630 = ( n285 & n720 ) | ( n285 & n6627 ) | ( n720 & n6627 ) ;
  assign n6631 = n1730 | n6630 ;
  assign n6632 = ( ~n1731 & n6629 ) | ( ~n1731 & n6631 ) | ( n6629 & n6631 ) ;
  assign n6633 = ( n3912 & ~n5135 ) | ( n3912 & n6299 ) | ( ~n5135 & n6299 ) ;
  buffer buf_n6634( .i (n6633), .o (n6634) );
  buffer buf_n6635( .i (n6634), .o (n6635) );
  buffer buf_n6636( .i (n6635), .o (n6636) );
  buffer buf_n6637( .i (n6636), .o (n6637) );
  buffer buf_n6638( .i (n6299), .o (n6638) );
  buffer buf_n6639( .i (n6349), .o (n6639) );
  assign n6640 = ( n3913 & n6638 ) | ( n3913 & ~n6639 ) | ( n6638 & ~n6639 ) ;
  assign n6641 = n6634 & n6640 ;
  buffer buf_n6642( .i (n6641), .o (n6642) );
  buffer buf_n6643( .i (n6642), .o (n6643) );
  buffer buf_n6644( .i (n5742), .o (n6644) );
  assign n6645 = n6642 | n6644 ;
  assign n6646 = ( ~n6637 & n6643 ) | ( ~n6637 & n6645 ) | ( n6643 & n6645 ) ;
  buffer buf_n6647( .i (n6646), .o (n6647) );
  buffer buf_n6648( .i (n6647), .o (n6648) );
  buffer buf_n6649( .i (n6509), .o (n6649) );
  buffer buf_n6650( .i (n6649), .o (n6650) );
  assign n6651 = ( ~n6386 & n6647 ) | ( ~n6386 & n6650 ) | ( n6647 & n6650 ) ;
  assign n6652 = ( n3826 & n4119 ) | ( n3826 & n6164 ) | ( n4119 & n6164 ) ;
  assign n6653 = ~n4120 & n6652 ;
  assign n6654 = n6650 & n6653 ;
  assign n6655 = ( ~n6648 & n6651 ) | ( ~n6648 & n6654 ) | ( n6651 & n6654 ) ;
  buffer buf_n6656( .i (n6655), .o (n6656) );
  buffer buf_n6657( .i (n6656), .o (n6657) );
  buffer buf_n6658( .i (n6657), .o (n6658) );
  buffer buf_n5817( .i (n5816), .o (n5817) );
  buffer buf_n5818( .i (n5817), .o (n5818) );
  buffer buf_n5819( .i (n5818), .o (n5819) );
  buffer buf_n5820( .i (n5819), .o (n5820) );
  buffer buf_n5821( .i (n5820), .o (n5821) );
  buffer buf_n5822( .i (n5821), .o (n5822) );
  buffer buf_n5823( .i (n5822), .o (n5823) );
  assign n6659 = n5820 & ~n6507 ;
  buffer buf_n6660( .i (n6659), .o (n6660) );
  buffer buf_n6661( .i (n6660), .o (n6661) );
  buffer buf_n6662( .i (n6386), .o (n6662) );
  assign n6663 = ( n6426 & ~n6660 ) | ( n6426 & n6662 ) | ( ~n6660 & n6662 ) ;
  assign n6664 = ( n5823 & n6661 ) | ( n5823 & ~n6663 ) | ( n6661 & ~n6663 ) ;
  assign n6665 = ( ~n6570 & n6656 ) | ( ~n6570 & n6664 ) | ( n6656 & n6664 ) ;
  buffer buf_n6666( .i (n6346), .o (n6666) );
  assign n6667 = ~n6665 & n6666 ;
  assign n6668 = ( n148 & n6658 ) | ( n148 & ~n6667 ) | ( n6658 & ~n6667 ) ;
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  assign n6669 = ( n6273 & n6518 ) | ( n6273 & ~n6618 ) | ( n6518 & ~n6618 ) ;
  assign n6670 = ~n1167 & n6669 ;
  buffer buf_n6671( .i (n6469), .o (n6671) );
  buffer buf_n6672( .i (n6671), .o (n6672) );
  assign n6673 = n6670 & ~n6672 ;
  buffer buf_n6674( .i (n6276), .o (n6674) );
  assign n6675 = ( n6569 & n6673 ) | ( n6569 & ~n6674 ) | ( n6673 & ~n6674 ) ;
  assign n6676 = ~n6570 & n6675 ;
  buffer buf_n6677( .i (n6676), .o (n6677) );
  buffer buf_n6678( .i (n6677), .o (n6678) );
  buffer buf_n6679( .i (n5194), .o (n6679) );
  assign n6680 = n6677 | n6679 ;
  assign n6681 = ( n6668 & n6678 ) | ( n6668 & n6680 ) | ( n6678 & n6680 ) ;
  buffer buf_n6682( .i (n6436), .o (n6682) );
  assign n6683 = n6681 | n6682 ;
  buffer buf_n5449( .i (n5448), .o (n5449) );
  buffer buf_n5450( .i (n5449), .o (n5450) );
  buffer buf_n5451( .i (n5450), .o (n5451) );
  buffer buf_n6684( .i (n6672), .o (n6684) );
  assign n6685 = ( n4873 & n6427 ) | ( n4873 & n6684 ) | ( n6427 & n6684 ) ;
  assign n6686 = n5451 & ~n6685 ;
  assign n6687 = ( ~n5482 & n6601 ) | ( ~n5482 & n6686 ) | ( n6601 & n6686 ) ;
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  assign n6688 = n431 & n6684 ;
  assign n6689 = n879 & n6688 ;
  assign n6690 = ~n5482 & n6689 ;
  assign n6691 = ( ~n4895 & n6687 ) | ( ~n4895 & n6690 ) | ( n6687 & n6690 ) ;
  assign n6692 = ~n6248 & n6691 ;
  assign n6693 = n6682 & ~n6692 ;
  assign n6694 = n6683 & ~n6693 ;
  buffer buf_n4028( .i (n4027), .o (n4028) );
  buffer buf_n4029( .i (n4028), .o (n4029) );
  buffer buf_n4030( .i (n4029), .o (n4030) );
  buffer buf_n4031( .i (n4030), .o (n4031) );
  buffer buf_n4032( .i (n4031), .o (n4032) );
  buffer buf_n4033( .i (n4032), .o (n4033) );
  assign n6695 = ( n4696 & ~n6638 ) | ( n4696 & n6639 ) | ( ~n6638 & n6639 ) ;
  buffer buf_n6696( .i (n6695), .o (n6696) );
  buffer buf_n6697( .i (n6696), .o (n6697) );
  buffer buf_n6698( .i (n6697), .o (n6698) );
  buffer buf_n6699( .i (n6698), .o (n6699) );
  assign n6700 = ( n5735 & n6395 ) | ( n5735 & n6696 ) | ( n6395 & n6696 ) ;
  buffer buf_n6701( .i (n6700), .o (n6701) );
  buffer buf_n6702( .i (n6701), .o (n6702) );
  assign n6703 = ~n4700 & n6701 ;
  assign n6704 = ( ~n6699 & n6702 ) | ( ~n6699 & n6703 ) | ( n6702 & n6703 ) ;
  assign n6705 = n6671 & n6704 ;
  assign n6706 = ~n6568 & n6705 ;
  buffer buf_n6707( .i (n6706), .o (n6707) );
  buffer buf_n6708( .i (n6707), .o (n6708) );
  buffer buf_n6709( .i (n6708), .o (n6709) );
  buffer buf_n6710( .i (n6684), .o (n6710) );
  assign n6711 = ( n879 & n6707 ) | ( n879 & ~n6710 ) | ( n6707 & ~n6710 ) ;
  assign n6712 = n4032 & ~n6711 ;
  assign n6713 = ( n4033 & n6709 ) | ( n4033 & ~n6712 ) | ( n6709 & ~n6712 ) ;
  assign n6714 = ~n1506 & n2785 ;
  assign n6715 = ( ~n726 & n4878 ) | ( ~n726 & n5742 ) | ( n4878 & n5742 ) ;
  assign n6716 = n727 & n6715 ;
  assign n6717 = ( n4974 & n5365 ) | ( n4974 & ~n5899 ) | ( n5365 & ~n5899 ) ;
  buffer buf_n6718( .i (n6717), .o (n6718) );
  assign n6722 = ( n6223 & n6363 ) | ( n6223 & n6718 ) | ( n6363 & n6718 ) ;
  buffer buf_n6723( .i (n6722), .o (n6723) );
  buffer buf_n6724( .i (n6723), .o (n6724) );
  buffer buf_n6725( .i (n6724), .o (n6725) );
  buffer buf_n6719( .i (n6718), .o (n6719) );
  buffer buf_n6720( .i (n6719), .o (n6720) );
  buffer buf_n6721( .i (n6720), .o (n6721) );
  assign n6726 = ( n6330 & n6349 ) | ( n6330 & ~n6723 ) | ( n6349 & ~n6723 ) ;
  assign n6727 = n6721 | n6726 ;
  assign n6728 = ( n6335 & ~n6725 ) | ( n6335 & n6727 ) | ( ~n6725 & n6727 ) ;
  assign n6729 = ( n3915 & ~n6114 ) | ( n3915 & n6728 ) | ( ~n6114 & n6728 ) ;
  assign n6730 = ( n4692 & n5298 ) | ( n4692 & ~n5972 ) | ( n5298 & ~n5972 ) ;
  buffer buf_n6731( .i (n6730), .o (n6731) );
  buffer buf_n6734( .i (n5299), .o (n6734) );
  assign n6735 = ~n6731 & n6734 ;
  buffer buf_n6736( .i (n6735), .o (n6736) );
  buffer buf_n6737( .i (n6736), .o (n6737) );
  buffer buf_n6732( .i (n6731), .o (n6732) );
  buffer buf_n6733( .i (n6732), .o (n6733) );
  assign n6738 = n6733 | n6736 ;
  assign n6739 = ( ~n6311 & n6737 ) | ( ~n6311 & n6738 ) | ( n6737 & n6738 ) ;
  buffer buf_n6740( .i (n3914), .o (n6740) );
  buffer buf_n6741( .i (n6113), .o (n6741) );
  assign n6742 = ( ~n6739 & n6740 ) | ( ~n6739 & n6741 ) | ( n6740 & n6741 ) ;
  assign n6743 = n6729 | n6742 ;
  assign n6744 = ~n6716 & n6743 ;
  assign n6745 = ~n6714 & n6744 ;
  assign n6746 = ~n6650 & n6745 ;
  assign n6747 = ( n5165 & n6326 ) | ( n5165 & ~n6329 ) | ( n6326 & ~n6329 ) ;
  buffer buf_n6748( .i (n6747), .o (n6748) );
  buffer buf_n6749( .i (n6748), .o (n6749) );
  buffer buf_n6750( .i (n6749), .o (n6750) );
  buffer buf_n6751( .i (n6326), .o (n6751) );
  buffer buf_n6752( .i (n6751), .o (n6752) );
  assign n6753 = ( n6603 & n6748 ) | ( n6603 & ~n6752 ) | ( n6748 & ~n6752 ) ;
  assign n6754 = ( n6259 & ~n6311 ) | ( n6259 & n6753 ) | ( ~n6311 & n6753 ) ;
  assign n6755 = ( ~n441 & n6750 ) | ( ~n441 & n6754 ) | ( n6750 & n6754 ) ;
  assign n6756 = ~n6464 & n6755 ;
  assign n6757 = n633 & n872 ;
  assign n6758 = n6464 & ~n6757 ;
  assign n6759 = n6756 | n6758 ;
  assign n6760 = n4863 | n6759 ;
  assign n6761 = n6650 & n6760 ;
  assign n6762 = n6746 | n6761 ;
  buffer buf_n6763( .i (n5655), .o (n6763) );
  assign n6764 = n6762 & n6763 ;
  buffer buf_n6765( .i (n6638), .o (n6765) );
  buffer buf_n6766( .i (n6639), .o (n6766) );
  assign n6767 = ( n1609 & ~n6765 ) | ( n1609 & n6766 ) | ( ~n6765 & n6766 ) ;
  buffer buf_n6768( .i (n5135), .o (n6768) );
  assign n6769 = ( ~n1608 & n6639 ) | ( ~n1608 & n6768 ) | ( n6639 & n6768 ) ;
  buffer buf_n6770( .i (n6603), .o (n6770) );
  assign n6771 = ( ~n6765 & n6769 ) | ( ~n6765 & n6770 ) | ( n6769 & n6770 ) ;
  assign n6772 = ~n6767 & n6771 ;
  assign n6773 = n6399 & n6772 ;
  buffer buf_n6774( .i (n5298), .o (n6774) );
  assign n6775 = ( ~n4552 & n6223 ) | ( ~n4552 & n6774 ) | ( n6223 & n6774 ) ;
  buffer buf_n6776( .i (n6775), .o (n6776) );
  buffer buf_n6777( .i (n6776), .o (n6777) );
  buffer buf_n6778( .i (n6777), .o (n6778) );
  buffer buf_n6779( .i (n6778), .o (n6779) );
  buffer buf_n6780( .i (n4635), .o (n6780) );
  assign n6781 = ( ~n6330 & n6776 ) | ( ~n6330 & n6780 ) | ( n6776 & n6780 ) ;
  buffer buf_n6782( .i (n6781), .o (n6782) );
  buffer buf_n6783( .i (n6782), .o (n6783) );
  assign n6784 = n4556 & n6782 ;
  assign n6785 = ( ~n6779 & n6783 ) | ( ~n6779 & n6784 ) | ( n6783 & n6784 ) ;
  assign n6786 = n6399 | n6785 ;
  assign n6787 = ( ~n6340 & n6773 ) | ( ~n6340 & n6786 ) | ( n6773 & n6786 ) ;
  assign n6788 = n6649 & ~n6787 ;
  assign n6789 = ~n395 & n5735 ;
  assign n6790 = ( ~n2630 & n2719 ) | ( ~n2630 & n6789 ) | ( n2719 & n6789 ) ;
  assign n6791 = n6340 & ~n6790 ;
  assign n6792 = n6649 | n6791 ;
  assign n6793 = ~n6788 & n6792 ;
  assign n6794 = ~n6568 & n6793 ;
  assign n6795 = n6763 | n6794 ;
  assign n6796 = ~n6764 & n6795 ;
  buffer buf_n6797( .i (n6796), .o (n6797) );
  buffer buf_n6798( .i (n6797), .o (n6798) );
  assign n6799 = n2707 & ~n6797 ;
  assign n6800 = ( n6713 & n6798 ) | ( n6713 & ~n6799 ) | ( n6798 & ~n6799 ) ;
  assign n6801 = n5597 | n6800 ;
  buffer buf_n6802( .i (n606), .o (n6802) );
  assign n6803 = n557 | n6802 ;
  assign n6804 = ( n513 & n558 ) | ( n513 & n6803 ) | ( n558 & n6803 ) ;
  assign n6805 = n6340 & ~n6804 ;
  assign n6806 = n2134 & n6644 ;
  buffer buf_n6807( .i (n6395), .o (n6807) );
  buffer buf_n6808( .i (n6807), .o (n6808) );
  assign n6809 = n6806 | n6808 ;
  assign n6810 = ~n6805 & n6809 ;
  buffer buf_n6811( .i (n6810), .o (n6811) );
  buffer buf_n6812( .i (n6811), .o (n6812) );
  buffer buf_n6813( .i (n6812), .o (n6813) );
  buffer buf_n6814( .i (n6291), .o (n6814) );
  assign n6815 = ( n6388 & n6504 ) | ( n6388 & ~n6814 ) | ( n6504 & ~n6814 ) ;
  buffer buf_n6816( .i (n6815), .o (n6816) );
  buffer buf_n6817( .i (n6816), .o (n6817) );
  buffer buf_n6818( .i (n6506), .o (n6818) );
  assign n6819 = ( n6649 & n6817 ) | ( n6649 & ~n6818 ) | ( n6817 & ~n6818 ) ;
  assign n6820 = ~n6808 & n6816 ;
  assign n6821 = ( ~n6420 & n6817 ) | ( ~n6420 & n6820 ) | ( n6817 & n6820 ) ;
  assign n6822 = n6819 | n6821 ;
  assign n6823 = ( n6426 & n6811 ) | ( n6426 & ~n6822 ) | ( n6811 & ~n6822 ) ;
  buffer buf_n6824( .i (n6424), .o (n6824) );
  assign n6825 = ~n6823 & n6824 ;
  assign n6826 = ( n5692 & n6813 ) | ( n5692 & ~n6825 ) | ( n6813 & ~n6825 ) ;
  assign n6827 = ~n6666 & n6826 ;
  assign n6828 = ( ~n606 & n6335 ) | ( ~n606 & n6766 ) | ( n6335 & n6766 ) ;
  buffer buf_n6829( .i (n6828), .o (n6829) );
  buffer buf_n6830( .i (n6829), .o (n6830) );
  buffer buf_n6831( .i (n6830), .o (n6831) );
  buffer buf_n6832( .i (n6770), .o (n6832) );
  buffer buf_n6833( .i (n6832), .o (n6833) );
  assign n6834 = ( ~n6807 & n6829 ) | ( ~n6807 & n6833 ) | ( n6829 & n6833 ) ;
  assign n6835 = ( n6442 & ~n6517 ) | ( n6442 & n6834 ) | ( ~n6517 & n6834 ) ;
  assign n6836 = n6831 & n6835 ;
  buffer buf_n6837( .i (n6836), .o (n6837) );
  buffer buf_n6838( .i (n6837), .o (n6838) );
  assign n6839 = ( n6276 & ~n6547 ) | ( n6276 & n6837 ) | ( ~n6547 & n6837 ) ;
  assign n6840 = ( n2313 & n6807 ) | ( n2313 & n6833 ) | ( n6807 & n6833 ) ;
  buffer buf_n6841( .i (n6840), .o (n6841) );
  assign n6842 = ( ~n6618 & n6818 ) | ( ~n6618 & n6841 ) | ( n6818 & n6841 ) ;
  assign n6843 = ( n6195 & n6818 ) | ( n6195 & ~n6841 ) | ( n6818 & ~n6841 ) ;
  assign n6844 = n6842 & ~n6843 ;
  assign n6845 = ~n6276 & n6844 ;
  assign n6846 = ( n6838 & ~n6839 ) | ( n6838 & n6845 ) | ( ~n6839 & n6845 ) ;
  assign n6847 = ( n6326 & n6327 ) | ( n6326 & n6329 ) | ( n6327 & n6329 ) ;
  buffer buf_n6848( .i (n6847), .o (n6848) );
  assign n6854 = ( n6583 & ~n6638 ) | ( n6583 & n6848 ) | ( ~n6638 & n6848 ) ;
  buffer buf_n6855( .i (n6854), .o (n6855) );
  assign n6858 = n6388 & ~n6855 ;
  buffer buf_n6859( .i (n6858), .o (n6859) );
  buffer buf_n6860( .i (n6859), .o (n6860) );
  buffer buf_n6856( .i (n6855), .o (n6856) );
  buffer buf_n6857( .i (n6856), .o (n6857) );
  assign n6861 = n6857 | n6859 ;
  buffer buf_n6862( .i (n6442), .o (n6862) );
  assign n6863 = ( n6860 & n6861 ) | ( n6860 & ~n6862 ) | ( n6861 & ~n6862 ) ;
  buffer buf_n6864( .i (n6863), .o (n6864) );
  buffer buf_n6865( .i (n6864), .o (n6865) );
  buffer buf_n6866( .i (n6509), .o (n6866) );
  buffer buf_n6867( .i (n6866), .o (n6867) );
  buffer buf_n6868( .i (n6867), .o (n6868) );
  assign n6869 = ( n6426 & ~n6864 ) | ( n6426 & n6868 ) | ( ~n6864 & n6868 ) ;
  assign n6870 = ( ~n4467 & n6807 ) | ( ~n4467 & n6833 ) | ( n6807 & n6833 ) ;
  buffer buf_n6871( .i (n6870), .o (n6871) );
  buffer buf_n6872( .i (n6871), .o (n6872) );
  assign n6873 = n6195 & ~n6871 ;
  assign n6874 = ( n6422 & ~n6872 ) | ( n6422 & n6873 ) | ( ~n6872 & n6873 ) ;
  assign n6875 = n6868 & n6874 ;
  assign n6876 = ( n6865 & n6869 ) | ( n6865 & n6875 ) | ( n6869 & n6875 ) ;
  assign n6877 = n6846 | n6876 ;
  assign n6878 = n6666 & n6877 ;
  assign n6879 = n6827 | n6878 ;
  assign n6880 = ~n6248 & n6879 ;
  assign n6881 = n5597 & ~n6880 ;
  assign n6882 = n6801 & ~n6881 ;
  assign n6883 = n6694 | n6882 ;
  assign n6884 = ( ~n6581 & n6632 ) | ( ~n6581 & n6883 ) | ( n6632 & n6883 ) ;
  assign n6885 = n6582 | n6884 ;
  buffer buf_n239( .i (n238), .o (n239) );
  assign n6886 = n1748 & ~n6546 ;
  assign n6887 = n707 & ~n6886 ;
  assign n6888 = n728 & n6164 ;
  assign n6889 = ( n6818 & n6862 ) | ( n6818 & n6888 ) | ( n6862 & n6888 ) ;
  assign n6890 = ~n6149 & n6889 ;
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2306( .i (n2305), .o (n2306) );
  buffer buf_n2307( .i (n2306), .o (n2307) );
  buffer buf_n6891( .i (n6584), .o (n6891) );
  buffer buf_n6892( .i (n6891), .o (n6892) );
  assign n6893 = ( ~n4376 & n5983 ) | ( ~n4376 & n6892 ) | ( n5983 & n6892 ) ;
  assign n6894 = ( ~n4376 & n5983 ) | ( ~n4376 & n6644 ) | ( n5983 & n6644 ) ;
  assign n6895 = ( n2307 & n6893 ) | ( n2307 & ~n6894 ) | ( n6893 & ~n6894 ) ;
  buffer buf_n6896( .i (n6740), .o (n6896) );
  buffer buf_n6897( .i (n6896), .o (n6897) );
  buffer buf_n6898( .i (n6897), .o (n6898) );
  buffer buf_n6899( .i (n6506), .o (n6899) );
  assign n6900 = ( n6895 & ~n6898 ) | ( n6895 & n6899 ) | ( ~n6898 & n6899 ) ;
  buffer buf_n6901( .i (n6223), .o (n6901) );
  buffer buf_n6902( .i (n6901), .o (n6902) );
  assign n6903 = ( n5393 & n6751 ) | ( n5393 & ~n6902 ) | ( n6751 & ~n6902 ) ;
  buffer buf_n6904( .i (n6903), .o (n6904) );
  buffer buf_n6905( .i (n6904), .o (n6905) );
  buffer buf_n6906( .i (n6905), .o (n6906) );
  buffer buf_n6907( .i (n6906), .o (n6907) );
  buffer buf_n6909( .i (n6752), .o (n6909) );
  assign n6910 = n6904 & ~n6909 ;
  buffer buf_n6911( .i (n6910), .o (n6911) );
  buffer buf_n6912( .i (n6911), .o (n6912) );
  buffer buf_n6913( .i (n5717), .o (n6913) );
  assign n6914 = ( n6892 & ~n6911 ) | ( n6892 & n6913 ) | ( ~n6911 & n6913 ) ;
  assign n6915 = ( n6907 & n6912 ) | ( n6907 & ~n6914 ) | ( n6912 & ~n6914 ) ;
  assign n6916 = ( n6898 & n6899 ) | ( n6898 & ~n6915 ) | ( n6899 & ~n6915 ) ;
  assign n6917 = n6900 & ~n6916 ;
  assign n6918 = n6890 | n6917 ;
  assign n6919 = ( n708 & ~n6887 ) | ( n708 & n6918 ) | ( ~n6887 & n6918 ) ;
  assign n6920 = n6710 & n6919 ;
  buffer buf_n6921( .i (n5972), .o (n6921) );
  assign n6922 = ( n20 & n6364 ) | ( n20 & n6921 ) | ( n6364 & n6921 ) ;
  buffer buf_n6923( .i (n6922), .o (n6923) );
  assign n6928 = ( ~n3912 & n6299 ) | ( ~n3912 & n6923 ) | ( n6299 & n6923 ) ;
  buffer buf_n6929( .i (n6928), .o (n6929) );
  buffer buf_n6930( .i (n6929), .o (n6930) );
  buffer buf_n6931( .i (n6930), .o (n6931) );
  buffer buf_n6932( .i (n6931), .o (n6932) );
  assign n6933 = ( n6584 & n6766 ) | ( n6584 & n6929 ) | ( n6766 & n6929 ) ;
  buffer buf_n6934( .i (n6933), .o (n6934) );
  buffer buf_n6935( .i (n6934), .o (n6935) );
  buffer buf_n6924( .i (n6923), .o (n6924) );
  buffer buf_n6925( .i (n6924), .o (n6925) );
  buffer buf_n6926( .i (n6925), .o (n6926) );
  buffer buf_n6927( .i (n6926), .o (n6927) );
  assign n6936 = n6927 & ~n6934 ;
  assign n6937 = ( n6932 & ~n6935 ) | ( n6932 & n6936 ) | ( ~n6935 & n6936 ) ;
  buffer buf_n6938( .i (n6937), .o (n6938) );
  buffer buf_n6939( .i (n6938), .o (n6939) );
  buffer buf_n6940( .i (n6808), .o (n6940) );
  buffer buf_n6941( .i (n6940), .o (n6941) );
  buffer buf_n6942( .i (n6273), .o (n6942) );
  assign n6943 = ( n6938 & n6941 ) | ( n6938 & n6942 ) | ( n6941 & n6942 ) ;
  assign n6944 = n729 & ~n6561 ;
  assign n6945 = ~n6942 & n6944 ;
  assign n6946 = ( n6939 & ~n6943 ) | ( n6939 & n6945 ) | ( ~n6943 & n6945 ) ;
  buffer buf_n4474( .i (n4473), .o (n4474) );
  buffer buf_n4475( .i (n4474), .o (n4475) );
  buffer buf_n4476( .i (n4475), .o (n4476) );
  buffer buf_n4477( .i (n4476), .o (n4477) );
  buffer buf_n4478( .i (n4477), .o (n4478) );
  buffer buf_n4479( .i (n4478), .o (n4479) );
  buffer buf_n4480( .i (n4479), .o (n4480) );
  buffer buf_n4481( .i (n4480), .o (n4481) );
  assign n6947 = ( ~n754 & n4481 ) | ( ~n754 & n6484 ) | ( n4481 & n6484 ) ;
  assign n6948 = n755 & n6947 ;
  assign n6949 = n6946 | n6948 ;
  assign n6950 = ~n6710 & n6949 ;
  assign n6951 = n6920 | n6950 ;
  assign n6952 = ( n3855 & n6679 ) | ( n3855 & ~n6951 ) | ( n6679 & ~n6951 ) ;
  buffer buf_n6953( .i (n6952), .o (n6953) );
  buffer buf_n6954( .i (n6953), .o (n6954) );
  assign n6955 = n208 & ~n6953 ;
  assign n6956 = ( n239 & ~n6954 ) | ( n239 & n6955 ) | ( ~n6954 & n6955 ) ;
  buffer buf_n6957( .i (n6956), .o (n6957) );
  buffer buf_n6958( .i (n6957), .o (n6958) );
  assign n6959 = ~n6833 & n6896 ;
  assign n6960 = n6165 & ~n6959 ;
  assign n6961 = ( n610 & n2497 ) | ( n610 & ~n6960 ) | ( n2497 & ~n6960 ) ;
  assign n6962 = n6867 & ~n6961 ;
  assign n6963 = n3014 | n6898 ;
  assign n6964 = ~n6867 & n6963 ;
  assign n6965 = n6962 | n6964 ;
  buffer buf_n6966( .i (n6547), .o (n6966) );
  assign n6967 = n6965 & ~n6966 ;
  assign n6968 = n1186 & ~n6892 ;
  buffer buf_n6969( .i (n6968), .o (n6969) );
  buffer buf_n6970( .i (n6969), .o (n6970) );
  assign n6971 = ( ~n1187 & n6442 ) | ( ~n1187 & n6509 ) | ( n6442 & n6509 ) ;
  assign n6972 = n6969 | n6971 ;
  assign n6973 = ( n6149 & n6970 ) | ( n6149 & n6972 ) | ( n6970 & n6972 ) ;
  assign n6974 = n6568 | n6973 ;
  assign n6975 = n6966 & n6974 ;
  assign n6976 = n6967 | n6975 ;
  assign n6977 = ~n6601 & n6976 ;
  assign n6978 = ( n4586 & ~n6618 ) | ( n4586 & n6862 ) | ( ~n6618 & n6862 ) ;
  buffer buf_n6979( .i (n4585), .o (n6979) );
  assign n6980 = ( ~n6469 & n6862 ) | ( ~n6469 & n6979 ) | ( n6862 & n6979 ) ;
  assign n6981 = ( n659 & ~n6978 ) | ( n659 & n6980 ) | ( ~n6978 & n6980 ) ;
  assign n6982 = n6868 | n6981 ;
  assign n6983 = n350 & ~n6671 ;
  assign n6984 = n6868 & ~n6983 ;
  assign n6985 = n6982 & ~n6984 ;
  buffer buf_n6986( .i (n6569), .o (n6986) );
  assign n6987 = n6985 & ~n6986 ;
  buffer buf_n6988( .i (n6552), .o (n6988) );
  assign n6989 = ~n6987 & n6988 ;
  assign n6990 = n6977 | n6989 ;
  buffer buf_n6991( .i (n6435), .o (n6991) );
  assign n6992 = n6990 & ~n6991 ;
  buffer buf_n6993( .i (n6734), .o (n6993) );
  buffer buf_n6994( .i (n6993), .o (n6994) );
  assign n6995 = ( n6392 & n6603 ) | ( n6392 & n6994 ) | ( n6603 & n6994 ) ;
  buffer buf_n6996( .i (n6995), .o (n6996) );
  assign n7000 = ( n6504 & n6891 ) | ( n6504 & ~n6996 ) | ( n6891 & ~n6996 ) ;
  buffer buf_n7001( .i (n7000), .o (n7001) );
  buffer buf_n7002( .i (n7001), .o (n7002) );
  buffer buf_n7003( .i (n7002), .o (n7003) );
  buffer buf_n6997( .i (n6996), .o (n6997) );
  buffer buf_n6998( .i (n6997), .o (n6998) );
  buffer buf_n6999( .i (n6998), .o (n6999) );
  buffer buf_n7004( .i (n5891), .o (n7004) );
  assign n7005 = ( ~n6506 & n7001 ) | ( ~n6506 & n7004 ) | ( n7001 & n7004 ) ;
  assign n7006 = n6999 | n7005 ;
  buffer buf_n7007( .i (n6892), .o (n7007) );
  buffer buf_n7008( .i (n7007), .o (n7008) );
  buffer buf_n7009( .i (n7008), .o (n7009) );
  assign n7010 = ( n7003 & n7006 ) | ( n7003 & ~n7009 ) | ( n7006 & ~n7009 ) ;
  assign n7011 = n6672 & ~n7010 ;
  assign n7012 = ( ~n1760 & n4785 ) | ( ~n1760 & n6546 ) | ( n4785 & n6546 ) ;
  assign n7013 = n6672 | n7012 ;
  assign n7014 = ( ~n6684 & n7011 ) | ( ~n6684 & n7013 ) | ( n7011 & n7013 ) ;
  buffer buf_n7015( .i (n6202), .o (n7015) );
  assign n7016 = n7014 & n7015 ;
  buffer buf_n7017( .i (n6891), .o (n7017) );
  assign n7018 = ~n925 & n7017 ;
  buffer buf_n7019( .i (n7018), .o (n7019) );
  assign n7020 = ~n6866 & n7019 ;
  assign n7021 = ( ~n927 & n6899 ) | ( ~n927 & n7019 ) | ( n6899 & n7019 ) ;
  assign n7022 = ( ~n6422 & n7020 ) | ( ~n6422 & n7021 ) | ( n7020 & n7021 ) ;
  buffer buf_n7023( .i (n6671), .o (n7023) );
  assign n7024 = ~n7022 & n7023 ;
  buffer buf_n7025( .i (n6832), .o (n7025) );
  assign n7026 = ( n2699 & n6505 ) | ( n2699 & n7025 ) | ( n6505 & n7025 ) ;
  buffer buf_n7027( .i (n7026), .o (n7027) );
  buffer buf_n7028( .i (n7027), .o (n7028) );
  assign n7029 = n6899 & ~n7027 ;
  buffer buf_n7030( .i (n7025), .o (n7030) );
  buffer buf_n7031( .i (n7030), .o (n7031) );
  buffer buf_n7032( .i (n7031), .o (n7032) );
  assign n7033 = ( ~n7028 & n7029 ) | ( ~n7028 & n7032 ) | ( n7029 & n7032 ) ;
  assign n7034 = ~n7023 & n7033 ;
  buffer buf_n7035( .i (n7023), .o (n7035) );
  assign n7036 = ( ~n7024 & n7034 ) | ( ~n7024 & n7035 ) | ( n7034 & n7035 ) ;
  assign n7037 = n7015 | n7036 ;
  assign n7038 = ( ~n6988 & n7016 ) | ( ~n6988 & n7037 ) | ( n7016 & n7037 ) ;
  buffer buf_n7039( .i (n6624), .o (n7039) );
  assign n7040 = n7038 & ~n7039 ;
  assign n7041 = n6991 & ~n7040 ;
  assign n7042 = n6992 | n7041 ;
  buffer buf_n7043( .i (n180), .o (n7043) );
  assign n7044 = n7042 & n7043 ;
  buffer buf_n7045( .i (n6504), .o (n7045) );
  buffer buf_n7046( .i (n7045), .o (n7046) );
  buffer buf_n7047( .i (n7046), .o (n7047) );
  assign n7048 = ( n6866 & ~n6940 ) | ( n6866 & n7047 ) | ( ~n6940 & n7047 ) ;
  buffer buf_n7049( .i (n7048), .o (n7049) );
  buffer buf_n7050( .i (n7049), .o (n7050) );
  buffer buf_n7051( .i (n7050), .o (n7051) );
  assign n7052 = n6596 & n7050 ;
  assign n7053 = ( ~n4230 & n7051 ) | ( ~n4230 & n7052 ) | ( n7051 & n7052 ) ;
  assign n7054 = n6392 | n6994 ;
  buffer buf_n7055( .i (n7054), .o (n7055) );
  buffer buf_n7058( .i (n6765), .o (n7058) );
  assign n7059 = ( n6832 & n7055 ) | ( n6832 & ~n7058 ) | ( n7055 & ~n7058 ) ;
  assign n7060 = ( n6832 & n6891 ) | ( n6832 & n7055 ) | ( n6891 & n7055 ) ;
  assign n7061 = ( n6045 & n7059 ) | ( n6045 & ~n7060 ) | ( n7059 & ~n7060 ) ;
  buffer buf_n7062( .i (n6913), .o (n7062) );
  assign n7063 = n7061 & n7062 ;
  assign n7064 = n1236 & n7045 ;
  assign n7065 = n7062 | n7064 ;
  assign n7066 = ~n7063 & n7065 ;
  assign n7067 = n6941 & ~n7066 ;
  buffer buf_n7056( .i (n7055), .o (n7056) );
  buffer buf_n7057( .i (n7056), .o (n7057) );
  assign n7068 = ~n2933 & n7025 ;
  assign n7069 = ( ~n2121 & n7057 ) | ( ~n2121 & n7068 ) | ( n7057 & n7068 ) ;
  assign n7070 = n7008 | n7069 ;
  assign n7071 = ~n6941 & n7070 ;
  assign n7072 = n7067 | n7071 ;
  buffer buf_n7073( .i (n7072), .o (n7073) );
  buffer buf_n7074( .i (n7073), .o (n7074) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n5067( .i (n5066), .o (n5067) );
  buffer buf_n5068( .i (n5067), .o (n5068) );
  assign n7075 = ( n280 & n1750 ) | ( n280 & ~n5068 ) | ( n1750 & ~n5068 ) ;
  assign n7076 = n7073 & ~n7075 ;
  assign n7077 = ( ~n7053 & n7074 ) | ( ~n7053 & n7076 ) | ( n7074 & n7076 ) ;
  buffer buf_n7078( .i (n6666), .o (n7078) );
  assign n7079 = ~n7077 & n7078 ;
  buffer buf_n7080( .i (n6584), .o (n7080) );
  assign n7081 = ( n5027 & ~n6814 ) | ( n5027 & n7080 ) | ( ~n6814 & n7080 ) ;
  buffer buf_n7082( .i (n7081), .o (n7082) );
  assign n7085 = n7007 & ~n7082 ;
  buffer buf_n7086( .i (n7085), .o (n7086) );
  buffer buf_n7087( .i (n7086), .o (n7087) );
  buffer buf_n7083( .i (n7082), .o (n7083) );
  buffer buf_n7084( .i (n7083), .o (n7084) );
  assign n7088 = n7084 | n7086 ;
  assign n7089 = ( ~n5655 & n7087 ) | ( ~n5655 & n7088 ) | ( n7087 & n7088 ) ;
  assign n7090 = ( ~n6596 & n6966 ) | ( ~n6596 & n7089 ) | ( n6966 & n7089 ) ;
  buffer buf_n6110( .i (n6109), .o (n6110) );
  buffer buf_n6111( .i (n6110), .o (n6111) );
  buffer buf_n6112( .i (n6111), .o (n6112) );
  assign n7091 = ( n928 & n2572 ) | ( n928 & ~n6112 ) | ( n2572 & ~n6112 ) ;
  buffer buf_n7092( .i (n928), .o (n7092) );
  assign n7093 = ( n6424 & n7091 ) | ( n6424 & n7092 ) | ( n7091 & n7092 ) ;
  buffer buf_n7094( .i (n6595), .o (n7094) );
  assign n7095 = ( n6966 & n7093 ) | ( n6966 & n7094 ) | ( n7093 & n7094 ) ;
  assign n7096 = n7090 & n7095 ;
  buffer buf_n7097( .i (n6546), .o (n7097) );
  assign n7098 = n1761 | n7097 ;
  buffer buf_n7099( .i (n6662), .o (n7099) );
  assign n7100 = ( n7094 & ~n7098 ) | ( n7094 & n7099 ) | ( ~n7098 & n7099 ) ;
  assign n7101 = ~n6489 & n7100 ;
  assign n7102 = n7096 | n7101 ;
  assign n7103 = ~n7078 & n7102 ;
  assign n7104 = n7079 | n7103 ;
  assign n7105 = ~n5847 & n7104 ;
  assign n7106 = n7043 | n7105 ;
  assign n7107 = ~n7044 & n7106 ;
  assign n7108 = ( n1000 & n3913 ) | ( n1000 & n6768 ) | ( n3913 & n6768 ) ;
  buffer buf_n7109( .i (n7108), .o (n7109) );
  buffer buf_n7110( .i (n7109), .o (n7110) );
  buffer buf_n7111( .i (n7110), .o (n7111) );
  buffer buf_n7112( .i (n6770), .o (n7112) );
  assign n7113 = ( n6741 & ~n7109 ) | ( n6741 & n7112 ) | ( ~n7109 & n7112 ) ;
  assign n7114 = ( ~n6644 & n6896 ) | ( ~n6644 & n7113 ) | ( n6896 & n7113 ) ;
  assign n7115 = ~n7111 & n7114 ;
  assign n7116 = n6940 | n7115 ;
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  assign n7117 = n1639 & ~n6897 ;
  assign n7118 = n6940 & ~n7117 ;
  assign n7119 = n7116 & ~n7118 ;
  assign n7120 = n6662 | n7119 ;
  assign n7121 = ( n3370 & n6165 ) | ( n3370 & ~n6808 ) | ( n6165 & ~n6808 ) ;
  buffer buf_n7122( .i (n6741), .o (n7122) );
  buffer buf_n7123( .i (n7122), .o (n7123) );
  assign n7124 = ( n3370 & n6517 ) | ( n3370 & ~n7123 ) | ( n6517 & ~n7123 ) ;
  assign n7125 = n7121 & n7124 ;
  assign n7126 = ~n6567 & n7125 ;
  assign n7127 = n6662 & ~n7126 ;
  assign n7128 = n7120 & ~n7127 ;
  assign n7129 = n6475 | n7128 ;
  buffer buf_n7130( .i (n6909), .o (n7130) );
  assign n7131 = ( n2670 & ~n5717 ) | ( n2670 & n7130 ) | ( ~n5717 & n7130 ) ;
  buffer buf_n7132( .i (n5824), .o (n7132) );
  assign n7133 = ( n5138 & n7130 ) | ( n5138 & n7132 ) | ( n7130 & n7132 ) ;
  assign n7134 = ~n7131 & n7133 ;
  buffer buf_n7135( .i (n7134), .o (n7135) );
  buffer buf_n7136( .i (n7135), .o (n7136) );
  buffer buf_n7137( .i (n7136), .o (n7137) );
  buffer buf_n7138( .i (n7123), .o (n7138) );
  assign n7139 = ( n1005 & n7135 ) | ( n1005 & ~n7138 ) | ( n7135 & ~n7138 ) ;
  assign n7140 = n1948 & ~n7139 ;
  assign n7141 = ( n1949 & n7137 ) | ( n1949 & ~n7140 ) | ( n7137 & ~n7140 ) ;
  assign n7142 = ~n6569 & n7141 ;
  assign n7143 = n6475 & ~n7142 ;
  assign n7144 = n7129 & ~n7143 ;
  assign n7145 = ( n3855 & n6190 ) | ( n3855 & ~n7144 ) | ( n6190 & ~n7144 ) ;
  buffer buf_n7146( .i (n7145), .o (n7146) );
  buffer buf_n7147( .i (n7146), .o (n7147) );
  buffer buf_n7148( .i (n5774), .o (n7148) );
  buffer buf_n7149( .i (n7148), .o (n7149) );
  buffer buf_n7150( .i (n7149), .o (n7150) );
  buffer buf_n7151( .i (n7150), .o (n7151) );
  assign n7152 = ~n7146 & n7151 ;
  assign n7153 = ( n267 & ~n7147 ) | ( n267 & n7152 ) | ( ~n7147 & n7152 ) ;
  assign n7154 = ( n3913 & n5929 ) | ( n3913 & ~n6752 ) | ( n5929 & ~n6752 ) ;
  buffer buf_n7155( .i (n7154), .o (n7155) );
  buffer buf_n7160( .i (n6766), .o (n7160) );
  assign n7161 = ( n7130 & n7155 ) | ( n7130 & ~n7160 ) | ( n7155 & ~n7160 ) ;
  buffer buf_n7162( .i (n7161), .o (n7162) );
  buffer buf_n7163( .i (n7162), .o (n7163) );
  buffer buf_n7164( .i (n7163), .o (n7164) );
  buffer buf_n7165( .i (n7164), .o (n7165) );
  assign n7166 = ( n6897 & n7062 ) | ( n6897 & n7162 ) | ( n7062 & n7162 ) ;
  buffer buf_n7167( .i (n7166), .o (n7167) );
  buffer buf_n7168( .i (n7167), .o (n7168) );
  buffer buf_n7156( .i (n7155), .o (n7156) );
  buffer buf_n7157( .i (n7156), .o (n7157) );
  buffer buf_n7158( .i (n7157), .o (n7158) );
  buffer buf_n7159( .i (n7158), .o (n7159) );
  assign n7169 = n7159 & ~n7167 ;
  assign n7170 = ( n7165 & ~n7168 ) | ( n7165 & n7169 ) | ( ~n7168 & n7169 ) ;
  assign n7171 = ( n6824 & ~n7035 ) | ( n6824 & n7170 ) | ( ~n7035 & n7170 ) ;
  buffer buf_n7172( .i (n7171), .o (n7172) );
  assign n7173 = ( ~n5194 & n7148 ) | ( ~n5194 & n7172 ) | ( n7148 & n7172 ) ;
  buffer buf_n7174( .i (n6710), .o (n7174) );
  assign n7175 = ( ~n7148 & n7172 ) | ( ~n7148 & n7174 ) | ( n7172 & n7174 ) ;
  assign n7176 = n7173 & n7175 ;
  assign n7177 = ( ~n2631 & n7004 ) | ( ~n2631 & n7062 ) | ( n7004 & n7062 ) ;
  buffer buf_n7178( .i (n7177), .o (n7178) );
  buffer buf_n7179( .i (n7178), .o (n7179) );
  buffer buf_n7180( .i (n7179), .o (n7180) );
  assign n7181 = ( n6484 & ~n6942 ) | ( n6484 & n7178 ) | ( ~n6942 & n7178 ) ;
  buffer buf_n7182( .i (n6867), .o (n7182) );
  assign n7183 = ( n6424 & n7181 ) | ( n6424 & ~n7182 ) | ( n7181 & ~n7182 ) ;
  assign n7184 = n7180 & n7183 ;
  buffer buf_n7185( .i (n7184), .o (n7185) );
  buffer buf_n7186( .i (n7185), .o (n7186) );
  buffer buf_n7187( .i (n733), .o (n7187) );
  assign n7188 = ( n7174 & n7185 ) | ( n7174 & ~n7187 ) | ( n7185 & ~n7187 ) ;
  assign n7189 = n7186 & ~n7188 ;
  assign n7190 = n7176 | n7189 ;
  assign n7191 = n120 | n7190 ;
  assign n7192 = ~n2010 & n7032 ;
  assign n7193 = ( ~n2124 & n3870 ) | ( ~n2124 & n7192 ) | ( n3870 & n7192 ) ;
  assign n7194 = n7094 & ~n7193 ;
  buffer buf_n7195( .i (n7138), .o (n7195) );
  buffer buf_n7196( .i (n2041), .o (n7196) );
  assign n7197 = ( n6942 & ~n7195 ) | ( n6942 & n7196 ) | ( ~n7195 & n7196 ) ;
  buffer buf_n7198( .i (n2040), .o (n7198) );
  assign n7199 = ( n6866 & n7138 ) | ( n6866 & n7198 ) | ( n7138 & n7198 ) ;
  buffer buf_n7200( .i (n6913), .o (n7200) );
  buffer buf_n7201( .i (n7200), .o (n7201) );
  buffer buf_n7202( .i (n7201), .o (n7202) );
  assign n7203 = ( n7032 & ~n7199 ) | ( n7032 & n7202 ) | ( ~n7199 & n7202 ) ;
  assign n7204 = ~n7197 & n7203 ;
  assign n7205 = n7094 | n7204 ;
  assign n7206 = ( ~n6489 & n7194 ) | ( ~n6489 & n7205 ) | ( n7194 & n7205 ) ;
  assign n7207 = n5284 | n7206 ;
  assign n7208 = n6595 & n7182 ;
  buffer buf_n7209( .i (n7032), .o (n7209) );
  assign n7210 = n542 | n7209 ;
  assign n7211 = ( ~n2099 & n7208 ) | ( ~n2099 & n7210 ) | ( n7208 & n7210 ) ;
  buffer buf_n7212( .i (n7035), .o (n7212) );
  assign n7213 = n7211 & ~n7212 ;
  buffer buf_n7214( .i (n6480), .o (n7214) );
  assign n7215 = ~n7213 & n7214 ;
  assign n7216 = n7207 & ~n7215 ;
  assign n7217 = ~n6248 & n7216 ;
  buffer buf_n7218( .i (n6178), .o (n7218) );
  buffer buf_n7219( .i (n7218), .o (n7219) );
  assign n7220 = ~n7217 & n7219 ;
  assign n7221 = n7191 & ~n7220 ;
  assign n7222 = n7153 | n7221 ;
  assign n7223 = ( ~n6957 & n7107 ) | ( ~n6957 & n7222 ) | ( n7107 & n7222 ) ;
  assign n7224 = n6958 | n7223 ;
  buffer buf_n4932( .i (n4931), .o (n4932) );
  buffer buf_n4933( .i (n4932), .o (n4933) );
  buffer buf_n4934( .i (n4933), .o (n4934) );
  buffer buf_n4935( .i (n4934), .o (n4935) );
  buffer buf_n4936( .i (n4935), .o (n4936) );
  buffer buf_n4626( .i (n4625), .o (n4626) );
  buffer buf_n4627( .i (n4626), .o (n4627) );
  buffer buf_n4628( .i (n4627), .o (n4628) );
  buffer buf_n4629( .i (n4628), .o (n4629) );
  buffer buf_n4630( .i (n4629), .o (n4630) );
  assign n7225 = ( n760 & n4630 ) | ( n760 & ~n4935 ) | ( n4630 & ~n4935 ) ;
  buffer buf_n5069( .i (n5068), .o (n5069) );
  buffer buf_n7226( .i (n6941), .o (n7226) );
  buffer buf_n7227( .i (n7226), .o (n7227) );
  buffer buf_n7228( .i (n7227), .o (n7228) );
  assign n7229 = ( n5069 & ~n6475 ) | ( n5069 & n7228 ) | ( ~n6475 & n7228 ) ;
  assign n7230 = ~n6527 & n7229 ;
  assign n7231 = n7039 & n7230 ;
  assign n7232 = n4630 & n7231 ;
  assign n7233 = ( n4936 & n7225 ) | ( n4936 & n7232 ) | ( n7225 & n7232 ) ;
  buffer buf_n7234( .i (n7233), .o (n7234) );
  buffer buf_n7235( .i (n7234), .o (n7235) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  assign n7236 = n573 & ~n6191 ;
  buffer buf_n7237( .i (n6189), .o (n7237) );
  assign n7238 = n7236 & n7237 ;
  buffer buf_n7239( .i (n6363), .o (n7239) );
  assign n7240 = ( n6734 & n6901 ) | ( n6734 & ~n7239 ) | ( n6901 & ~n7239 ) ;
  buffer buf_n7241( .i (n7240), .o (n7241) );
  buffer buf_n7246( .i (n6902), .o (n7246) );
  assign n7247 = ( n6583 & ~n7241 ) | ( n6583 & n7246 ) | ( ~n7241 & n7246 ) ;
  buffer buf_n7248( .i (n7247), .o (n7248) );
  buffer buf_n7249( .i (n7248), .o (n7249) );
  buffer buf_n7250( .i (n7249), .o (n7250) );
  buffer buf_n7251( .i (n7250), .o (n7251) );
  assign n7252 = ( ~n7058 & n7130 ) | ( ~n7058 & n7248 ) | ( n7130 & n7248 ) ;
  buffer buf_n7253( .i (n7252), .o (n7253) );
  buffer buf_n7254( .i (n7253), .o (n7254) );
  buffer buf_n7242( .i (n7241), .o (n7242) );
  buffer buf_n7243( .i (n7242), .o (n7243) );
  buffer buf_n7244( .i (n7243), .o (n7244) );
  buffer buf_n7245( .i (n7244), .o (n7245) );
  assign n7255 = n7245 & n7253 ;
  assign n7256 = ( ~n7251 & n7254 ) | ( ~n7251 & n7255 ) | ( n7254 & n7255 ) ;
  assign n7257 = ~n7195 & n7256 ;
  buffer buf_n7258( .i (n6567), .o (n7258) );
  assign n7259 = n7257 & ~n7258 ;
  buffer buf_n7260( .i (n7259), .o (n7260) );
  buffer buf_n7261( .i (n7260), .o (n7261) );
  buffer buf_n4499( .i (n4498), .o (n4499) );
  buffer buf_n4500( .i (n4499), .o (n4500) );
  buffer buf_n4501( .i (n4500), .o (n4501) );
  assign n7262 = n4501 | n7260 ;
  assign n7263 = ( n4032 & n7261 ) | ( n4032 & n7262 ) | ( n7261 & n7262 ) ;
  assign n7264 = ~n4895 & n7263 ;
  buffer buf_n7265( .i (n7264), .o (n7265) );
  buffer buf_n7266( .i (n7265), .o (n7266) );
  assign n7267 = n761 | n7265 ;
  assign n7268 = ( n7238 & n7266 ) | ( n7238 & n7267 ) | ( n7266 & n7267 ) ;
  buffer buf_n7269( .i (n4559), .o (n7269) );
  assign n7270 = ( n3911 & ~n6327 ) | ( n3911 & n7269 ) | ( ~n6327 & n7269 ) ;
  buffer buf_n7271( .i (n7270), .o (n7271) );
  buffer buf_n7276( .i (n6370), .o (n7276) );
  assign n7277 = ( n6768 & n7271 ) | ( n6768 & ~n7276 ) | ( n7271 & ~n7276 ) ;
  buffer buf_n7278( .i (n7277), .o (n7278) );
  buffer buf_n7279( .i (n7278), .o (n7279) );
  buffer buf_n7280( .i (n7279), .o (n7280) );
  buffer buf_n7281( .i (n7280), .o (n7281) );
  assign n7282 = ( n6740 & ~n7080 ) | ( n6740 & n7278 ) | ( ~n7080 & n7278 ) ;
  buffer buf_n7283( .i (n7282), .o (n7283) );
  buffer buf_n7284( .i (n7283), .o (n7284) );
  buffer buf_n7272( .i (n7271), .o (n7272) );
  buffer buf_n7273( .i (n7272), .o (n7273) );
  buffer buf_n7274( .i (n7273), .o (n7274) );
  buffer buf_n7275( .i (n7274), .o (n7275) );
  assign n7285 = ~n7275 & n7283 ;
  assign n7286 = ( ~n7281 & n7284 ) | ( ~n7281 & n7285 ) | ( n7284 & n7285 ) ;
  assign n7287 = n7202 | n7286 ;
  assign n7288 = n3121 & n7123 ;
  assign n7289 = ~n6898 & n7288 ;
  assign n7290 = n7202 & ~n7289 ;
  assign n7291 = n7287 & ~n7290 ;
  assign n7292 = n7227 | n7291 ;
  buffer buf_n7293( .i (n6583), .o (n7293) );
  assign n7294 = n5824 & n7293 ;
  assign n7295 = ( n6741 & n6814 ) | ( n6741 & n7294 ) | ( n6814 & n7294 ) ;
  buffer buf_n7296( .i (n7295), .o (n7296) );
  buffer buf_n7297( .i (n7296), .o (n7297) );
  buffer buf_n7298( .i (n7297), .o (n7298) );
  assign n7299 = ( n7004 & n7007 ) | ( n7004 & ~n7296 ) | ( n7007 & ~n7296 ) ;
  assign n7300 = ( n7138 & n7201 ) | ( n7138 & n7299 ) | ( n7201 & n7299 ) ;
  assign n7301 = ~n7298 & n7300 ;
  assign n7302 = ~n7258 & n7301 ;
  assign n7303 = n7227 & ~n7302 ;
  assign n7304 = n7292 & ~n7303 ;
  assign n7305 = n7214 | n7304 ;
  buffer buf_n7306( .i (n5300), .o (n7306) );
  assign n7307 = ( n5924 & n7269 ) | ( n5924 & n7306 ) | ( n7269 & n7306 ) ;
  buffer buf_n7308( .i (n7307), .o (n7308) );
  buffer buf_n7309( .i (n7308), .o (n7309) );
  buffer buf_n7310( .i (n7309), .o (n7310) );
  buffer buf_n7311( .i (n7310), .o (n7311) );
  buffer buf_n7312( .i (n7311), .o (n7312) );
  buffer buf_n7313( .i (n7312), .o (n7313) );
  buffer buf_n7314( .i (n7313), .o (n7314) );
  buffer buf_n7315( .i (n7314), .o (n7315) );
  buffer buf_n7316( .i (n7123), .o (n7316) );
  buffer buf_n7317( .i (n7004), .o (n7317) );
  assign n7318 = ( ~n7313 & n7316 ) | ( ~n7313 & n7317 ) | ( n7316 & n7317 ) ;
  buffer buf_n7319( .i (n6909), .o (n7319) );
  buffer buf_n7320( .i (n7319), .o (n7320) );
  buffer buf_n7321( .i (n7320), .o (n7321) );
  buffer buf_n7322( .i (n7321), .o (n7322) );
  buffer buf_n7323( .i (n7322), .o (n7323) );
  assign n7324 = ( n7195 & n7318 ) | ( n7195 & n7323 ) | ( n7318 & n7323 ) ;
  assign n7325 = ( n1949 & n7315 ) | ( n1949 & ~n7324 ) | ( n7315 & ~n7324 ) ;
  assign n7326 = n746 & n1766 ;
  buffer buf_n7327( .i (n7326), .o (n7327) );
  buffer buf_n7328( .i (n7327), .o (n7328) );
  assign n7329 = n5655 | n7327 ;
  assign n7330 = ( n7325 & n7328 ) | ( n7325 & n7329 ) | ( n7328 & n7329 ) ;
  assign n7331 = ~n6986 & n7330 ;
  assign n7332 = n7214 & ~n7331 ;
  assign n7333 = n7305 & ~n7332 ;
  assign n7334 = n7218 | n7333 ;
  buffer buf_n4330( .i (n4329), .o (n4330) );
  buffer buf_n4331( .i (n4330), .o (n4331) );
  assign n7335 = ( n2212 & ~n7008 ) | ( n2212 & n7317 ) | ( ~n7008 & n7317 ) ;
  assign n7336 = ( n2212 & n7317 ) | ( n2212 & n7322 ) | ( n7317 & n7322 ) ;
  assign n7337 = ( n4331 & n7335 ) | ( n4331 & ~n7336 ) | ( n7335 & ~n7336 ) ;
  assign n7338 = n7023 & n7337 ;
  assign n7339 = ( n5393 & ~n6370 ) | ( n5393 & n6751 ) | ( ~n6370 & n6751 ) ;
  buffer buf_n7340( .i (n7339), .o (n7340) );
  buffer buf_n7346( .i (n7246), .o (n7346) );
  assign n7347 = ( n7293 & n7340 ) | ( n7293 & ~n7346 ) | ( n7340 & ~n7346 ) ;
  buffer buf_n7348( .i (n7347), .o (n7348) );
  assign n7351 = n7017 & ~n7348 ;
  buffer buf_n7352( .i (n7351), .o (n7352) );
  buffer buf_n7353( .i (n7352), .o (n7353) );
  buffer buf_n7349( .i (n7348), .o (n7349) );
  buffer buf_n7350( .i (n7349), .o (n7350) );
  assign n7354 = n7350 | n7352 ;
  assign n7355 = ( ~n7009 & n7353 ) | ( ~n7009 & n7354 ) | ( n7353 & n7354 ) ;
  buffer buf_n7356( .i (n7195), .o (n7356) );
  assign n7357 = n7355 | n7356 ;
  assign n7358 = ( ~n7035 & n7338 ) | ( ~n7035 & n7357 ) | ( n7338 & n7357 ) ;
  assign n7359 = n7015 & n7358 ;
  assign n7360 = ( n6291 & ~n6904 ) | ( n6291 & n6909 ) | ( ~n6904 & n6909 ) ;
  buffer buf_n7361( .i (n7360), .o (n7361) );
  buffer buf_n7362( .i (n7361), .o (n7362) );
  buffer buf_n7363( .i (n7362), .o (n7363) );
  buffer buf_n7364( .i (n7363), .o (n7364) );
  buffer buf_n7365( .i (n7160), .o (n7365) );
  assign n7366 = ( ~n7017 & n7361 ) | ( ~n7017 & n7365 ) | ( n7361 & n7365 ) ;
  buffer buf_n7367( .i (n7366), .o (n7367) );
  buffer buf_n7368( .i (n7367), .o (n7368) );
  buffer buf_n6908( .i (n6907), .o (n6908) );
  assign n7369 = n6908 & n7367 ;
  assign n7370 = ( ~n7364 & n7368 ) | ( ~n7364 & n7369 ) | ( n7368 & n7369 ) ;
  assign n7371 = n7356 & ~n7370 ;
  buffer buf_n3615( .i (n3614), .o (n3615) );
  assign n7372 = n3615 | n4421 ;
  assign n7373 = ~n7323 & n7372 ;
  assign n7374 = n7356 | n7373 ;
  assign n7375 = ~n7371 & n7374 ;
  assign n7376 = n7015 | n7375 ;
  assign n7377 = ( ~n6988 & n7359 ) | ( ~n6988 & n7376 ) | ( n7359 & n7376 ) ;
  assign n7378 = ~n7039 & n7377 ;
  assign n7379 = n7218 & ~n7378 ;
  assign n7380 = n7334 & ~n7379 ;
  assign n7381 = n1399 & n2611 ;
  assign n7382 = n445 & n7381 ;
  buffer buf_n7383( .i (n7382), .o (n7383) );
  buffer buf_n7384( .i (n7383), .o (n7384) );
  buffer buf_n7385( .i (n7384), .o (n7385) );
  buffer buf_n7386( .i (n6814), .o (n7386) );
  buffer buf_n7387( .i (n7386), .o (n7387) );
  assign n7388 = ( n2211 & ~n7321 ) | ( n2211 & n7387 ) | ( ~n7321 & n7387 ) ;
  assign n7389 = ( ~n2210 & n7017 ) | ( ~n2210 & n7386 ) | ( n7017 & n7386 ) ;
  assign n7390 = ( n6517 & ~n7321 ) | ( n6517 & n7389 ) | ( ~n7321 & n7389 ) ;
  assign n7391 = ~n7388 & n7390 ;
  buffer buf_n7392( .i (n7047), .o (n7392) );
  assign n7393 = n7391 | n7392 ;
  assign n7394 = n3281 | n7322 ;
  assign n7395 = n7392 & n7394 ;
  assign n7396 = n7393 & ~n7395 ;
  buffer buf_n7397( .i (n7258), .o (n7397) );
  assign n7398 = ( n7383 & n7396 ) | ( n7383 & ~n7397 ) | ( n7396 & ~n7397 ) ;
  buffer buf_n7399( .i (n7099), .o (n7399) );
  assign n7400 = ~n7398 & n7399 ;
  assign n7401 = ( n6988 & n7385 ) | ( n6988 & ~n7400 ) | ( n7385 & ~n7400 ) ;
  buffer buf_n7402( .i (n7401), .o (n7402) );
  buffer buf_n7403( .i (n7402), .o (n7403) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  assign n7404 = n1202 & n7402 ;
  buffer buf_n4539( .i (n4538), .o (n4539) );
  buffer buf_n4540( .i (n4539), .o (n4540) );
  assign n7405 = n4540 & ~n6816 ;
  buffer buf_n7406( .i (n7405), .o (n7406) );
  buffer buf_n7407( .i (n7406), .o (n7407) );
  assign n7408 = n794 & n7269 ;
  buffer buf_n7409( .i (n7269), .o (n7409) );
  assign n7410 = ( n2882 & ~n7408 ) | ( n2882 & n7409 ) | ( ~n7408 & n7409 ) ;
  buffer buf_n7411( .i (n6327), .o (n7411) );
  buffer buf_n7412( .i (n7411), .o (n7412) );
  assign n7413 = ( n6994 & n7410 ) | ( n6994 & ~n7412 ) | ( n7410 & ~n7412 ) ;
  buffer buf_n7414( .i (n7413), .o (n7414) );
  assign n7415 = ( n7080 & ~n7112 ) | ( n7080 & n7414 ) | ( ~n7112 & n7414 ) ;
  assign n7416 = ( ~n7058 & n7112 ) | ( ~n7058 & n7414 ) | ( n7112 & n7414 ) ;
  assign n7417 = n7415 | n7416 ;
  buffer buf_n7418( .i (n7417), .o (n7418) );
  buffer buf_n7419( .i (n7418), .o (n7419) );
  buffer buf_n7420( .i (n7419), .o (n7420) );
  assign n7421 = ( n6518 & n7316 ) | ( n6518 & n7418 ) | ( n7316 & n7418 ) ;
  assign n7422 = n7406 & n7421 ;
  assign n7423 = ( ~n7407 & n7420 ) | ( ~n7407 & n7422 ) | ( n7420 & n7422 ) ;
  assign n7424 = n7099 & ~n7423 ;
  buffer buf_n2285( .i (n2284), .o (n2285) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n7425( .i (n7276), .o (n7425) );
  buffer buf_n7426( .i (n7425), .o (n7426) );
  assign n7427 = ( ~n7112 & n7160 ) | ( ~n7112 & n7426 ) | ( n7160 & n7426 ) ;
  buffer buf_n7428( .i (n7080), .o (n7428) );
  assign n7429 = n7427 | n7428 ;
  assign n7430 = ~n2287 & n7429 ;
  assign n7431 = ( n7047 & ~n7316 ) | ( n7047 & n7430 ) | ( ~n7316 & n7430 ) ;
  assign n7432 = ( n491 & n922 ) | ( n491 & n7246 ) | ( n922 & n7246 ) ;
  buffer buf_n7433( .i (n7432), .o (n7433) );
  buffer buf_n7434( .i (n7433), .o (n7434) );
  buffer buf_n7435( .i (n7434), .o (n7435) );
  buffer buf_n7436( .i (n6770), .o (n7436) );
  assign n7437 = ( ~n7160 & n7433 ) | ( ~n7160 & n7436 ) | ( n7433 & n7436 ) ;
  assign n7438 = ( n494 & ~n7428 ) | ( n494 & n7437 ) | ( ~n7428 & n7437 ) ;
  assign n7439 = ( ~n495 & n7435 ) | ( ~n495 & n7438 ) | ( n7435 & n7438 ) ;
  assign n7440 = ( n7047 & n7316 ) | ( n7047 & ~n7439 ) | ( n7316 & ~n7439 ) ;
  assign n7441 = n7431 & ~n7440 ;
  assign n7442 = ( n1502 & n7276 ) | ( n1502 & n7412 ) | ( n7276 & n7412 ) ;
  buffer buf_n7443( .i (n7442), .o (n7443) );
  buffer buf_n7444( .i (n7443), .o (n7444) );
  buffer buf_n7445( .i (n7444), .o (n7445) );
  buffer buf_n7446( .i (n7346), .o (n7446) );
  assign n7447 = ( n7426 & ~n7443 ) | ( n7426 & n7446 ) | ( ~n7443 & n7446 ) ;
  assign n7448 = ( n7025 & n7428 ) | ( n7025 & n7447 ) | ( n7428 & n7447 ) ;
  assign n7449 = n7445 & ~n7448 ;
  buffer buf_n7450( .i (n7046), .o (n7450) );
  buffer buf_n7451( .i (n7122), .o (n7451) );
  buffer buf_n7452( .i (n7451), .o (n7452) );
  assign n7453 = ( n7449 & ~n7450 ) | ( n7449 & n7452 ) | ( ~n7450 & n7452 ) ;
  buffer buf_n7454( .i (n7436), .o (n7454) );
  assign n7455 = ( n2260 & n7428 ) | ( n2260 & n7454 ) | ( n7428 & n7454 ) ;
  buffer buf_n7456( .i (n7293), .o (n7456) );
  buffer buf_n7457( .i (n7456), .o (n7457) );
  assign n7458 = ( n2260 & n7365 ) | ( n2260 & n7457 ) | ( n7365 & n7457 ) ;
  assign n7459 = ( n874 & n7455 ) | ( n874 & ~n7458 ) | ( n7455 & ~n7458 ) ;
  assign n7460 = ( n7450 & n7452 ) | ( n7450 & n7459 ) | ( n7452 & n7459 ) ;
  assign n7461 = n7453 & n7460 ;
  assign n7462 = n7441 | n7461 ;
  assign n7463 = ~n7099 & n7462 ;
  assign n7464 = n7424 | n7463 ;
  assign n7465 = ( n6527 & ~n6624 ) | ( n6527 & n7464 ) | ( ~n6624 & n7464 ) ;
  assign n7466 = n394 & n2175 ;
  buffer buf_n7467( .i (n7466), .o (n7467) );
  buffer buf_n7468( .i (n7467), .o (n7468) );
  assign n7469 = n4752 | n7425 ;
  assign n7470 = ( n4752 & ~n7293 ) | ( n4752 & n7425 ) | ( ~n7293 & n7425 ) ;
  assign n7471 = ( n7456 & ~n7469 ) | ( n7456 & n7470 ) | ( ~n7469 & n7470 ) ;
  assign n7472 = n7467 | n7471 ;
  assign n7473 = ( ~n7030 & n7468 ) | ( ~n7030 & n7472 ) | ( n7468 & n7472 ) ;
  assign n7474 = n7201 | n7473 ;
  assign n7475 = n1118 & ~n7412 ;
  buffer buf_n7476( .i (n7475), .o (n7476) );
  buffer buf_n7477( .i (n7476), .o (n7477) );
  buffer buf_n7478( .i (n6113), .o (n7478) );
  assign n7479 = ( n7058 & ~n7476 ) | ( n7058 & n7478 ) | ( ~n7476 & n7478 ) ;
  assign n7480 = ( n1121 & n7477 ) | ( n1121 & ~n7479 ) | ( n7477 & ~n7479 ) ;
  assign n7481 = n7387 & n7480 ;
  assign n7482 = n7201 & ~n7481 ;
  assign n7483 = n7474 & ~n7482 ;
  assign n7484 = ( n4751 & n6768 ) | ( n4751 & ~n7276 ) | ( n6768 & ~n7276 ) ;
  buffer buf_n7485( .i (n7484), .o (n7485) );
  assign n7488 = n7478 & ~n7485 ;
  buffer buf_n7489( .i (n7488), .o (n7489) );
  buffer buf_n7490( .i (n7489), .o (n7490) );
  buffer buf_n7486( .i (n7485), .o (n7486) );
  buffer buf_n7487( .i (n7486), .o (n7487) );
  assign n7491 = n7487 | n7489 ;
  assign n7492 = ( ~n7452 & n7490 ) | ( ~n7452 & n7491 ) | ( n7490 & n7491 ) ;
  buffer buf_n7493( .i (n7031), .o (n7493) );
  assign n7494 = ( ~n7202 & n7492 ) | ( ~n7202 & n7493 ) | ( n7492 & n7493 ) ;
  assign n7495 = ( ~n5067 & n7483 ) | ( ~n5067 & n7494 ) | ( n7483 & n7494 ) ;
  buffer buf_n7496( .i (n6484), .o (n7496) );
  buffer buf_n7497( .i (n7496), .o (n7497) );
  assign n7498 = n7495 & ~n7497 ;
  buffer buf_n7499( .i (n6765), .o (n7499) );
  assign n7500 = ( n5242 & ~n7436 ) | ( n5242 & n7499 ) | ( ~n7436 & n7499 ) ;
  buffer buf_n7501( .i (n5929), .o (n7501) );
  assign n7502 = ~n5241 & n7501 ;
  assign n7503 = ( ~n5242 & n7456 ) | ( ~n5242 & n7502 ) | ( n7456 & n7502 ) ;
  assign n7504 = n7500 & ~n7503 ;
  assign n7505 = n7387 | n7504 ;
  buffer buf_n7506( .i (n6329), .o (n7506) );
  buffer buf_n7507( .i (n7506), .o (n7507) );
  buffer buf_n7508( .i (n7507), .o (n7508) );
  assign n7509 = n5026 | n7508 ;
  assign n7510 = ( n5027 & ~n7132 ) | ( n5027 & n7509 ) | ( ~n7132 & n7509 ) ;
  assign n7511 = n7045 & ~n7510 ;
  assign n7512 = n7387 & ~n7511 ;
  assign n7513 = n7505 & ~n7512 ;
  buffer buf_n7514( .i (n7452), .o (n7514) );
  assign n7515 = n7513 & n7514 ;
  assign n7516 = n1253 & n7317 ;
  assign n7517 = n611 & n7516 ;
  assign n7518 = n7515 | n7517 ;
  assign n7519 = n7497 & n7518 ;
  assign n7520 = n7498 | n7519 ;
  assign n7521 = ( n6527 & n6624 ) | ( n6527 & ~n7520 ) | ( n6624 & ~n7520 ) ;
  assign n7522 = n7465 & ~n7521 ;
  buffer buf_n7523( .i (n7409), .o (n7523) );
  assign n7524 = ( n7308 & n7507 ) | ( n7308 & ~n7523 ) | ( n7507 & ~n7523 ) ;
  buffer buf_n7525( .i (n7524), .o (n7525) );
  buffer buf_n7526( .i (n7525), .o (n7526) );
  buffer buf_n7527( .i (n7526), .o (n7527) );
  buffer buf_n7528( .i (n7527), .o (n7528) );
  assign n7529 = ( n7132 & n7478 ) | ( n7132 & n7525 ) | ( n7478 & n7525 ) ;
  buffer buf_n7530( .i (n7529), .o (n7530) );
  buffer buf_n7531( .i (n7530), .o (n7531) );
  assign n7532 = n7312 & ~n7530 ;
  assign n7533 = ( n7528 & ~n7531 ) | ( n7528 & n7532 ) | ( ~n7531 & n7532 ) ;
  buffer buf_n7534( .i (n7533), .o (n7534) );
  buffer buf_n7535( .i (n7534), .o (n7535) );
  buffer buf_n4379( .i (n4378), .o (n4379) );
  buffer buf_n4380( .i (n4379), .o (n4380) );
  assign n7536 = ( n4380 & n7097 ) | ( n4380 & n7534 ) | ( n7097 & n7534 ) ;
  assign n7537 = n7535 & ~n7536 ;
  buffer buf_n7538( .i (n7537), .o (n7538) );
  buffer buf_n7539( .i (n7538), .o (n7539) );
  buffer buf_n7540( .i (n6994), .o (n7540) );
  assign n7541 = ( n6113 & n7425 ) | ( n6113 & n7540 ) | ( n7425 & n7540 ) ;
  buffer buf_n7542( .i (n7541), .o (n7542) );
  assign n7543 = ( n7045 & n7457 ) | ( n7045 & ~n7542 ) | ( n7457 & ~n7542 ) ;
  assign n7544 = ( ~n7386 & n7457 ) | ( ~n7386 & n7542 ) | ( n7457 & n7542 ) ;
  assign n7545 = ~n7543 & n7544 ;
  buffer buf_n7546( .i (n7200), .o (n7546) );
  assign n7547 = ~n7545 & n7546 ;
  assign n7548 = n4108 & ~n7046 ;
  assign n7549 = n7546 | n7548 ;
  assign n7550 = ~n7547 & n7549 ;
  buffer buf_n7551( .i (n7550), .o (n7551) );
  buffer buf_n7552( .i (n7551), .o (n7552) );
  assign n7553 = ( n6824 & ~n7227 ) | ( n6824 & n7551 ) | ( ~n7227 & n7551 ) ;
  buffer buf_n7554( .i (n7451), .o (n7554) );
  assign n7555 = n277 & ~n7554 ;
  buffer buf_n7556( .i (n7546), .o (n7556) );
  assign n7557 = ( n7392 & n7555 ) | ( n7392 & n7556 ) | ( n7555 & n7556 ) ;
  buffer buf_n7558( .i (n7556), .o (n7558) );
  assign n7559 = n7557 & ~n7558 ;
  buffer buf_n7560( .i (n7226), .o (n7560) );
  assign n7561 = n7559 & n7560 ;
  assign n7562 = ( n7552 & ~n7553 ) | ( n7552 & n7561 ) | ( ~n7553 & n7561 ) ;
  assign n7563 = n278 & n713 ;
  assign n7564 = ( n7182 & n7356 ) | ( n7182 & n7563 ) | ( n7356 & n7563 ) ;
  assign n7565 = ~n6674 & n7564 ;
  buffer buf_n7566( .i (n7565), .o (n7566) );
  assign n7567 = ( ~n7538 & n7562 ) | ( ~n7538 & n7566 ) | ( n7562 & n7566 ) ;
  buffer buf_n7568( .i (n6986), .o (n7568) );
  assign n7569 = ~n7566 & n7568 ;
  assign n7570 = ( n7539 & n7567 ) | ( n7539 & ~n7569 ) | ( n7567 & ~n7569 ) ;
  assign n7571 = n7522 | n7570 ;
  assign n7572 = ( n7403 & ~n7404 ) | ( n7403 & n7571 ) | ( ~n7404 & n7571 ) ;
  assign n7573 = n7380 | n7572 ;
  assign n7574 = ( ~n7234 & n7268 ) | ( ~n7234 & n7573 ) | ( n7268 & n7573 ) ;
  assign n7575 = n7235 | n7574 ;
  buffer buf_n7576( .i (n7575), .o (n7576) );
  buffer buf_n6058( .i (n6057), .o (n6058) );
  buffer buf_n6059( .i (n6058), .o (n6059) );
  buffer buf_n6060( .i (n6059), .o (n6060) );
  buffer buf_n6061( .i (n6060), .o (n6061) );
  buffer buf_n6062( .i (n6061), .o (n6062) );
  buffer buf_n6063( .i (n6062), .o (n6063) );
  buffer buf_n6064( .i (n6063), .o (n6064) );
  buffer buf_n6065( .i (n6064), .o (n6065) );
  buffer buf_n6066( .i (n6065), .o (n6066) );
  buffer buf_n6067( .i (n6066), .o (n6067) );
  buffer buf_n7577( .i (n7365), .o (n7577) );
  buffer buf_n7578( .i (n7577), .o (n7578) );
  assign n7579 = n1974 & ~n7578 ;
  buffer buf_n7580( .i (n7579), .o (n7580) );
  buffer buf_n7581( .i (n7580), .o (n7581) );
  assign n7582 = ( ~n7097 & n7558 ) | ( ~n7097 & n7580 ) | ( n7558 & n7580 ) ;
  assign n7583 = ( n1977 & n7581 ) | ( n1977 & n7582 ) | ( n7581 & n7582 ) ;
  assign n7584 = n7228 & n7583 ;
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n4165( .i (n4164), .o (n4165) );
  buffer buf_n4166( .i (n4165), .o (n4166) );
  buffer buf_n4167( .i (n4166), .o (n4167) );
  buffer buf_n4168( .i (n4167), .o (n4168) );
  buffer buf_n4169( .i (n4168), .o (n4169) );
  buffer buf_n4170( .i (n4169), .o (n4170) );
  buffer buf_n4171( .i (n4170), .o (n4171) );
  buffer buf_n4172( .i (n4171), .o (n4172) );
  assign n7585 = ( n4170 & n7514 ) | ( n4170 & ~n7556 ) | ( n7514 & ~n7556 ) ;
  assign n7586 = ( n7496 & n7558 ) | ( n7496 & ~n7585 ) | ( n7558 & ~n7585 ) ;
  assign n7587 = ( n447 & n4172 ) | ( n447 & ~n7586 ) | ( n4172 & ~n7586 ) ;
  assign n7588 = n7228 | n7587 ;
  buffer buf_n7589( .i (n7228), .o (n7589) );
  assign n7590 = ( n7584 & n7588 ) | ( n7584 & ~n7589 ) | ( n7588 & ~n7589 ) ;
  assign n7591 = n6190 & ~n7590 ;
  buffer buf_n7592( .i (n7578), .o (n7592) );
  assign n7593 = n7323 | n7592 ;
  buffer buf_n7594( .i (n7593), .o (n7594) );
  buffer buf_n7595( .i (n7097), .o (n7595) );
  assign n7596 = ( n7497 & ~n7594 ) | ( n7497 & n7595 ) | ( ~n7594 & n7595 ) ;
  buffer buf_n7597( .i (n7558), .o (n7597) );
  assign n7598 = ( ~n7594 & n7595 ) | ( ~n7594 & n7597 ) | ( n7595 & n7597 ) ;
  assign n7599 = ( n964 & n7596 ) | ( n964 & ~n7598 ) | ( n7596 & ~n7598 ) ;
  assign n7600 = ~n7174 & n7599 ;
  buffer buf_n7601( .i (n6184), .o (n7601) );
  assign n7602 = n7600 | n7601 ;
  assign n7603 = ~n7591 & n7602 ;
  assign n7604 = ( n5847 & ~n6067 ) | ( n5847 & n7603 ) | ( ~n6067 & n7603 ) ;
  buffer buf_n6500( .i (n6499), .o (n6500) );
  buffer buf_n6501( .i (n6500), .o (n6501) );
  buffer buf_n6502( .i (n6501), .o (n6502) );
  buffer buf_n6503( .i (n6502), .o (n6503) );
  assign n7605 = n6503 & n7212 ;
  buffer buf_n7606( .i (n7595), .o (n7606) );
  assign n7607 = ( n6503 & n7212 ) | ( n6503 & ~n7606 ) | ( n7212 & ~n7606 ) ;
  assign n7608 = ( n6242 & ~n7605 ) | ( n6242 & n7607 ) | ( ~n7605 & n7607 ) ;
  assign n7609 = n6435 | n7608 ;
  assign n7610 = n4896 | n7609 ;
  buffer buf_n7611( .i (n7039), .o (n7611) );
  buffer buf_n7612( .i (n7611), .o (n7612) );
  assign n7613 = ( n6067 & n7610 ) | ( n6067 & n7612 ) | ( n7610 & n7612 ) ;
  assign n7614 = n7604 & ~n7613 ;
  buffer buf_n7615( .i (n7614), .o (n7615) );
  buffer buf_n7616( .i (n7615), .o (n7616) );
  buffer buf_n2677( .i (n2676), .o (n2677) );
  buffer buf_n2937( .i (n2936), .o (n2937) );
  buffer buf_n2938( .i (n2937), .o (n2938) );
  assign n7617 = ( n2676 & n2938 ) | ( n2676 & n7560 ) | ( n2938 & n7560 ) ;
  assign n7618 = ~n2677 & n7617 ;
  buffer buf_n7619( .i (n7618), .o (n7619) );
  buffer buf_n7620( .i (n7619), .o (n7620) );
  buffer buf_n5144( .i (n5143), .o (n5144) );
  assign n7621 = n5144 & ~n7595 ;
  buffer buf_n7622( .i (n7560), .o (n7622) );
  assign n7623 = ( n7399 & n7621 ) | ( n7399 & n7622 ) | ( n7621 & n7622 ) ;
  assign n7624 = ~n7589 & n7623 ;
  assign n7625 = n1402 & ~n1510 ;
  assign n7626 = n402 & n7625 ;
  buffer buf_n7627( .i (n7626), .o (n7627) );
  assign n7628 = ( ~n7619 & n7624 ) | ( ~n7619 & n7627 ) | ( n7624 & n7627 ) ;
  buffer buf_n7629( .i (n7568), .o (n7629) );
  assign n7630 = ~n7627 & n7629 ;
  assign n7631 = ( n7620 & n7628 ) | ( n7620 & ~n7630 ) | ( n7628 & ~n7630 ) ;
  buffer buf_n7632( .i (n7631), .o (n7632) );
  buffer buf_n7633( .i (n7632), .o (n7633) );
  assign n7634 = n2710 & n7632 ;
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n5945( .i (n5944), .o (n5945) );
  buffer buf_n5946( .i (n5945), .o (n5946) );
  buffer buf_n5947( .i (n5946), .o (n5947) );
  buffer buf_n5948( .i (n5947), .o (n5948) );
  buffer buf_n5949( .i (n5948), .o (n5949) );
  buffer buf_n5950( .i (n5949), .o (n5950) );
  buffer buf_n5951( .i (n5950), .o (n5951) );
  buffer buf_n5952( .i (n5951), .o (n5952) );
  buffer buf_n5953( .i (n5952), .o (n5953) );
  buffer buf_n5954( .i (n5953), .o (n5954) );
  assign n7635 = ( ~n719 & n808 ) | ( ~n719 & n5954 ) | ( n808 & n5954 ) ;
  assign n7636 = n720 & n7635 ;
  buffer buf_n4122( .i (n4121), .o (n4122) );
  buffer buf_n4123( .i (n4122), .o (n4123) );
  buffer buf_n4124( .i (n4123), .o (n4124) );
  buffer buf_n4125( .i (n4124), .o (n4125) );
  assign n7637 = ( n5929 & n7507 ) | ( n5929 & n7523 ) | ( n7507 & n7523 ) ;
  buffer buf_n7638( .i (n7637), .o (n7638) );
  assign n7639 = ( n7132 & n7456 ) | ( n7132 & ~n7638 ) | ( n7456 & ~n7638 ) ;
  buffer buf_n7640( .i (n7412), .o (n7640) );
  buffer buf_n7641( .i (n7640), .o (n7641) );
  assign n7642 = ( ~n7436 & n7638 ) | ( ~n7436 & n7641 ) | ( n7638 & n7641 ) ;
  assign n7643 = ~n7639 & n7642 ;
  assign n7644 = n7321 | n7643 ;
  assign n7645 = n2177 & n6913 ;
  buffer buf_n7646( .i (n7320), .o (n7646) );
  assign n7647 = ~n7645 & n7646 ;
  assign n7648 = n7644 & ~n7647 ;
  assign n7649 = n7514 & n7648 ;
  buffer buf_n7650( .i (n7649), .o (n7650) );
  buffer buf_n7651( .i (n7650), .o (n7651) );
  buffer buf_n7652( .i (n7386), .o (n7652) );
  buffer buf_n7653( .i (n7652), .o (n7653) );
  buffer buf_n7654( .i (n7653), .o (n7654) );
  assign n7655 = ( n350 & ~n2010 ) | ( n350 & n7654 ) | ( ~n2010 & n7654 ) ;
  assign n7656 = n351 & ~n7655 ;
  assign n7657 = n7650 | n7656 ;
  assign n7658 = ( n7622 & n7651 ) | ( n7622 & n7657 ) | ( n7651 & n7657 ) ;
  assign n7659 = ~n4125 & n7658 ;
  buffer buf_n7660( .i (n7659), .o (n7660) );
  buffer buf_n7661( .i (n7660), .o (n7661) );
  buffer buf_n3267( .i (n3266), .o (n3267) );
  assign n7662 = ~n3264 & n7346 ;
  buffer buf_n7663( .i (n7662), .o (n7663) );
  buffer buf_n7664( .i (n7663), .o (n7664) );
  buffer buf_n7665( .i (n7499), .o (n7665) );
  assign n7666 = ( n7122 & n7663 ) | ( n7122 & ~n7665 ) | ( n7663 & ~n7665 ) ;
  assign n7667 = ( ~n3267 & n7664 ) | ( ~n3267 & n7666 ) | ( n7664 & n7666 ) ;
  assign n7668 = n7031 & n7667 ;
  assign n7669 = ( n1048 & ~n7478 ) | ( n1048 & n7499 ) | ( ~n7478 & n7499 ) ;
  assign n7670 = ( n396 & ~n7365 ) | ( n396 & n7669 ) | ( ~n7365 & n7669 ) ;
  assign n7671 = ( ~n4496 & n7577 ) | ( ~n4496 & n7670 ) | ( n7577 & n7670 ) ;
  assign n7672 = ~n7031 & n7671 ;
  assign n7673 = ( n7493 & ~n7668 ) | ( n7493 & n7672 ) | ( ~n7668 & n7672 ) ;
  buffer buf_n7674( .i (n7556), .o (n7674) );
  assign n7675 = n7673 | n7674 ;
  assign n7676 = n926 & ~n7577 ;
  assign n7677 = n566 & n7676 ;
  assign n7678 = n398 & n1140 ;
  assign n7679 = n7677 | n7678 ;
  assign n7680 = n7674 & n7679 ;
  assign n7681 = n7675 & ~n7680 ;
  assign n7682 = ( ~n5774 & n7622 ) | ( ~n5774 & n7681 ) | ( n7622 & n7681 ) ;
  buffer buf_n1142( .i (n1141), .o (n1142) );
  assign n7683 = n407 & ~n1142 ;
  assign n7684 = ( n1861 & n6993 ) | ( n1861 & n7411 ) | ( n6993 & n7411 ) ;
  buffer buf_n7685( .i (n7684), .o (n7685) );
  buffer buf_n7686( .i (n7685), .o (n7686) );
  buffer buf_n7687( .i (n7686), .o (n7687) );
  assign n7688 = ( n7508 & n7640 ) | ( n7508 & ~n7685 ) | ( n7640 & ~n7685 ) ;
  assign n7689 = n1864 & n7688 ;
  assign n7690 = ( n7665 & ~n7687 ) | ( n7665 & n7689 ) | ( ~n7687 & n7689 ) ;
  buffer buf_n7691( .i (n7690), .o (n7691) );
  buffer buf_n7692( .i (n7691), .o (n7692) );
  assign n7693 = ( n7554 & n7578 ) | ( n7554 & n7691 ) | ( n7578 & n7691 ) ;
  assign n7694 = ( ~n347 & n1081 ) | ( ~n347 & n7665 ) | ( n1081 & n7665 ) ;
  assign n7695 = n348 & n7694 ;
  assign n7696 = ~n7578 & n7695 ;
  assign n7697 = ( n7692 & ~n7693 ) | ( n7692 & n7696 ) | ( ~n7693 & n7696 ) ;
  buffer buf_n7698( .i (n7501), .o (n7698) );
  buffer buf_n7699( .i (n7698), .o (n7699) );
  assign n7700 = ~n426 & n7699 ;
  buffer buf_n7701( .i (n7700), .o (n7701) );
  assign n7702 = n1306 & n7701 ;
  assign n7703 = ( n289 & ~n428 ) | ( n289 & n7701 ) | ( ~n428 & n7701 ) ;
  assign n7704 = ( n7392 & n7702 ) | ( n7392 & n7703 ) | ( n7702 & n7703 ) ;
  assign n7705 = n7697 | n7704 ;
  assign n7706 = ( n408 & ~n7683 ) | ( n408 & n7705 ) | ( ~n7683 & n7705 ) ;
  assign n7707 = ( n5774 & n7622 ) | ( n5774 & n7706 ) | ( n7622 & n7706 ) ;
  assign n7708 = ~n7682 & n7707 ;
  assign n7709 = ~n1135 & n7322 ;
  buffer buf_n7710( .i (n7646), .o (n7710) );
  assign n7711 = n1546 | n7710 ;
  assign n7712 = ~n7709 & n7711 ;
  buffer buf_n7713( .i (n7514), .o (n7713) );
  assign n7714 = ~n7712 & n7713 ;
  assign n7715 = ( n1170 & n7446 ) | ( n1170 & n7499 ) | ( n7446 & n7499 ) ;
  buffer buf_n7716( .i (n7715), .o (n7716) );
  buffer buf_n7717( .i (n7716), .o (n7717) );
  assign n7718 = n1165 & ~n7716 ;
  assign n7719 = ( n1173 & ~n7717 ) | ( n1173 & n7718 ) | ( ~n7717 & n7718 ) ;
  assign n7720 = ~n7323 & n7719 ;
  assign n7721 = n7713 | n7720 ;
  assign n7722 = ~n7714 & n7721 ;
  buffer buf_n7723( .i (n6674), .o (n7723) );
  assign n7724 = ( n7399 & n7722 ) | ( n7399 & ~n7723 ) | ( n7722 & ~n7723 ) ;
  assign n7725 = ( n2069 & n6780 ) | ( n2069 & ~n7411 ) | ( n6780 & ~n7411 ) ;
  buffer buf_n7726( .i (n7725), .o (n7726) );
  buffer buf_n7729( .i (n6780), .o (n7729) );
  buffer buf_n7730( .i (n7729), .o (n7730) );
  assign n7731 = ~n7726 & n7730 ;
  buffer buf_n7732( .i (n7731), .o (n7732) );
  buffer buf_n7733( .i (n7732), .o (n7733) );
  buffer buf_n7727( .i (n7726), .o (n7727) );
  buffer buf_n7728( .i (n7727), .o (n7728) );
  assign n7734 = n7728 | n7732 ;
  assign n7735 = ( ~n7451 & n7733 ) | ( ~n7451 & n7734 ) | ( n7733 & n7734 ) ;
  assign n7736 = n7710 & ~n7735 ;
  assign n7737 = n1211 & ~n7451 ;
  assign n7738 = n7710 | n7737 ;
  assign n7739 = ~n7736 & n7738 ;
  buffer buf_n7740( .i (n7450), .o (n7740) );
  buffer buf_n7741( .i (n7740), .o (n7741) );
  assign n7742 = n7739 | n7741 ;
  buffer buf_n6849( .i (n6848), .o (n6849) );
  buffer buf_n6850( .i (n6849), .o (n6850) );
  buffer buf_n6851( .i (n6850), .o (n6851) );
  buffer buf_n6852( .i (n6851), .o (n6852) );
  buffer buf_n6853( .i (n6852), .o (n6853) );
  buffer buf_n7743( .i (n7122), .o (n7743) );
  assign n7744 = ( n7007 & ~n7646 ) | ( n7007 & n7743 ) | ( ~n7646 & n7743 ) ;
  assign n7745 = n6853 & n7744 ;
  assign n7746 = ~n7592 & n7745 ;
  assign n7747 = n7741 & ~n7746 ;
  assign n7748 = n7742 & ~n7747 ;
  assign n7749 = ( n7399 & n7723 ) | ( n7399 & ~n7748 ) | ( n7723 & ~n7748 ) ;
  assign n7750 = n7724 & ~n7749 ;
  assign n7751 = ( ~n7629 & n7708 ) | ( ~n7629 & n7750 ) | ( n7708 & n7750 ) ;
  assign n7752 = ~n7660 & n7751 ;
  assign n7753 = ( ~n7612 & n7661 ) | ( ~n7612 & n7752 ) | ( n7661 & n7752 ) ;
  assign n7754 = n7636 | n7753 ;
  assign n7755 = ( n7633 & ~n7634 ) | ( n7633 & n7754 ) | ( ~n7634 & n7754 ) ;
  buffer buf_n4069( .i (n4068), .o (n4069) );
  buffer buf_n7756( .i (n7710), .o (n7756) );
  assign n7757 = ( ~n589 & n4069 ) | ( ~n589 & n7756 ) | ( n4069 & n7756 ) ;
  assign n7758 = ~n7226 & n7757 ;
  buffer buf_n7759( .i (n7758), .o (n7759) );
  buffer buf_n7760( .i (n7759), .o (n7760) );
  buffer buf_n7761( .i (n7760), .o (n7761) );
  buffer buf_n5078( .i (n5077), .o (n5078) );
  buffer buf_n5079( .i (n5078), .o (n5079) );
  buffer buf_n5080( .i (n5079), .o (n5080) );
  assign n7762 = ( n5080 & n7496 ) | ( n5080 & ~n7741 ) | ( n7496 & ~n7741 ) ;
  assign n7763 = ( n5079 & ~n7592 ) | ( n5079 & n7756 ) | ( ~n7592 & n7756 ) ;
  assign n7764 = ( ~n7182 & n7741 ) | ( ~n7182 & n7763 ) | ( n7741 & n7763 ) ;
  assign n7765 = n7762 | n7764 ;
  buffer buf_n7766( .i (n7597), .o (n7766) );
  assign n7767 = ( n7759 & ~n7765 ) | ( n7759 & n7766 ) | ( ~n7765 & n7766 ) ;
  assign n7768 = n7174 & ~n7767 ;
  assign n7769 = ( n7078 & n7761 ) | ( n7078 & ~n7768 ) | ( n7761 & ~n7768 ) ;
  buffer buf_n7770( .i (n7769), .o (n7770) );
  buffer buf_n7771( .i (n7770), .o (n7771) );
  assign n7772 = ( n357 & n7612 ) | ( n357 & n7770 ) | ( n7612 & n7770 ) ;
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  assign n7773 = ( n1411 & n6188 ) | ( n1411 & n7149 ) | ( n6188 & n7149 ) ;
  assign n7774 = ~n7150 & n7773 ;
  assign n7775 = ~n357 & n7774 ;
  assign n7776 = ( n7771 & ~n7772 ) | ( n7771 & n7775 ) | ( ~n7772 & n7775 ) ;
  assign n7777 = ( ~n6780 & n7411 ) | ( ~n6780 & n7506 ) | ( n7411 & n7506 ) ;
  buffer buf_n7778( .i (n7777), .o (n7778) );
  assign n7783 = ( n3914 & n7640 ) | ( n3914 & ~n7778 ) | ( n7640 & ~n7778 ) ;
  buffer buf_n7784( .i (n7783), .o (n7784) );
  buffer buf_n7785( .i (n7784), .o (n7785) );
  buffer buf_n7786( .i (n7785), .o (n7786) );
  buffer buf_n7787( .i (n7786), .o (n7787) );
  buffer buf_n7788( .i (n7730), .o (n7788) );
  buffer buf_n7789( .i (n7788), .o (n7789) );
  assign n7790 = ( ~n7454 & n7784 ) | ( ~n7454 & n7789 ) | ( n7784 & n7789 ) ;
  buffer buf_n7791( .i (n7790), .o (n7791) );
  buffer buf_n7792( .i (n7791), .o (n7792) );
  buffer buf_n7779( .i (n7778), .o (n7779) );
  buffer buf_n7780( .i (n7779), .o (n7780) );
  buffer buf_n7781( .i (n7780), .o (n7781) );
  buffer buf_n7782( .i (n7781), .o (n7782) );
  assign n7793 = n7782 & n7791 ;
  assign n7794 = ( ~n7787 & n7792 ) | ( ~n7787 & n7793 ) | ( n7792 & n7793 ) ;
  assign n7795 = n7226 | n7794 ;
  assign n7796 = ~n1332 & n7743 ;
  buffer buf_n7797( .i (n7030), .o (n7797) );
  assign n7798 = ( ~n1333 & n7796 ) | ( ~n1333 & n7797 ) | ( n7796 & n7797 ) ;
  assign n7799 = ~n6567 & n7798 ;
  buffer buf_n7800( .i (n7756), .o (n7800) );
  assign n7801 = ~n7799 & n7800 ;
  assign n7802 = n7795 & ~n7801 ;
  assign n7803 = n7766 | n7802 ;
  buffer buf_n7804( .i (n7554), .o (n7804) );
  assign n7805 = ( ~n7009 & n7493 ) | ( ~n7009 & n7804 ) | ( n7493 & n7804 ) ;
  assign n7806 = ( n7009 & n7493 ) | ( n7009 & ~n7756 ) | ( n7493 & ~n7756 ) ;
  assign n7807 = n7805 | n7806 ;
  assign n7808 = n7397 | n7807 ;
  assign n7809 = n7766 & n7808 ;
  assign n7810 = n7803 & ~n7809 ;
  assign n7811 = n6178 | n7810 ;
  assign n7812 = ( ~n3950 & n7454 ) | ( ~n3950 & n7789 ) | ( n7454 & n7789 ) ;
  buffer buf_n7813( .i (n7812), .o (n7813) );
  buffer buf_n7814( .i (n7813), .o (n7814) );
  buffer buf_n7815( .i (n7814), .o (n7815) );
  buffer buf_n7816( .i (n7815), .o (n7816) );
  buffer buf_n7817( .i (n7646), .o (n7817) );
  assign n7818 = ( n7546 & ~n7813 ) | ( n7546 & n7817 ) | ( ~n7813 & n7817 ) ;
  buffer buf_n7819( .i (n7818), .o (n7819) );
  buffer buf_n7820( .i (n7819), .o (n7820) );
  assign n7821 = ~n3954 & n7819 ;
  assign n7822 = ( n7816 & n7820 ) | ( n7816 & n7821 ) | ( n7820 & n7821 ) ;
  assign n7823 = n927 & n7554 ;
  buffer buf_n7824( .i (n310), .o (n7824) );
  assign n7825 = n7823 & ~n7824 ;
  buffer buf_n7826( .i (n7825), .o (n7826) );
  buffer buf_n7827( .i (n7826), .o (n7827) );
  assign n7828 = n6763 & ~n7826 ;
  assign n7829 = ( n7822 & n7827 ) | ( n7822 & ~n7828 ) | ( n7827 & ~n7828 ) ;
  assign n7830 = ~n7568 & n7829 ;
  assign n7831 = n6178 & ~n7830 ;
  assign n7832 = n7811 & ~n7831 ;
  assign n7833 = n7151 & n7832 ;
  assign n7834 = ~n341 & n572 ;
  buffer buf_n7835( .i (n6752), .o (n7835) );
  assign n7836 = ( n3914 & ~n7730 ) | ( n3914 & n7835 ) | ( ~n7730 & n7835 ) ;
  buffer buf_n7837( .i (n7836), .o (n7837) );
  buffer buf_n7838( .i (n7837), .o (n7838) );
  buffer buf_n7839( .i (n7838), .o (n7839) );
  buffer buf_n7840( .i (n7839), .o (n7840) );
  assign n7841 = n6896 & ~n7837 ;
  buffer buf_n7842( .i (n7841), .o (n7842) );
  buffer buf_n7843( .i (n7842), .o (n7843) );
  assign n7844 = ( ~n7008 & n7817 ) | ( ~n7008 & n7842 ) | ( n7817 & n7842 ) ;
  assign n7845 = ( ~n7840 & n7843 ) | ( ~n7840 & n7844 ) | ( n7843 & n7844 ) ;
  buffer buf_n7846( .i (n7740), .o (n7846) );
  assign n7847 = ( n7209 & n7845 ) | ( n7209 & n7846 ) | ( n7845 & n7846 ) ;
  buffer buf_n7848( .i (n7743), .o (n7848) );
  assign n7849 = ( n729 & n4480 ) | ( n729 & n7848 ) | ( n4480 & n7848 ) ;
  assign n7850 = ~n7804 & n7849 ;
  assign n7851 = n7209 & n7850 ;
  buffer buf_n7852( .i (n7846), .o (n7852) );
  assign n7853 = ( n7847 & n7851 ) | ( n7847 & ~n7852 ) | ( n7851 & ~n7852 ) ;
  assign n7854 = ~n7766 & n7853 ;
  buffer buf_n7855( .i (n7854), .o (n7855) );
  buffer buf_n7856( .i (n7855), .o (n7856) );
  assign n7857 = n759 | n7855 ;
  assign n7858 = ( n7834 & n7856 ) | ( n7834 & n7857 ) | ( n7856 & n7857 ) ;
  assign n7859 = n7151 | n7858 ;
  assign n7860 = ( ~n209 & n7833 ) | ( ~n209 & n7859 ) | ( n7833 & n7859 ) ;
  assign n7861 = n7776 | n7860 ;
  assign n7862 = ( ~n7615 & n7755 ) | ( ~n7615 & n7861 ) | ( n7755 & n7861 ) ;
  assign n7863 = n7616 | n7862 ;
  assign n7864 = n7258 & ~n7674 ;
  buffer buf_n7865( .i (n6897), .o (n7865) );
  buffer buf_n7866( .i (n7865), .o (n7866) );
  buffer buf_n7867( .i (n7866), .o (n7867) );
  assign n7868 = ( n4847 & n7674 ) | ( n4847 & ~n7867 ) | ( n7674 & ~n7867 ) ;
  assign n7869 = n4847 & n7800 ;
  assign n7870 = ( n7864 & n7868 ) | ( n7864 & ~n7869 ) | ( n7868 & ~n7869 ) ;
  assign n7871 = ~n4721 & n7870 ;
  buffer buf_n7872( .i (n7871), .o (n7872) );
  buffer buf_n7873( .i (n7872), .o (n7873) );
  buffer buf_n3704( .i (n3703), .o (n3704) );
  buffer buf_n3705( .i (n3704), .o (n3705) );
  buffer buf_n3706( .i (n3705), .o (n3706) );
  buffer buf_n3707( .i (n3706), .o (n3707) );
  buffer buf_n3708( .i (n3707), .o (n3708) );
  buffer buf_n3709( .i (n3708), .o (n3709) );
  buffer buf_n3710( .i (n3709), .o (n3710) );
  buffer buf_n3711( .i (n3710), .o (n3711) );
  buffer buf_n4848( .i (n4847), .o (n4848) );
  buffer buf_n4849( .i (n4848), .o (n4849) );
  buffer buf_n4850( .i (n4849), .o (n4850) );
  assign n7874 = n3711 & n4850 ;
  assign n7875 = n7872 | n7874 ;
  assign n7876 = ( ~n7611 & n7873 ) | ( ~n7611 & n7875 ) | ( n7873 & n7875 ) ;
  assign n7877 = n7219 | n7876 ;
  buffer buf_n3712( .i (n3711), .o (n3712) );
  assign n7878 = n3709 & ~n6763 ;
  buffer buf_n7879( .i (n7878), .o (n7879) );
  buffer buf_n7880( .i (n7879), .o (n7880) );
  buffer buf_n7881( .i (n7597), .o (n7881) );
  buffer buf_n7882( .i (n7881), .o (n7882) );
  assign n7883 = ( n7589 & n7879 ) | ( n7589 & ~n7882 ) | ( n7879 & ~n7882 ) ;
  assign n7884 = ( n3712 & n7880 ) | ( n3712 & n7883 ) | ( n7880 & n7883 ) ;
  assign n7885 = ~n7611 & n7884 ;
  assign n7886 = n7219 & ~n7885 ;
  assign n7887 = n7877 & ~n7886 ;
  buffer buf_n7888( .i (n7887), .o (n7888) );
  buffer buf_n7889( .i (n7888), .o (n7889) );
  buffer buf_n2678( .i (n2677), .o (n2678) );
  buffer buf_n2679( .i (n2678), .o (n2679) );
  buffer buf_n2680( .i (n2679), .o (n2680) );
  buffer buf_n2681( .i (n2680), .o (n2681) );
  buffer buf_n2682( .i (n2681), .o (n2682) );
  buffer buf_n2683( .i (n2682), .o (n2683) );
  buffer buf_n2684( .i (n2683), .o (n2684) );
  assign n7890 = n2684 & n7888 ;
  buffer buf_n4275( .i (n4274), .o (n4275) );
  buffer buf_n4276( .i (n4275), .o (n4276) );
  buffer buf_n4277( .i (n4276), .o (n4277) );
  buffer buf_n4278( .i (n4277), .o (n4278) );
  buffer buf_n4279( .i (n4278), .o (n4279) );
  buffer buf_n4280( .i (n4279), .o (n4280) );
  buffer buf_n4281( .i (n4280), .o (n4281) );
  buffer buf_n4282( .i (n4281), .o (n4282) );
  buffer buf_n4283( .i (n4282), .o (n4283) );
  buffer buf_n4284( .i (n4283), .o (n4284) );
  buffer buf_n5804( .i (n5803), .o (n5804) );
  buffer buf_n5805( .i (n5804), .o (n5805) );
  buffer buf_n5806( .i (n5805), .o (n5806) );
  buffer buf_n7891( .i (n7457), .o (n7891) );
  buffer buf_n7892( .i (n7891), .o (n7892) );
  buffer buf_n7893( .i (n7892), .o (n7893) );
  buffer buf_n7894( .i (n7893), .o (n7894) );
  assign n7895 = ( n4284 & ~n5806 ) | ( n4284 & n7894 ) | ( ~n5806 & n7894 ) ;
  assign n7896 = n7597 & ~n7895 ;
  buffer buf_n7341( .i (n7340), .o (n7341) );
  buffer buf_n7342( .i (n7341), .o (n7342) );
  buffer buf_n7343( .i (n7342), .o (n7343) );
  buffer buf_n7344( .i (n7343), .o (n7344) );
  buffer buf_n7345( .i (n7344), .o (n7345) );
  assign n7897 = ~n7345 & n7740 ;
  assign n7898 = n7049 & ~n7897 ;
  buffer buf_n7899( .i (n7200), .o (n7899) );
  buffer buf_n7900( .i (n7899), .o (n7900) );
  buffer buf_n7901( .i (n7900), .o (n7901) );
  buffer buf_n7902( .i (n7901), .o (n7902) );
  assign n7903 = n7898 | n7902 ;
  assign n7904 = ( ~n7881 & n7896 ) | ( ~n7881 & n7903 ) | ( n7896 & n7903 ) ;
  assign n7905 = n7568 | n7904 ;
  buffer buf_n7906( .i (n7560), .o (n7906) );
  assign n7907 = n592 | n7906 ;
  buffer buf_n7908( .i (n6986), .o (n7908) );
  assign n7909 = n7907 & n7908 ;
  assign n7910 = n7905 & ~n7909 ;
  assign n7911 = ( n237 & n6189 ) | ( n237 & n7910 ) | ( n6189 & n7910 ) ;
  buffer buf_n7912( .i (n7911), .o (n7912) );
  assign n7913 = ( n151 & ~n7043 ) | ( n151 & n7912 ) | ( ~n7043 & n7912 ) ;
  buffer buf_n7914( .i (n150), .o (n7914) );
  assign n7915 = ( n239 & ~n7912 ) | ( n239 & n7914 ) | ( ~n7912 & n7914 ) ;
  assign n7916 = n7913 & ~n7915 ;
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  assign n7917 = n934 & ~n7150 ;
  assign n7918 = n602 & n7917 ;
  assign n7919 = n721 & ~n7918 ;
  buffer buf_n7920( .i (n6751), .o (n7920) );
  assign n7921 = ( n1000 & n7523 ) | ( n1000 & n7920 ) | ( n7523 & n7920 ) ;
  buffer buf_n7922( .i (n7921), .o (n7922) );
  buffer buf_n7923( .i (n7922), .o (n7923) );
  buffer buf_n7924( .i (n7923), .o (n7924) );
  buffer buf_n7925( .i (n7508), .o (n7925) );
  assign n7926 = ( n7426 & ~n7922 ) | ( n7426 & n7925 ) | ( ~n7922 & n7925 ) ;
  buffer buf_n7927( .i (n7446), .o (n7927) );
  assign n7928 = ( n7320 & n7926 ) | ( n7320 & ~n7927 ) | ( n7926 & ~n7927 ) ;
  assign n7929 = ~n7924 & n7928 ;
  assign n7930 = n7450 | n7929 ;
  buffer buf_n7931( .i (n7320), .o (n7931) );
  assign n7932 = n2056 & n7931 ;
  buffer buf_n7933( .i (n7046), .o (n7933) );
  assign n7934 = ~n7932 & n7933 ;
  assign n7935 = n7930 & ~n7934 ;
  assign n7936 = n7901 & n7935 ;
  buffer buf_n7937( .i (n7540), .o (n7937) );
  assign n7938 = ( n1002 & n7426 ) | ( n1002 & n7937 ) | ( n7426 & n7937 ) ;
  buffer buf_n7939( .i (n7523), .o (n7939) );
  assign n7940 = ( n1001 & n7346 ) | ( n1001 & ~n7939 ) | ( n7346 & ~n7939 ) ;
  assign n7941 = ( n7925 & n7937 ) | ( n7925 & ~n7940 ) | ( n7937 & ~n7940 ) ;
  assign n7942 = ~n7938 & n7941 ;
  assign n7943 = n7931 | n7942 ;
  assign n7944 = n2834 & ~n7665 ;
  assign n7945 = n7931 & ~n7944 ;
  assign n7946 = n7943 & ~n7945 ;
  buffer buf_n7947( .i (n7937), .o (n7947) );
  buffer buf_n7948( .i (n7947), .o (n7948) );
  buffer buf_n7949( .i (n2120), .o (n7949) );
  assign n7950 = ( n7931 & ~n7948 ) | ( n7931 & n7949 ) | ( ~n7948 & n7949 ) ;
  buffer buf_n7951( .i (n7939), .o (n7951) );
  buffer buf_n7952( .i (n7951), .o (n7952) );
  assign n7953 = ( n2120 & n7947 ) | ( n2120 & ~n7952 ) | ( n7947 & ~n7952 ) ;
  buffer buf_n7954( .i (n7319), .o (n7954) );
  buffer buf_n7955( .i (n7954), .o (n7955) );
  assign n7956 = ( n7030 & ~n7953 ) | ( n7030 & n7955 ) | ( ~n7953 & n7955 ) ;
  assign n7957 = ~n7950 & n7956 ;
  assign n7958 = n7946 | n7957 ;
  assign n7959 = ~n7901 & n7958 ;
  assign n7960 = n7936 | n7959 ;
  assign n7961 = ~n7212 & n7960 ;
  assign n7962 = n5410 & ~n7454 ;
  assign n7963 = ( ~n5409 & n7319 ) | ( ~n5409 & n7698 ) | ( n7319 & n7698 ) ;
  buffer buf_n7964( .i (n7925), .o (n7964) );
  assign n7965 = ( n744 & ~n7963 ) | ( n744 & n7964 ) | ( ~n7963 & n7964 ) ;
  buffer buf_n7966( .i (n7964), .o (n7966) );
  assign n7967 = ( n7962 & ~n7965 ) | ( n7962 & n7966 ) | ( ~n7965 & n7966 ) ;
  buffer buf_n7968( .i (n7967), .o (n7968) );
  buffer buf_n7969( .i (n7968), .o (n7969) );
  assign n7970 = ( n7654 & n7740 ) | ( n7654 & n7968 ) | ( n7740 & n7968 ) ;
  assign n7971 = ( ~n745 & n4880 ) | ( ~n745 & n7577 ) | ( n4880 & n7577 ) ;
  assign n7972 = n746 & n7971 ;
  assign n7973 = ~n7654 & n7972 ;
  assign n7974 = ( n7969 & ~n7970 ) | ( n7969 & n7973 ) | ( ~n7970 & n7973 ) ;
  buffer buf_n7975( .i (n5881), .o (n7975) );
  assign n7976 = ( ~n3733 & n6363 ) | ( ~n3733 & n7975 ) | ( n6363 & n7975 ) ;
  buffer buf_n7977( .i (n7976), .o (n7977) );
  assign n7982 = ( n6993 & ~n7506 ) | ( n6993 & n7977 ) | ( ~n7506 & n7977 ) ;
  buffer buf_n7983( .i (n7982), .o (n7983) );
  buffer buf_n7984( .i (n7983), .o (n7984) );
  buffer buf_n7985( .i (n7984), .o (n7985) );
  buffer buf_n7986( .i (n7985), .o (n7986) );
  assign n7987 = ( ~n7501 & n7835 ) | ( ~n7501 & n7983 ) | ( n7835 & n7983 ) ;
  buffer buf_n7988( .i (n7987), .o (n7988) );
  buffer buf_n7989( .i (n7988), .o (n7989) );
  buffer buf_n7978( .i (n7977), .o (n7978) );
  buffer buf_n7979( .i (n7978), .o (n7979) );
  buffer buf_n7980( .i (n7979), .o (n7980) );
  buffer buf_n7981( .i (n7980), .o (n7981) );
  assign n7990 = ~n7981 & n7988 ;
  assign n7991 = ( ~n7986 & n7989 ) | ( ~n7986 & n7990 ) | ( n7989 & n7990 ) ;
  buffer buf_n7992( .i (n7991), .o (n7992) );
  buffer buf_n7993( .i (n7992), .o (n7993) );
  assign n7994 = ( n7592 & n7654 ) | ( n7592 & ~n7992 ) | ( n7654 & ~n7992 ) ;
  assign n7995 = ( n5924 & ~n6734 ) | ( n5924 & n6901 ) | ( ~n6734 & n6901 ) ;
  buffer buf_n7996( .i (n7995), .o (n7996) );
  assign n8001 = ( ~n7246 & n7507 ) | ( ~n7246 & n7996 ) | ( n7507 & n7996 ) ;
  buffer buf_n8002( .i (n8001), .o (n8002) );
  buffer buf_n8003( .i (n8002), .o (n8003) );
  buffer buf_n8004( .i (n8003), .o (n8004) );
  buffer buf_n8005( .i (n8004), .o (n8005) );
  assign n8006 = ( n7698 & ~n7937 ) | ( n7698 & n8002 ) | ( ~n7937 & n8002 ) ;
  buffer buf_n8007( .i (n8006), .o (n8007) );
  buffer buf_n8008( .i (n8007), .o (n8008) );
  buffer buf_n7997( .i (n7996), .o (n7997) );
  buffer buf_n7998( .i (n7997), .o (n7998) );
  buffer buf_n7999( .i (n7998), .o (n7999) );
  buffer buf_n8000( .i (n7999), .o (n8000) );
  assign n8009 = ~n8000 & n8007 ;
  assign n8010 = ( ~n8005 & n8008 ) | ( ~n8005 & n8009 ) | ( n8008 & n8009 ) ;
  buffer buf_n8011( .i (n7653), .o (n8011) );
  assign n8012 = n8010 & n8011 ;
  assign n8013 = ( n7993 & n7994 ) | ( n7993 & n8012 ) | ( n7994 & n8012 ) ;
  assign n8014 = n7974 | n8013 ;
  buffer buf_n8015( .i (n7713), .o (n8015) );
  buffer buf_n8016( .i (n8015), .o (n8016) );
  assign n8017 = n8014 & n8016 ;
  assign n8018 = n7961 | n8017 ;
  buffer buf_n8019( .i (n8018), .o (n8019) );
  buffer buf_n8020( .i (n8019), .o (n8020) );
  assign n8021 = ( ~n6191 & n7611 ) | ( ~n6191 & n8019 ) | ( n7611 & n8019 ) ;
  assign n8022 = n314 | n2202 ;
  assign n8023 = ( n282 & n694 ) | ( n282 & n8022 ) | ( n694 & n8022 ) ;
  assign n8024 = n283 & ~n8023 ;
  buffer buf_n8025( .i (n7629), .o (n8025) );
  assign n8026 = n8024 & ~n8025 ;
  assign n8027 = ( n8020 & ~n8021 ) | ( n8020 & n8026 ) | ( ~n8021 & n8026 ) ;
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  assign n8028 = ( ~n745 & n4225 ) | ( ~n745 & n7743 ) | ( n4225 & n7743 ) ;
  assign n8029 = n746 & n8028 ;
  assign n8030 = ~n7893 & n8029 ;
  buffer buf_n8031( .i (n8030), .o (n8031) );
  buffer buf_n8032( .i (n8031), .o (n8032) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  assign n8033 = ( n7319 & n7698 ) | ( n7319 & ~n7951 ) | ( n7698 & ~n7951 ) ;
  buffer buf_n8034( .i (n8033), .o (n8034) );
  buffer buf_n8035( .i (n8034), .o (n8035) );
  buffer buf_n8036( .i (n8035), .o (n8036) );
  assign n8037 = ( ~n7200 & n7652 ) | ( ~n7200 & n8034 ) | ( n7652 & n8034 ) ;
  assign n8038 = ( n7848 & n7899 ) | ( n7848 & ~n8037 ) | ( n7899 & ~n8037 ) ;
  assign n8039 = ( n1496 & n8036 ) | ( n1496 & ~n8038 ) | ( n8036 & ~n8038 ) ;
  buffer buf_n8040( .i (n8039), .o (n8040) );
  buffer buf_n8041( .i (n8040), .o (n8041) );
  buffer buf_n8042( .i (n7894), .o (n8042) );
  assign n8043 = ( n7852 & n8040 ) | ( n7852 & n8042 ) | ( n8040 & n8042 ) ;
  assign n8044 = ( n8032 & n8041 ) | ( n8032 & ~n8043 ) | ( n8041 & ~n8043 ) ;
  assign n8045 = ~n7214 & n8044 ;
  buffer buf_n8046( .i (n7789), .o (n8046) );
  assign n8047 = n4281 & n8046 ;
  assign n8048 = ( n4225 & ~n7955 ) | ( n4225 & n8046 ) | ( ~n7955 & n8046 ) ;
  assign n8049 = ~n4225 & n7955 ;
  assign n8050 = ( ~n8047 & n8048 ) | ( ~n8047 & n8049 ) | ( n8048 & n8049 ) ;
  buffer buf_n8051( .i (n8050), .o (n8051) );
  buffer buf_n8052( .i (n8051), .o (n8052) );
  assign n8053 = ( n7894 & n7901 ) | ( n7894 & ~n8051 ) | ( n7901 & ~n8051 ) ;
  assign n8054 = ( ~n8031 & n8052 ) | ( ~n8031 & n8053 ) | ( n8052 & n8053 ) ;
  assign n8055 = ( n1384 & n2610 ) | ( n1384 & ~n6110 ) | ( n2610 & ~n6110 ) ;
  assign n8056 = ( n7817 & n7848 ) | ( n7817 & ~n8055 ) | ( n7848 & ~n8055 ) ;
  buffer buf_n8057( .i (n8056), .o (n8057) );
  assign n8058 = ( ~n7713 & n7846 ) | ( ~n7713 & n8057 ) | ( n7846 & n8057 ) ;
  assign n8059 = ( n7800 & n7846 ) | ( n7800 & ~n8057 ) | ( n7846 & ~n8057 ) ;
  assign n8060 = n8058 & ~n8059 ;
  assign n8061 = n8054 & ~n8060 ;
  buffer buf_n8062( .i (n6480), .o (n8062) );
  assign n8063 = ~n8061 & n8062 ;
  assign n8064 = n8045 | n8063 ;
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n2158( .i (n2157), .o (n2158) );
  buffer buf_n8065( .i (n8011), .o (n8065) );
  assign n8066 = n7800 | n8065 ;
  assign n8067 = ( n597 & n2158 ) | ( n597 & n8066 ) | ( n2158 & n8066 ) ;
  assign n8068 = ( n598 & ~n8016 ) | ( n598 & n8067 ) | ( ~n8016 & n8067 ) ;
  buffer buf_n4422( .i (n4421), .o (n4422) );
  assign n8069 = n4422 & ~n7804 ;
  buffer buf_n8070( .i (n7817), .o (n8070) );
  buffer buf_n8071( .i (n8070), .o (n8071) );
  assign n8072 = n8069 & n8071 ;
  buffer buf_n8073( .i (n8072), .o (n8073) );
  buffer buf_n8074( .i (n8073), .o (n8074) );
  buffer buf_n8075( .i (n8042), .o (n8075) );
  assign n8076 = n8073 | n8075 ;
  assign n8077 = ( n8068 & n8074 ) | ( n8068 & n8076 ) | ( n8074 & n8076 ) ;
  buffer buf_n8078( .i (n6242), .o (n8078) );
  assign n8079 = ( n4895 & n8077 ) | ( n4895 & n8078 ) | ( n8077 & n8078 ) ;
  assign n8080 = ( ~n435 & n8064 ) | ( ~n435 & n8079 ) | ( n8064 & n8079 ) ;
  assign n8081 = ( n7501 & n7835 ) | ( n7501 & n7939 ) | ( n7835 & n7939 ) ;
  buffer buf_n8082( .i (n8081), .o (n8082) );
  assign n8083 = ( n7947 & n7954 ) | ( n7947 & ~n8082 ) | ( n7954 & ~n8082 ) ;
  assign n8084 = ( ~n7699 & n7947 ) | ( ~n7699 & n8082 ) | ( n7947 & n8082 ) ;
  assign n8085 = ~n8083 & n8084 ;
  assign n8086 = n7865 | n8085 ;
  buffer buf_n8087( .i (n7540), .o (n8087) );
  buffer buf_n8088( .i (n8087), .o (n8088) );
  assign n8089 = n3866 | n8088 ;
  assign n8090 = n7955 | n8089 ;
  assign n8091 = n7865 & n8090 ;
  assign n8092 = n8086 & ~n8091 ;
  buffer buf_n8093( .i (n7804), .o (n8093) );
  assign n8094 = ( n7894 & n8092 ) | ( n7894 & n8093 ) | ( n8092 & n8093 ) ;
  buffer buf_n8095( .i (n8094), .o (n8095) );
  buffer buf_n8096( .i (n7497), .o (n8096) );
  assign n8097 = ( ~n8075 & n8095 ) | ( ~n8075 & n8096 ) | ( n8095 & n8096 ) ;
  assign n8098 = ( n8016 & ~n8095 ) | ( n8016 & n8096 ) | ( ~n8095 & n8096 ) ;
  assign n8099 = n8097 & ~n8098 ;
  buffer buf_n8100( .i (n8099), .o (n8100) );
  buffer buf_n8101( .i (n8100), .o (n8101) );
  assign n8102 = n8025 & ~n8100 ;
  assign n8103 = ( n8080 & n8101 ) | ( n8080 & ~n8102 ) | ( n8101 & ~n8102 ) ;
  assign n8104 = n8027 | n8103 ;
  assign n8105 = ( n722 & ~n7919 ) | ( n722 & n8104 ) | ( ~n7919 & n8104 ) ;
  assign n8106 = n7916 | n8105 ;
  assign n8107 = ( n7889 & ~n7890 ) | ( n7889 & n8106 ) | ( ~n7890 & n8106 ) ;
  assign y0 = n421 ;
  assign y1 = n767 ;
  assign y2 = n1099 ;
  assign y3 = n1422 ;
  assign y4 = n1960 ;
  assign y5 = n2625 ;
  assign y6 = n3116 ;
  assign y7 = n3493 ;
  assign y8 = n3862 ;
  assign y9 = n4367 ;
  assign y10 = n4799 ;
  assign y11 = n5162 ;
  assign y12 = n5561 ;
  assign y13 = n5852 ;
  assign y14 = n6214 ;
  assign y15 = n6535 ;
  assign y16 = n6885 ;
  assign y17 = n7224 ;
  assign y18 = n7576 ;
  assign y19 = n7863 ;
  assign y20 = n8107 ;
endmodule
