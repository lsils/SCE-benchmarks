module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G6 , G7 , G8 , G9 , G3519 , G3520 , G3521 , G3522 , G3523 , G3524 , G3525 , G3526 , G3527 , G3528 , G3529 , G3530 , G3531 , G3532 , G3533 , G3534 , G3535 , G3536 , G3537 , G3538 , G3539 , G3540 );
  input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G6 , G7 , G8 , G9 ;
  output G3519 , G3520 , G3521 , G3522 , G3523 , G3524 , G3525 , G3526 , G3527 , G3528 , G3529 , G3530 , G3531 , G3532 , G3533 , G3534 , G3535 , G3536 , G3537 , G3538 , G3539 , G3540 ;
  wire n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 ;
  assign n51 = G8 | G9 ;
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  assign n77 = G10 | G7 ;
  buffer buf_n78( .i (n77), .o (n78) );
  assign n79 = n76 | n78 ;
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  inverter inv_n93( .i (n92), .o (n93) );
  assign n94 = G12 | G13 ;
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  assign n142 = ~G11 | ~n141 ;
  assign n143 = G1 | G3 ;
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  assign n171 = G32 & ~G9 ;
  assign n172 = G31 & ~G8 ;
  assign n173 = n171 | n172 ;
  assign n174 = ~G13 & G36 ;
  assign n175 = ~G14 & G37 ;
  assign n176 = n174 | n175 ;
  assign n177 = n173 | n176 ;
  assign n178 = ~G11 & G34 ;
  assign n179 = ~G12 & G35 ;
  assign n180 = n178 | n179 ;
  assign n181 = ~G10 & G33 ;
  assign n182 = G30 & ~G7 ;
  assign n183 = n181 | n182 ;
  assign n184 = n180 | n183 ;
  assign n185 = n177 | n184 ;
  assign n186 = n170 & n185 ;
  assign n187 = ~G1 & G2 ;
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  assign n223 = ~G3 & n222 ;
  buffer buf_n224( .i (n223), .o (n224) );
  assign n225 = ~G7 & n75 ;
  buffer buf_n226( .i (n225), .o (n226) );
  assign n227 = n224 & n226 ;
  assign n228 = G2 | n144 ;
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  assign n253 = G35 | G36 ;
  assign n254 = G34 & n253 ;
  assign n255 = ~n252 & n254 ;
  assign n256 = n227 | n255 ;
  assign n257 = n186 | n256 ;
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  inverter inv_n268( .i (n267), .o (n268) );
  assign n269 = G36 | G37 ;
  assign n270 = G36 & G37 ;
  assign n271 = n269 & ~n270 ;
  buffer buf_n272( .i (n271), .o (n272) );
  assign n273 = G34 & ~G35 ;
  assign n274 = ~G34 & G35 ;
  assign n275 = n273 | n274 ;
  buffer buf_n276( .i (n275), .o (n276) );
  assign n277 = n272 | n276 ;
  assign n278 = n272 & n276 ;
  assign n279 = n277 & ~n278 ;
  buffer buf_n280( .i (n279), .o (n280) );
  assign n281 = G30 & ~G31 ;
  assign n282 = ~G30 & G31 ;
  assign n283 = n281 | n282 ;
  buffer buf_n284( .i (n283), .o (n284) );
  assign n285 = G32 | G33 ;
  assign n286 = G32 & G33 ;
  assign n287 = n285 & ~n286 ;
  buffer buf_n288( .i (n287), .o (n288) );
  assign n289 = n284 | n288 ;
  assign n290 = n284 & n288 ;
  assign n291 = n289 & ~n290 ;
  buffer buf_n292( .i (n291), .o (n292) );
  assign n293 = n280 | n292 ;
  assign n294 = n280 & n292 ;
  assign n295 = n293 & ~n294 ;
  assign n296 = G8 & G9 ;
  assign n297 = n52 & ~n296 ;
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  assign n323 = G10 & G7 ;
  assign n324 = n78 & ~n323 ;
  buffer buf_n325( .i (n324), .o (n325) );
  assign n326 = ~n322 & n325 ;
  assign n327 = n322 & ~n325 ;
  assign n328 = n326 | n327 ;
  buffer buf_n329( .i (n328), .o (n329) );
  assign n330 = ~G11 & G13 ;
  assign n331 = G11 & ~G13 ;
  assign n332 = n330 | n331 ;
  buffer buf_n333( .i (n332), .o (n333) );
  assign n334 = G12 | G14 ;
  assign n335 = G12 & G14 ;
  assign n336 = n334 & ~n335 ;
  buffer buf_n337( .i (n336), .o (n337) );
  assign n338 = n333 & ~n337 ;
  assign n339 = ~n333 & n337 ;
  assign n340 = n338 | n339 ;
  buffer buf_n341( .i (n340), .o (n341) );
  assign n342 = n329 & n341 ;
  assign n343 = n329 | n341 ;
  assign n344 = ~n342 & n343 ;
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  assign n353 = G3 & n188 ;
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  assign n367 = G7 | n366 ;
  assign n368 = ~G1 & G3 ;
  buffer buf_n369( .i (n368), .o (n369) );
  assign n370 = G1 & G2 ;
  buffer buf_n371( .i (n370), .o (n371) );
  assign n375 = G1 & G3 ;
  assign n376 = G4 & n375 ;
  assign n377 = n371 | n376 ;
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  assign n392 = n369 | n386 ;
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  assign n396 = G7 & n395 ;
  assign n397 = n367 & ~n396 ;
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  assign n398 = G7 | n53 ;
  assign n399 = G3 & n398 ;
  assign n400 = G3 | G4 ;
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  assign n411 = G21 & ~n410 ;
  assign n412 = ~G3 & G4 ;
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  assign n442 = ~G8 & n422 ;
  assign n443 = n411 | n442 ;
  assign n444 = n399 | n443 ;
  assign n445 = n391 & n444 ;
  assign n446 = n397 | n445 ;
  buffer buf_n447( .i (n446), .o (n447) );
  assign n457 = G25 | G26 ;
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  assign n472 = G5 | G6 ;
  assign n473 = ~G1 & n472 ;
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  assign n477 = G4 & G5 ;
  buffer buf_n478( .i (n477), .o (n478) );
  assign n509 = n371 & ~n478 ;
  buffer buf_n510( .i (n509), .o (n510) );
  assign n523 = G38 & ~n510 ;
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  assign n532 = n475 & n531 ;
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n476( .i (n475), .o (n476) );
  assign n536 = G30 & ~n476 ;
  assign n537 = G4 | G49 ;
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  assign n548 = G28 & ~n547 ;
  assign n549 = G10 & ~G4 ;
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  assign n558 = G29 & G4 ;
  assign n559 = n557 | n558 ;
  assign n560 = n548 | n559 ;
  assign n561 = n536 | n560 ;
  assign n562 = ~n522 & n561 ;
  assign n563 = n535 | n562 ;
  buffer buf_n564( .i (n563), .o (n564) );
  assign n565 = n467 & ~n564 ;
  assign n566 = n447 | n565 ;
  buffer buf_n567( .i (n566), .o (n567) );
  assign n572 = G23 | G24 ;
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  assign n583 = ~n564 & n582 ;
  assign n584 = n447 & n583 ;
  buffer buf_n585( .i (n584), .o (n585) );
  assign n591 = n567 & ~n585 ;
  buffer buf_n592( .i (n591), .o (n592) );
  assign n600 = G8 & n395 ;
  assign n601 = G8 | n366 ;
  assign n602 = ~n600 & n601 ;
  assign n603 = G3 & n298 ;
  assign n604 = ~G9 & n422 ;
  assign n605 = G22 & ~G3 ;
  buffer buf_n606( .i (n605), .o (n606) );
  assign n625 = ~G4 & n606 ;
  assign n626 = n604 | n625 ;
  assign n627 = n603 | n626 ;
  assign n628 = n391 & n627 ;
  assign n629 = n602 | n628 ;
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n468( .i (n467), .o (n468) );
  assign n635 = G31 & ~n476 ;
  assign n636 = G29 & ~n547 ;
  assign n637 = G11 | G4 ;
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  assign n644 = ~G30 & G4 ;
  assign n645 = n643 & ~n644 ;
  assign n646 = n636 | n645 ;
  assign n647 = n635 | n646 ;
  assign n648 = ~n522 & n647 ;
  assign n649 = n535 | n648 ;
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  assign n652 = n468 & ~n651 ;
  assign n653 = n631 | n652 ;
  assign n654 = n582 & ~n650 ;
  assign n655 = n630 & n654 ;
  buffer buf_n656( .i (n655), .o (n656) );
  assign n666 = n653 & ~n656 ;
  buffer buf_n667( .i (n666), .o (n667) );
  assign n670 = n592 & n667 ;
  buffer buf_n671( .i (n670), .o (n671) );
  assign n673 = G3 & n379 ;
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  assign n682 = n393 & ~n681 ;
  assign n683 = G10 & ~n682 ;
  assign n684 = ~G10 & n364 ;
  assign n685 = G8 | n408 ;
  assign n686 = ~G11 & n420 ;
  assign n687 = n685 & ~n686 ;
  assign n688 = n388 & ~n687 ;
  assign n689 = n684 | n688 ;
  assign n690 = n683 | n689 ;
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  assign n694 = G33 & ~n474 ;
  assign n695 = G31 & ~n545 ;
  assign n696 = G13 | G4 ;
  assign n697 = ~G32 & G4 ;
  assign n698 = n696 & ~n697 ;
  assign n699 = n695 | n698 ;
  assign n700 = n694 | n699 ;
  assign n701 = ~n520 & n700 ;
  assign n702 = n533 | n701 ;
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  assign n705 = n466 & ~n704 ;
  assign n706 = n692 | n705 ;
  assign n707 = n580 & ~n703 ;
  assign n708 = n691 & n707 ;
  buffer buf_n709( .i (n708), .o (n709) );
  assign n715 = n706 & ~n709 ;
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  assign n730 = n358 | n675 ;
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  assign n737 = ~G9 & n736 ;
  assign n738 = G7 & ~n408 ;
  assign n739 = G10 & n420 ;
  assign n740 = n738 | n739 ;
  assign n741 = n388 & n740 ;
  assign n742 = G9 & ~n393 ;
  assign n743 = n741 | n742 ;
  assign n744 = n737 | n743 ;
  buffer buf_n745( .i (n744), .o (n745) );
  assign n748 = G32 & ~n474 ;
  assign n749 = G30 & ~n545 ;
  assign n750 = G12 | G4 ;
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  assign n753 = ~G31 & G4 ;
  assign n754 = n752 & ~n753 ;
  assign n755 = n749 | n754 ;
  assign n756 = n748 | n755 ;
  assign n757 = ~n520 & n756 ;
  assign n758 = n533 | n757 ;
  buffer buf_n759( .i (n758), .o (n759) );
  assign n760 = n465 & ~n759 ;
  assign n761 = n745 | n760 ;
  buffer buf_n762( .i (n761), .o (n762) );
  assign n768 = n580 & ~n759 ;
  assign n769 = n745 & n768 ;
  buffer buf_n770( .i (n769), .o (n770) );
  assign n777 = n762 & ~n770 ;
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  assign n782 = n719 & n781 ;
  assign n783 = n671 & n782 ;
  buffer buf_n784( .i (n783), .o (n784) );
  assign n791 = G11 | n95 ;
  assign n792 = G3 & n791 ;
  assign n793 = G9 | n401 ;
  assign n794 = ~G12 & n413 ;
  assign n795 = n793 & ~n794 ;
  assign n796 = ~n792 & n795 ;
  assign n797 = n382 & ~n796 ;
  assign n798 = ~G1 & G4 ;
  assign n799 = n354 | n798 ;
  assign n800 = n379 | n799 ;
  buffer buf_n801( .i (n800), .o (n801) );
  assign n806 = G11 & ~n801 ;
  assign n807 = ~G11 & n357 ;
  assign n808 = n806 | n807 ;
  assign n809 = n797 | n808 ;
  buffer buf_n810( .i (n809), .o (n810) );
  assign n827 = G32 & ~n539 ;
  assign n828 = G14 | G4 ;
  assign n829 = ~G33 & G4 ;
  assign n830 = n828 & ~n829 ;
  assign n831 = n827 | n830 ;
  assign n832 = G1 | G6 ;
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  assign n843 = G38 | n835 ;
  assign n844 = ~G34 & n835 ;
  assign n845 = n843 & ~n844 ;
  assign n846 = n831 | n845 ;
  assign n847 = ~n514 & n846 ;
  buffer buf_n848( .i (n847), .o (n848) );
  assign n856 = n573 & ~n848 ;
  assign n857 = n810 & n856 ;
  buffer buf_n858( .i (n857), .o (n858) );
  assign n864 = n458 & ~n848 ;
  assign n865 = n810 | n864 ;
  buffer buf_n866( .i (n865), .o (n866) );
  assign n871 = ~n858 & n866 ;
  buffer buf_n872( .i (n871), .o (n872) );
  assign n887 = G12 | n357 ;
  assign n888 = G12 & n801 ;
  assign n889 = n887 & ~n888 ;
  assign n890 = G12 & G13 ;
  assign n891 = n95 & ~n890 ;
  buffer buf_n892( .i (n891), .o (n892) );
  assign n925 = n674 & n892 ;
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  assign n926 = ~G3 & n374 ;
  buffer buf_n927( .i (n926), .o (n927) );
  assign n932 = G13 & G4 ;
  assign n933 = n550 | n932 ;
  assign n934 = n927 & n933 ;
  assign n935 = n925 | n934 ;
  assign n936 = n889 | n935 ;
  buffer buf_n937( .i (n936), .o (n937) );
  assign n948 = G5 | n833 ;
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  assign n953 = n524 & ~n950 ;
  buffer buf_n954( .i (n953), .o (n954) );
  assign n959 = G35 & n949 ;
  assign n960 = G33 & ~n538 ;
  assign n961 = G39 | G4 ;
  assign n962 = ~G34 & G4 ;
  assign n963 = n961 & ~n962 ;
  assign n964 = n960 | n963 ;
  assign n965 = n959 | n964 ;
  assign n966 = ~n513 & n965 ;
  assign n967 = n954 | n966 ;
  buffer buf_n968( .i (n967), .o (n968) );
  assign n978 = n573 & ~n968 ;
  assign n979 = n937 & n978 ;
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n969( .i (n968), .o (n969) );
  assign n997 = n459 & ~n969 ;
  assign n998 = n938 | n997 ;
  assign n999 = ~n980 & n998 ;
  buffer buf_n1000( .i (n999), .o (n1000) );
  assign n1009 = n872 & n1000 ;
  buffer buf_n1010( .i (n1009), .o (n1010) );
  assign n1012 = ~G13 & n731 ;
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  assign n1013 = G13 & ~n803 ;
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  assign n1014 = G14 & G4 ;
  assign n1015 = n638 & ~n1014 ;
  assign n1016 = n929 & ~n1015 ;
  assign n1017 = n1013 | n1016 ;
  assign n1018 = n1012 | n1017 ;
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  assign n1024 = G36 & n950 ;
  assign n1025 = G35 & G4 ;
  assign n1026 = ~G4 & G40 ;
  assign n1027 = n1025 | n1026 ;
  assign n1028 = G34 & ~n539 ;
  assign n1029 = n1027 | n1028 ;
  assign n1030 = n1024 | n1029 ;
  assign n1031 = ~n514 & n1030 ;
  buffer buf_n1032( .i (n1031), .o (n1032) );
  assign n1040 = n956 | n1032 ;
  buffer buf_n1041( .i (n1040), .o (n1041) );
  assign n1048 = n575 & ~n1041 ;
  assign n1049 = n1019 & n1048 ;
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  assign n1059 = n461 & ~n1042 ;
  assign n1060 = n1020 | n1059 ;
  assign n1061 = ~n1050 & n1060 ;
  buffer buf_n1062( .i (n1061), .o (n1062) );
  assign n1072 = n1010 & n1062 ;
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  assign n1074 = ~n678 & n805 ;
  assign n1075 = G14 & ~n1074 ;
  assign n1076 = ~G14 & n361 ;
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  assign n1077 = G39 & G4 ;
  assign n1078 = n751 & ~n1077 ;
  assign n1079 = n931 & ~n1078 ;
  assign n1080 = n1076 | n1079 ;
  assign n1081 = n1075 | n1080 ;
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  assign n1090 = G37 & n952 ;
  assign n1091 = G36 & G4 ;
  assign n1092 = ~G4 & G41 ;
  assign n1093 = n1091 | n1092 ;
  assign n1094 = G35 & ~n541 ;
  assign n1095 = n1093 | n1094 ;
  assign n1096 = n1090 | n1095 ;
  assign n1097 = ~n516 & n1096 ;
  buffer buf_n1098( .i (n1097), .o (n1098) );
  assign n1104 = n958 | n1098 ;
  buffer buf_n1105( .i (n1104), .o (n1105) );
  assign n1110 = n577 & ~n1105 ;
  assign n1111 = n1082 & n1110 ;
  buffer buf_n1112( .i (n1111), .o (n1112) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  assign n1116 = n463 & ~n1106 ;
  assign n1117 = n1083 | n1116 ;
  assign n1118 = ~n1112 & n1117 ;
  buffer buf_n1119( .i (n1118), .o (n1119) );
  assign n1125 = n1073 & n1119 ;
  buffer buf_n1126( .i (n1125), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n1133( .i (n1132), .o (n1133) );
  assign n1134 = n784 & n1133 ;
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  assign n1158 = n1073 & n1114 ;
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1053( .i (n1052), .o (n1053) );
  assign n1159 = n1011 & n1053 ;
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  assign n1160 = n870 & n984 ;
  assign n1161 = n863 | n1160 ;
  assign n1162 = n1159 | n1161 ;
  assign n1163 = n1158 | n1162 ;
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  assign n1172 = n785 & n1171 ;
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  assign n1173 = n714 & n767 ;
  assign n1174 = n776 | n1173 ;
  assign n1175 = n672 & n1174 ;
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  assign n1176 = n571 & n660 ;
  assign n1177 = n590 | n1176 ;
  assign n1178 = n1175 | n1177 ;
  buffer buf_n1179( .i (n1178), .o (n1179) );
  assign n1180 = n1172 | n1179 ;
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  assign n1202 = G27 & G48 ;
  buffer buf_n1203( .i (n1202), .o (n1203) );
  assign n1236 = ~n229 & n1203 ;
  buffer buf_n1237( .i (n1236), .o (n1237) );
  assign n1250 = n1023 & n1237 ;
  buffer buf_n1251( .i (n1250), .o (n1251) );
  assign n1252 = n1064 | n1251 ;
  assign n1253 = n1064 & n1251 ;
  assign n1254 = n1252 & ~n1253 ;
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  assign n1269 = n1089 & n1242 ;
  buffer buf_n1270( .i (n1269), .o (n1270) );
  assign n1271 = n1124 | n1270 ;
  assign n1272 = n1124 & n1270 ;
  assign n1273 = n1271 & ~n1272 ;
  buffer buf_n1274( .i (n1273), .o (n1274) );
  assign n1284 = G47 & n1274 ;
  assign n1285 = ~n1261 & n1284 ;
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1304( .i (n1303), .o (n1304) );
  buffer buf_n1305( .i (n1304), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  assign n1309 = G5 & ~n245 ;
  buffer buf_n1310( .i (n1309), .o (n1310) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  buffer buf_n1313( .i (n1312), .o (n1313) );
  buffer buf_n1314( .i (n1313), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  assign n1316 = n226 & ~n1315 ;
  assign n1317 = n1164 & ~n1242 ;
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  assign n1333 = ~G1 & n1332 ;
  assign n1334 = n1316 | n1333 ;
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n1280( .i (n1279), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  assign n1347 = ~G2 & n441 ;
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  assign n1350 = n1283 & n1349 ;
  assign n1351 = ~G6 & n1310 ;
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  assign n1357 = ~G23 & G3 ;
  assign n1358 = n218 & ~n1357 ;
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  assign n1364 = G25 & G3 ;
  buffer buf_n1365( .i (n1364), .o (n1365) );
  assign n1366 = G24 & G3 ;
  buffer buf_n1367( .i (n1366), .o (n1367) );
  assign n1368 = G26 & ~n1367 ;
  buffer buf_n1369( .i (n1368), .o (n1369) );
  assign n1370 = n1365 & n1369 ;
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1373( .i (n1372), .o (n1373) );
  buffer buf_n1374( .i (n1373), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  assign n1379 = G39 | G43 ;
  buffer buf_n1380( .i (n1379), .o (n1380) );
  assign n1381 = ~n1375 & n1380 ;
  assign n1382 = ~G3 & G41 ;
  assign n1383 = G4 & ~n1382 ;
  assign n1384 = ~n1381 & n1383 ;
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  assign n1385 = G24 | n471 ;
  assign n1386 = G3 & n1385 ;
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  buffer buf_n1390( .i (n1389), .o (n1390) );
  buffer buf_n1391( .i (n1390), .o (n1391) );
  assign n1395 = G40 & n1391 ;
  assign n1396 = G26 | n1367 ;
  buffer buf_n1397( .i (n1396), .o (n1397) );
  assign n1398 = n1365 | n1397 ;
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  assign n1407 = G44 & n1402 ;
  assign n1408 = n1395 | n1407 ;
  assign n1409 = ~n1365 & n1369 ;
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  assign n1417 = G41 | G45 ;
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  assign n1420 = ~n1413 & n1419 ;
  assign n1421 = n1365 & ~n1397 ;
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  assign n1429 = G42 | G46 ;
  assign n1430 = ~n1425 & n1429 ;
  assign n1431 = n1420 | n1430 ;
  assign n1432 = n1408 | n1431 ;
  assign n1433 = n1384 & ~n1432 ;
  assign n1434 = G3 & n1410 ;
  buffer buf_n1435( .i (n1434), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  assign n1441 = G11 | n1436 ;
  buffer buf_n1442( .i (n1441), .o (n1442) );
  assign n1444 = G13 | n1373 ;
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  assign n1447 = n1442 & n1446 ;
  assign n1448 = G9 | n1372 ;
  buffer buf_n1449( .i (n1448), .o (n1449) );
  assign n1451 = G7 | n1412 ;
  assign n1452 = n1449 & n1451 ;
  assign n1453 = G10 | n1424 ;
  assign n1454 = ~G8 & n1401 ;
  assign n1455 = n1453 & ~n1454 ;
  assign n1456 = n1452 & n1455 ;
  assign n1457 = G22 & ~n1423 ;
  assign n1458 = G4 | n1457 ;
  buffer buf_n1459( .i (n1458), .o (n1459) );
  assign n1463 = ~G12 & n1390 ;
  buffer buf_n1464( .i (n1463), .o (n1464) );
  assign n1468 = n1459 | n1464 ;
  assign n1469 = n1456 & ~n1468 ;
  assign n1470 = n1447 & n1469 ;
  assign n1471 = n1433 | n1470 ;
  assign n1472 = ~n1360 & n1471 ;
  assign n1473 = n1353 & ~n1472 ;
  assign n1474 = ~n1350 & n1473 ;
  assign n1475 = G47 & ~n1274 ;
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  assign n1485 = ~G47 & n1282 ;
  assign n1486 = n1353 | n1485 ;
  assign n1487 = n1484 | n1486 ;
  assign n1488 = ~n1474 & n1487 ;
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  inverter inv_n1501( .i (n1500), .o (n1501) );
  buffer buf_n693( .i (n692), .o (n693) );
  assign n1502 = n693 & n1240 ;
  buffer buf_n1503( .i (n1502), .o (n1503) );
  assign n1504 = n716 | n1503 ;
  assign n1505 = n716 & n1503 ;
  assign n1506 = n1504 & ~n1505 ;
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  assign n1522 = ~G2 & G4 ;
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  assign n1526 = n1521 & n1525 ;
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  assign n1527 = G20 & n1406 ;
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  assign n1528 = ~G8 & n1394 ;
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  assign n1529 = G19 & ~n1416 ;
  assign n1530 = n1528 | n1529 ;
  assign n1531 = n1527 | n1530 ;
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  assign n1532 = G7 | n1440 ;
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n1461( .i (n1460), .o (n1461) );
  buffer buf_n1462( .i (n1461), .o (n1462) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  assign n1533 = G18 & ~n1427 ;
  buffer buf_n1376( .i (n1375), .o (n1376) );
  assign n1534 = ~G21 & G9 ;
  assign n1535 = n1376 | n1534 ;
  assign n1536 = ~n1533 & n1535 ;
  assign n1537 = ~n1462 & n1536 ;
  assign n1538 = n1532 & n1537 ;
  assign n1539 = ~n1531 & n1538 ;
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  assign n1540 = G40 & n1405 ;
  assign n1541 = n1467 | n1540 ;
  assign n1542 = G41 & ~n1416 ;
  buffer buf_n1377( .i (n1376), .o (n1377) );
  assign n1543 = G11 & ~G39 ;
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  assign n1546 = n1377 | n1545 ;
  assign n1547 = ~n1542 & n1546 ;
  assign n1548 = ~n1541 & n1547 ;
  assign n1549 = G13 | n1440 ;
  buffer buf_n1428( .i (n1427), .o (n1428) );
  assign n1550 = G14 & ~G42 ;
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  assign n1556 = n1428 | n1555 ;
  assign n1557 = G4 & n1556 ;
  assign n1558 = n1549 & n1557 ;
  assign n1559 = n1548 & n1558 ;
  assign n1560 = n1539 | n1559 ;
  assign n1561 = ~n1363 & n1560 ;
  assign n1562 = n1356 & ~n1561 ;
  assign n1563 = ~n1526 & n1562 ;
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1038( .i (n1037), .o (n1038) );
  buffer buf_n1039( .i (n1038), .o (n1039) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  assign n1564 = n1039 | n1103 ;
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  assign n1565 = G24 | n855 ;
  assign n1566 = n1564 | n1565 ;
  assign n1567 = n977 | n1566 ;
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n1109( .i (n1108), .o (n1109) );
  assign n1568 = n1047 & n1109 ;
  assign n1569 = G24 & n855 ;
  assign n1570 = n976 & n1569 ;
  assign n1571 = n1568 & n1570 ;
  assign n1572 = n1567 & ~n1571 ;
  assign n1573 = n1241 | n1572 ;
  assign n1574 = n1126 & n1241 ;
  assign n1575 = n1573 & ~n1574 ;
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  assign n1589 = G47 & ~n1588 ;
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  assign n1592 = ~n1321 & n1509 ;
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  assign n1601 = ~n729 & n1329 ;
  assign n1602 = n1600 | n1601 ;
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  assign n1605 = n1591 | n1604 ;
  assign n1606 = n1590 & n1603 ;
  assign n1607 = n1356 | n1606 ;
  assign n1608 = n1605 & ~n1607 ;
  assign n1609 = n1563 | n1608 ;
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  assign n1620 = G47 & n1576 ;
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  assign n1632 = n747 & n1240 ;
  buffer buf_n1633( .i (n1632), .o (n1633) );
  assign n1634 = n778 & ~n1633 ;
  assign n1635 = ~n778 & n1633 ;
  assign n1636 = n1634 | n1635 ;
  buffer buf_n1637( .i (n1636), .o (n1637) );
  assign n1651 = n1507 & n1637 ;
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  assign n1655 = G27 & ~n236 ;
  buffer buf_n1656( .i (n1655), .o (n1656) );
  assign n1664 = n634 & n1656 ;
  buffer buf_n1665( .i (n1664), .o (n1665) );
  assign n1666 = n669 | n1665 ;
  assign n1667 = n669 & n1665 ;
  assign n1668 = n1666 & ~n1667 ;
  buffer buf_n1669( .i (n1668), .o (n1669) );
  assign n1678 = n1654 & n1669 ;
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  assign n1683 = n790 & n1682 ;
  assign n1684 = n790 | n1682 ;
  assign n1685 = ~n1683 & n1684 ;
  assign n1686 = n1631 & ~n1685 ;
  buffer buf_n1687( .i (n1686), .o (n1687) );
  assign n1688 = n785 | n1323 ;
  assign n1689 = ~n1179 & n1688 ;
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  assign n1694 = n776 & ~n1246 ;
  buffer buf_n1638( .i (n1637), .o (n1638) );
  assign n1695 = n713 & ~n1244 ;
  buffer buf_n1696( .i (n1695), .o (n1696) );
  assign n1700 = n1638 & ~n1696 ;
  assign n1701 = n1694 | n1700 ;
  buffer buf_n1702( .i (n1701), .o (n1702) );
  assign n1704 = n1669 & n1702 ;
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  buffer buf_n1658( .i (n1657), .o (n1658) );
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  assign n1707 = n665 & ~n1663 ;
  assign n1708 = n1706 | n1707 ;
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1710( .i (n1709), .o (n1710) );
  assign n1711 = n1693 & n1710 ;
  assign n1712 = n1693 | n1710 ;
  assign n1713 = ~n1711 & n1712 ;
  buffer buf_n1714( .i (n1713), .o (n1714) );
  assign n1715 = n1687 & n1714 ;
  assign n1716 = n1687 | n1714 ;
  assign n1717 = ~n1715 & n1716 ;
  assign n1718 = G1 | G2 ;
  buffer buf_n1719( .i (n1718), .o (n1719) );
  assign n1720 = n170 & n1719 ;
  assign n1721 = ~n1717 & n1720 ;
  assign n1722 = G7 & ~G9 ;
  assign n1723 = n78 | n320 ;
  assign n1724 = ~n1722 & n1723 ;
  assign n1725 = n1719 | n1724 ;
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  assign n1726 = ~G14 & n224 ;
  assign n1727 = ~n924 & n1726 ;
  assign n1728 = n1725 & ~n1727 ;
  assign n1729 = ~n1721 & n1728 ;
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n1732( .i (n1731), .o (n1732) );
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n1734( .i (n1733), .o (n1734) );
  buffer buf_n1735( .i (n1734), .o (n1735) );
  buffer buf_n1736( .i (n1735), .o (n1736) );
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  inverter inv_n1739( .i (n1738), .o (n1739) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  assign n1740 = ~n369 & n842 ;
  assign n1741 = ~n199 & n1740 ;
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  assign n1767 = n1115 & ~n1240 ;
  buffer buf_n1768( .i (n1767), .o (n1768) );
  assign n1773 = n1255 | n1768 ;
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  assign n1778 = n1071 & n1772 ;
  assign n1779 = n1777 & ~n1778 ;
  buffer buf_n1780( .i (n1779), .o (n1780) );
  assign n1781 = n1476 | n1780 ;
  assign n1782 = n1476 & n1780 ;
  assign n1783 = n1781 & ~n1782 ;
  buffer buf_n1784( .i (n1783), .o (n1784) );
  assign n1789 = n1326 & n1784 ;
  assign n1790 = n1310 | n1789 ;
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  assign n1794 = n947 & n1241 ;
  buffer buf_n1795( .i (n1794), .o (n1795) );
  assign n1796 = n1008 | n1795 ;
  assign n1797 = n1008 & n1795 ;
  assign n1798 = n1796 & ~n1797 ;
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  assign n1809 = n1058 & ~n1243 ;
  assign n1810 = n1774 & ~n1809 ;
  buffer buf_n1811( .i (n1810), .o (n1811) );
  assign n1813 = n1799 | n1811 ;
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1800( .i (n1799), .o (n1800) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  assign n1817 = n1800 & n1812 ;
  assign n1818 = n1814 & ~n1817 ;
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  assign n1821 = ~n1287 & n1820 ;
  assign n1822 = n1286 & ~n1819 ;
  buffer buf_n1823( .i (n1822), .o (n1823) );
  assign n1827 = n1821 | n1823 ;
  buffer buf_n1828( .i (n1827), .o (n1828) );
  assign n1832 = n1328 & ~n1828 ;
  assign n1833 = n1791 | n1832 ;
  assign n1834 = ~n1763 & n1833 ;
  buffer buf_n1824( .i (n1823), .o (n1824) );
  buffer buf_n1825( .i (n1824), .o (n1825) );
  buffer buf_n1826( .i (n1825), .o (n1826) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n1247( .i (n1246), .o (n1247) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  assign n1835 = n996 & ~n1249 ;
  assign n1836 = n1816 & ~n1835 ;
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  assign n1838 = n826 & n1247 ;
  buffer buf_n1839( .i (n1838), .o (n1839) );
  assign n1840 = n886 | n1839 ;
  assign n1841 = n886 & n1839 ;
  assign n1842 = n1840 & ~n1841 ;
  buffer buf_n1843( .i (n1842), .o (n1843) );
  assign n1848 = n1837 & ~n1843 ;
  assign n1849 = ~n1837 & n1843 ;
  assign n1850 = n1848 | n1849 ;
  buffer buf_n1851( .i (n1850), .o (n1851) );
  assign n1852 = n1826 & ~n1851 ;
  assign n1853 = ~n1826 & n1851 ;
  assign n1854 = n1852 | n1853 ;
  assign n1855 = ~n1834 & n1854 ;
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  buffer buf_n1846( .i (n1845), .o (n1846) );
  buffer buf_n1847( .i (n1846), .o (n1847) );
  assign n1856 = n1349 & n1847 ;
  assign n1857 = ~G19 & G7 ;
  buffer buf_n1858( .i (n1857), .o (n1858) );
  assign n1859 = n1425 | n1858 ;
  assign n1860 = G21 & n1401 ;
  assign n1861 = G20 & ~n1412 ;
  assign n1862 = n1860 | n1861 ;
  assign n1863 = n1859 & ~n1862 ;
  assign n1864 = G10 & ~G22 ;
  assign n1865 = n1375 | n1864 ;
  assign n1866 = n1863 & n1865 ;
  assign n1867 = ~G9 & n1390 ;
  buffer buf_n1868( .i (n1867), .o (n1868) );
  assign n1870 = G8 | n1436 ;
  assign n1871 = ~n1868 & n1870 ;
  assign n1872 = ~G4 & n1871 ;
  assign n1873 = n1866 & n1872 ;
  assign n1874 = n1380 & ~n1426 ;
  assign n1875 = G12 & ~G40 ;
  buffer buf_n1876( .i (n1875), .o (n1876) );
  assign n1878 = n1375 | n1876 ;
  assign n1879 = ~n1874 & n1878 ;
  assign n1880 = G42 & ~n1413 ;
  assign n1881 = G41 & n1402 ;
  assign n1882 = n1880 | n1881 ;
  assign n1883 = G14 | n1436 ;
  assign n1884 = ~G13 & n1390 ;
  assign n1885 = G4 & ~n1884 ;
  assign n1886 = n1883 & n1885 ;
  assign n1887 = ~n1882 & n1886 ;
  assign n1888 = n1879 & n1887 ;
  assign n1889 = n1873 | n1888 ;
  assign n1890 = ~n1360 & n1889 ;
  assign n1891 = n1353 & ~n1890 ;
  assign n1892 = ~n1856 & n1891 ;
  assign n1893 = n1855 | n1892 ;
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1895( .i (n1894), .o (n1895) );
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1897( .i (n1896), .o (n1897) );
  buffer buf_n1898( .i (n1897), .o (n1898) );
  buffer buf_n1899( .i (n1898), .o (n1899) );
  buffer buf_n1900( .i (n1899), .o (n1900) );
  buffer buf_n1901( .i (n1900), .o (n1901) );
  buffer buf_n1902( .i (n1901), .o (n1902) );
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1904( .i (n1903), .o (n1904) );
  buffer buf_n1905( .i (n1904), .o (n1905) );
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  assign n1907 = n1326 | n1784 ;
  buffer buf_n1908( .i (n1907), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  assign n1912 = ~n1793 & n1911 ;
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  assign n1913 = n1763 & ~n1788 ;
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  assign n1914 = n1268 & n1348 ;
  buffer buf_n1915( .i (n1389), .o (n1915) );
  assign n1916 = G39 & n1915 ;
  assign n1917 = G44 & ~n1412 ;
  assign n1918 = n1916 | n1917 ;
  assign n1919 = n1418 & ~n1424 ;
  assign n1920 = G43 & n1401 ;
  assign n1921 = n1919 | n1920 ;
  assign n1922 = n1918 | n1921 ;
  buffer buf_n1923( .i (n1435), .o (n1923) );
  assign n1924 = G40 & ~n1923 ;
  assign n1925 = n1373 | n1551 ;
  assign n1926 = G4 & n1925 ;
  assign n1927 = ~n1924 & n1926 ;
  assign n1928 = ~n1922 & n1927 ;
  buffer buf_n1929( .i (n1400), .o (n1929) );
  assign n1930 = ~G7 & n1929 ;
  buffer buf_n1931( .i (n1411), .o (n1931) );
  assign n1932 = G22 & ~n1931 ;
  assign n1933 = n1930 | n1932 ;
  assign n1934 = G12 | n1372 ;
  buffer buf_n1935( .i (n1934), .o (n1935) );
  assign n1938 = G9 | n1424 ;
  assign n1939 = n1935 & n1938 ;
  assign n1940 = ~n1933 & n1939 ;
  assign n1941 = G10 | n1435 ;
  buffer buf_n1942( .i (n1941), .o (n1942) );
  assign n1946 = G8 | n1371 ;
  assign n1947 = ~G4 & n1946 ;
  buffer buf_n1948( .i (n1947), .o (n1948) );
  assign n1953 = ~G11 & n1388 ;
  buffer buf_n1954( .i (n1953), .o (n1954) );
  assign n1959 = G21 & ~n1422 ;
  buffer buf_n1960( .i (n1959), .o (n1960) );
  assign n1965 = n1954 | n1960 ;
  assign n1966 = n1948 & ~n1965 ;
  assign n1967 = n1942 & n1966 ;
  assign n1968 = n1940 & n1967 ;
  assign n1969 = n1928 | n1968 ;
  assign n1970 = ~n1359 & n1969 ;
  assign n1971 = n1352 & ~n1970 ;
  assign n1972 = ~n1914 & n1971 ;
  assign n1973 = n1913 | n1972 ;
  assign n1974 = n1912 | n1973 ;
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  buffer buf_n1978( .i (n1977), .o (n1978) );
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  buffer buf_n1981( .i (n1980), .o (n1981) );
  buffer buf_n1982( .i (n1981), .o (n1982) );
  buffer buf_n1983( .i (n1982), .o (n1983) );
  buffer buf_n1984( .i (n1983), .o (n1984) );
  buffer buf_n1985( .i (n1984), .o (n1985) );
  buffer buf_n1986( .i (n1985), .o (n1986) );
  buffer buf_n1987( .i (n1986), .o (n1987) );
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  assign n1988 = ~n1313 & n1910 ;
  assign n1989 = ~n1831 & n1988 ;
  buffer buf_n1801( .i (n1800), .o (n1801) );
  buffer buf_n1802( .i (n1801), .o (n1802) );
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  assign n1990 = n1348 & n1808 ;
  assign n1991 = G21 & ~n1413 ;
  buffer buf_n1992( .i (n1423), .o (n1992) );
  assign n1993 = G8 | n1992 ;
  assign n1994 = G11 & G7 ;
  assign n1995 = n1373 | n1994 ;
  assign n1996 = n1993 & n1995 ;
  assign n1997 = ~n1991 & n1996 ;
  assign n1998 = G9 | n1923 ;
  assign n1999 = G20 & ~n1422 ;
  assign n2000 = G4 | n1999 ;
  buffer buf_n2001( .i (n2000), .o (n2001) );
  assign n2005 = ~G10 & n1388 ;
  buffer buf_n2006( .i (n2005), .o (n2006) );
  assign n2009 = G22 & n1400 ;
  assign n2010 = n2006 | n2009 ;
  assign n2011 = n2001 | n2010 ;
  assign n2012 = n1998 & ~n2011 ;
  assign n2013 = n1997 & n2012 ;
  assign n2014 = G42 & n1929 ;
  assign n2015 = G40 | G44 ;
  assign n2016 = ~n1992 & n2015 ;
  assign n2017 = n2014 | n2016 ;
  assign n2018 = G43 & ~n1931 ;
  assign n2019 = ~G14 & n1915 ;
  assign n2020 = n2018 | n2019 ;
  assign n2021 = n2017 | n2020 ;
  assign n2022 = G39 & ~n1923 ;
  assign n2023 = G13 & ~G41 ;
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2028( .i (n1372), .o (n2028) );
  assign n2029 = n2024 | n2028 ;
  assign n2030 = G4 & n2029 ;
  assign n2031 = ~n2022 & n2030 ;
  assign n2032 = ~n2021 & n2031 ;
  assign n2033 = n2013 | n2032 ;
  assign n2034 = ~n1359 & n2033 ;
  assign n2035 = n1352 & ~n2034 ;
  assign n2036 = ~n1990 & n2035 ;
  assign n2037 = n1311 | n1908 ;
  assign n2038 = ~n1762 & n2037 ;
  assign n2039 = n1830 & ~n2038 ;
  assign n2040 = n2036 | n2039 ;
  assign n2041 = n1989 | n2040 ;
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  assign n2055 = n1626 & n1679 ;
  buffer buf_n2056( .i (n2055), .o (n2056) );
  assign n2061 = n1622 & n1652 ;
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  buffer buf_n2064( .i (n2063), .o (n2064) );
  buffer buf_n2065( .i (n2064), .o (n2065) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  assign n2066 = n1670 | n1703 ;
  assign n2067 = ~n1705 & n2066 ;
  assign n2068 = ~n2065 & n2067 ;
  assign n2069 = n2056 | n2068 ;
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n2073( .i (n2072), .o (n2073) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  assign n2075 = n1593 | n1699 ;
  buffer buf_n2076( .i (n2075), .o (n2076) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  assign n2077 = n1509 & n1622 ;
  assign n2078 = n1640 | n2077 ;
  assign n2079 = ~n2062 & n2078 ;
  buffer buf_n2080( .i (n2079), .o (n2080) );
  assign n2081 = n2076 | n2080 ;
  assign n2082 = n2076 & n2080 ;
  assign n2083 = n2081 & ~n2082 ;
  buffer buf_n2084( .i (n2083), .o (n2084) );
  assign n2090 = n1627 & ~n1690 ;
  buffer buf_n2091( .i (n2090), .o (n2091) );
  assign n2093 = n2084 | n2091 ;
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  assign n2096 = n1314 | n2095 ;
  assign n2097 = ~n1765 & n2096 ;
  assign n2098 = n2074 & ~n2097 ;
  assign n2099 = ~n1313 & n2094 ;
  buffer buf_n2100( .i (n2099), .o (n2100) );
  assign n2103 = ~n2073 & n2100 ;
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  assign n2104 = n1523 & n1677 ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1877( .i (n1876), .o (n1877) );
  assign n2105 = n1427 | n1877 ;
  assign n2106 = n1443 & n2105 ;
  assign n2107 = ~G14 & n1403 ;
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n2007( .i (n2006), .o (n2007) );
  buffer buf_n2008( .i (n2007), .o (n2008) );
  assign n2108 = n1450 & ~n2008 ;
  assign n2109 = ~n2107 & n2108 ;
  assign n2110 = G39 & ~n1414 ;
  assign n2111 = G4 & n1445 ;
  assign n2112 = ~n2110 & n2111 ;
  assign n2113 = n2109 & n2112 ;
  assign n2114 = n2106 & n2113 ;
  assign n2115 = G16 & ~n1427 ;
  assign n2116 = G17 & ~n1414 ;
  assign n2117 = G22 & n1392 ;
  assign n2118 = n2116 | n2117 ;
  assign n2119 = n2115 | n2118 ;
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n2003), .o (n2004) );
  assign n2120 = G21 & ~n1437 ;
  assign n2121 = G18 & n1402 ;
  assign n2122 = n1374 | n1858 ;
  assign n2123 = ~n2121 & n2122 ;
  assign n2124 = ~n2120 & n2123 ;
  assign n2125 = ~n2004 & n2124 ;
  assign n2126 = ~n2119 & n2125 ;
  assign n2127 = n2114 | n2126 ;
  assign n2128 = ~n1361 & n2127 ;
  assign n2129 = n1354 & ~n2128 ;
  assign n2130 = ~n2104 & n2129 ;
  assign n2131 = n2103 | n2130 ;
  assign n2132 = n2098 | n2131 ;
  buffer buf_n2133( .i (n2132), .o (n2133) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  buffer buf_n2136( .i (n2135), .o (n2136) );
  buffer buf_n2137( .i (n2136), .o (n2137) );
  buffer buf_n2138( .i (n2137), .o (n2138) );
  buffer buf_n2139( .i (n2138), .o (n2139) );
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n2143( .i (n2142), .o (n2143) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  assign n2144 = n456 & n1661 ;
  buffer buf_n2145( .i (n2144), .o (n2145) );
  assign n2146 = n599 | n2145 ;
  assign n2147 = n599 & n2145 ;
  assign n2148 = n2146 & ~n2147 ;
  buffer buf_n2149( .i (n2148), .o (n2149) );
  buffer buf_n2150( .i (n2149), .o (n2150) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  buffer buf_n2152( .i (n2151), .o (n2152) );
  buffer buf_n2153( .i (n2152), .o (n2153) );
  assign n2154 = n1524 & n2153 ;
  buffer buf_n1378( .i (n1377), .o (n1378) );
  assign n2155 = G18 | G22 ;
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n2158( .i (n2157), .o (n2158) );
  buffer buf_n2159( .i (n2158), .o (n2159) );
  assign n2160 = ~n1378 & n2159 ;
  assign n2161 = G16 & ~n1415 ;
  assign n2162 = G20 & ~n1438 ;
  assign n2163 = n2161 | n2162 ;
  assign n2164 = G17 & n1403 ;
  assign n2165 = G15 | G19 ;
  assign n2166 = ~n1426 & n2165 ;
  assign n2167 = n2164 | n2166 ;
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  assign n2168 = G21 & n1392 ;
  assign n2169 = n508 & ~n2168 ;
  assign n2170 = ~n2167 & n2169 ;
  assign n2171 = ~n2163 & n2170 ;
  assign n2172 = ~n2160 & n2171 ;
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  assign n2173 = G5 & n1945 ;
  buffer buf_n1869( .i (n1868), .o (n1869) );
  assign n2174 = G14 | n1414 ;
  assign n2175 = ~n1869 & n2174 ;
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  assign n2176 = ~G13 & n1403 ;
  assign n2177 = n1937 & ~n2176 ;
  assign n2178 = n2175 & n2177 ;
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n2179( .i (n1426), .o (n2179) );
  assign n2180 = n1544 | n2179 ;
  assign n2181 = n1951 & n2180 ;
  assign n2182 = n2178 & n2181 ;
  assign n2183 = n2173 & n2182 ;
  assign n2184 = n2172 | n2183 ;
  assign n2185 = ~n1362 & n2184 ;
  assign n2186 = n1355 & ~n2185 ;
  assign n2187 = ~n2154 & n2186 ;
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  assign n2188 = n2085 & n2092 ;
  buffer buf_n2189( .i (n2188), .o (n2189) );
  assign n2193 = ~n2070 & n2092 ;
  assign n2194 = n1313 | n2193 ;
  assign n2195 = n2189 | n2194 ;
  assign n2196 = ~n1765 & n2195 ;
  buffer buf_n2057( .i (n2056), .o (n2057) );
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  assign n2197 = n1709 & ~n2149 ;
  assign n2198 = ~n1709 & n2149 ;
  assign n2199 = n2197 | n2198 ;
  buffer buf_n2200( .i (n2199), .o (n2200) );
  assign n2201 = n2060 & ~n2200 ;
  assign n2202 = ~n2060 & n2200 ;
  assign n2203 = n2201 | n2202 ;
  assign n2204 = ~n2196 & n2203 ;
  assign n2205 = n2187 | n2204 ;
  buffer buf_n2206( .i (n2205), .o (n2206) );
  buffer buf_n2207( .i (n2206), .o (n2207) );
  buffer buf_n2208( .i (n2207), .o (n2208) );
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n2211( .i (n2210), .o (n2211) );
  buffer buf_n2212( .i (n2211), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  buffer buf_n2214( .i (n2213), .o (n2214) );
  buffer buf_n2215( .i (n2214), .o (n2215) );
  buffer buf_n2216( .i (n2215), .o (n2216) );
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n2102( .i (n2101), .o (n2102) );
  buffer buf_n2190( .i (n2189), .o (n2190) );
  buffer buf_n2191( .i (n2190), .o (n2191) );
  buffer buf_n2192( .i (n2191), .o (n2192) );
  assign n2217 = n2102 & ~n2192 ;
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  buffer buf_n1644( .i (n1643), .o (n1644) );
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  assign n2218 = n1524 & n1650 ;
  assign n2219 = G39 & n1404 ;
  assign n2220 = G40 & ~n1415 ;
  assign n2221 = n2219 | n2220 ;
  buffer buf_n1955( .i (n1954), .o (n1955) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  assign n2222 = G10 & G14 ;
  assign n2223 = n1376 | n2222 ;
  assign n2224 = ~n1958 & n2223 ;
  assign n2225 = ~n2221 & n2224 ;
  assign n2226 = G12 | n1439 ;
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  assign n2227 = n2027 | n2179 ;
  assign n2228 = G4 & n2227 ;
  assign n2229 = n2226 & n2228 ;
  assign n2230 = n2225 & n2229 ;
  assign n2231 = G17 & ~n1428 ;
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  assign n2232 = G19 & n1404 ;
  assign n2233 = n1964 | n2232 ;
  assign n2234 = n2231 | n2233 ;
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n622( .i (n621), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n2235( .i (n1931), .o (n2235) );
  buffer buf_n2236( .i (n2235), .o (n2236) );
  assign n2237 = n2156 & ~n2236 ;
  assign n2238 = n624 | n2237 ;
  assign n2239 = ~G7 & n1392 ;
  buffer buf_n2240( .i (n1374), .o (n2240) );
  assign n2241 = G20 & ~n2240 ;
  assign n2242 = n2239 | n2241 ;
  assign n2243 = n2238 | n2242 ;
  assign n2244 = n1952 & ~n2243 ;
  assign n2245 = ~n2234 & n2244 ;
  assign n2246 = n2230 | n2245 ;
  assign n2247 = ~n1362 & n2246 ;
  assign n2248 = n1355 & ~n2247 ;
  assign n2249 = ~n2218 & n2248 ;
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2089( .i (n2088), .o (n2089) );
  assign n2250 = n1766 & ~n2089 ;
  assign n2251 = n2249 | n2250 ;
  assign n2252 = n2217 | n2251 ;
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  assign n2263 = n2133 | n2206 ;
  buffer buf_n2264( .i (n2263), .o (n2264) );
  buffer buf_n2265( .i (n2264), .o (n2265) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  assign n2269 = n1610 | n2253 ;
  buffer buf_n2270( .i (n2269), .o (n2270) );
  assign n2271 = n1894 | n2042 ;
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2273( .i (n2272), .o (n2273) );
  buffer buf_n2274( .i (n2273), .o (n2274) );
  assign n2275 = n1489 & ~n1975 ;
  buffer buf_n2276( .i (n2275), .o (n2276) );
  buffer buf_n2277( .i (n2276), .o (n2277) );
  buffer buf_n2278( .i (n2277), .o (n2278) );
  assign n2279 = ~n2274 & n2278 ;
  assign n2280 = ~n2270 & n2279 ;
  assign n2281 = ~n2266 & n2280 ;
  buffer buf_n2282( .i (n2281), .o (n2282) );
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  inverter inv_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2267( .i (n2266), .o (n2267) );
  buffer buf_n2268( .i (n2267), .o (n2268) );
  assign n2287 = G48 & ~n2268 ;
  assign n2288 = G27 & ~n2282 ;
  assign n2289 = ~n2287 & n2288 ;
  buffer buf_n2290( .i (n2289), .o (n2290) );
  inverter inv_n2291( .i (n2290), .o (n2291) );
  assign n2292 = n1611 & n2254 ;
  assign n2293 = n2270 & ~n2292 ;
  buffer buf_n2294( .i (n2293), .o (n2294) );
  assign n2295 = ~n1490 & n1976 ;
  assign n2296 = n2276 | n2295 ;
  buffer buf_n2297( .i (n2296), .o (n2297) );
  assign n2298 = n1895 & n2043 ;
  assign n2299 = n2272 & ~n2298 ;
  buffer buf_n2300( .i (n2299), .o (n2300) );
  assign n2301 = n2297 | n2300 ;
  assign n2302 = n2297 & n2300 ;
  assign n2303 = n2301 & ~n2302 ;
  buffer buf_n2304( .i (n2303), .o (n2304) );
  assign n2305 = n2294 & n2304 ;
  assign n2306 = n2294 | n2304 ;
  assign n2307 = ~n2305 & n2306 ;
  buffer buf_n2308( .i (n2307), .o (n2308) );
  assign n2309 = n2134 & n2207 ;
  assign n2310 = n2264 & ~n2309 ;
  buffer buf_n2311( .i (n2310), .o (n2311) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  assign n2316 = G50 & n2312 ;
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  assign n2317 = G50 | n2311 ;
  assign n2318 = ~n1235 & n2317 ;
  assign n2319 = ~n2316 & n2318 ;
  buffer buf_n2320( .i (n2319), .o (n2320) );
  assign n2321 = n2308 & n2320 ;
  assign n2322 = n2308 | n2320 ;
  assign n2323 = n2321 | ~n2322 ;
  buffer buf_n2313( .i (n2312), .o (n2313) );
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2315( .i (n2314), .o (n2315) );
  assign n2324 = n2308 | n2315 ;
  assign n2325 = n2308 & n2315 ;
  assign n2326 = n2324 & ~n2325 ;
  assign G3519 = n93 ;
  assign G3520 = n142 ;
  assign G3521 = n268 ;
  assign G3522 = n295 ;
  assign G3523 = n352 ;
  assign G3524 = n1157 ;
  assign G3525 = n1201 ;
  assign G3526 = n1308 ;
  assign G3527 = n1346 ;
  assign G3528 = n1501 ;
  assign G3529 = n1619 ;
  assign G3530 = n1739 ;
  assign G3531 = n1906 ;
  assign G3532 = n1987 ;
  assign G3533 = n2054 ;
  assign G3534 = n2143 ;
  assign G3535 = n2216 ;
  assign G3536 = n2262 ;
  assign G3537 = n2286 ;
  assign G3538 = n2291 ;
  assign G3539 = n2323 ;
  assign G3540 = n2326 ;
endmodule
