module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 ;
  wire n2 , n3 , n4 , n5 , n6 , n8 , n9 , n10 , n12 , n13 , n15 , n16 , n17 , n18 , n19 , n20 , n22 , n23 , n24 , n25 , n26 , n28 , n29 , n31 , n32 , n33 , n34 , n36 , n37 , n38 , n39 , n40 , n42 , n43 , n44 , n45 , n46 , n47 , n49 , n50 , n51 , n52 , n54 , n55 , n57 , n58 , n59 , n60 , n62 , n63 , n64 , n65 , n67 , n68 , n69 , n70 , n71 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n111 , n112 , n113 , n114 , n116 , n117 , n118 , n119 , n121 , n122 , n123 , n124 , n126 , n127 , n128 , n129 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 ;
  buffer buf_n15( .i (x3), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n36( .i (x7), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n22( .i (x4), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  assign n143 = n25 | n39 ;
  buffer buf_n81( .i (x15), .o (n81) );
  buffer buf_n92( .i (x16), .o (n92) );
  assign n144 = n81 & n92 ;
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n73( .i (x14), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n111( .i (x18), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  assign n148 = n74 & n112 ;
  assign n149 = n145 & n148 ;
  buffer buf_n150( .i (n149), .o (n150) );
  assign n151 = ( n40 & n143 ) | ( n40 & ~n150 ) | ( n143 & ~n150 ) ;
  assign n152 = n20 & n151 ;
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n12( .i (x2), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n28( .i (x5), .o (n28) );
  buffer buf_n67( .i (x13), .o (n67) );
  assign n155 = n28 & n67 ;
  assign n156 = n13 & n155 ;
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n8( .i (x1), .o (n8) );
  assign n161 = ~n2 & n8 ;
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n101( .i (x17), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n113( .i (n112), .o (n113) );
  assign n166 = ~n103 & n113 ;
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  assign n169 = n165 & ~n168 ;
  assign n170 = n160 & n169 ;
  buffer buf_n171( .i (n170), .o (n171) );
  assign n172 = n154 & n171 ;
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n49( .i (x9), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  assign n175 = n16 & ~n50 ;
  buffer buf_n9( .i (n8), .o (n9) );
  assign n176 = n9 | n13 ;
  assign n177 = n175 & ~n176 ;
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  assign n180 = n40 & n71 ;
  assign n181 = n179 & n180 ;
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n131( .i (x22), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n121( .i (x20), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n126( .i (x21), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n116( .i (x19), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  assign n185 = n69 | n118 ;
  assign n186 = ( n124 & n129 ) | ( n124 & ~n185 ) | ( n129 & ~n185 ) ;
  assign n187 = ~n127 & n132 ;
  buffer buf_n188( .i (n187), .o (n188) );
  assign n189 = ( n124 & n129 ) | ( n124 & n188 ) | ( n129 & n188 ) ;
  assign n190 = n186 & ~n189 ;
  buffer buf_n191( .i (n190), .o (n191) );
  assign n195 = n137 & n191 ;
  assign n196 = n182 | n195 ;
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n82( .i (n81), .o (n82) );
  assign n199 = ~n29 & n82 ;
  buffer buf_n200( .i (n199), .o (n200) );
  assign n204 = n24 & n69 ;
  assign n205 = n200 & n204 ;
  buffer buf_n206( .i (n205), .o (n206) );
  assign n207 = ~n168 & n206 ;
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  assign n210 = n25 & n84 ;
  assign n211 = ~n167 & n210 ;
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  assign n212 = n75 & n94 ;
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  assign n215 = n211 & ~n214 ;
  buffer buf_n216( .i (n215), .o (n216) );
  assign n217 = ~n29 & n68 ;
  buffer buf_n218( .i (n217), .o (n218) );
  assign n219 = n24 & ~n113 ;
  assign n220 = n218 & n219 ;
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  assign n224 = ( n208 & ~n216 ) | ( n208 & n223 ) | ( ~n216 & n223 ) ;
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n54( .i (x10), .o (n54) );
  buffer buf_n57( .i (x11), .o (n57) );
  assign n227 = n54 & n57 ;
  assign n228 = ~n13 & n227 ;
  assign n229 = n162 & n228 ;
  buffer buf_n230( .i (n229), .o (n230) );
  assign n236 = n178 | n230 ;
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  assign n241 = n225 & ~n240 ;
  assign n242 = ( n198 & n226 ) | ( n198 & ~n241 ) | ( n226 & ~n241 ) ;
  assign n243 = n174 | n242 ;
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  assign n244 = n77 & n147 ;
  assign n245 = n221 & ~n244 ;
  assign n246 = n237 & n245 ;
  buffer buf_n247( .i (n246), .o (n247) );
  assign n249 = ~n8 & n12 ;
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n55( .i (n54), .o (n55) );
  assign n255 = ~n3 & n55 ;
  assign n256 = n250 & n255 ;
  buffer buf_n257( .i (n256), .o (n257) );
  assign n259 = n12 | n15 ;
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n10( .i (n9), .o (n10) );
  assign n262 = n4 & ~n10 ;
  assign n263 = ~n261 & n262 ;
  assign n264 = n257 | n263 ;
  buffer buf_n265( .i (n264), .o (n265) );
  assign n266 = n25 & n218 ;
  buffer buf_n267( .i (n266), .o (n267) );
  assign n268 = n147 | n213 ;
  assign n269 = n267 & ~n268 ;
  assign n270 = n265 & n269 ;
  buffer buf_n271( .i (n270), .o (n271) );
  assign n272 = n247 | n271 ;
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n183( .i (n182), .o (n183) );
  assign n275 = n4 & ~n260 ;
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  assign n278 = ~n9 & n68 ;
  buffer buf_n279( .i (n278), .o (n279) );
  assign n281 = n52 & n279 ;
  assign n282 = n276 & n281 ;
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n31( .i (x6), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  assign n290 = n34 & n279 ;
  assign n291 = n276 & n290 ;
  buffer buf_n292( .i (n291), .o (n292) );
  assign n294 = n283 | n292 ;
  buffer buf_n295( .i (n294), .o (n295) );
  assign n296 = n183 | n295 ;
  buffer buf_n297( .i (n296), .o (n297) );
  assign n298 = n273 | n297 ;
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  assign n299 = ~n79 & n265 ;
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  assign n300 = n78 & n179 ;
  assign n301 = ( n79 & n232 ) | ( n79 & n300 ) | ( n232 & n300 ) ;
  assign n302 = ( n99 & n299 ) | ( n99 & n301 ) | ( n299 & n301 ) ;
  assign n303 = n209 & n302 ;
  buffer buf_n304( .i (n303), .o (n304) );
  assign n305 = n157 & n163 ;
  buffer buf_n306( .i (n305), .o (n306) );
  assign n309 = n16 & ~n37 ;
  assign n310 = n16 | n32 ;
  assign n311 = ~n309 & n310 ;
  buffer buf_n312( .i (n311), .o (n312) );
  assign n315 = ( ~n15 & n73 ) | ( ~n15 & n81 ) | ( n73 & n81 ) ;
  buffer buf_n316( .i (n315), .o (n316) );
  assign n318 = n23 & ~n93 ;
  assign n319 = ( n24 & ~n316 ) | ( n24 & n318 ) | ( ~n316 & n318 ) ;
  buffer buf_n320( .i (n319), .o (n320) );
  assign n323 = n312 | n320 ;
  assign n324 = n306 & n323 ;
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n114( .i (n113), .o (n114) );
  assign n327 = n104 | n114 ;
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  assign n332 = n84 & n104 ;
  buffer buf_n333( .i (n332), .o (n333) );
  assign n334 = n328 & ~n333 ;
  assign n335 = ( ~n314 & n329 ) | ( ~n314 & n334 ) | ( n329 & n334 ) ;
  assign n336 = n325 & ~n335 ;
  buffer buf_n337( .i (n336), .o (n337) );
  assign n339 = ~n18 & n76 ;
  assign n340 = n150 | n339 ;
  buffer buf_n317( .i (n316), .o (n317) );
  assign n341 = n95 & n317 ;
  buffer buf_n342( .i (n341), .o (n342) );
  assign n346 = ~n340 & n342 ;
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n119( .i (n118), .o (n119) );
  assign n349 = ( n70 & n119 ) | ( n70 & ~n124 ) | ( n119 & ~n124 ) ;
  assign n350 = ( n119 & ~n124 ) | ( n119 & n188 ) | ( ~n124 & n188 ) ;
  assign n351 = ~n349 & n350 ;
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n26( .i (n25), .o (n26) );
  assign n355 = n26 & n164 ;
  assign n356 = n159 & n355 ;
  buffer buf_n357( .i (n356), .o (n357) );
  assign n358 = n353 | n357 ;
  assign n359 = ( n348 & n354 ) | ( n348 & n358 ) | ( n354 & n358 ) ;
  assign n360 = n337 | n359 ;
  assign n361 = n304 | n360 ;
  assign n362 = n298 | n361 ;
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  assign n363 = n313 & ~n333 ;
  assign n364 = n322 | n363 ;
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  assign n367 = n171 | n193 ;
  assign n368 = ( n194 & n366 ) | ( n194 & n367 ) | ( n366 & n367 ) ;
  assign n369 = n297 | n368 ;
  assign n370 = n274 | n369 ;
  assign n371 = ( ~n69 & n123 ) | ( ~n69 & n133 ) | ( n123 & n133 ) ;
  assign n372 = n117 & n127 ;
  assign n373 = ( n123 & n133 ) | ( n123 & ~n372 ) | ( n133 & ~n372 ) ;
  assign n374 = n371 & ~n373 ;
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n42( .i (x8), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n378( .i (n68), .o (n378) );
  assign n379 = n44 & n378 ;
  buffer buf_n380( .i (n379), .o (n380) );
  assign n382 = n6 & n380 ;
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  assign n384 = n18 & n60 ;
  assign n385 = n252 & n384 ;
  buffer buf_n386( .i (n385), .o (n386) );
  assign n387 = n383 & n386 ;
  assign n388 = n377 | n387 ;
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n326( .i (n325), .o (n326) );
  assign n391 = n109 & n326 ;
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  assign n393 = n90 & ~n389 ;
  assign n394 = ( n390 & n392 ) | ( n390 & ~n393 ) | ( n392 & ~n393 ) ;
  buffer buf_n338( .i (n337), .o (n338) );
  assign n395 = n347 & n357 ;
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  assign n398 = n338 | n397 ;
  assign n399 = n394 | n398 ;
  assign n400 = ( n97 & n214 ) | ( n97 & n328 ) | ( n214 & n328 ) ;
  assign n401 = n265 & ~n400 ;
  assign n402 = n94 & n103 ;
  assign n403 = n75 | n113 ;
  assign n404 = ( n114 & n402 ) | ( n114 & n403 ) | ( n402 & n403 ) ;
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  assign n407 = n179 & ~n405 ;
  assign n408 = ( n232 & ~n406 ) | ( n232 & n407 ) | ( ~n406 & n407 ) ;
  assign n409 = n401 | n408 ;
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  assign n412 = n304 & ~n411 ;
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n62( .i (x12), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  assign n413 = n65 & n114 ;
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  assign n419 = n271 | n417 ;
  assign n420 = n248 | n419 ;
  buffer buf_n421( .i (n420), .o (n421) );
  assign n422 = n412 | n421 ;
  buffer buf_n418( .i (n417), .o (n418) );
  assign n423 = n206 | n414 ;
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  assign n427 = ( n410 & n418 ) | ( n410 & n426 ) | ( n418 & n426 ) ;
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  assign n430 = n216 & n308 ;
  buffer buf_n431( .i (n430), .o (n431) );
  assign n432 = n396 | n431 ;
  assign n433 = n304 | n432 ;
  assign n434 = n428 | n433 ;
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n280( .i (n279), .o (n280) );
  assign n435 = n276 & n280 ;
  assign n436 = n47 & n435 ;
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  assign n439 = n295 | n438 ;
  assign n440 = n184 | n439 ;
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n381( .i (n380), .o (n381) );
  assign n443 = n277 & n381 ;
  buffer buf_n444( .i (n443), .o (n444) );
  assign n445 = n293 | n444 ;
  assign n446 = n183 | n445 ;
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n139( .i (x23), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  assign n447 = ~n114 & n142 ;
  buffer buf_n448( .i (n447), .o (n448) );
  assign n449 = n165 & n448 ;
  assign n450 = n160 & n449 ;
  buffer buf_n451( .i (n450), .o (n451) );
  assign n452 = ~n345 & n451 ;
  assign n453 = n446 | n452 ;
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  assign n455 = n326 & ~n331 ;
  buffer buf_n456( .i (n455), .o (n456) );
  assign n457 = n273 | n456 ;
  assign n458 = n454 | n457 ;
  assign n459 = n304 | n397 ;
  assign n460 = n348 & n451 ;
  buffer buf_n461( .i (n460), .o (n461) );
  assign n462 = n392 | n461 ;
  assign n463 = n459 | n462 ;
  assign n464 = ~n214 & n267 ;
  buffer buf_n258( .i (n257), .o (n258) );
  assign n465 = n147 & n167 ;
  assign n466 = n258 & ~n465 ;
  assign n467 = n464 & n466 ;
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  assign n471 = n225 & n235 ;
  assign n472 = n470 | n471 ;
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  assign n474 = n254 & n383 ;
  assign n475 = n444 | n474 ;
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  assign n480 = n203 & ~n329 ;
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  assign y0 = n243 ;
  assign y1 = n362 ;
  assign y2 = n370 ;
  assign y3 = n399 ;
  assign y4 = n422 ;
  assign y5 = n434 ;
  assign y6 = n442 ;
  assign y7 = n429 ;
  assign y8 = n458 ;
  assign y9 = n463 ;
  assign y10 = n473 ;
  assign y11 = n289 ;
  assign y12 = n479 ;
  assign y13 = n485 ;
endmodule
