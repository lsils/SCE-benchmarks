module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 ;
  buffer buf_n22( .i (x2), .o (n22) );
  buffer buf_n61( .i (x6), .o (n61) );
  assign n78 = n22 & n61 ;
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n41( .i (x4), .o (n41) );
  assign n85 = n2 | n41 ;
  buffer buf_n86( .i (n85), .o (n86) );
  assign n94 = n79 & ~n86 ;
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n42( .i (n41), .o (n42) );
  assign n99 = n3 & n42 ;
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n62( .i (n61), .o (n62) );
  assign n107 = n23 | n62 ;
  buffer buf_n108( .i (n107), .o (n108) );
  assign n114 = n100 & ~n108 ;
  assign n115 = n95 | n114 ;
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n12( .i (x1), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n70( .i (x7), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  assign n118 = n14 & ~n72 ;
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n30( .i (x3), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n51( .i (x5), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  assign n122 = ~n31 & n52 ;
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  assign n127 = ~n101 & n124 ;
  assign n128 = n120 & n127 ;
  assign n129 = n13 & n52 ;
  buffer buf_n130( .i (n129), .o (n130) );
  assign n134 = n100 & n130 ;
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n32( .i (n31), .o (n32) );
  assign n139 = n32 & n72 ;
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  assign n143 = n135 & n141 ;
  assign n144 = n128 | n143 ;
  assign n145 = ~n117 & n144 ;
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n63( .i (n62), .o (n63) );
  assign n148 = n32 | n63 ;
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n43( .i (n42), .o (n43) );
  assign n152 = n24 & ~n43 ;
  buffer buf_n153( .i (n152), .o (n153) );
  assign n155 = n149 & n153 ;
  buffer buf_n156( .i (n155), .o (n156) );
  assign n158 = n8 & ~n156 ;
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  assign n159 = ~n34 & n45 ;
  assign n160 = ( n46 & ~n82 ) | ( n46 & n159 ) | ( ~n82 & n159 ) ;
  assign n161 = n18 | n160 ;
  assign n162 = n158 & n161 ;
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  assign n164 = n110 & n132 ;
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n53( .i (n52), .o (n53) );
  assign n167 = n14 | n53 ;
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  assign n173 = ~n98 & n171 ;
  assign n174 = ~n166 & n173 ;
  assign n175 = n163 | n174 ;
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  assign n176 = n56 & n82 ;
  assign n177 = n16 & n45 ;
  assign n178 = ( n46 & ~n110 ) | ( n46 & n177 ) | ( ~n110 & n177 ) ;
  assign n179 = ~n176 & n178 ;
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n157( .i (n156), .o (n157) );
  assign n181 = ~n17 & n56 ;
  assign n182 = n8 & n181 ;
  assign n183 = ~n157 & n182 ;
  assign n184 = n180 | n183 ;
  assign n185 = ~n146 & n184 ;
  assign n186 = ( n147 & n175 ) | ( n147 & ~n185 ) | ( n175 & ~n185 ) ;
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n73( .i (n72), .o (n73) );
  assign n188 = n33 | n73 ;
  assign n189 = n168 | n188 ;
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  assign n193 = ( n17 & n56 ) | ( n17 & n141 ) | ( n56 & n141 ) ;
  assign n194 = n116 & ~n193 ;
  assign n195 = n43 & n53 ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n199 = ~n6 & n196 ;
  buffer buf_n64( .i (n63), .o (n64) );
  assign n200 = ( n64 & n73 ) | ( n64 & n80 ) | ( n73 & n80 ) ;
  buffer buf_n201( .i (n200), .o (n201) );
  assign n205 = n199 & ~n201 ;
  assign n206 = n190 & n205 ;
  assign n207 = ( n191 & n194 ) | ( n191 & n206 ) | ( n194 & n206 ) ;
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  assign n211 = n44 & n73 ;
  buffer buf_n212( .i (n211), .o (n212) );
  assign n214 = n17 | n212 ;
  assign n215 = ( n8 & n198 ) | ( n8 & n214 ) | ( n198 & n214 ) ;
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  assign n218 = ~n208 & n217 ;
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  assign n221 = n138 & n216 ;
  assign n222 = ~n208 & n221 ;
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  assign n225 = ( ~n187 & n220 ) | ( ~n187 & n224 ) | ( n220 & n224 ) ;
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  assign n226 = n81 & n140 ;
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  assign n229 = n171 & n228 ;
  assign n230 = n91 | n165 ;
  assign n231 = n229 | n230 ;
  assign n232 = ( n93 & ~n146 ) | ( n93 & n231 ) | ( ~n146 & n231 ) ;
  buffer buf_n233( .i (n232), .o (n233) );
  assign n234 = ~n219 & n233 ;
  assign n235 = ~n223 & n233 ;
  assign n236 = ( n187 & n234 ) | ( n187 & n235 ) | ( n234 & n235 ) ;
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n74( .i (n73), .o (n74) );
  assign n237 = n65 & ~n74 ;
  assign n238 = n169 | n237 ;
  buffer buf_n239( .i (n72), .o (n239) );
  assign n240 = n15 | n239 ;
  buffer buf_n241( .i (n240), .o (n241) );
  assign n243 = n110 & n241 ;
  buffer buf_n25( .i (n24), .o (n25) );
  assign n244 = n25 & n54 ;
  buffer buf_n245( .i (n244), .o (n245) );
  assign n247 = n241 | n245 ;
  assign n248 = ( n238 & n243 ) | ( n238 & ~n247 ) | ( n243 & ~n247 ) ;
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n172( .i (n171), .o (n172) );
  assign n251 = n105 & ~n172 ;
  assign n252 = n250 & n251 ;
  assign n253 = ~n131 & n168 ;
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  assign n258 = ~n9 & n48 ;
  assign n259 = n204 & n258 ;
  assign n260 = n257 & n259 ;
  assign n261 = n252 | n260 ;
  assign n262 = n210 | n261 ;
  assign n263 = n187 | n262 ;
  buffer buf_n142( .i (n141), .o (n142) );
  assign n264 = n116 & ~n142 ;
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n192( .i (n191), .o (n192) );
  assign n269 = n192 & ~n256 ;
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n106( .i (n105), .o (n106) );
  assign n272 = n34 & n81 ;
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  assign n277 = n106 & n276 ;
  assign n278 = ~n270 & n277 ;
  assign n279 = ( n268 & ~n271 ) | ( n268 & n278 ) | ( ~n271 & n278 ) ;
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  assign n280 = ~n32 & n63 ;
  buffer buf_n281( .i (n280), .o (n281) );
  assign n284 = ( ~n65 & n149 ) | ( ~n65 & n281 ) | ( n149 & n281 ) ;
  buffer buf_n285( .i (n284), .o (n285) );
  assign n286 = n126 | n285 ;
  assign n287 = n47 & n254 ;
  assign n288 = ( n48 & ~n286 ) | ( n48 & n287 ) | ( ~n286 & n287 ) ;
  assign n289 = n13 & ~n42 ;
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n35( .i (n34), .o (n35) );
  assign n294 = n27 | n35 ;
  assign n295 = n293 & ~n294 ;
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  assign n296 = ~n26 & n55 ;
  buffer buf_n297( .i (n296), .o (n297) );
  assign n299 = ( n57 & ~n151 ) | ( n57 & n297 ) | ( ~n151 & n297 ) ;
  buffer buf_n28( .i (n27), .o (n28) );
  assign n300 = n28 & ~n57 ;
  assign n301 = ( ~n295 & n299 ) | ( ~n295 & n300 ) | ( n299 & n300 ) ;
  assign n302 = ~n288 & n301 ;
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  assign n303 = n57 & ~n76 ;
  buffer buf_n304( .i (n303), .o (n304) );
  assign n305 = n180 & n304 ;
  assign n306 = n302 | n305 ;
  assign n307 = n23 & n71 ;
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  assign n312 = n46 & ~n169 ;
  assign n313 = n290 & ~n308 ;
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  assign n316 = ( ~n311 & n312 ) | ( ~n311 & n315 ) | ( n312 & n315 ) ;
  assign n317 = n45 | n124 ;
  buffer buf_n318( .i (n317), .o (n318) );
  assign n320 = n202 & n318 ;
  assign n321 = n316 & n320 ;
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n10( .i (n9), .o (n10) );
  assign n324 = n44 & n64 ;
  buffer buf_n325( .i (n324), .o (n325) );
  assign n327 = n310 & n325 ;
  assign n328 = n254 & n327 ;
  buffer buf_n329( .i (n328), .o (n329) );
  assign n330 = n10 & ~n329 ;
  assign n331 = ~n322 & n330 ;
  assign n332 = ~n306 & n331 ;
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n333( .i (n16), .o (n333) );
  assign n334 = n154 | n333 ;
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n83( .i (n82), .o (n83) );
  assign n337 = ( n83 & ~n198 ) | ( n83 & n273 ) | ( ~n198 & n273 ) ;
  assign n338 = n335 & n337 ;
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n77( .i (n76), .o (n77) );
  assign n339 = ~n43 & n63 ;
  buffer buf_n340( .i (n339), .o (n340) );
  assign n344 = ~n124 & n340 ;
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  assign n347 = ( n68 & n77 ) | ( n68 & n346 ) | ( n77 & n346 ) ;
  assign n348 = ( n336 & n338 ) | ( n336 & n347 ) | ( n338 & n347 ) ;
  assign n349 = n28 & ~n126 ;
  buffer buf_n121( .i (n120), .o (n121) );
  assign n350 = n47 & n121 ;
  assign n351 = ~n15 & n239 ;
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  assign n355 = ~n47 & n353 ;
  assign n356 = ( n349 & n350 ) | ( n349 & n355 ) | ( n350 & n355 ) ;
  buffer buf_n357( .i (n62), .o (n357) );
  assign n358 = n24 & ~n357 ;
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n362( .i (n123), .o (n362) );
  assign n363 = n359 & n362 ;
  assign n364 = n314 & n363 ;
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n213( .i (n212), .o (n213) );
  assign n367 = n66 | n333 ;
  assign n368 = ( n67 & n213 ) | ( n67 & n367 ) | ( n213 & n367 ) ;
  assign n369 = n365 | n368 ;
  assign n370 = n356 | n369 ;
  assign n371 = ~n348 & n370 ;
  buffer buf_n111( .i (n110), .o (n111) );
  assign n372 = ~n111 & n126 ;
  assign n373 = n9 & ~n372 ;
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n374( .i (n55), .o (n374) );
  assign n375 = n27 | n374 ;
  assign n376 = n142 & ~n375 ;
  assign n377 = n343 & n376 ;
  assign n378 = n373 | n377 ;
  buffer buf_n49( .i (n48), .o (n49) );
  assign n379 = n111 & ~n227 ;
  assign n380 = ~n55 & n359 ;
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n133( .i (n132), .o (n133) );
  assign n383 = n133 | n381 ;
  assign n384 = ( ~n379 & n382 ) | ( ~n379 & n383 ) | ( n382 & n383 ) ;
  assign n385 = ~n49 & n384 ;
  assign n386 = n378 | n385 ;
  assign n387 = n371 | n386 ;
  assign n388 = ~n332 & n387 ;
  assign n389 = n279 | n388 ;
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n84( .i (n83), .o (n84) );
  assign n390 = ( n19 & ~n84 ) | ( n19 & n191 ) | ( ~n84 & n191 ) ;
  assign n391 = n329 | n390 ;
  assign n392 = n163 & ~n391 ;
  assign n393 = ~n323 & n392 ;
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n326( .i (n325), .o (n326) );
  assign n394 = n121 & ~n326 ;
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n395( .i (n7), .o (n395) );
  assign n396 = n361 | n395 ;
  assign n397 = ( ~n104 & n394 ) | ( ~n104 & n396 ) | ( n394 & n396 ) ;
  assign n398 = ~n59 & n397 ;
  assign n399 = n88 & ~n119 ;
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  assign n403 = n37 & n343 ;
  assign n404 = n402 & n403 ;
  assign n405 = ( n39 & n398 ) | ( n39 & n404 ) | ( n398 & n404 ) ;
  assign n406 = ~n345 & n395 ;
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n409( .i (n44), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  assign n412 = n142 & ~n411 ;
  assign n413 = n298 & n412 ;
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n246( .i (n245), .o (n246) );
  assign n414 = ~n242 & n246 ;
  assign n415 = ~n319 & n414 ;
  assign n416 = n413 | n415 ;
  buffer buf_n354( .i (n353), .o (n354) );
  assign n417 = ~n75 & n410 ;
  assign n418 = ( n27 & ~n75 ) | ( n27 & n410 ) | ( ~n75 & n410 ) ;
  assign n419 = ( ~n126 & n417 ) | ( ~n126 & n418 ) | ( n417 & n418 ) ;
  buffer buf_n420( .i (n26), .o (n420) );
  assign n421 = ( n75 & n333 ) | ( n75 & ~n420 ) | ( n333 & ~n420 ) ;
  buffer buf_n422( .i (n125), .o (n422) );
  assign n423 = ( n242 & n421 ) | ( n242 & n422 ) | ( n421 & n422 ) ;
  assign n424 = ( n354 & n419 ) | ( n354 & n423 ) | ( n419 & n423 ) ;
  assign n425 = ~n407 & n424 ;
  assign n426 = ( ~n408 & n416 ) | ( ~n408 & n425 ) | ( n416 & n425 ) ;
  assign n427 = n405 | n426 ;
  assign n428 = n393 | n427 ;
  assign n429 = n7 & n212 ;
  buffer buf_n430( .i (n74), .o (n430) );
  assign n431 = n89 | n430 ;
  assign n432 = ~n429 & n431 ;
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  assign n435 = n283 & n297 ;
  assign n436 = n274 | n435 ;
  assign n437 = n20 & n436 ;
  assign n438 = n36 & ~n111 ;
  assign n439 = ~n171 & n438 ;
  assign n440 = ~n433 & n439 ;
  assign n441 = ( ~n434 & n437 ) | ( ~n434 & n440 ) | ( n437 & n440 ) ;
  buffer buf_n366( .i (n365), .o (n366) );
  assign n442 = ~n36 & n213 ;
  assign n443 = n382 & n442 ;
  assign n444 = n366 | n443 ;
  buffer buf_n445( .i (n374), .o (n445) );
  assign n446 = n103 & ~n445 ;
  assign n447 = ~n76 & n170 ;
  assign n448 = ( n354 & ~n446 ) | ( n354 & n447 ) | ( ~n446 & n447 ) ;
  assign n449 = ~n374 & n430 ;
  buffer buf_n450( .i (n449), .o (n450) );
  assign n453 = n285 & ~n400 ;
  assign n454 = ( n28 & ~n76 ) | ( n28 & n445 ) | ( ~n76 & n445 ) ;
  assign n455 = ( n450 & n453 ) | ( n450 & n454 ) | ( n453 & n454 ) ;
  assign n456 = ~n448 & n455 ;
  assign n457 = n444 | n456 ;
  assign n458 = n441 | n457 ;
  assign n459 = n38 & n249 ;
  assign n460 = ( ~n19 & n37 ) | ( ~n19 & n104 ) | ( n37 & n104 ) ;
  assign n461 = n249 | n460 ;
  assign n462 = ( n106 & n459 ) | ( n106 & ~n461 ) | ( n459 & ~n461 ) ;
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  assign n463 = n352 | n420 ;
  assign n464 = n65 | n409 ;
  assign n465 = ( ~n120 & n410 ) | ( ~n120 & n464 ) | ( n410 & n464 ) ;
  assign n466 = ~n16 & n26 ;
  assign n467 = ( ~n212 & n420 ) | ( ~n212 & n466 ) | ( n420 & n466 ) ;
  assign n468 = ( ~n463 & n465 ) | ( ~n463 & n467 ) | ( n465 & n467 ) ;
  assign n469 = n395 & n422 ;
  assign n470 = ~n468 & n469 ;
  buffer buf_n471( .i (n470), .o (n471) );
  assign n472 = n452 | n471 ;
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  assign n473 = ( n19 & ~n58 ) | ( n19 & n77 ) | ( ~n58 & n77 ) ;
  assign n474 = ( n113 & n304 ) | ( n113 & ~n473 ) | ( n304 & ~n473 ) ;
  assign n475 = n471 | n474 ;
  assign n476 = ( n462 & n472 ) | ( n462 & n475 ) | ( n472 & n475 ) ;
  assign n477 = n458 | n476 ;
  assign n478 = n428 | n477 ;
  assign y0 = n225 ;
  assign y1 = n236 ;
  assign y2 = n263 ;
  assign y3 = n389 ;
  assign y4 = n478 ;
endmodule
