module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n204 , n205 , n207 , n208 , n209 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n258 , n259 , n260 , n261 , n262 , n263 , n265 , n266 , n267 , n268 , n269 , n270 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n348 , n349 , n350 , n351 , n352 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n519 , n520 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 ;
  buffer buf_n613( .i (x48), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n624( .i (x49), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  assign n634 = n615 | n626 ;
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n28( .i (x1), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n601( .i (x47), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  assign n640 = n34 | n607 ;
  buffer buf_n641( .i (n640), .o (n641) );
  assign n642 = n639 | n641 ;
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n39( .i (x2), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n50( .i (x3), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n61( .i (x4), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  assign n685 = n52 | n63 ;
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  assign n688 = n44 & n687 ;
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n272( .i (x22), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n136( .i (x11), .o (n136) );
  assign n734 = ~n2 & n136 ;
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  buffer buf_n738( .i (n737), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  assign n742 = ~n279 & n740 ;
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n608( .i (n607), .o (n608) );
  assign n744 = ~n608 & n638 ;
  buffer buf_n745( .i (n744), .o (n745) );
  assign n761 = n743 & n745 ;
  buffer buf_n315( .i (x27), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n324( .i (x28), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n332( .i (x29), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  assign n762 = n330 | n338 ;
  assign n763 = n322 & n762 ;
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  assign n765 = n7 | n277 ;
  buffer buf_n766( .i (n765), .o (n766) );
  assign n770 = n143 | n766 ;
  buffer buf_n771( .i (n770), .o (n771) );
  assign n775 = n764 & ~n771 ;
  assign n776 = n761 | n775 ;
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  assign n777 = ~n56 & n330 ;
  buffer buf_n45( .i (n44), .o (n45) );
  assign n778 = ~n45 & n321 ;
  assign n779 = n777 | n778 ;
  buffer buf_n283( .i (x23), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  assign n780 = n289 & ~n607 ;
  buffer buf_n307( .i (x26), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  assign n781 = ~n34 & n313 ;
  assign n782 = n780 | n781 ;
  assign n783 = n779 | n782 ;
  buffer buf_n299( .i (x25), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  assign n784 = n305 & ~n630 ;
  buffer buf_n291( .i (x24), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  assign n785 = n297 & ~n619 ;
  assign n786 = n784 | n785 ;
  buffer buf_n73( .i (x5), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n340( .i (x30), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  assign n787 = ~n79 & n346 ;
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  assign n788 = ~n67 & n338 ;
  assign n789 = n787 | n788 ;
  assign n790 = n786 | n789 ;
  assign n791 = n783 | n790 ;
  assign n792 = n769 & n791 ;
  assign n793 = n776 | n792 ;
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  assign n833 = n321 & ~n330 ;
  assign n834 = ~n321 & n330 ;
  assign n835 = n833 | n834 ;
  buffer buf_n836( .i (n835), .o (n836) );
  assign n837 = n338 | n346 ;
  assign n838 = n338 & n346 ;
  assign n839 = n837 & ~n838 ;
  buffer buf_n840( .i (n839), .o (n840) );
  assign n841 = n836 | n840 ;
  assign n842 = n836 & n840 ;
  assign n843 = n841 & ~n842 ;
  buffer buf_n844( .i (n843), .o (n844) );
  assign n845 = n289 & ~n297 ;
  assign n846 = ~n289 & n297 ;
  assign n847 = n845 | n846 ;
  buffer buf_n848( .i (n847), .o (n848) );
  assign n849 = n305 | n313 ;
  assign n850 = n305 & n313 ;
  assign n851 = n849 & ~n850 ;
  buffer buf_n852( .i (n851), .o (n852) );
  assign n853 = n848 | n852 ;
  assign n854 = n848 & n852 ;
  assign n855 = n853 & ~n854 ;
  buffer buf_n856( .i (n855), .o (n856) );
  assign n857 = n844 & n856 ;
  assign n858 = n844 | n856 ;
  assign n859 = ~n857 & n858 ;
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  buffer buf_n886( .i (n885), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  assign n897 = ~n48 & n70 ;
  assign n898 = n48 & ~n70 ;
  assign n899 = n897 | n898 ;
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  assign n901 = n59 & n82 ;
  assign n902 = n59 | n82 ;
  assign n903 = ~n901 & n902 ;
  buffer buf_n904( .i (n903), .o (n904) );
  assign n905 = ~n900 & n904 ;
  assign n906 = n900 & ~n904 ;
  assign n907 = n905 | n906 ;
  buffer buf_n908( .i (n907), .o (n908) );
  assign n909 = n616 & n627 ;
  assign n910 = n635 & ~n909 ;
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n35( .i (n34), .o (n35) );
  assign n916 = n35 & n608 ;
  assign n917 = n641 & ~n916 ;
  buffer buf_n918( .i (n917), .o (n918) );
  assign n919 = ~n915 & n918 ;
  assign n920 = n915 & ~n918 ;
  assign n921 = n919 | n920 ;
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  assign n925 = n908 | n924 ;
  assign n926 = n908 & n924 ;
  assign n927 = n925 & ~n926 ;
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  assign n962 = n2 & n136 ;
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n365( .i (x33), .o (n365) );
  buffer buf_n522( .i (x44), .o (n522) );
  assign n965 = n365 & n522 ;
  buffer buf_n966( .i (n965), .o (n966) );
  assign n974 = n963 & ~n966 ;
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n584( .i (x46), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  assign n980 = n3 | n585 ;
  buffer buf_n981( .i (n980), .o (n981) );
  assign n984 = n525 | n981 ;
  buffer buf_n985( .i (n984), .o (n985) );
  assign n987 = n337 & n985 ;
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n519( .i (x43), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  assign n988 = n366 | n520 ;
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  assign n992 = n319 & ~n990 ;
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n378( .i (x34), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  assign n993 = ~n368 & n381 ;
  assign n994 = n327 & n368 ;
  assign n995 = n993 | n994 ;
  assign n996 = n992 | n995 ;
  assign n997 = n987 | n996 ;
  assign n998 = ~n978 & n997 ;
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n348( .i (x31), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  assign n1000 = n352 & ~n975 ;
  buffer buf_n1001( .i (n1000), .o (n1001) );
  assign n1002 = ~n986 & n1001 ;
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  assign n1005 = n999 | n1004 ;
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n183( .i (x15), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n192( .i (x16), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  assign n1007 = n190 | n199 ;
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  assign n1011 = ~n1006 & n1010 ;
  assign n1012 = n274 & n735 ;
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n964( .i (n963), .o (n964) );
  assign n1017 = n3 & n273 ;
  assign n1018 = n367 & n1017 ;
  assign n1019 = n964 | n1018 ;
  buffer buf_n1020( .i (n1019), .o (n1020) );
  assign n1024 = n277 & n1020 ;
  buffer buf_n1025( .i (n1024), .o (n1025) );
  assign n1026 = n1016 | n1025 ;
  buffer buf_n1027( .i (n1026), .o (n1027) );
  assign n1028 = ~n70 & n1027 ;
  assign n1029 = ~n5 & n368 ;
  assign n1030 = n1013 | n1029 ;
  assign n1031 = n1020 | n1030 ;
  buffer buf_n1032( .i (n1031), .o (n1032) );
  assign n1033 = n68 & ~n1032 ;
  assign n1034 = ~n275 & n964 ;
  buffer buf_n1035( .i (n1034), .o (n1035) );
  assign n1036 = n41 | n367 ;
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n1039( .i (n367), .o (n1039) );
  assign n1040 = n76 & n1039 ;
  assign n1041 = n1037 & ~n1040 ;
  assign n1042 = n1035 & ~n1041 ;
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  assign n1045 = n1033 | n1044 ;
  buffer buf_n1046( .i (n1045), .o (n1046) );
  assign n1047 = n1028 | n1046 ;
  buffer buf_n1048( .i (n1047), .o (n1048) );
  assign n1051 = n1011 & n1048 ;
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n204( .i (x17), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n207( .i (x18), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  assign n1058 = n205 | n208 ;
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  buffer buf_n1061( .i (n1060), .o (n1061) );
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  assign n1069 = ~n1006 & n1067 ;
  buffer buf_n1070( .i (n1069), .o (n1070) );
  assign n1071 = n1049 | n1070 ;
  assign n1072 = ~n1052 & n1071 ;
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  assign n1077 = n57 | n1016 ;
  assign n1078 = n57 & n1032 ;
  assign n1079 = n1077 & ~n1078 ;
  buffer buf_n1080( .i (n366), .o (n1080) );
  assign n1081 = n30 & ~n1080 ;
  buffer buf_n1082( .i (n1081), .o (n1082) );
  assign n1083 = n64 & n1039 ;
  assign n1084 = n1082 | n1083 ;
  assign n1085 = n1035 & n1084 ;
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  assign n1088 = n54 & n65 ;
  assign n1089 = n687 & ~n1088 ;
  buffer buf_n1090( .i (n1089), .o (n1090) );
  assign n1094 = n1025 & n1090 ;
  assign n1095 = n1087 | n1094 ;
  assign n1096 = n1079 | n1095 ;
  buffer buf_n1097( .i (n1096), .o (n1097) );
  assign n1100 = n329 & n985 ;
  buffer buf_n354( .i (x32), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  assign n1101 = n357 | n1039 ;
  assign n1102 = ~n318 & n1039 ;
  assign n1103 = n1101 & ~n1102 ;
  assign n1104 = n311 & ~n990 ;
  assign n1105 = n1103 | n1104 ;
  assign n1106 = n1100 | n1105 ;
  assign n1107 = ~n978 & n1106 ;
  assign n1108 = n1003 | n1107 ;
  buffer buf_n1109( .i (n1108), .o (n1109) );
  assign n1111 = n1009 & ~n1109 ;
  assign n1112 = n1097 & n1111 ;
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  buffer buf_n1110( .i (n1109), .o (n1110) );
  assign n1122 = n1067 & ~n1110 ;
  assign n1123 = n1098 | n1122 ;
  assign n1124 = ~n1113 & n1123 ;
  buffer buf_n1125( .i (n1124), .o (n1125) );
  assign n1126 = n46 & ~n1032 ;
  assign n1127 = ~n46 & n1016 ;
  assign n1128 = n1126 | n1127 ;
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  assign n1129 = n274 | n1080 ;
  buffer buf_n1130( .i (n1129), .o (n1130) );
  assign n1132 = n628 | n1130 ;
  assign n1133 = ~n274 & n1080 ;
  buffer buf_n1134( .i (n1133), .o (n1134) );
  assign n1142 = ~n54 & n1134 ;
  assign n1143 = n1132 & ~n1142 ;
  assign n1144 = n43 | n686 ;
  assign n1145 = n277 & n1144 ;
  assign n1146 = n1143 & ~n1145 ;
  assign n1147 = n1022 & ~n1146 ;
  buffer buf_n1148( .i (n1147), .o (n1148) );
  assign n1149 = n1128 | n1148 ;
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1153( .i (n1080), .o (n1153) );
  assign n1154 = ~n310 & n1153 ;
  assign n1155 = n76 | n1153 ;
  assign n1156 = ~n1154 & n1155 ;
  assign n1157 = n303 & ~n990 ;
  assign n1158 = n1156 | n1157 ;
  buffer buf_n982( .i (n981), .o (n982) );
  assign n1159 = n352 | n982 ;
  assign n1160 = ~n319 & n982 ;
  assign n1161 = n1159 & ~n1160 ;
  assign n1162 = n1158 | n1161 ;
  assign n1163 = ~n978 & n1162 ;
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  assign n1166 = n1009 & ~n1165 ;
  assign n1167 = n1150 & n1166 ;
  buffer buf_n1168( .i (n1167), .o (n1168) );
  assign n1170 = n1066 & ~n1165 ;
  assign n1171 = n1150 | n1170 ;
  buffer buf_n1172( .i (n1171), .o (n1172) );
  assign n1173 = ~n1168 & n1172 ;
  buffer buf_n1174( .i (n1173), .o (n1174) );
  assign n1175 = n1125 & n1174 ;
  buffer buf_n1176( .i (n1175), .o (n1176) );
  assign n1177 = n1074 & n1176 ;
  buffer buf_n1178( .i (n1177), .o (n1178) );
  assign n1179 = n345 & n985 ;
  buffer buf_n1180( .i (n989), .o (n1180) );
  assign n1181 = n328 & ~n1180 ;
  assign n1182 = n335 & n1153 ;
  buffer buf_n389( .i (x35), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  assign n1183 = n392 & ~n1153 ;
  assign n1184 = n1182 | n1183 ;
  assign n1185 = n1181 | n1184 ;
  assign n1186 = n1179 | n1185 ;
  buffer buf_n1187( .i (n977), .o (n1187) );
  assign n1188 = n1186 & ~n1187 ;
  buffer buf_n1189( .i (n1188), .o (n1189) );
  assign n1190 = n1004 | n1189 ;
  buffer buf_n1191( .i (n1190), .o (n1191) );
  assign n1193 = n1010 & ~n1191 ;
  buffer buf_n1194( .i (n366), .o (n1194) );
  assign n1195 = n52 | n1194 ;
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1194), .o (n1197) );
  assign n1198 = n357 & n1197 ;
  assign n1199 = n1196 & ~n1198 ;
  assign n1200 = n1035 & ~n1199 ;
  buffer buf_n1201( .i (n1200), .o (n1201) );
  assign n1202 = ~n79 & n1015 ;
  assign n1203 = n1201 | n1202 ;
  buffer buf_n1204( .i (n1203), .o (n1204) );
  assign n1205 = ~n1025 & n1032 ;
  assign n1206 = n81 & ~n1205 ;
  assign n1207 = n1204 | n1206 ;
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  assign n1212 = n1193 & n1209 ;
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  assign n1219 = n1068 & ~n1192 ;
  assign n1220 = n1210 | n1219 ;
  assign n1221 = ~n1213 & n1220 ;
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  assign n1226 = n1178 & n1225 ;
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n1228( .i (n1227), .o (n1228) );
  buffer buf_n1229( .i (n1228), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  assign n1232 = ~n5 & n275 ;
  buffer buf_n1233( .i (n1232), .o (n1233) );
  assign n1234 = n1020 | n1233 ;
  buffer buf_n1235( .i (n1234), .o (n1235) );
  assign n1236 = n608 & n1235 ;
  buffer buf_n1237( .i (n607), .o (n1237) );
  assign n1238 = n1016 | n1237 ;
  assign n1239 = ~n1236 & n1238 ;
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1135( .i (n1134), .o (n1135) );
  assign n1240 = ~n618 & n1135 ;
  buffer buf_n160( .i (x13), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  assign n1241 = n165 & ~n1131 ;
  assign n1242 = n1240 | n1241 ;
  assign n1243 = n606 | n636 ;
  assign n1244 = n278 & n1243 ;
  assign n1245 = n1242 | n1244 ;
  assign n1246 = n1023 & n1245 ;
  assign n1247 = n1239 | n1246 ;
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n586( .i (n585), .o (n586) );
  assign n1252 = n524 | n586 ;
  assign n1253 = ~n5 & n1252 ;
  buffer buf_n1254( .i (n1253), .o (n1254) );
  buffer buf_n1255( .i (n1254), .o (n1255) );
  assign n1256 = n1001 & n1255 ;
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n979( .i (n978), .o (n979) );
  assign n1259 = n289 & ~n1255 ;
  buffer buf_n265( .i (x21), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  assign n1260 = n268 & n1197 ;
  assign n1261 = n1082 | n1260 ;
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n258( .i (x20), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n991( .i (n990), .o (n991) );
  assign n1263 = n263 & ~n991 ;
  assign n1264 = n1262 | n1263 ;
  assign n1265 = n1259 | n1264 ;
  assign n1266 = ~n979 & n1265 ;
  assign n1267 = n1258 | n1266 ;
  buffer buf_n1268( .i (n1267), .o (n1268) );
  assign n1269 = n1010 & ~n1268 ;
  assign n1270 = n1249 & n1269 ;
  buffer buf_n1271( .i (n1270), .o (n1271) );
  assign n1273 = n1067 & ~n1268 ;
  assign n1274 = n1249 | n1273 ;
  buffer buf_n1275( .i (n1274), .o (n1275) );
  assign n1276 = ~n1271 & n1275 ;
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n1278( .i (n1015), .o (n1278) );
  assign n1279 = n620 | n1278 ;
  assign n1280 = n620 & n1235 ;
  assign n1281 = n1279 & ~n1280 ;
  assign n1282 = ~n629 & n1135 ;
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n172( .i (x14), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  assign n1283 = n175 & ~n275 ;
  buffer buf_n1284( .i (n1283), .o (n1284) );
  assign n1288 = ~n370 & n1284 ;
  assign n1289 = n1282 | n1288 ;
  assign n1290 = n278 & n911 ;
  assign n1291 = n1289 | n1290 ;
  assign n1292 = n1023 & n1291 ;
  assign n1293 = n1281 | n1292 ;
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  assign n1298 = n297 & ~n1255 ;
  buffer buf_n1038( .i (n1037), .o (n1038) );
  assign n1299 = ~n287 & n369 ;
  assign n1300 = n1038 & ~n1299 ;
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  assign n1301 = n270 & ~n991 ;
  assign n1302 = n1300 | n1301 ;
  assign n1303 = n1298 | n1302 ;
  assign n1304 = ~n979 & n1303 ;
  assign n1305 = n1258 | n1304 ;
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1066), .o (n1307) );
  assign n1308 = ~n1306 & n1307 ;
  buffer buf_n1309( .i (n1308), .o (n1309) );
  assign n1310 = n1296 | n1309 ;
  assign n1311 = n1010 & ~n1306 ;
  assign n1312 = n1295 & n1311 ;
  buffer buf_n1313( .i (n1312), .o (n1313) );
  assign n1314 = n1310 & ~n1313 ;
  buffer buf_n1315( .i (n1314), .o (n1315) );
  assign n1316 = n1277 & n1315 ;
  buffer buf_n1317( .i (n1316), .o (n1317) );
  assign n1318 = ~n35 & n1278 ;
  assign n1319 = n618 | n1131 ;
  assign n1320 = ~n44 & n1135 ;
  assign n1321 = n1319 & ~n1320 ;
  assign n1322 = n1022 & ~n1321 ;
  assign n1323 = n1318 | n1322 ;
  buffer buf_n36( .i (n35), .o (n36) );
  assign n1324 = ~n1025 & n1235 ;
  assign n1325 = n36 & ~n1324 ;
  assign n1326 = n1323 | n1325 ;
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  assign n1331 = n313 & ~n1255 ;
  assign n1332 = n65 | n369 ;
  assign n1333 = ~n303 & n369 ;
  assign n1334 = n1332 & ~n1333 ;
  assign n1335 = n296 & ~n991 ;
  assign n1336 = n1334 | n1335 ;
  assign n1337 = n1331 | n1336 ;
  assign n1338 = ~n979 & n1337 ;
  assign n1339 = n1258 | n1338 ;
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1342( .i (n1009), .o (n1342) );
  assign n1343 = ~n1340 & n1342 ;
  assign n1344 = n1328 & n1343 ;
  buffer buf_n1345( .i (n1344), .o (n1345) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  assign n1349 = n1068 & ~n1341 ;
  assign n1350 = n1329 | n1349 ;
  assign n1351 = ~n1345 & n1350 ;
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  assign n1362 = ~n294 & n1197 ;
  assign n1363 = n1196 & ~n1362 ;
  assign n1364 = n287 & ~n1180 ;
  assign n1365 = n1363 | n1364 ;
  assign n1366 = n304 & ~n1254 ;
  assign n1367 = n1365 | n1366 ;
  assign n1368 = ~n1187 & n1367 ;
  buffer buf_n1369( .i (n1368), .o (n1369) );
  assign n1370 = n1258 | n1369 ;
  buffer buf_n1371( .i (n1370), .o (n1371) );
  assign n1372 = n1307 & ~n1371 ;
  buffer buf_n631( .i (n630), .o (n631) );
  assign n1373 = n631 & ~n1235 ;
  buffer buf_n1374( .i (n1134), .o (n1374) );
  assign n1375 = n33 & n1374 ;
  assign n1376 = n606 & ~n1131 ;
  assign n1377 = n1375 | n1376 ;
  assign n1378 = n1022 & n1377 ;
  assign n1379 = n1373 | n1378 ;
  buffer buf_n1380( .i (n1379), .o (n1380) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  assign n1381 = ~n633 & n1027 ;
  assign n1382 = n1380 | n1381 ;
  buffer buf_n1383( .i (n1382), .o (n1383) );
  assign n1385 = n1372 | n1383 ;
  buffer buf_n1386( .i (n1385), .o (n1386) );
  assign n1389 = n1342 & ~n1371 ;
  assign n1390 = n1383 & n1389 ;
  buffer buf_n1391( .i (n1390), .o (n1391) );
  assign n1397 = n1386 & ~n1391 ;
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  assign n1400 = n1353 & n1399 ;
  assign n1401 = n1317 & n1400 ;
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  assign n1408 = n1231 & n1407 ;
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  buffer buf_n1414( .i (n1413), .o (n1414) );
  buffer buf_n1415( .i (n1414), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  assign n1434 = n1275 & n1313 ;
  assign n1435 = n1272 | n1434 ;
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1392( .i (n1391), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1346( .i (n1345), .o (n1346) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  assign n1439 = n1347 & n1388 ;
  assign n1440 = n1394 | n1439 ;
  assign n1441 = n1317 & n1440 ;
  assign n1442 = n1438 | n1441 ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  assign n1448 = n1178 & n1218 ;
  buffer buf_n1053( .i (n1052), .o (n1053) );
  buffer buf_n1054( .i (n1053), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  assign n1449 = n1055 & n1176 ;
  buffer buf_n1169( .i (n1168), .o (n1169) );
  assign n1450 = n1113 & n1172 ;
  assign n1451 = n1169 | n1450 ;
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  assign n1455 = n1449 | n1454 ;
  buffer buf_n1456( .i (n1455), .o (n1456) );
  assign n1457 = n1448 | n1456 ;
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  assign n1461 = n1406 & n1460 ;
  assign n1462 = n1447 | n1461 ;
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n211( .i (x19), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n474( .i (x42), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  assign n1488 = n220 & n483 ;
  buffer buf_n1489( .i (n1488), .o (n1489) );
  assign n1525 = ~n773 & n1489 ;
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  assign n1536 = n1050 & n1527 ;
  buffer buf_n1537( .i (n1536), .o (n1537) );
  assign n1538 = n1073 | n1537 ;
  assign n1539 = n1073 & n1537 ;
  assign n1540 = n1538 & ~n1539 ;
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n448( .i (x41), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  assign n1545 = n1211 & n1527 ;
  buffer buf_n1546( .i (n1545), .o (n1546) );
  assign n1547 = n1222 & n1546 ;
  assign n1548 = n1222 | n1546 ;
  assign n1549 = ~n1547 & n1548 ;
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  assign n1553 = n469 & n1552 ;
  assign n1554 = ~n1544 & n1553 ;
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n1556( .i (n1555), .o (n1556) );
  buffer buf_n1557( .i (n1556), .o (n1557) );
  buffer buf_n1558( .i (n1557), .o (n1558) );
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n1575( .i (n1574), .o (n1575) );
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n774( .i (n773), .o (n774) );
  assign n1583 = n534 & ~n774 ;
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  assign n1606 = n760 & ~n1594 ;
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  buffer buf_n1534( .i (n1533), .o (n1534) );
  buffer buf_n1535( .i (n1534), .o (n1535) );
  assign n1607 = n1458 & ~n1535 ;
  buffer buf_n1608( .i (n1607), .o (n1608) );
  assign n1616 = ~n26 & n1608 ;
  assign n1617 = n1606 | n1616 ;
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n1621( .i (n1620), .o (n1621) );
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n1633( .i (n1632), .o (n1633) );
  buffer buf_n1634( .i (n1633), .o (n1634) );
  buffer buf_n1635( .i (n1634), .o (n1635) );
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n1637( .i (n1636), .o (n1637) );
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  assign n1643 = ~n469 & n1552 ;
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  assign n1644 = ~n599 & n1585 ;
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  assign n1658 = n1643 | n1650 ;
  assign n1659 = n469 & ~n1552 ;
  buffer buf_n1660( .i (n1659), .o (n1660) );
  assign n1661 = n1658 | n1660 ;
  buffer buf_n400( .i (x36), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n438( .i (x40), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  assign n1662 = n408 | n446 ;
  buffer buf_n209( .i (n208), .o (n209) );
  assign n1663 = n192 & n272 ;
  buffer buf_n1664( .i (n1663), .o (n1664) );
  assign n1665 = n209 | n1664 ;
  buffer buf_n1666( .i (n1665), .o (n1666) );
  assign n1667 = n205 & n273 ;
  buffer buf_n1668( .i (n1667), .o (n1668) );
  buffer buf_n1669( .i (n1668), .o (n1669) );
  assign n1670 = ~n1666 & n1669 ;
  buffer buf_n1671( .i (n1670), .o (n1671) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  assign n1676 = n1662 & ~n1674 ;
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n430( .i (x39), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  assign n1677 = n395 | n436 ;
  buffer buf_n1678( .i (n1677), .o (n1678) );
  assign n1679 = n209 & ~n1664 ;
  buffer buf_n1680( .i (n1679), .o (n1680) );
  assign n1681 = ~n1669 & n1680 ;
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  assign n1686 = n1678 & ~n1684 ;
  buffer buf_n1687( .i (n1686), .o (n1687) );
  assign n1688 = n1676 | n1687 ;
  buffer buf_n420( .i (x38), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  assign n1689 = n1666 | n1669 ;
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n1691( .i (n1690), .o (n1691) );
  buffer buf_n1692( .i (n1691), .o (n1692) );
  assign n1694 = n428 & n1692 ;
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  assign n1695 = n195 | n1059 ;
  assign n1696 = n276 & n1695 ;
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  assign n1701 = n386 & n1699 ;
  assign n1702 = n1694 | n1701 ;
  buffer buf_n1703( .i (n1702), .o (n1703) );
  assign n1704 = n1688 | n1703 ;
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  assign n1705 = ~n281 & n398 ;
  assign n1706 = n375 & ~n1705 ;
  assign n1707 = n1669 & n1680 ;
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1710( .i (n1709), .o (n1710) );
  buffer buf_n1711( .i (n1710), .o (n1711) );
  buffer buf_n1712( .i (n1711), .o (n1712) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n410( .i (x37), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  assign n1713 = n362 | n418 ;
  buffer buf_n1714( .i (n1713), .o (n1714) );
  assign n1715 = ~n1712 & n1714 ;
  assign n1716 = n1706 & ~n1715 ;
  assign n1717 = ~n1704 & n1716 ;
  assign n1718 = n69 | n1710 ;
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  assign n1721 = n278 & n1682 ;
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  assign n1725 = n48 | n1723 ;
  buffer buf_n1726( .i (n1725), .o (n1726) );
  assign n1727 = n1720 & n1726 ;
  assign n1728 = ~n58 & n1699 ;
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  assign n1730 = n179 & ~n1672 ;
  assign n1731 = n373 | n1730 ;
  buffer buf_n1732( .i (n1731), .o (n1732) );
  assign n1733 = n1729 | n1732 ;
  buffer buf_n609( .i (n608), .o (n609) );
  assign n1734 = n609 | n1684 ;
  assign n1735 = n631 | n1709 ;
  buffer buf_n1736( .i (n1735), .o (n1736) );
  assign n1737 = n1734 & n1736 ;
  assign n1738 = n36 | n1673 ;
  buffer buf_n621( .i (n620), .o (n621) );
  assign n1739 = ~n621 & n1692 ;
  assign n1740 = n1738 & ~n1739 ;
  assign n1741 = n1737 & n1740 ;
  assign n1742 = ~n1733 & n1741 ;
  assign n1743 = n1727 & n1742 ;
  assign n1744 = n1717 | n1743 ;
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n741( .i (n740), .o (n741) );
  assign n1746 = ~n190 & n279 ;
  assign n1747 = n741 & ~n1746 ;
  buffer buf_n1748( .i (n1747), .o (n1748) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  assign n1755 = n1745 & ~n1753 ;
  buffer buf_n1756( .i (n1755), .o (n1756) );
  buffer buf_n1757( .i (n1756), .o (n1757) );
  assign n1758 = n1646 & ~n1757 ;
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n1139( .i (n1138), .o (n1139) );
  buffer buf_n1140( .i (n1139), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  assign n1760 = ~n147 & n1141 ;
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  assign n1768 = n1550 & n1767 ;
  assign n1769 = n1759 & ~n1768 ;
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  assign n1773 = n1661 & ~n1772 ;
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n1775( .i (n1774), .o (n1775) );
  buffer buf_n1776( .i (n1775), .o (n1776) );
  buffer buf_n1777( .i (n1776), .o (n1777) );
  buffer buf_n1778( .i (n1777), .o (n1778) );
  buffer buf_n1779( .i (n1778), .o (n1779) );
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n1799( .i (n1798), .o (n1799) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  assign n1800 = n1330 & n1527 ;
  buffer buf_n1801( .i (n1800), .o (n1801) );
  assign n1802 = n1352 | n1801 ;
  assign n1803 = n1352 & n1801 ;
  assign n1804 = n1802 & ~n1803 ;
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n376( .i (n375), .o (n376) );
  assign n1813 = ~n147 & n376 ;
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  assign n1821 = n1805 & n1820 ;
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  assign n1822 = n387 & n1693 ;
  assign n1823 = n1729 | n1822 ;
  assign n1824 = n46 & ~n361 ;
  buffer buf_n1825( .i (n1824), .o (n1825) );
  assign n1826 = n1711 | n1825 ;
  buffer buf_n1685( .i (n1684), .o (n1685) );
  assign n1827 = n398 & ~n1685 ;
  assign n1828 = n1826 & ~n1827 ;
  assign n1829 = ~n1823 & n1828 ;
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  assign n1830 = n71 | n1724 ;
  assign n1831 = n79 & ~n406 ;
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  assign n1834 = n1674 | n1833 ;
  assign n1835 = n375 & n1834 ;
  assign n1836 = n1830 & n1835 ;
  assign n1837 = n1829 & n1836 ;
  buffer buf_n126( .i (x10), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  assign n1838 = n134 & ~n1684 ;
  assign n1839 = ~n621 & n1699 ;
  assign n1840 = n1838 | n1839 ;
  buffer buf_n149( .i (x12), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  assign n1841 = n158 & n1693 ;
  assign n1842 = n1840 | n1841 ;
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  assign n1844 = ~n167 & n631 ;
  assign n1845 = n1710 | n1844 ;
  buffer buf_n116( .i (x9), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  assign n1846 = n124 & ~n1673 ;
  assign n1847 = n1845 & ~n1846 ;
  assign n1848 = ~n1732 & n1847 ;
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  assign n1849 = n611 | n1724 ;
  assign n1850 = n1848 & n1849 ;
  assign n1851 = ~n1843 & n1850 ;
  assign n1852 = n1837 | n1851 ;
  assign n1853 = ~n1752 & n1852 ;
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  assign n1858 = n1647 & ~n1857 ;
  assign n1859 = ~n1821 & n1858 ;
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  assign n1870 = n1227 & n1534 ;
  assign n1871 = n999 | n1189 ;
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  assign n1872 = n201 | n1164 ;
  assign n1873 = n1871 | n1872 ;
  assign n1874 = n1110 | n1873 ;
  buffer buf_n1875( .i (n1874), .o (n1875) );
  assign n1876 = n1006 & n1191 ;
  buffer buf_n202( .i (n201), .o (n202) );
  assign n1877 = n202 & n1165 ;
  assign n1878 = n1110 & n1877 ;
  assign n1879 = n1876 & n1878 ;
  assign n1880 = n1875 & ~n1879 ;
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n1883( .i (n1882), .o (n1883) );
  buffer buf_n1884( .i (n1883), .o (n1884) );
  buffer buf_n1885( .i (n1884), .o (n1885) );
  buffer buf_n1886( .i (n1885), .o (n1886) );
  buffer buf_n1887( .i (n1886), .o (n1887) );
  assign n1888 = n1534 | n1887 ;
  assign n1889 = ~n1870 & n1888 ;
  buffer buf_n1890( .i (n1889), .o (n1890) );
  assign n1891 = n472 & ~n1890 ;
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  buffer buf_n1894( .i (n1893), .o (n1894) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  assign n1895 = ~n1608 & n1810 ;
  buffer buf_n1896( .i (n1895), .o (n1896) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  assign n1897 = ~n1361 & n1609 ;
  assign n1898 = n1896 | n1897 ;
  buffer buf_n1899( .i (n1898), .o (n1899) );
  assign n1900 = n1894 & n1899 ;
  assign n1901 = n1657 | n1900 ;
  assign n1902 = n1894 | n1899 ;
  buffer buf_n1903( .i (n1902), .o (n1903) );
  assign n1904 = ~n1901 & n1903 ;
  assign n1905 = n1869 | n1904 ;
  buffer buf_n1906( .i (n1905), .o (n1906) );
  buffer buf_n1907( .i (n1906), .o (n1907) );
  buffer buf_n1908( .i (n1907), .o (n1908) );
  buffer buf_n1909( .i (n1908), .o (n1909) );
  buffer buf_n1910( .i (n1909), .o (n1910) );
  buffer buf_n1911( .i (n1910), .o (n1911) );
  buffer buf_n1912( .i (n1911), .o (n1912) );
  buffer buf_n1913( .i (n1912), .o (n1913) );
  buffer buf_n1914( .i (n1913), .o (n1914) );
  buffer buf_n1915( .i (n1914), .o (n1915) );
  buffer buf_n1916( .i (n1915), .o (n1916) );
  buffer buf_n1917( .i (n1916), .o (n1917) );
  buffer buf_n1918( .i (n1917), .o (n1918) );
  buffer buf_n1919( .i (n1918), .o (n1919) );
  buffer buf_n1920( .i (n1919), .o (n1920) );
  buffer buf_n1921( .i (n1920), .o (n1921) );
  buffer buf_n1922( .i (n1921), .o (n1922) );
  buffer buf_n1923( .i (n1922), .o (n1923) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n1384( .i (n1383), .o (n1384) );
  assign n1925 = n1384 & n1526 ;
  buffer buf_n1926( .i (n1925), .o (n1926) );
  buffer buf_n1927( .i (n1926), .o (n1927) );
  assign n1928 = n1398 & ~n1927 ;
  assign n1929 = ~n1398 & n1927 ;
  assign n1930 = n1928 | n1929 ;
  buffer buf_n1931( .i (n1930), .o (n1931) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  assign n1940 = n1348 & ~n1530 ;
  buffer buf_n1941( .i (n1940), .o (n1941) );
  assign n1949 = n1931 & ~n1941 ;
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  assign n1950 = n1396 & ~n1532 ;
  assign n1951 = n1949 | n1950 ;
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  assign n1954 = n223 & ~n774 ;
  buffer buf_n1955( .i (n1954), .o (n1955) );
  assign n1956 = n1297 & n1955 ;
  buffer buf_n1957( .i (n1956), .o (n1957) );
  assign n1958 = n1315 & n1957 ;
  assign n1959 = n1315 | n1957 ;
  assign n1960 = ~n1958 & n1959 ;
  buffer buf_n1961( .i (n1960), .o (n1961) );
  buffer buf_n1962( .i (n1961), .o (n1962) );
  buffer buf_n1963( .i (n1962), .o (n1963) );
  buffer buf_n1964( .i (n1963), .o (n1964) );
  assign n1966 = n1952 & n1964 ;
  buffer buf_n1967( .i (n1966), .o (n1967) );
  assign n1968 = n1313 & ~n1955 ;
  buffer buf_n1969( .i (n1968), .o (n1969) );
  buffer buf_n1970( .i (n1969), .o (n1970) );
  buffer buf_n1971( .i (n1970), .o (n1971) );
  buffer buf_n1972( .i (n1971), .o (n1972) );
  buffer buf_n1973( .i (n1972), .o (n1973) );
  buffer buf_n1974( .i (n1973), .o (n1974) );
  buffer buf_n1975( .i (n1974), .o (n1975) );
  buffer buf_n1976( .i (n1975), .o (n1976) );
  buffer buf_n1977( .i (n1976), .o (n1977) );
  assign n1978 = n1967 | n1977 ;
  buffer buf_n1979( .i (n1978), .o (n1979) );
  buffer buf_n1980( .i (n1979), .o (n1980) );
  assign n1981 = n1406 | n1608 ;
  assign n1982 = ~n1447 & n1981 ;
  buffer buf_n1983( .i (n1982), .o (n1983) );
  assign n1984 = n1980 & n1983 ;
  assign n1985 = n1980 | n1983 ;
  assign n1986 = ~n1984 & n1985 ;
  buffer buf_n1987( .i (n1986), .o (n1987) );
  buffer buf_n1965( .i (n1964), .o (n1965) );
  buffer buf_n1932( .i (n1931), .o (n1932) );
  buffer buf_n1933( .i (n1932), .o (n1933) );
  assign n1988 = n1807 & n1933 ;
  buffer buf_n1989( .i (n1988), .o (n1989) );
  assign n1993 = n1965 & n1989 ;
  buffer buf_n1994( .i (n1993), .o (n1994) );
  assign n1996 = n1407 | n1994 ;
  assign n1997 = n1407 & n1994 ;
  assign n1998 = n1996 & ~n1997 ;
  assign n1999 = n472 & n1890 ;
  buffer buf_n2000( .i (n1999), .o (n2000) );
  buffer buf_n2001( .i (n2000), .o (n2001) );
  assign n2002 = ~n1998 & n2001 ;
  buffer buf_n2003( .i (n2002), .o (n2003) );
  buffer buf_n2004( .i (n2003), .o (n2004) );
  assign n2005 = n1987 | n2004 ;
  assign n2006 = n1987 & n2004 ;
  assign n2007 = n2005 & ~n2006 ;
  assign n2008 = n10 | n144 ;
  buffer buf_n2009( .i (n2008), .o (n2009) );
  assign n2010 = n769 & n2009 ;
  buffer buf_n2011( .i (n2010), .o (n2011) );
  buffer buf_n2012( .i (n2011), .o (n2012) );
  buffer buf_n2013( .i (n2012), .o (n2013) );
  buffer buf_n2014( .i (n2013), .o (n2014) );
  buffer buf_n2015( .i (n2014), .o (n2015) );
  buffer buf_n2016( .i (n2015), .o (n2016) );
  buffer buf_n2017( .i (n2016), .o (n2017) );
  buffer buf_n2018( .i (n2017), .o (n2018) );
  buffer buf_n2019( .i (n2018), .o (n2019) );
  buffer buf_n2020( .i (n2019), .o (n2020) );
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  buffer buf_n2024( .i (n2023), .o (n2024) );
  buffer buf_n2025( .i (n2024), .o (n2025) );
  buffer buf_n2026( .i (n2025), .o (n2026) );
  buffer buf_n2027( .i (n2026), .o (n2027) );
  buffer buf_n2028( .i (n2027), .o (n2028) );
  buffer buf_n2029( .i (n2028), .o (n2029) );
  buffer buf_n2030( .i (n2029), .o (n2030) );
  buffer buf_n2031( .i (n2030), .o (n2031) );
  assign n2032 = ~n2007 & n2031 ;
  assign n2033 = n641 | n913 ;
  assign n2034 = n609 & ~n632 ;
  assign n2035 = n2033 & ~n2034 ;
  assign n2036 = n2009 | n2035 ;
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  assign n2037 = ~n82 & n743 ;
  assign n2038 = ~n1093 & n2037 ;
  assign n2039 = n2036 & ~n2038 ;
  buffer buf_n2040( .i (n2039), .o (n2040) );
  buffer buf_n2041( .i (n2040), .o (n2041) );
  buffer buf_n2042( .i (n2041), .o (n2042) );
  buffer buf_n2043( .i (n2042), .o (n2043) );
  buffer buf_n2044( .i (n2043), .o (n2044) );
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n2046( .i (n2045), .o (n2046) );
  buffer buf_n2047( .i (n2046), .o (n2047) );
  buffer buf_n2048( .i (n2047), .o (n2048) );
  buffer buf_n2049( .i (n2048), .o (n2049) );
  buffer buf_n2050( .i (n2049), .o (n2050) );
  buffer buf_n2051( .i (n2050), .o (n2051) );
  buffer buf_n2052( .i (n2051), .o (n2052) );
  buffer buf_n2053( .i (n2052), .o (n2053) );
  buffer buf_n2054( .i (n2053), .o (n2054) );
  buffer buf_n2055( .i (n2054), .o (n2055) );
  buffer buf_n2056( .i (n2055), .o (n2056) );
  buffer buf_n2057( .i (n2056), .o (n2057) );
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  assign n2061 = ~n2032 & n2060 ;
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  buffer buf_n2064( .i (n2063), .o (n2064) );
  buffer buf_n2065( .i (n2064), .o (n2065) );
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n2070( .i (n2069), .o (n2070) );
  buffer buf_n2071( .i (n2070), .o (n2071) );
  buffer buf_n2072( .i (n2071), .o (n2072) );
  buffer buf_n2073( .i (n2072), .o (n2073) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n2075( .i (n2074), .o (n2075) );
  buffer buf_n2076( .i (n2075), .o (n2076) );
  buffer buf_n2077( .i (n2076), .o (n2077) );
  buffer buf_n2078( .i (n2077), .o (n2078) );
  buffer buf_n983( .i (n982), .o (n983) );
  assign n2079 = n983 & ~n1233 ;
  buffer buf_n2080( .i (n2079), .o (n2080) );
  buffer buf_n2081( .i (n2080), .o (n2081) );
  assign n2082 = ~n741 & n2081 ;
  buffer buf_n2083( .i (n2082), .o (n2083) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n2085( .i (n2084), .o (n2085) );
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2089( .i (n2088), .o (n2089) );
  buffer buf_n2090( .i (n2089), .o (n2090) );
  buffer buf_n2091( .i (n2090), .o (n2091) );
  buffer buf_n2092( .i (n2091), .o (n2092) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n2099( .i (n2098), .o (n2099) );
  buffer buf_n2100( .i (n2099), .o (n2100) );
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n2102( .i (n2101), .o (n2102) );
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n2106( .i (n2105), .o (n2106) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  assign n2110 = n1057 & ~n1532 ;
  buffer buf_n2111( .i (n2110), .o (n2111) );
  assign n2112 = n1216 & ~n1530 ;
  buffer buf_n2113( .i (n2112), .o (n2113) );
  assign n2114 = n1541 | n2113 ;
  buffer buf_n2115( .i (n2114), .o (n2115) );
  assign n2116 = ~n2111 & n2115 ;
  buffer buf_n2117( .i (n2116), .o (n2117) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  assign n2118 = n1099 & n1526 ;
  buffer buf_n2119( .i (n2118), .o (n2119) );
  assign n2120 = n1125 & n2119 ;
  assign n2121 = n1125 | n2119 ;
  assign n2122 = ~n2120 & n2121 ;
  buffer buf_n2123( .i (n2122), .o (n2123) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  buffer buf_n2128( .i (n2127), .o (n2128) );
  assign n2129 = n2117 & n2128 ;
  buffer buf_n2130( .i (n2129), .o (n2130) );
  assign n2131 = n2117 | n2128 ;
  buffer buf_n2132( .i (n2131), .o (n2132) );
  assign n2133 = ~n2130 & n2132 ;
  buffer buf_n2134( .i (n2133), .o (n2134) );
  assign n2136 = n1558 & ~n2134 ;
  buffer buf_n2137( .i (n2136), .o (n2137) );
  buffer buf_n2135( .i (n2134), .o (n2135) );
  assign n2139 = ~n1559 & n2135 ;
  assign n2140 = n2137 | n2139 ;
  buffer buf_n2141( .i (n2140), .o (n2141) );
  assign n2142 = n1615 & ~n2141 ;
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  assign n2143 = n1076 & n2113 ;
  buffer buf_n2144( .i (n2143), .o (n2144) );
  assign n2145 = n2115 & ~n2144 ;
  buffer buf_n2146( .i (n2145), .o (n2146) );
  assign n2147 = n1660 & n2146 ;
  assign n2148 = n1660 | n2146 ;
  assign n2149 = ~n2147 & n2148 ;
  buffer buf_n2150( .i (n2149), .o (n2150) );
  assign n2152 = n1610 & n2150 ;
  assign n2153 = n1597 | n2152 ;
  buffer buf_n2154( .i (n2153), .o (n2154) );
  buffer buf_n2155( .i (n2154), .o (n2155) );
  buffer buf_n2156( .i (n2155), .o (n2156) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  assign n2158 = n2142 | n2157 ;
  assign n2159 = ~n2106 & n2158 ;
  buffer buf_n2138( .i (n2137), .o (n2138) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  assign n2160 = n1152 & n1526 ;
  buffer buf_n2161( .i (n2160), .o (n2161) );
  assign n2162 = n1174 & n2161 ;
  assign n2163 = n1174 | n2161 ;
  assign n2164 = ~n2162 & n2163 ;
  buffer buf_n2165( .i (n2164), .o (n2165) );
  buffer buf_n2166( .i (n2165), .o (n2166) );
  buffer buf_n2167( .i (n2166), .o (n2167) );
  buffer buf_n2168( .i (n2167), .o (n2168) );
  buffer buf_n2169( .i (n2168), .o (n2169) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  buffer buf_n2171( .i (n2170), .o (n2171) );
  buffer buf_n2172( .i (n2171), .o (n2172) );
  buffer buf_n2173( .i (n2172), .o (n2173) );
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  assign n2175 = n1121 & ~n1534 ;
  buffer buf_n2176( .i (n2175), .o (n2176) );
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n2177), .o (n2178) );
  assign n2179 = n2132 & ~n2178 ;
  buffer buf_n2180( .i (n2179), .o (n2180) );
  assign n2181 = ~n2174 & n2180 ;
  assign n2182 = n2174 & ~n2180 ;
  assign n2183 = n2181 | n2182 ;
  buffer buf_n2184( .i (n2183), .o (n2184) );
  assign n2185 = ~n2138 & n2184 ;
  assign n2186 = n2138 & ~n2184 ;
  assign n2187 = n2185 | n2186 ;
  buffer buf_n2188( .i (n2187), .o (n2188) );
  buffer buf_n2189( .i (n2188), .o (n2189) );
  assign n2190 = ~n2159 & n2189 ;
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  assign n2191 = n37 & ~n181 ;
  assign n2192 = n1712 | n2191 ;
  buffer buf_n2193( .i (n1683), .o (n2193) );
  assign n2194 = n157 & ~n2193 ;
  buffer buf_n168( .i (n167), .o (n168) );
  assign n2195 = n168 & n1692 ;
  assign n2196 = n2194 | n2195 ;
  assign n2197 = ~n133 & n1237 ;
  buffer buf_n2198( .i (n2197), .o (n2198) );
  assign n2199 = n1674 | n2198 ;
  assign n2200 = ~n2196 & n2199 ;
  assign n2201 = n2192 & n2200 ;
  buffer buf_n622( .i (n621), .o (n622) );
  assign n2202 = n622 | n1723 ;
  buffer buf_n2203( .i (n630), .o (n2203) );
  assign n2204 = n1698 & ~n2203 ;
  buffer buf_n2205( .i (n2204), .o (n2205) );
  buffer buf_n2206( .i (n2205), .o (n2206) );
  assign n2207 = n2202 & ~n2206 ;
  assign n2208 = ~n376 & n2207 ;
  assign n2209 = n2201 & n2208 ;
  assign n2210 = n58 & ~n386 ;
  buffer buf_n2211( .i (n2210), .o (n2211) );
  assign n2212 = n1712 | n2211 ;
  buffer buf_n1675( .i (n1674), .o (n1675) );
  assign n2213 = ~n1675 & n1714 ;
  assign n2214 = n2212 & ~n2213 ;
  assign n2215 = n408 & ~n2193 ;
  buffer buf_n2216( .i (n2215), .o (n2216) );
  assign n2217 = n398 & n1693 ;
  assign n2218 = n2216 | n2217 ;
  assign n2219 = n82 | n1723 ;
  buffer buf_n2220( .i (n1698), .o (n2220) );
  assign n2221 = ~n69 & n2220 ;
  assign n2222 = n374 & ~n2221 ;
  assign n2223 = n2219 & n2222 ;
  assign n2224 = ~n2218 & n2223 ;
  assign n2225 = n2214 & n2224 ;
  assign n2226 = n2209 | n2225 ;
  buffer buf_n2227( .i (n2226), .o (n2227) );
  assign n2228 = ~n1753 & n2227 ;
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  assign n2231 = n1646 & ~n2230 ;
  buffer buf_n2232( .i (n2231), .o (n2232) );
  assign n2233 = n1767 & n2166 ;
  assign n2234 = n2232 & ~n2233 ;
  buffer buf_n2235( .i (n2234), .o (n2235) );
  buffer buf_n2236( .i (n2235), .o (n2236) );
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  buffer buf_n2241( .i (n2240), .o (n2241) );
  buffer buf_n2242( .i (n2241), .o (n2242) );
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n2244( .i (n2243), .o (n2244) );
  buffer buf_n2245( .i (n2244), .o (n2245) );
  buffer buf_n2246( .i (n2245), .o (n2246) );
  buffer buf_n2247( .i (n2246), .o (n2247) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  assign n2249 = n2190 | n2248 ;
  buffer buf_n2250( .i (n2249), .o (n2250) );
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  buffer buf_n2257( .i (n2256), .o (n2257) );
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  buffer buf_n2263( .i (n2262), .o (n2263) );
  buffer buf_n2264( .i (n2263), .o (n2264) );
  assign n2265 = n2099 & ~n2150 ;
  assign n2266 = n36 | n1722 ;
  buffer buf_n2267( .i (n2266), .o (n2267) );
  assign n2269 = n619 | n1708 ;
  assign n2270 = ~n372 & n2269 ;
  buffer buf_n2271( .i (n2270), .o (n2271) );
  assign n2273 = n166 & ~n1671 ;
  buffer buf_n2274( .i (n2273), .o (n2274) );
  assign n2276 = ~n45 & n1697 ;
  buffer buf_n2277( .i (n2276), .o (n2277) );
  assign n2279 = n2274 | n2277 ;
  assign n2280 = n2271 & ~n2279 ;
  assign n2281 = n2267 & n2280 ;
  assign n2282 = n632 | n1673 ;
  assign n2283 = n57 | n1709 ;
  buffer buf_n2284( .i (n2283), .o (n2284) );
  assign n2285 = n2282 & n2284 ;
  buffer buf_n2286( .i (n1691), .o (n2286) );
  assign n2287 = ~n609 & n2286 ;
  assign n2288 = n180 & ~n2193 ;
  assign n2289 = n2287 | n2288 ;
  assign n2290 = n2285 & ~n2289 ;
  assign n2291 = n2281 & n2290 ;
  buffer buf_n2292( .i (n1672), .o (n2292) );
  assign n2293 = n1678 & ~n2292 ;
  assign n2294 = n418 & n2286 ;
  assign n2295 = n2293 | n2294 ;
  assign n2296 = n362 & n2220 ;
  assign n2297 = n428 & ~n2193 ;
  assign n2298 = n2296 | n2297 ;
  assign n2299 = n2295 | n2298 ;
  buffer buf_n2300( .i (n1722), .o (n2300) );
  assign n2301 = n387 & ~n2300 ;
  assign n2302 = n1710 | n1832 ;
  assign n2303 = n374 & n2302 ;
  assign n2304 = ~n2301 & n2303 ;
  assign n2305 = ~n2299 & n2304 ;
  assign n2306 = n2291 | n2305 ;
  buffer buf_n2307( .i (n2306), .o (n2307) );
  assign n2308 = ~n1752 & n2307 ;
  buffer buf_n2309( .i (n2308), .o (n2309) );
  buffer buf_n2310( .i (n2309), .o (n2310) );
  assign n2311 = n1645 & ~n2310 ;
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  assign n2314 = n1541 & n1767 ;
  assign n2315 = n2313 & ~n2314 ;
  buffer buf_n2316( .i (n2315), .o (n2316) );
  buffer buf_n2317( .i (n2316), .o (n2317) );
  buffer buf_n2318( .i (n2317), .o (n2318) );
  buffer buf_n2319( .i (n2318), .o (n2319) );
  buffer buf_n2320( .i (n2319), .o (n2320) );
  buffer buf_n2321( .i (n2320), .o (n2321) );
  assign n2322 = n2265 | n2321 ;
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2151( .i (n2150), .o (n2151) );
  assign n2325 = n1611 | n2151 ;
  buffer buf_n2326( .i (n2325), .o (n2326) );
  assign n2327 = ~n2154 & n2326 ;
  assign n2328 = n2324 | n2327 ;
  buffer buf_n2329( .i (n2328), .o (n2329) );
  buffer buf_n2330( .i (n2329), .o (n2330) );
  buffer buf_n2331( .i (n2330), .o (n2331) );
  buffer buf_n2332( .i (n2331), .o (n2332) );
  buffer buf_n2333( .i (n2332), .o (n2333) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n2335( .i (n2334), .o (n2335) );
  buffer buf_n2336( .i (n2335), .o (n2336) );
  buffer buf_n2337( .i (n2336), .o (n2337) );
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  buffer buf_n2340( .i (n2339), .o (n2340) );
  buffer buf_n2341( .i (n2340), .o (n2341) );
  buffer buf_n2342( .i (n2341), .o (n2342) );
  buffer buf_n2343( .i (n2342), .o (n2343) );
  buffer buf_n2344( .i (n2343), .o (n2344) );
  buffer buf_n2345( .i (n2344), .o (n2345) );
  buffer buf_n2346( .i (n2345), .o (n2346) );
  buffer buf_n2347( .i (n2346), .o (n2347) );
  buffer buf_n2348( .i (n2347), .o (n2348) );
  buffer buf_n1598( .i (n1597), .o (n1598) );
  buffer buf_n1599( .i (n1598), .o (n1599) );
  assign n2349 = n1599 | n2326 ;
  assign n2350 = ~n2103 & n2349 ;
  assign n2351 = n2141 & ~n2350 ;
  assign n2352 = n1767 & n2124 ;
  assign n2353 = n633 | n2300 ;
  assign n2354 = n179 & n1691 ;
  assign n2355 = ~n34 & n1697 ;
  buffer buf_n2356( .i (n2355), .o (n2356) );
  assign n2358 = n2354 | n2356 ;
  assign n2359 = n155 & ~n1671 ;
  assign n2360 = n372 | n2359 ;
  buffer buf_n2361( .i (n2360), .o (n2361) );
  assign n2365 = n2358 | n2361 ;
  assign n2366 = n2353 & ~n2365 ;
  buffer buf_n169( .i (n168), .o (n169) );
  assign n2367 = n169 & ~n1685 ;
  assign n2368 = n621 | n2292 ;
  buffer buf_n2369( .i (n45), .o (n2369) );
  assign n2370 = n1237 & n2369 ;
  buffer buf_n2371( .i (n1709), .o (n2371) );
  assign n2372 = n2370 | n2371 ;
  assign n2373 = n2368 & n2372 ;
  assign n2374 = ~n2367 & n2373 ;
  assign n2375 = n2366 & n2374 ;
  assign n2376 = ~n81 & n2220 ;
  buffer buf_n2377( .i (n1683), .o (n2377) );
  assign n2378 = n418 & ~n2377 ;
  assign n2379 = n2376 | n2378 ;
  assign n2380 = n385 | n427 ;
  assign n2381 = ~n2292 & n2380 ;
  assign n2382 = n408 & n2286 ;
  assign n2383 = n2381 | n2382 ;
  assign n2384 = n2379 | n2383 ;
  assign n2385 = n67 & ~n395 ;
  buffer buf_n2386( .i (n2385), .o (n2386) );
  assign n2387 = n2371 | n2386 ;
  assign n2388 = n374 & n2387 ;
  buffer buf_n363( .i (n362), .o (n363) );
  assign n2389 = n363 & ~n2300 ;
  assign n2390 = n2388 & ~n2389 ;
  assign n2391 = ~n2384 & n2390 ;
  assign n2392 = n2375 | n2391 ;
  buffer buf_n2393( .i (n2392), .o (n2393) );
  assign n2394 = ~n1752 & n2393 ;
  buffer buf_n2395( .i (n2394), .o (n2395) );
  buffer buf_n2396( .i (n2395), .o (n2396) );
  assign n2397 = n1645 & ~n2396 ;
  buffer buf_n2398( .i (n2397), .o (n2398) );
  buffer buf_n2399( .i (n2398), .o (n2399) );
  assign n2400 = ~n2352 & n2399 ;
  buffer buf_n2401( .i (n2400), .o (n2401) );
  buffer buf_n2402( .i (n2401), .o (n2402) );
  buffer buf_n2403( .i (n2402), .o (n2403) );
  buffer buf_n2404( .i (n2403), .o (n2404) );
  buffer buf_n2405( .i (n2404), .o (n2405) );
  buffer buf_n2406( .i (n2405), .o (n2406) );
  buffer buf_n2407( .i (n2406), .o (n2407) );
  buffer buf_n2408( .i (n2407), .o (n2408) );
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n2410( .i (n2409), .o (n2410) );
  buffer buf_n2411( .i (n2410), .o (n2411) );
  assign n2412 = n2351 | n2411 ;
  assign n2413 = ~n1599 & n2326 ;
  buffer buf_n2414( .i (n2413), .o (n2414) );
  assign n2415 = ~n2141 & n2414 ;
  buffer buf_n2416( .i (n2415), .o (n2416) );
  assign n2417 = n2412 | n2416 ;
  buffer buf_n2418( .i (n2417), .o (n2418) );
  buffer buf_n2419( .i (n2418), .o (n2419) );
  buffer buf_n2420( .i (n2419), .o (n2420) );
  buffer buf_n2421( .i (n2420), .o (n2421) );
  buffer buf_n2422( .i (n2421), .o (n2422) );
  buffer buf_n2423( .i (n2422), .o (n2423) );
  buffer buf_n2424( .i (n2423), .o (n2424) );
  buffer buf_n2425( .i (n2424), .o (n2425) );
  buffer buf_n2426( .i (n2425), .o (n2426) );
  buffer buf_n2427( .i (n2426), .o (n2427) );
  buffer buf_n2428( .i (n2427), .o (n2428) );
  buffer buf_n2429( .i (n2428), .o (n2429) );
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  buffer buf_n2432( .i (n2431), .o (n2432) );
  buffer buf_n2433( .i (n2432), .o (n2433) );
  buffer buf_n2434( .i (n2433), .o (n2434) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1990( .i (n1989), .o (n1990) );
  buffer buf_n1991( .i (n1990), .o (n1991) );
  buffer buf_n1992( .i (n1991), .o (n1992) );
  assign n2435 = n1992 & n2000 ;
  buffer buf_n2436( .i (n2435), .o (n2436) );
  buffer buf_n1934( .i (n1933), .o (n1934) );
  buffer buf_n1935( .i (n1934), .o (n1935) );
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1937( .i (n1936), .o (n1937) );
  buffer buf_n1938( .i (n1937), .o (n1938) );
  buffer buf_n1939( .i (n1938), .o (n1939) );
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  assign n2437 = n1812 & n2000 ;
  assign n2438 = n1939 | n2437 ;
  assign n2439 = ~n2436 & n2438 ;
  buffer buf_n2440( .i (n2439), .o (n2440) );
  buffer buf_n1942( .i (n1941), .o (n1942) );
  buffer buf_n1943( .i (n1942), .o (n1943) );
  buffer buf_n1944( .i (n1943), .o (n1944) );
  buffer buf_n1945( .i (n1944), .o (n1945) );
  buffer buf_n1946( .i (n1945), .o (n1946) );
  buffer buf_n1947( .i (n1946), .o (n1947) );
  buffer buf_n1948( .i (n1947), .o (n1948) );
  assign n2441 = n1896 | n1948 ;
  buffer buf_n2442( .i (n2441), .o (n2442) );
  buffer buf_n2443( .i (n2442), .o (n2443) );
  buffer buf_n2444( .i (n2443), .o (n2444) );
  assign n2445 = n2440 | n2444 ;
  assign n2446 = n2440 & n2444 ;
  assign n2447 = n2445 & ~n2446 ;
  buffer buf_n2448( .i (n2447), .o (n2448) );
  assign n2449 = ~n1983 & n2001 ;
  buffer buf_n2450( .i (n2449), .o (n2450) );
  buffer buf_n2451( .i (n2450), .o (n2451) );
  buffer buf_n2452( .i (n2451), .o (n2452) );
  buffer buf_n2453( .i (n2452), .o (n2453) );
  buffer buf_n2454( .i (n2453), .o (n2454) );
  assign n2455 = n2448 | n2454 ;
  buffer buf_n2456( .i (n2455), .o (n2456) );
  assign n2457 = ~n1605 & n2456 ;
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  assign n2459 = n1953 | n1965 ;
  assign n2460 = ~n1967 & n2459 ;
  buffer buf_n2461( .i (n2460), .o (n2461) );
  buffer buf_n2462( .i (n2461), .o (n2462) );
  buffer buf_n2463( .i (n2462), .o (n2463) );
  assign n2464 = ~n2436 & n2463 ;
  buffer buf_n1995( .i (n1994), .o (n1995) );
  assign n2465 = n1995 & n2000 ;
  buffer buf_n2466( .i (n2465), .o (n2466) );
  buffer buf_n2467( .i (n2466), .o (n2467) );
  assign n2468 = n2464 | n2467 ;
  buffer buf_n2469( .i (n2468), .o (n2469) );
  buffer buf_n2470( .i (n2469), .o (n2470) );
  buffer buf_n2471( .i (n2470), .o (n2471) );
  buffer buf_n2472( .i (n2471), .o (n2472) );
  buffer buf_n2473( .i (n2472), .o (n2473) );
  buffer buf_n2474( .i (n2473), .o (n2474) );
  buffer buf_n2475( .i (n2474), .o (n2475) );
  assign n2476 = n2458 & ~n2475 ;
  assign n2477 = n1820 & n1961 ;
  buffer buf_n1754( .i (n1753), .o (n1754) );
  assign n2478 = n363 & ~n1685 ;
  buffer buf_n2479( .i (n2478), .o (n2479) );
  assign n2480 = n375 & n1719 ;
  assign n2481 = ~n2479 & n2480 ;
  buffer buf_n2482( .i (n81), .o (n2482) );
  assign n2483 = n1693 & ~n2482 ;
  buffer buf_n2357( .i (n2356), .o (n2357) );
  assign n2484 = n1736 & ~n2357 ;
  assign n2485 = ~n2483 & n2484 ;
  buffer buf_n2486( .i (n2485), .o (n2486) );
  assign n2487 = n2481 & n2486 ;
  assign n2488 = n1675 | n2211 ;
  assign n2489 = n1726 & n2488 ;
  buffer buf_n2490( .i (n2489), .o (n2490) );
  assign n2491 = n2487 & n2490 ;
  buffer buf_n2362( .i (n2361), .o (n2362) );
  buffer buf_n2363( .i (n2362), .o (n2363) );
  buffer buf_n2364( .i (n2363), .o (n2364) );
  assign n2492 = n1711 | n2198 ;
  assign n2493 = n124 & n2286 ;
  buffer buf_n2494( .i (n2493), .o (n2494) );
  assign n2495 = n2492 & ~n2494 ;
  buffer buf_n170( .i (n169), .o (n170) );
  assign n2496 = n170 & ~n1724 ;
  assign n2497 = n2495 & ~n2496 ;
  assign n2498 = ~n2364 & n2497 ;
  buffer buf_n93( .i (x7), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  assign n2499 = n103 & ~n1675 ;
  buffer buf_n105( .i (x8), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  assign n2500 = n114 & ~n1685 ;
  buffer buf_n1700( .i (n1699), .o (n1700) );
  assign n2501 = n181 & n1700 ;
  assign n2502 = n2500 | n2501 ;
  assign n2503 = n2499 | n2502 ;
  buffer buf_n2504( .i (n2503), .o (n2504) );
  assign n2505 = n2498 & ~n2504 ;
  assign n2506 = n2491 | n2505 ;
  buffer buf_n2507( .i (n2506), .o (n2507) );
  assign n2508 = ~n1754 & n2507 ;
  buffer buf_n2509( .i (n2508), .o (n2509) );
  buffer buf_n2510( .i (n2509), .o (n2510) );
  assign n2511 = n1647 & ~n2510 ;
  assign n2512 = ~n2477 & n2511 ;
  buffer buf_n2513( .i (n2512), .o (n2513) );
  buffer buf_n2514( .i (n2513), .o (n2514) );
  buffer buf_n2515( .i (n2514), .o (n2515) );
  buffer buf_n2516( .i (n2515), .o (n2516) );
  buffer buf_n2517( .i (n2516), .o (n2517) );
  buffer buf_n2518( .i (n2517), .o (n2518) );
  buffer buf_n2519( .i (n2518), .o (n2519) );
  buffer buf_n2520( .i (n2519), .o (n2520) );
  buffer buf_n2521( .i (n2520), .o (n2521) );
  buffer buf_n2522( .i (n2521), .o (n2522) );
  buffer buf_n2523( .i (n2522), .o (n2523) );
  buffer buf_n2524( .i (n2523), .o (n2524) );
  buffer buf_n2525( .i (n2524), .o (n2525) );
  buffer buf_n2526( .i (n2525), .o (n2526) );
  buffer buf_n2527( .i (n2526), .o (n2527) );
  buffer buf_n2528( .i (n2527), .o (n2528) );
  buffer buf_n2529( .i (n2528), .o (n2529) );
  assign n2530 = n2476 | n2529 ;
  buffer buf_n2107( .i (n2106), .o (n2107) );
  buffer buf_n2108( .i (n2107), .o (n2108) );
  buffer buf_n2109( .i (n2108), .o (n2109) );
  assign n2531 = n1605 | n2456 ;
  assign n2532 = ~n2109 & n2531 ;
  assign n2533 = n2475 & ~n2532 ;
  buffer buf_n2534( .i (n2533), .o (n2534) );
  assign n2535 = n2530 | n2534 ;
  buffer buf_n2536( .i (n2535), .o (n2536) );
  buffer buf_n2537( .i (n2536), .o (n2537) );
  buffer buf_n2538( .i (n2537), .o (n2538) );
  buffer buf_n2539( .i (n2538), .o (n2539) );
  buffer buf_n2540( .i (n2539), .o (n2540) );
  buffer buf_n2541( .i (n2540), .o (n2541) );
  buffer buf_n2542( .i (n2541), .o (n2542) );
  buffer buf_n2543( .i (n2542), .o (n2543) );
  buffer buf_n2544( .i (n2543), .o (n2544) );
  buffer buf_n2545( .i (n2544), .o (n2545) );
  buffer buf_n2546( .i (n2545), .o (n2546) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  assign n2547 = n1251 & n1955 ;
  buffer buf_n2548( .i (n2547), .o (n2548) );
  assign n2549 = n1277 | n2548 ;
  assign n2550 = n1277 & n2548 ;
  assign n2551 = n2549 & ~n2550 ;
  buffer buf_n2552( .i (n2551), .o (n2552) );
  buffer buf_n2553( .i (n2552), .o (n2553) );
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2555( .i (n2554), .o (n2555) );
  buffer buf_n2556( .i (n2555), .o (n2556) );
  buffer buf_n2557( .i (n2556), .o (n2557) );
  buffer buf_n2558( .i (n2557), .o (n2558) );
  buffer buf_n2559( .i (n2558), .o (n2559) );
  assign n2560 = n1979 & ~n2559 ;
  assign n2561 = ~n1979 & n2559 ;
  assign n2562 = n2560 | n2561 ;
  buffer buf_n2563( .i (n2562), .o (n2563) );
  assign n2564 = n2467 & ~n2563 ;
  assign n2565 = ~n2467 & n2563 ;
  assign n2566 = n2564 | n2565 ;
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n2568( .i (n2567), .o (n2568) );
  buffer buf_n2569( .i (n2568), .o (n2569) );
  buffer buf_n2570( .i (n2569), .o (n2570) );
  buffer buf_n2571( .i (n2570), .o (n2571) );
  buffer buf_n2572( .i (n2571), .o (n2572) );
  assign n2573 = n2448 & n2454 ;
  buffer buf_n2574( .i (n2573), .o (n2574) );
  assign n2577 = n2454 & ~n2471 ;
  assign n2578 = n1604 | n2577 ;
  assign n2579 = n2574 | n2578 ;
  assign n2580 = ~n2109 & n2579 ;
  assign n2581 = n2572 & ~n2580 ;
  assign n2582 = n1820 & n2552 ;
  buffer buf_n2583( .i (n1691), .o (n2583) );
  assign n2584 = n113 & n2583 ;
  buffer buf_n84( .i (x6), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  assign n2585 = n91 | n133 ;
  assign n2586 = ~n2292 & n2585 ;
  assign n2587 = n2584 | n2586 ;
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  assign n2588 = n168 & n2220 ;
  assign n2589 = n973 & ~n2588 ;
  assign n2590 = ~n2587 & n2589 ;
  assign n2591 = n158 & ~n2300 ;
  buffer buf_n2592( .i (n2377), .o (n2592) );
  assign n2593 = n102 & ~n2592 ;
  assign n2594 = n2591 | n2593 ;
  assign n2595 = n2590 & ~n2594 ;
  assign n2596 = n121 | n177 ;
  buffer buf_n2597( .i (n2596), .o (n2597) );
  buffer buf_n2598( .i (n1708), .o (n2598) );
  assign n2599 = n2597 & ~n2598 ;
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  buffer buf_n2602( .i (n2601), .o (n2602) );
  buffer buf_n2603( .i (n2602), .o (n2603) );
  assign n2604 = n2595 & ~n2603 ;
  buffer buf_n2268( .i (n2267), .o (n2268) );
  assign n2605 = n533 & n2268 ;
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2606( .i (n1672), .o (n2606) );
  buffer buf_n2607( .i (n2606), .o (n2607) );
  assign n2608 = n1825 | n2607 ;
  assign n2609 = n2272 & n2608 ;
  assign n2610 = ~n69 & n2583 ;
  assign n2611 = n2284 & ~n2610 ;
  buffer buf_n2612( .i (n80), .o (n2612) );
  assign n2613 = n2377 | n2612 ;
  assign n2614 = ~n2205 & n2613 ;
  assign n2615 = n2611 & n2614 ;
  assign n2616 = n2609 & n2615 ;
  assign n2617 = n2605 & n2616 ;
  assign n2618 = n2604 | n2617 ;
  buffer buf_n2619( .i (n2618), .o (n2619) );
  buffer buf_n2620( .i (n2619), .o (n2620) );
  assign n2621 = ~n1754 & n2620 ;
  buffer buf_n2622( .i (n2621), .o (n2622) );
  buffer buf_n2623( .i (n2622), .o (n2623) );
  assign n2624 = n1647 & ~n2623 ;
  assign n2625 = ~n2582 & n2624 ;
  buffer buf_n2626( .i (n2625), .o (n2626) );
  buffer buf_n2627( .i (n2626), .o (n2627) );
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  buffer buf_n2631( .i (n2630), .o (n2631) );
  buffer buf_n2632( .i (n2631), .o (n2632) );
  buffer buf_n2633( .i (n2632), .o (n2633) );
  buffer buf_n2634( .i (n2633), .o (n2634) );
  buffer buf_n2635( .i (n2634), .o (n2635) );
  buffer buf_n2636( .i (n2635), .o (n2636) );
  buffer buf_n2637( .i (n2636), .o (n2637) );
  buffer buf_n2638( .i (n2637), .o (n2638) );
  buffer buf_n2639( .i (n2638), .o (n2639) );
  buffer buf_n2640( .i (n2639), .o (n2640) );
  buffer buf_n2641( .i (n2640), .o (n2641) );
  buffer buf_n2642( .i (n2641), .o (n2642) );
  assign n2643 = n2581 | n2642 ;
  buffer buf_n2644( .i (n2643), .o (n2644) );
  buffer buf_n2645( .i (n2644), .o (n2645) );
  buffer buf_n2646( .i (n2645), .o (n2646) );
  buffer buf_n2647( .i (n2646), .o (n2647) );
  buffer buf_n2648( .i (n2647), .o (n2648) );
  buffer buf_n2649( .i (n2648), .o (n2649) );
  buffer buf_n2650( .i (n2649), .o (n2650) );
  buffer buf_n2651( .i (n2650), .o (n2651) );
  buffer buf_n2652( .i (n2651), .o (n2652) );
  buffer buf_n2653( .i (n2652), .o (n2653) );
  buffer buf_n2654( .i (n2653), .o (n2654) );
  buffer buf_n2655( .i (n2654), .o (n2655) );
  assign n2656 = n2106 & ~n2448 ;
  assign n2657 = n362 & n2583 ;
  assign n2658 = n386 & ~n2377 ;
  assign n2659 = n2657 | n2658 ;
  buffer buf_n2278( .i (n2277), .o (n2278) );
  assign n2660 = n35 & n80 ;
  assign n2661 = n2371 | n2660 ;
  assign n2662 = ~n2278 & n2661 ;
  assign n2663 = ~n2659 & n2662 ;
  buffer buf_n2664( .i (n1722), .o (n2664) );
  assign n2665 = n59 | n2664 ;
  assign n2666 = n2386 | n2606 ;
  buffer buf_n2667( .i (n373), .o (n2667) );
  assign n2668 = n2666 & n2667 ;
  assign n2669 = n2665 & n2668 ;
  assign n2670 = n2663 & n2669 ;
  assign n2671 = n114 & ~n2607 ;
  buffer buf_n2275( .i (n2274), .o (n2275) );
  assign n2672 = n134 & n2583 ;
  assign n2673 = n2275 | n2672 ;
  assign n2674 = n2671 | n2673 ;
  assign n2675 = n156 & ~n2598 ;
  assign n2676 = ~n1237 & n1698 ;
  assign n2677 = n2675 | n2676 ;
  buffer buf_n1285( .i (n1284), .o (n1285) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  assign n2678 = ~n1683 & n2597 ;
  assign n2679 = n1287 | n2678 ;
  assign n2680 = n2677 | n2679 ;
  assign n2681 = n2272 & ~n2680 ;
  assign n2682 = ~n2674 & n2681 ;
  assign n2683 = n2670 | n2682 ;
  buffer buf_n2684( .i (n2683), .o (n2684) );
  buffer buf_n2685( .i (n2684), .o (n2685) );
  buffer buf_n2686( .i (n2685), .o (n2686) );
  assign n2687 = ~n1754 & n2686 ;
  buffer buf_n2688( .i (n2687), .o (n2688) );
  assign n2689 = n1646 & ~n2688 ;
  buffer buf_n2690( .i (n2689), .o (n2690) );
  assign n2691 = n1820 & n1931 ;
  assign n2692 = n2690 & ~n2691 ;
  buffer buf_n2693( .i (n2692), .o (n2693) );
  buffer buf_n2694( .i (n2693), .o (n2694) );
  buffer buf_n2695( .i (n2694), .o (n2695) );
  buffer buf_n2696( .i (n2695), .o (n2696) );
  buffer buf_n2697( .i (n2696), .o (n2697) );
  buffer buf_n2698( .i (n2697), .o (n2698) );
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n2700( .i (n2699), .o (n2700) );
  buffer buf_n2701( .i (n2700), .o (n2701) );
  buffer buf_n2702( .i (n2701), .o (n2702) );
  buffer buf_n2703( .i (n2702), .o (n2703) );
  buffer buf_n2704( .i (n2703), .o (n2704) );
  buffer buf_n2705( .i (n2704), .o (n2705) );
  assign n2706 = n2656 | n2705 ;
  buffer buf_n2707( .i (n2706), .o (n2707) );
  buffer buf_n2708( .i (n2707), .o (n2708) );
  buffer buf_n2709( .i (n2708), .o (n2709) );
  buffer buf_n2575( .i (n2574), .o (n2575) );
  buffer buf_n2576( .i (n2575), .o (n2576) );
  assign n2710 = n2458 & ~n2576 ;
  assign n2711 = n2709 | n2710 ;
  buffer buf_n2712( .i (n2711), .o (n2712) );
  buffer buf_n2713( .i (n2712), .o (n2713) );
  buffer buf_n2714( .i (n2713), .o (n2714) );
  buffer buf_n2715( .i (n2714), .o (n2715) );
  buffer buf_n2716( .i (n2715), .o (n2716) );
  buffer buf_n2717( .i (n2716), .o (n2717) );
  buffer buf_n2718( .i (n2717), .o (n2718) );
  buffer buf_n2719( .i (n2718), .o (n2719) );
  buffer buf_n2720( .i (n2719), .o (n2720) );
  buffer buf_n2721( .i (n2720), .o (n2721) );
  buffer buf_n2722( .i (n2721), .o (n2722) );
  buffer buf_n2723( .i (n2722), .o (n2723) );
  assign n2724 = n2536 | n2645 ;
  buffer buf_n2725( .i (n2724), .o (n2725) );
  assign n2726 = n1787 & ~n2336 ;
  buffer buf_n2727( .i (n2726), .o (n2727) );
  assign n2728 = n2252 | n2422 ;
  buffer buf_n2729( .i (n2728), .o (n2729) );
  assign n2730 = n2727 & ~n2729 ;
  assign n2731 = n1913 | n2712 ;
  buffer buf_n2732( .i (n2731), .o (n2732) );
  assign n2735 = n2730 & ~n2732 ;
  assign n2736 = ~n2725 & n2735 ;
  buffer buf_n2737( .i (n2736), .o (n2737) );
  buffer buf_n2738( .i (n2737), .o (n2738) );
  buffer buf_n2739( .i (n2738), .o (n2739) );
  buffer buf_n2740( .i (n2739), .o (n2740) );
  buffer buf_n2741( .i (n2740), .o (n2741) );
  buffer buf_n2742( .i (n2741), .o (n2742) );
  buffer buf_n2743( .i (n2742), .o (n2743) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  buffer buf_n245( .i (n244), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  assign n2744 = n256 & ~n2737 ;
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  assign n2745 = n517 & ~n2725 ;
  buffer buf_n2746( .i (n2745), .o (n2746) );
  buffer buf_n2747( .i (n2746), .o (n2747) );
  assign n2748 = n2744 & ~n2747 ;
  buffer buf_n2749( .i (n2748), .o (n2749) );
  buffer buf_n2750( .i (n2749), .o (n2750) );
  buffer buf_n2751( .i (n2750), .o (n2751) );
  buffer buf_n2752( .i (n2751), .o (n2752) );
  buffer buf_n536( .i (x45), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  assign n2753 = n2537 & n2646 ;
  assign n2754 = n2725 & ~n2753 ;
  buffer buf_n2755( .i (n2754), .o (n2755) );
  buffer buf_n2756( .i (n2755), .o (n2756) );
  assign n2760 = n582 & n2756 ;
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  buffer buf_n1505( .i (n1504), .o (n1505) );
  buffer buf_n1506( .i (n1505), .o (n1506) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1518( .i (n1517), .o (n1518) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n1522( .i (n1521), .o (n1522) );
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  assign n2761 = n581 | n2755 ;
  assign n2762 = ~n1524 & n2761 ;
  assign n2763 = ~n2760 & n2762 ;
  buffer buf_n2764( .i (n2763), .o (n2764) );
  buffer buf_n2733( .i (n2732), .o (n2733) );
  buffer buf_n2734( .i (n2733), .o (n2734) );
  assign n2765 = n1916 & n2715 ;
  assign n2766 = n2734 & ~n2765 ;
  buffer buf_n2767( .i (n2766), .o (n2767) );
  assign n2768 = ~n1788 & n2337 ;
  assign n2769 = n2727 | n2768 ;
  buffer buf_n2770( .i (n2769), .o (n2770) );
  assign n2771 = n2253 & n2423 ;
  assign n2772 = n2729 & ~n2771 ;
  buffer buf_n2773( .i (n2772), .o (n2773) );
  assign n2774 = n2770 | n2773 ;
  assign n2775 = n2770 & n2773 ;
  assign n2776 = n2774 & ~n2775 ;
  buffer buf_n2777( .i (n2776), .o (n2777) );
  assign n2778 = n2767 | n2777 ;
  assign n2779 = n2767 & n2777 ;
  assign n2780 = n2778 & ~n2779 ;
  buffer buf_n2781( .i (n2780), .o (n2781) );
  assign n2782 = n2764 & n2781 ;
  assign n2783 = n2764 | n2781 ;
  assign n2784 = ~n2782 & n2783 ;
  buffer buf_n2757( .i (n2756), .o (n2757) );
  buffer buf_n2758( .i (n2757), .o (n2758) );
  buffer buf_n2759( .i (n2758), .o (n2759) );
  assign n2785 = n2759 & n2781 ;
  assign n2786 = n2759 | n2781 ;
  assign n2787 = ~n2785 & n2786 ;
  assign y0 = ~n684 ;
  assign y1 = ~n733 ;
  assign y2 = ~n832 ;
  assign y3 = n896 ;
  assign y4 = n961 ;
  assign y5 = n1433 ;
  assign y6 = n1487 ;
  assign y7 = n1582 ;
  assign y8 = n1642 ;
  assign y9 = ~n1799 ;
  assign y10 = n1924 ;
  assign y11 = ~n2078 ;
  assign y12 = n2264 ;
  assign y13 = n2348 ;
  assign y14 = n2434 ;
  assign y15 = n2546 ;
  assign y16 = n2655 ;
  assign y17 = n2723 ;
  assign y18 = ~n2743 ;
  assign y19 = ~n2752 ;
  assign y20 = ~n2784 ;
  assign y21 = n2787 ;
endmodule
