module top( N1 , N101 , N105 , N109 , N113 , N117 , N121 , N125 , N129 , N13 , N130 , N131 , N132 , N133 , N134 , N135 , N136 , N137 , N17 , N21 , N25 , N29 , N33 , N37 , N41 , N45 , N49 , N5 , N53 , N57 , N61 , N65 , N69 , N73 , N77 , N81 , N85 , N89 , N9 , N93 , N97 , N724 , N725 , N726 , N727 , N728 , N729 , N730 , N731 , N732 , N733 , N734 , N735 , N736 , N737 , N738 , N739 , N740 , N741 , N742 , N743 , N744 , N745 , N746 , N747 , N748 , N749 , N750 , N751 , N752 , N753 , N754 , N755 );
  input N1 , N101 , N105 , N109 , N113 , N117 , N121 , N125 , N129 , N13 , N130 , N131 , N132 , N133 , N134 , N135 , N136 , N137 , N17 , N21 , N25 , N29 , N33 , N37 , N41 , N45 , N49 , N5 , N53 , N57 , N61 , N65 , N69 , N73 , N77 , N81 , N85 , N89 , N9 , N93 , N97 ;
  output N724 , N725 , N726 , N727 , N728 , N729 , N730 , N731 , N732 , N733 , N734 , N735 , N736 , N737 , N738 , N739 , N740 , N741 , N742 , N743 , N744 , N745 , N746 , N747 , N748 , N749 , N750 , N751 , N752 , N753 , N754 , N755 ;
  wire n1028 , n1029 , n1030 , n1032 , n1034 , n1035 , n1036 , n1038 , n1039 , n1040 , n1042 , n1043 , n1044 , n1046 , n1047 , n1048 , n1050 , n1051 , n1052 , n1054 , n1055 , n1056 , n1059 , n1060 , n1061 , n1063 , n1064 , n1065 , n1067 , n1068 , n1069 , n1072 , n1073 , n1074 , n1076 , n1077 , n1078 , n1092 , n1094 , n1095 , n1096 , n1098 , n1099 , n1100 , n1102 , n1103 , n1104 , n1106 , n1107 , n1108 , n1110 , n1111 , n1112 , n1114 , n1115 , n1116 , n1118 , n1119 , n1120 , n1122 , n1123 , n1124 , n1126 , n1127 , n1128 , n1130 , n1131 , n1132 , n1134 , n1135 , n1136 , n1138 , n1139 , n1140 , n1153 , n1155 , n1156 , n1157 , n1159 , n1160 , n1161 , n1163 , n1164 , n1165 , n1167 , n1168 , n1169 , n1171 , n1172 , n1173 , n1175 , n1176 , n1177 , n1179 , n1180 , n1181 , n1183 , n1184 , n1185 , n1187 , n1188 , n1189 , n1191 , n1192 , n1193 , n1195 , n1196 , n1197 , n1199 , n1200 , n1201 , n1214 , n1222 , n1224 , n1227 , n1228 , n1230 , n1233 , n1234 , n1236 , n1237 , n1238 , n1240 , n1241 , n1242 , n1244 , n1245 , n1246 , n1248 , n1249 , n1250 , n1252 , n1253 , n1254 , n1257 , n1258 , n1259 , n1261 , n1262 , n1263 , n1276 , n1277 , n1278 , n1280 , n1282 , n1283 , n1284 , n1286 , n1287 , n1288 , n1290 , n1291 , n1292 , n1294 , n1295 , n1296 , n1298 , n1299 , n1300 , n1302 , n1303 , n1304 , n1307 , n1308 , n1309 , n1311 , n1312 , n1313 , n1327 , n1337 , n1345 , n1355 , n1363 , n1364 , n1366 , n1369 , n1370 , n1372 , n1375 , n1376 , n1378 , n1379 , n1380 , n1382 , n1383 , n1384 , n1386 , n1387 , n1388 , n1390 , n1391 , n1392 , n1405 , n1406 , n1412 , n1413 , n1414 , n1415 , n1416 , n1418 , n1419 , n1420 , n1422 , n1424 , n1425 , n1426 , n1428 , n1429 , n1430 , n1432 , n1433 , n1434 , n1436 , n1437 , n1438 , n1440 , n1441 , n1442 , n1455 , n1456 , n1457 , n1459 , n1461 , n1462 , n1463 , n1465 , n1466 , n1467 , n1469 , n1470 , n1471 , n1473 , n1474 , n1475 , n1477 , n1478 , n1479 , n1492 , n1498 , n1500 , n1502 , n1504 , n1505 , n1506 , n1507 , n1509 , n1510 , n1511 , n1512 , n1514 , n1515 , n1516 , n1517 , n1519 , n1520 , n1521 , n1522 , n1530 , n1532 , n1534 , n1535 , n1536 , n1537 , n1539 , n1540 , n1541 , n1542 , n1544 , n1545 , n1546 , n1547 , n1549 , n1550 , n1551 , n1552 , n1558 , n1560 , n1562 , n1564 , n1565 , n1566 , n1567 , n1569 , n1570 , n1571 , n1572 , n1574 , n1575 , n1576 , n1577 , n1579 , n1580 , n1581 , n1582 , n1584 , n1586 , n1587 , n1588 , n1589 , n1591 , n1592 , n1593 , n1594 , n1596 , n1597 , n1598 , n1599 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1612 , n1614 , n1616 , n1618 , n1619 , n1620 , n1621 , n1623 , n1624 , n1625 , n1626 , n1628 , n1629 , n1630 , n1631 , n1633 , n1634 , n1635 , n1636 , n1638 , n1640 , n1642 , n1643 , n1644 , n1645 , n1647 , n1648 , n1649 , n1650 , n1652 , n1653 , n1654 , n1655 , n1657 , n1658 , n1659 , n1660 , n1662 , n1664 , n1665 , n1666 , n1667 , n1669 , n1670 , n1671 , n1672 , n1674 , n1675 , n1676 , n1677 , n1679 , n1680 , n1681 , n1682 , n1684 , n1686 , n1687 , n1688 , n1689 , n1691 , n1692 , n1693 , n1694 , n1696 , n1697 , n1698 , n1699 , n1701 , n1702 , n1703 ;
  buffer buf_n42( .i (N1), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n477( .i (N33), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n593( .i (N49), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  buffer buf_n597( .i (n596), .o (n597) );
  buffer buf_n598( .i (n597), .o (n598) );
  assign n1028 = n482 & ~n598 ;
  assign n1029 = ~n482 & n598 ;
  assign n1030 = n1028 | n1029 ;
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n274( .i (N129), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n353( .i (N137), .o (n353) );
  buffer buf_n354( .i (n353), .o (n354) );
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  assign n1032 = n277 & n356 ;
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n361( .i (N17), .o (n361) );
  buffer buf_n362( .i (n361), .o (n362) );
  buffer buf_n363( .i (n362), .o (n363) );
  assign n1034 = n44 & ~n363 ;
  assign n1035 = ~n44 & n363 ;
  assign n1036 = n1034 | n1035 ;
  buffer buf_n1037( .i (n1036), .o (n1037) );
  assign n1038 = n1033 & ~n1037 ;
  assign n1039 = ~n1033 & n1037 ;
  assign n1040 = n1038 | n1039 ;
  buffer buf_n1041( .i (n1040), .o (n1041) );
  assign n1042 = n1031 | n1041 ;
  assign n1043 = n1031 & n1041 ;
  assign n1044 = n1042 & ~n1043 ;
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n796( .i (N73), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n798( .i (n797), .o (n798) );
  buffer buf_n825( .i (N77), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n827( .i (n826), .o (n827) );
  assign n1046 = n798 | n827 ;
  assign n1047 = n798 & n827 ;
  assign n1048 = n1046 & ~n1047 ;
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n738( .i (N65), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n767( .i (N69), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  assign n1050 = n740 & ~n769 ;
  assign n1051 = ~n740 & n769 ;
  assign n1052 = n1050 | n1051 ;
  buffer buf_n1053( .i (n1052), .o (n1053) );
  assign n1054 = ~n1049 & n1053 ;
  assign n1055 = n1049 & ~n1053 ;
  assign n1056 = n1054 | n1055 ;
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n912( .i (N89), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n970( .i (N93), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  assign n1059 = n914 | n972 ;
  assign n1060 = n914 & n972 ;
  assign n1061 = n1059 & ~n1060 ;
  buffer buf_n1062( .i (n1061), .o (n1062) );
  buffer buf_n854( .i (N81), .o (n854) );
  buffer buf_n855( .i (n854), .o (n855) );
  buffer buf_n856( .i (n855), .o (n856) );
  buffer buf_n883( .i (N85), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n885( .i (n884), .o (n885) );
  assign n1063 = n856 & ~n885 ;
  assign n1064 = ~n856 & n885 ;
  assign n1065 = n1063 | n1064 ;
  buffer buf_n1066( .i (n1065), .o (n1066) );
  assign n1067 = ~n1062 & n1066 ;
  assign n1068 = n1062 & ~n1066 ;
  assign n1069 = n1067 | n1068 ;
  buffer buf_n1070( .i (n1069), .o (n1070) );
  assign n1072 = n1057 & n1070 ;
  assign n1073 = n1057 | n1070 ;
  assign n1074 = ~n1072 & n1073 ;
  buffer buf_n1075( .i (n1074), .o (n1075) );
  assign n1076 = ~n1045 & n1075 ;
  assign n1077 = n1045 & ~n1075 ;
  assign n1078 = n1076 | n1077 ;
  buffer buf_n1079( .i (n1078), .o (n1079) );
  buffer buf_n1080( .i (n1079), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n1086( .i (n1085), .o (n1086) );
  buffer buf_n1087( .i (n1086), .o (n1087) );
  buffer buf_n1088( .i (n1087), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n337( .i (N135), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  assign n1092 = n344 & n360 ;
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n100( .i (N105), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n216( .i (N121), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  assign n1094 = n103 & ~n219 ;
  assign n1095 = ~n103 & n219 ;
  assign n1096 = n1094 | n1095 ;
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n799( .i (n798), .o (n799) );
  buffer buf_n915( .i (n914), .o (n915) );
  assign n1098 = n799 & ~n915 ;
  assign n1099 = ~n799 & n915 ;
  assign n1100 = n1098 | n1099 ;
  buffer buf_n1101( .i (n1100), .o (n1101) );
  assign n1102 = ~n1097 & n1101 ;
  assign n1103 = n1097 & ~n1101 ;
  assign n1104 = n1102 | n1103 ;
  buffer buf_n1105( .i (n1104), .o (n1105) );
  assign n1106 = n1093 & n1105 ;
  assign n1107 = n1093 | n1105 ;
  assign n1108 = ~n1106 & n1107 ;
  buffer buf_n1109( .i (n1108), .o (n1109) );
  buffer buf_n278( .i (N13), .o (n278) );
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n941( .i (N9), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  assign n1110 = n281 | n944 ;
  assign n1111 = n281 & n944 ;
  assign n1112 = n1110 & ~n1111 ;
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n622( .i (N5), .o (n622) );
  buffer buf_n623( .i (n622), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  assign n1114 = n45 & ~n625 ;
  assign n1115 = ~n45 & n625 ;
  assign n1116 = n1114 | n1115 ;
  buffer buf_n1117( .i (n1116), .o (n1117) );
  assign n1118 = ~n1113 & n1117 ;
  assign n1119 = n1113 & ~n1117 ;
  assign n1120 = n1118 | n1119 ;
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n535( .i (N41), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n564( .i (N45), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  assign n1122 = n538 | n567 ;
  assign n1123 = n538 & n567 ;
  assign n1124 = n1122 & ~n1123 ;
  buffer buf_n1125( .i (n1124), .o (n1125) );
  buffer buf_n506( .i (N37), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  assign n1126 = n480 & ~n509 ;
  assign n1127 = ~n480 & n509 ;
  assign n1128 = n1126 | n1127 ;
  buffer buf_n1129( .i (n1128), .o (n1129) );
  assign n1130 = ~n1125 & n1129 ;
  assign n1131 = n1125 & ~n1129 ;
  assign n1132 = n1130 | n1131 ;
  buffer buf_n1133( .i (n1132), .o (n1133) );
  assign n1134 = n1121 & n1133 ;
  assign n1135 = n1121 | n1133 ;
  assign n1136 = ~n1134 & n1135 ;
  buffer buf_n1137( .i (n1136), .o (n1137) );
  assign n1138 = ~n1109 & n1137 ;
  assign n1139 = n1109 & ~n1137 ;
  assign n1140 = n1138 | n1139 ;
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  buffer buf_n345( .i (N136), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  buffer buf_n350( .i (n349), .o (n350) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  assign n1153 = n352 & n360 ;
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n129( .i (N109), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n245( .i (N125), .o (n245) );
  buffer buf_n246( .i (n245), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  assign n1155 = n132 & ~n248 ;
  assign n1156 = ~n132 & n248 ;
  assign n1157 = n1155 | n1156 ;
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n828( .i (n827), .o (n828) );
  buffer buf_n973( .i (n972), .o (n973) );
  assign n1159 = n828 & ~n973 ;
  assign n1160 = ~n828 & n973 ;
  assign n1161 = n1159 | n1160 ;
  buffer buf_n1162( .i (n1161), .o (n1162) );
  assign n1163 = ~n1158 & n1162 ;
  assign n1164 = n1158 & ~n1162 ;
  assign n1165 = n1163 | n1164 ;
  buffer buf_n1166( .i (n1165), .o (n1166) );
  assign n1167 = n1154 & n1166 ;
  assign n1168 = n1154 | n1166 ;
  assign n1169 = ~n1167 & n1168 ;
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n419( .i (N25), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n448( .i (N29), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  assign n1171 = n422 | n451 ;
  assign n1172 = n422 & n451 ;
  assign n1173 = n1171 & ~n1172 ;
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n390( .i (N21), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  assign n1175 = n364 & ~n393 ;
  assign n1176 = ~n364 & n393 ;
  assign n1177 = n1175 | n1176 ;
  buffer buf_n1178( .i (n1177), .o (n1178) );
  assign n1179 = ~n1174 & n1178 ;
  assign n1180 = n1174 & ~n1178 ;
  assign n1181 = n1179 | n1180 ;
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n680( .i (N57), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n709( .i (N61), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n711( .i (n710), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  assign n1183 = n683 | n712 ;
  assign n1184 = n683 & n712 ;
  assign n1185 = n1183 & ~n1184 ;
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n651( .i (N53), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  assign n1187 = n596 & ~n654 ;
  assign n1188 = ~n596 & n654 ;
  assign n1189 = n1187 | n1188 ;
  buffer buf_n1190( .i (n1189), .o (n1190) );
  assign n1191 = ~n1186 & n1190 ;
  assign n1192 = n1186 & ~n1190 ;
  assign n1193 = n1191 | n1192 ;
  buffer buf_n1194( .i (n1193), .o (n1194) );
  assign n1195 = n1182 & n1194 ;
  assign n1196 = n1182 | n1194 ;
  assign n1197 = ~n1195 & n1196 ;
  buffer buf_n1198( .i (n1197), .o (n1198) );
  assign n1199 = ~n1170 & n1198 ;
  assign n1200 = n1170 & ~n1198 ;
  assign n1201 = n1199 | n1200 ;
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n1203( .i (n1202), .o (n1203) );
  assign n1214 = n1142 & ~n1203 ;
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n311( .i (N131), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  assign n1222 = n318 & n360 ;
  buffer buf_n1223( .i (n1222), .o (n1223) );
  assign n1224 = n538 & ~n683 ;
  buffer buf_n1225( .i (n537), .o (n1225) );
  buffer buf_n1226( .i (n682), .o (n1226) );
  assign n1227 = ~n1225 & n1226 ;
  assign n1228 = n1224 | n1227 ;
  buffer buf_n1229( .i (n1228), .o (n1229) );
  assign n1230 = ~n422 & n944 ;
  buffer buf_n1231( .i (n421), .o (n1231) );
  buffer buf_n1232( .i (n943), .o (n1232) );
  assign n1233 = n1231 & ~n1232 ;
  assign n1234 = n1230 | n1233 ;
  buffer buf_n1235( .i (n1234), .o (n1235) );
  assign n1236 = ~n1229 & n1235 ;
  assign n1237 = n1229 & ~n1235 ;
  assign n1238 = n1236 | n1237 ;
  buffer buf_n1239( .i (n1238), .o (n1239) );
  assign n1240 = n1223 & n1239 ;
  assign n1241 = n1223 | n1239 ;
  assign n1242 = ~n1240 & n1241 ;
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  assign n1244 = n102 | n131 ;
  assign n1245 = n102 & n131 ;
  assign n1246 = n1244 & ~n1245 ;
  buffer buf_n1247( .i (n1246), .o (n1247) );
  buffer buf_n71( .i (N101), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n999( .i (N97), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  assign n1248 = ~n73 & n1001 ;
  assign n1249 = n73 & ~n1001 ;
  assign n1250 = n1248 | n1249 ;
  buffer buf_n1251( .i (n1250), .o (n1251) );
  assign n1252 = ~n1247 & n1251 ;
  assign n1253 = n1247 & ~n1251 ;
  assign n1254 = n1252 | n1253 ;
  buffer buf_n1255( .i (n1254), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  assign n1257 = n1058 & n1256 ;
  assign n1258 = n1058 | n1256 ;
  assign n1259 = ~n1257 & n1258 ;
  buffer buf_n1260( .i (n1259), .o (n1260) );
  assign n1261 = ~n1243 & n1260 ;
  assign n1262 = n1243 & ~n1260 ;
  assign n1263 = n1261 | n1262 ;
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  assign n1276 = n511 & ~n656 ;
  assign n1277 = ~n511 & n656 ;
  assign n1278 = n1276 | n1277 ;
  buffer buf_n1279( .i (n1278), .o (n1279) );
  buffer buf_n307( .i (N130), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  assign n1280 = n310 & n356 ;
  buffer buf_n1281( .i (n1280), .o (n1281) );
  assign n1282 = ~n392 & n624 ;
  assign n1283 = n392 & ~n624 ;
  assign n1284 = n1282 | n1283 ;
  buffer buf_n1285( .i (n1284), .o (n1285) );
  assign n1286 = n1281 & ~n1285 ;
  assign n1287 = ~n1281 & n1285 ;
  assign n1288 = n1286 | n1287 ;
  buffer buf_n1289( .i (n1288), .o (n1289) );
  assign n1290 = n1279 | n1289 ;
  assign n1291 = n1279 & n1289 ;
  assign n1292 = n1290 & ~n1291 ;
  buffer buf_n1293( .i (n1292), .o (n1293) );
  assign n1294 = n218 | n247 ;
  assign n1295 = n218 & n247 ;
  assign n1296 = n1294 & ~n1295 ;
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n158( .i (N113), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n187( .i (N117), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  assign n1298 = n160 & ~n189 ;
  assign n1299 = ~n160 & n189 ;
  assign n1300 = n1298 | n1299 ;
  buffer buf_n1301( .i (n1300), .o (n1301) );
  assign n1302 = ~n1297 & n1301 ;
  assign n1303 = n1297 & ~n1301 ;
  assign n1304 = n1302 | n1303 ;
  buffer buf_n1305( .i (n1304), .o (n1305) );
  assign n1307 = n1255 & n1305 ;
  assign n1308 = n1255 | n1305 ;
  assign n1309 = ~n1307 & n1308 ;
  buffer buf_n1310( .i (n1309), .o (n1310) );
  assign n1311 = ~n1293 & n1310 ;
  assign n1312 = n1293 & ~n1310 ;
  assign n1313 = n1311 | n1312 ;
  buffer buf_n1314( .i (n1313), .o (n1314) );
  assign n1327 = ~n1079 & n1314 ;
  buffer buf_n1328( .i (n1327), .o (n1328) );
  assign n1337 = ~n1265 & n1328 ;
  buffer buf_n1338( .i (n1337), .o (n1338) );
  assign n1345 = n1079 & ~n1314 ;
  buffer buf_n1346( .i (n1345), .o (n1346) );
  assign n1355 = ~n1265 & n1346 ;
  buffer buf_n1356( .i (n1355), .o (n1356) );
  assign n1363 = n1338 | n1356 ;
  buffer buf_n319( .i (N132), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n321( .i (n320), .o (n321) );
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  assign n1364 = n326 & n360 ;
  buffer buf_n1365( .i (n1364), .o (n1365) );
  assign n1366 = n567 & ~n712 ;
  buffer buf_n1367( .i (n566), .o (n1367) );
  buffer buf_n1368( .i (n711), .o (n1368) );
  assign n1369 = ~n1367 & n1368 ;
  assign n1370 = n1366 | n1369 ;
  buffer buf_n1371( .i (n1370), .o (n1371) );
  assign n1372 = n281 & ~n451 ;
  buffer buf_n1373( .i (n280), .o (n1373) );
  buffer buf_n1374( .i (n450), .o (n1374) );
  assign n1375 = ~n1373 & n1374 ;
  assign n1376 = n1372 | n1375 ;
  buffer buf_n1377( .i (n1376), .o (n1377) );
  assign n1378 = ~n1371 & n1377 ;
  assign n1379 = n1371 & ~n1377 ;
  assign n1380 = n1378 | n1379 ;
  buffer buf_n1381( .i (n1380), .o (n1381) );
  assign n1382 = n1365 & n1381 ;
  assign n1383 = n1365 | n1381 ;
  assign n1384 = ~n1382 & n1383 ;
  buffer buf_n1385( .i (n1384), .o (n1385) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  assign n1386 = n1071 & n1306 ;
  assign n1387 = n1071 | n1306 ;
  assign n1388 = ~n1386 & n1387 ;
  buffer buf_n1389( .i (n1388), .o (n1389) );
  assign n1390 = ~n1385 & n1389 ;
  assign n1391 = n1385 & ~n1389 ;
  assign n1392 = n1390 | n1391 ;
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  buffer buf_n1397( .i (n1396), .o (n1397) );
  assign n1405 = n1363 & ~n1397 ;
  assign n1406 = n1265 & ~n1394 ;
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  assign n1412 = ~n1266 & n1395 ;
  assign n1413 = n1407 | n1412 ;
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  assign n1414 = n1083 | n1318 ;
  assign n1415 = n1413 & ~n1414 ;
  assign n1416 = n1405 | n1415 ;
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n1003( .i (n1002), .o (n1003) );
  buffer buf_n1004( .i (n1003), .o (n1004) );
  buffer buf_n1005( .i (n1004), .o (n1005) );
  assign n1418 = ~n164 & n1005 ;
  assign n1419 = n164 & ~n1005 ;
  assign n1420 = n1418 | n1419 ;
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n327( .i (N133), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  assign n1422 = n331 & n357 ;
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n741( .i (n740), .o (n741) );
  buffer buf_n857( .i (n856), .o (n857) );
  assign n1424 = n741 & ~n857 ;
  assign n1425 = ~n741 & n857 ;
  assign n1426 = n1424 | n1425 ;
  buffer buf_n1427( .i (n1426), .o (n1427) );
  assign n1428 = n1423 & ~n1427 ;
  assign n1429 = ~n1423 & n1427 ;
  assign n1430 = n1428 | n1429 ;
  buffer buf_n1431( .i (n1430), .o (n1431) );
  assign n1432 = n1421 | n1431 ;
  assign n1433 = n1421 & n1431 ;
  assign n1434 = n1432 & ~n1433 ;
  buffer buf_n1435( .i (n1434), .o (n1435) );
  assign n1436 = n1121 & n1182 ;
  assign n1437 = n1121 | n1182 ;
  assign n1438 = ~n1436 & n1437 ;
  buffer buf_n1439( .i (n1438), .o (n1439) );
  assign n1440 = ~n1435 & n1439 ;
  assign n1441 = n1435 & ~n1439 ;
  assign n1442 = n1440 | n1441 ;
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  assign n1455 = n77 & ~n193 ;
  assign n1456 = ~n77 & n193 ;
  assign n1457 = n1455 | n1456 ;
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n332( .i (N134), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  assign n1459 = n336 & n357 ;
  buffer buf_n1460( .i (n1459), .o (n1460) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n886( .i (n885), .o (n886) );
  assign n1461 = n770 & ~n886 ;
  assign n1462 = ~n770 & n886 ;
  assign n1463 = n1461 | n1462 ;
  buffer buf_n1464( .i (n1463), .o (n1464) );
  assign n1465 = n1460 & ~n1464 ;
  assign n1466 = ~n1460 & n1464 ;
  assign n1467 = n1465 | n1466 ;
  buffer buf_n1468( .i (n1467), .o (n1468) );
  assign n1469 = n1458 | n1468 ;
  assign n1470 = n1458 & n1468 ;
  assign n1471 = n1469 & ~n1470 ;
  buffer buf_n1472( .i (n1471), .o (n1472) );
  assign n1473 = n1133 & n1194 ;
  assign n1474 = n1133 | n1194 ;
  assign n1475 = ~n1473 & n1474 ;
  buffer buf_n1476( .i (n1475), .o (n1476) );
  assign n1477 = ~n1472 & n1476 ;
  assign n1478 = n1472 & ~n1476 ;
  assign n1479 = n1477 | n1478 ;
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  assign n1492 = n1444 & ~n1481 ;
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  assign n1498 = n1417 & n1497 ;
  buffer buf_n1499( .i (n1498), .o (n1499) );
  assign n1500 = n1221 & n1499 ;
  buffer buf_n1501( .i (n1500), .o (n1501) );
  assign n1502 = n1091 & n1501 ;
  buffer buf_n1503( .i (n1502), .o (n1503) );
  assign n1504 = n70 | n1503 ;
  assign n1505 = n70 & n1503 ;
  assign n1506 = n1504 & ~n1505 ;
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  buffer buf_n632( .i (n631), .o (n632) );
  buffer buf_n633( .i (n632), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  buffer buf_n636( .i (n635), .o (n636) );
  buffer buf_n637( .i (n636), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  buffer buf_n641( .i (n640), .o (n641) );
  buffer buf_n642( .i (n641), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  buffer buf_n649( .i (n648), .o (n649) );
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n1319( .i (n1318), .o (n1319) );
  buffer buf_n1320( .i (n1319), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  buffer buf_n1323( .i (n1322), .o (n1323) );
  buffer buf_n1324( .i (n1323), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  assign n1507 = n1326 & n1501 ;
  buffer buf_n1508( .i (n1507), .o (n1508) );
  assign n1509 = n650 | n1508 ;
  assign n1510 = n650 & n1508 ;
  assign n1511 = n1509 & ~n1510 ;
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n946( .i (n945), .o (n946) );
  buffer buf_n947( .i (n946), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n950( .i (n949), .o (n950) );
  buffer buf_n951( .i (n950), .o (n951) );
  buffer buf_n952( .i (n951), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  assign n1512 = n1275 & n1501 ;
  buffer buf_n1513( .i (n1512), .o (n1513) );
  assign n1514 = n969 & n1513 ;
  assign n1515 = n969 | n1513 ;
  assign n1516 = ~n1514 & n1515 ;
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  buffer buf_n284( .i (n283), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  buffer buf_n291( .i (n290), .o (n291) );
  buffer buf_n292( .i (n291), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n1398( .i (n1397), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  assign n1517 = n1404 & n1501 ;
  buffer buf_n1518( .i (n1517), .o (n1518) );
  assign n1519 = ~n306 & n1518 ;
  assign n1520 = n306 & ~n1518 ;
  assign n1521 = n1519 | n1520 ;
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  assign n1522 = ~n1142 & n1203 ;
  buffer buf_n1523( .i (n1522), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  assign n1530 = n1499 & n1529 ;
  buffer buf_n1531( .i (n1530), .o (n1531) );
  assign n1532 = n1091 & n1531 ;
  buffer buf_n1533( .i (n1532), .o (n1533) );
  assign n1534 = n389 | n1533 ;
  assign n1535 = n389 & n1533 ;
  assign n1536 = n1534 & ~n1535 ;
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  buffer buf_n401( .i (n400), .o (n401) );
  buffer buf_n402( .i (n401), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n407( .i (n406), .o (n407) );
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  assign n1537 = n1326 & n1531 ;
  buffer buf_n1538( .i (n1537), .o (n1538) );
  assign n1539 = n418 | n1538 ;
  assign n1540 = n418 & n1538 ;
  assign n1541 = n1539 & ~n1540 ;
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  assign n1542 = n1275 & n1531 ;
  buffer buf_n1543( .i (n1542), .o (n1543) );
  assign n1544 = n447 & n1543 ;
  assign n1545 = n447 | n1543 ;
  assign n1546 = ~n1544 & n1545 ;
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  assign n1547 = n1404 & n1531 ;
  buffer buf_n1548( .i (n1547), .o (n1548) );
  assign n1549 = ~n476 & n1548 ;
  assign n1550 = n476 & ~n1548 ;
  assign n1551 = n1549 | n1550 ;
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  assign n1552 = ~n1444 & n1481 ;
  buffer buf_n1553( .i (n1552), .o (n1553) );
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n1556( .i (n1555), .o (n1556) );
  buffer buf_n1557( .i (n1556), .o (n1557) );
  assign n1558 = n1417 & n1557 ;
  buffer buf_n1559( .i (n1558), .o (n1559) );
  assign n1560 = n1221 & n1559 ;
  buffer buf_n1561( .i (n1560), .o (n1561) );
  assign n1562 = n1091 & n1561 ;
  buffer buf_n1563( .i (n1562), .o (n1563) );
  assign n1564 = n505 | n1563 ;
  assign n1565 = n505 & n1563 ;
  assign n1566 = n1564 & ~n1565 ;
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  assign n1567 = n1326 & n1561 ;
  buffer buf_n1568( .i (n1567), .o (n1568) );
  assign n1569 = n534 | n1568 ;
  assign n1570 = n534 & n1568 ;
  assign n1571 = n1569 & ~n1570 ;
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  assign n1572 = n1275 & n1561 ;
  buffer buf_n1573( .i (n1572), .o (n1573) );
  assign n1574 = n563 & n1573 ;
  assign n1575 = n563 | n1573 ;
  assign n1576 = ~n1574 & n1575 ;
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  buffer buf_n579( .i (n578), .o (n579) );
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  buffer buf_n589( .i (n588), .o (n589) );
  buffer buf_n590( .i (n589), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  assign n1577 = n1404 & n1561 ;
  buffer buf_n1578( .i (n1577), .o (n1578) );
  assign n1579 = n592 | n1578 ;
  assign n1580 = n592 & n1578 ;
  assign n1581 = n1579 & ~n1580 ;
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  assign n1582 = n1529 & n1559 ;
  buffer buf_n1583( .i (n1582), .o (n1583) );
  assign n1584 = n1091 & n1583 ;
  buffer buf_n1585( .i (n1584), .o (n1585) );
  assign n1586 = n621 | n1585 ;
  assign n1587 = n621 & n1585 ;
  assign n1588 = n1586 & ~n1587 ;
  buffer buf_n657( .i (n656), .o (n657) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n659( .i (n658), .o (n659) );
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  assign n1589 = n1326 & n1583 ;
  buffer buf_n1590( .i (n1589), .o (n1590) );
  assign n1591 = n679 | n1590 ;
  assign n1592 = n679 & n1590 ;
  assign n1593 = n1591 & ~n1592 ;
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  buffer buf_n688( .i (n687), .o (n688) );
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n692( .i (n691), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  buffer buf_n702( .i (n701), .o (n702) );
  buffer buf_n703( .i (n702), .o (n703) );
  buffer buf_n704( .i (n703), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  assign n1594 = n1275 & n1583 ;
  buffer buf_n1595( .i (n1594), .o (n1595) );
  assign n1596 = n708 & n1595 ;
  assign n1597 = n708 | n1595 ;
  assign n1598 = ~n1596 & n1597 ;
  buffer buf_n713( .i (n712), .o (n713) );
  buffer buf_n714( .i (n713), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n718( .i (n717), .o (n718) );
  buffer buf_n719( .i (n718), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n722( .i (n721), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n732( .i (n731), .o (n732) );
  buffer buf_n733( .i (n732), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n737( .i (n736), .o (n737) );
  assign n1599 = n1404 & n1583 ;
  buffer buf_n1600( .i (n1599), .o (n1600) );
  assign n1601 = n737 & n1600 ;
  assign n1602 = n737 | n1600 ;
  assign n1603 = ~n1601 & n1602 ;
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n746( .i (n745), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  buffer buf_n748( .i (n747), .o (n748) );
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n1448( .i (n1447), .o (n1448) );
  buffer buf_n1449( .i (n1448), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  buffer buf_n1347( .i (n1346), .o (n1347) );
  buffer buf_n1348( .i (n1347), .o (n1348) );
  buffer buf_n1349( .i (n1348), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  assign n1604 = n1493 | n1553 ;
  buffer buf_n1143( .i (n1142), .o (n1143) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1204( .i (n1203), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  assign n1605 = n1144 | n1205 ;
  assign n1606 = n1604 & ~n1605 ;
  assign n1607 = n1215 | n1523 ;
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  assign n1608 = n1446 | n1483 ;
  assign n1609 = n1607 & ~n1608 ;
  assign n1610 = n1606 | n1609 ;
  buffer buf_n1611( .i (n1610), .o (n1611) );
  assign n1612 = n1411 & n1611 ;
  buffer buf_n1613( .i (n1612), .o (n1613) );
  assign n1614 = n1354 & n1613 ;
  buffer buf_n1615( .i (n1614), .o (n1615) );
  assign n1616 = n1454 & n1615 ;
  buffer buf_n1617( .i (n1616), .o (n1617) );
  assign n1618 = n766 | n1617 ;
  assign n1619 = n766 & n1617 ;
  assign n1620 = n1618 & ~n1619 ;
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n773( .i (n772), .o (n773) );
  buffer buf_n774( .i (n773), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n1484( .i (n1483), .o (n1484) );
  buffer buf_n1485( .i (n1484), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n1488( .i (n1487), .o (n1488) );
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  assign n1621 = n1491 & n1615 ;
  buffer buf_n1622( .i (n1621), .o (n1622) );
  assign n1623 = n795 | n1622 ;
  assign n1624 = n795 & n1622 ;
  assign n1625 = n1623 & ~n1624 ;
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  buffer buf_n804( .i (n803), .o (n804) );
  buffer buf_n805( .i (n804), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  buffer buf_n810( .i (n809), .o (n810) );
  buffer buf_n811( .i (n810), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n815( .i (n814), .o (n815) );
  buffer buf_n816( .i (n815), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n822( .i (n821), .o (n822) );
  buffer buf_n823( .i (n822), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n1151( .i (n1150), .o (n1151) );
  buffer buf_n1152( .i (n1151), .o (n1152) );
  assign n1626 = n1152 & n1615 ;
  buffer buf_n1627( .i (n1626), .o (n1627) );
  assign n1628 = ~n824 & n1627 ;
  assign n1629 = n824 & ~n1627 ;
  assign n1630 = n1628 | n1629 ;
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  buffer buf_n832( .i (n831), .o (n832) );
  buffer buf_n833( .i (n832), .o (n833) );
  buffer buf_n834( .i (n833), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n839( .i (n838), .o (n839) );
  buffer buf_n840( .i (n839), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  buffer buf_n844( .i (n843), .o (n844) );
  buffer buf_n845( .i (n844), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  assign n1631 = n1213 & n1615 ;
  buffer buf_n1632( .i (n1631), .o (n1632) );
  assign n1633 = n853 & n1632 ;
  assign n1634 = n853 | n1632 ;
  assign n1635 = ~n1633 & n1634 ;
  buffer buf_n858( .i (n857), .o (n858) );
  buffer buf_n859( .i (n858), .o (n859) );
  buffer buf_n860( .i (n859), .o (n860) );
  buffer buf_n861( .i (n860), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  assign n1636 = n1400 & n1611 ;
  buffer buf_n1637( .i (n1636), .o (n1637) );
  assign n1638 = n1362 & n1637 ;
  buffer buf_n1639( .i (n1638), .o (n1639) );
  assign n1640 = n1454 & n1639 ;
  buffer buf_n1641( .i (n1640), .o (n1641) );
  assign n1642 = n882 | n1641 ;
  assign n1643 = n882 & n1641 ;
  assign n1644 = n1642 & ~n1643 ;
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n891( .i (n890), .o (n891) );
  buffer buf_n892( .i (n891), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  assign n1645 = n1491 & n1639 ;
  buffer buf_n1646( .i (n1645), .o (n1646) );
  assign n1647 = n911 | n1646 ;
  assign n1648 = n911 & n1646 ;
  assign n1649 = n1647 & ~n1648 ;
  buffer buf_n916( .i (n915), .o (n916) );
  buffer buf_n917( .i (n916), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  buffer buf_n921( .i (n920), .o (n921) );
  buffer buf_n922( .i (n921), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  assign n1650 = n1152 & n1639 ;
  buffer buf_n1651( .i (n1650), .o (n1651) );
  assign n1652 = n940 & n1651 ;
  assign n1653 = n940 | n1651 ;
  assign n1654 = ~n1652 & n1653 ;
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n976( .i (n975), .o (n976) );
  buffer buf_n977( .i (n976), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  buffer buf_n985( .i (n984), .o (n985) );
  buffer buf_n986( .i (n985), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  buffer buf_n991( .i (n990), .o (n991) );
  buffer buf_n992( .i (n991), .o (n992) );
  buffer buf_n993( .i (n992), .o (n993) );
  buffer buf_n994( .i (n993), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  assign n1655 = n1213 & n1639 ;
  buffer buf_n1656( .i (n1655), .o (n1656) );
  assign n1657 = n998 | n1656 ;
  assign n1658 = n998 & n1656 ;
  assign n1659 = n1657 & ~n1658 ;
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n1017( .i (n1016), .o (n1017) );
  buffer buf_n1018( .i (n1017), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1027( .i (n1026), .o (n1027) );
  buffer buf_n1329( .i (n1328), .o (n1329) );
  buffer buf_n1330( .i (n1329), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  buffer buf_n1332( .i (n1331), .o (n1332) );
  buffer buf_n1333( .i (n1332), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  assign n1660 = n1336 & n1613 ;
  buffer buf_n1661( .i (n1660), .o (n1661) );
  assign n1662 = n1454 & n1661 ;
  buffer buf_n1663( .i (n1662), .o (n1663) );
  assign n1664 = n1027 | n1663 ;
  assign n1665 = n1027 & n1663 ;
  assign n1666 = n1664 & ~n1665 ;
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  assign n1667 = n1491 & n1661 ;
  buffer buf_n1668( .i (n1667), .o (n1668) );
  assign n1669 = n99 | n1668 ;
  assign n1670 = n99 & n1668 ;
  assign n1671 = n1669 & ~n1670 ;
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  assign n1672 = n1152 & n1661 ;
  buffer buf_n1673( .i (n1672), .o (n1673) );
  assign n1674 = ~n128 & n1673 ;
  assign n1675 = n128 & ~n1673 ;
  assign n1676 = n1674 | n1675 ;
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  assign n1677 = n1213 & n1661 ;
  buffer buf_n1678( .i (n1677), .o (n1678) );
  assign n1679 = n157 & n1678 ;
  assign n1680 = n157 | n1678 ;
  assign n1681 = ~n1679 & n1680 ;
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  buffer buf_n1342( .i (n1341), .o (n1342) );
  buffer buf_n1343( .i (n1342), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  assign n1682 = n1344 & n1637 ;
  buffer buf_n1683( .i (n1682), .o (n1683) );
  assign n1684 = n1454 & n1683 ;
  buffer buf_n1685( .i (n1684), .o (n1685) );
  assign n1686 = n186 | n1685 ;
  assign n1687 = n186 & n1685 ;
  assign n1688 = n1686 & ~n1687 ;
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  assign n1689 = n1491 & n1683 ;
  buffer buf_n1690( .i (n1689), .o (n1690) );
  assign n1691 = n215 | n1690 ;
  assign n1692 = n215 & n1690 ;
  assign n1693 = n1691 & ~n1692 ;
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  assign n1694 = n1152 & n1683 ;
  buffer buf_n1695( .i (n1694), .o (n1695) );
  assign n1696 = n244 & n1695 ;
  assign n1697 = n244 | n1695 ;
  assign n1698 = ~n1696 & n1697 ;
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  assign n1699 = n1213 & n1683 ;
  buffer buf_n1700( .i (n1699), .o (n1700) );
  assign n1701 = n273 | n1700 ;
  assign n1702 = n273 & n1700 ;
  assign n1703 = n1701 & ~n1702 ;
  assign N724 = n1506 ;
  assign N725 = n1511 ;
  assign N726 = n1516 ;
  assign N727 = n1521 ;
  assign N728 = n1536 ;
  assign N729 = n1541 ;
  assign N730 = n1546 ;
  assign N731 = n1551 ;
  assign N732 = n1566 ;
  assign N733 = n1571 ;
  assign N734 = n1576 ;
  assign N735 = n1581 ;
  assign N736 = n1588 ;
  assign N737 = n1593 ;
  assign N738 = n1598 ;
  assign N739 = n1603 ;
  assign N740 = n1620 ;
  assign N741 = n1625 ;
  assign N742 = n1630 ;
  assign N743 = n1635 ;
  assign N744 = n1644 ;
  assign N745 = n1649 ;
  assign N746 = n1654 ;
  assign N747 = n1659 ;
  assign N748 = n1666 ;
  assign N749 = n1671 ;
  assign N750 = n1676 ;
  assign N751 = n1681 ;
  assign N752 = n1688 ;
  assign N753 = n1693 ;
  assign N754 = n1698 ;
  assign N755 = n1703 ;
endmodule
