module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n113 , n114 , n115 , n116 , n117 , n118 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 ;
  buffer buf_n76( .i (x7), .o (n76) );
  buffer buf_n86( .i (x8), .o (n86) );
  assign n156 = n76 & n86 ;
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n102( .i (x9), .o (n102) );
  buffer buf_n113( .i (x10), .o (n113) );
  assign n158 = n102 & n113 ;
  buffer buf_n159( .i (n158), .o (n159) );
  assign n160 = n157 & n159 ;
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n137( .i (x12), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  assign n165 = n78 & ~n139 ;
  buffer buf_n166( .i (n165), .o (n166) );
  assign n168 = ~n161 & n166 ;
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  assign n170 = n89 | n116 ;
  buffer buf_n171( .i (n170), .o (n171) );
  assign n172 = n102 | n113 ;
  buffer buf_n173( .i (n172), .o (n173) );
  assign n175 = n157 & ~n173 ;
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n177( .i (n176), .o (n177) );
  assign n180 = n171 & ~n177 ;
  assign n181 = n169 & n180 ;
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n90( .i (n89), .o (n90) );
  assign n188 = ~n80 & n90 ;
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n120( .i (x11), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  assign n191 = ~n103 & n121 ;
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  assign n195 = n118 | n194 ;
  assign n196 = n189 & n195 ;
  buffer buf_n122( .i (n121), .o (n122) );
  assign n197 = n115 & n122 ;
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  assign n201 = n79 & n105 ;
  assign n202 = ~n198 & n201 ;
  buffer buf_n203( .i (n202), .o (n203) );
  assign n204 = ~n143 & n203 ;
  assign n205 = ( ~n144 & n196 ) | ( ~n144 & n204 ) | ( n196 & n204 ) ;
  assign n206 = n182 | n205 ;
  buffer buf_n207( .i (n206), .o (n207) );
  buffer buf_n208( .i (n207), .o (n208) );
  buffer buf_n209( .i (n208), .o (n209) );
  buffer buf_n44( .i (x4), .o (n44) );
  buffer buf_n45( .i (n44), .o (n45) );
  buffer buf_n46( .i (n45), .o (n46) );
  buffer buf_n47( .i (n46), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n19( .i (x2), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n33( .i (x3), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n146( .i (x13), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  buffer buf_n148( .i (n147), .o (n148) );
  assign n210 = n35 | n148 ;
  buffer buf_n211( .i (n210), .o (n211) );
  assign n212 = n23 & n211 ;
  buffer buf_n65( .i (x6), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  assign n213 = n20 | n34 ;
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  assign n222 = n69 | n215 ;
  assign n223 = ~n212 & n222 ;
  assign n224 = n50 & ~n223 ;
  buffer buf_n9( .i (x1), .o (n9) );
  assign n225 = ~n9 & n146 ;
  buffer buf_n226( .i (n225), .o (n226) );
  assign n230 = n21 & ~n226 ;
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n149( .i (n148), .o (n149) );
  assign n233 = n12 & n149 ;
  buffer buf_n234( .i (n233), .o (n234) );
  assign n236 = n232 | n234 ;
  buffer buf_n55( .i (x5), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  assign n237 = n67 & n148 ;
  buffer buf_n238( .i (n237), .o (n238) );
  assign n239 = n35 | n46 ;
  buffer buf_n240( .i (n239), .o (n240) );
  assign n244 = n238 & ~n240 ;
  assign n245 = n60 & ~n244 ;
  assign n246 = n236 & n245 ;
  assign n247 = ~n224 & n246 ;
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  assign n248 = ~n37 & n238 ;
  assign n249 = n232 & n248 ;
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  assign n252 = n247 | n251 ;
  buffer buf_n253( .i (n252), .o (n253) );
  assign n254 = n45 & ~n56 ;
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  assign n258 = n211 & n256 ;
  assign n259 = n232 & n258 ;
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  assign n264 = n253 | n263 ;
  buffer buf_n265( .i (n264), .o (n265) );
  assign n266 = n209 & n265 ;
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  assign n267 = n4 & n35 ;
  buffer buf_n268( .i (n267), .o (n268) );
  assign n269 = ( ~n13 & n48 ) | ( ~n13 & n268 ) | ( n48 & n268 ) ;
  assign n270 = ( n13 & n48 ) | ( n13 & n268 ) | ( n48 & n268 ) ;
  assign n271 = ~n269 & n270 ;
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n275( .i (n274), .o (n275) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  assign n278 = n69 & n80 ;
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  assign n281 = n77 | n114 ;
  buffer buf_n282( .i (n281), .o (n282) );
  buffer buf_n283( .i (n282), .o (n283) );
  assign n284 = n124 | n283 ;
  buffer buf_n285( .i (n284), .o (n285) );
  assign n286 = ~n279 & n285 ;
  buffer buf_n91( .i (n90), .o (n91) );
  assign n287 = n66 & n103 ;
  buffer buf_n288( .i (n287), .o (n288) );
  assign n289 = n77 & n114 ;
  buffer buf_n290( .i (n289), .o (n290) );
  assign n291 = ~n288 & n290 ;
  buffer buf_n292( .i (n291), .o (n292) );
  assign n295 = n91 & ~n292 ;
  assign n296 = ~n203 & n295 ;
  assign n297 = ~n286 & n296 ;
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n70( .i (n69), .o (n70) );
  assign n299 = n105 & ~n116 ;
  buffer buf_n300( .i (n299), .o (n300) );
  assign n302 = n69 | n80 ;
  assign n303 = ( n70 & ~n300 ) | ( n70 & n302 ) | ( ~n300 & n302 ) ;
  buffer buf_n125( .i (n124), .o (n125) );
  assign n304 = n76 | n86 ;
  buffer buf_n305( .i (n304), .o (n305) );
  assign n309 = n159 & ~n305 ;
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n174( .i (n173), .o (n174) );
  assign n315 = n123 | n174 ;
  buffer buf_n316( .i (n315), .o (n316) );
  assign n317 = ( n125 & ~n311 ) | ( n125 & n316 ) | ( ~n311 & n316 ) ;
  assign n318 = n303 & n317 ;
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n306( .i (n305), .o (n306) );
  assign n321 = n192 & ~n306 ;
  buffer buf_n322( .i (n321), .o (n322) );
  assign n323 = n138 & ~n147 ;
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  assign n329 = ~n322 & n326 ;
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  assign n332 = n319 & n331 ;
  assign n333 = ~n298 & n332 ;
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  assign n336 = n277 & n335 ;
  assign n337 = n266 | n336 ;
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  assign n340 = ~n20 & n34 ;
  buffer buf_n341( .i (n340), .o (n341) );
  assign n342 = n56 & ~n147 ;
  buffer buf_n343( .i (n342), .o (n343) );
  assign n344 = n341 & n343 ;
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  assign n348 = n260 | n347 ;
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  assign n349 = n20 & ~n45 ;
  buffer buf_n350( .i (n349), .o (n350) );
  assign n354 = n58 & n350 ;
  buffer buf_n355( .i (n354), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  assign n358 = n22 & n58 ;
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n241( .i (n240), .o (n241) );
  assign n362 = ~n234 & n241 ;
  assign n363 = n360 & n362 ;
  assign n364 = ( n153 & n357 ) | ( n153 & n363 ) | ( n357 & n363 ) ;
  assign n365 = n348 | n364 ;
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  assign n369 = n209 & n368 ;
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  assign n370 = n42 & n274 ;
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  assign n371 = n6 & ~n13 ;
  assign n372 = n355 & n371 ;
  assign n373 = n255 & n341 ;
  buffer buf_n374( .i (n373), .o (n374) );
  assign n375 = ~n10 & n45 ;
  buffer buf_n376( .i (n375), .o (n376) );
  assign n380 = n22 & ~n376 ;
  assign n381 = n268 & ~n380 ;
  assign n382 = ~n374 & n381 ;
  assign n383 = n372 | n382 ;
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  assign n387 = n370 | n386 ;
  buffer buf_n388( .i (n387), .o (n388) );
  assign n389 = n335 & n388 ;
  assign n390 = n369 | n389 ;
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  assign n393 = n56 | n66 ;
  buffer buf_n394( .i (n393), .o (n394) );
  assign n396 = ~n255 & n394 ;
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  assign n399 = ~n21 & n148 ;
  buffer buf_n400( .i (n399), .o (n400) );
  assign n402 = n231 | n400 ;
  buffer buf_n403( .i (n402), .o (n403) );
  assign n404 = n398 | n403 ;
  buffer buf_n257( .i (n256), .o (n257) );
  assign n405 = n215 | n256 ;
  assign n406 = ( ~n232 & n257 ) | ( ~n232 & n405 ) | ( n257 & n405 ) ;
  buffer buf_n401( .i (n400), .o (n401) );
  assign n407 = ~n68 & n214 ;
  buffer buf_n408( .i (n407), .o (n408) );
  buffer buf_n409( .i (n12), .o (n409) );
  assign n410 = n400 & ~n409 ;
  assign n411 = ( n401 & n408 ) | ( n401 & n410 ) | ( n408 & n410 ) ;
  assign n412 = n406 & ~n411 ;
  assign n413 = n404 & n412 ;
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  assign n416 = n253 | n415 ;
  buffer buf_n417( .i (n416), .o (n417) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  assign n418 = n25 | n50 ;
  buffer buf_n61( .i (n60), .o (n61) );
  assign n419 = n50 & n61 ;
  assign n420 = ( n25 & ~n61 ) | ( n25 & n152 ) | ( ~n61 & n152 ) ;
  assign n421 = ( ~n418 & n419 ) | ( ~n418 & n420 ) | ( n419 & n420 ) ;
  buffer buf_n422( .i (n421), .o (n422) );
  assign n423 = n53 | n422 ;
  assign n424 = n207 & n423 ;
  buffer buf_n425( .i (n424), .o (n425) );
  assign n426 = n417 & n425 ;
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n7( .i (n6), .o (n7) );
  assign n429 = n7 & ~n374 ;
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  assign n431 = ( ~n14 & n60 ) | ( ~n14 & n216 ) | ( n60 & n216 ) ;
  assign n432 = ~n217 & n431 ;
  assign n433 = ( n16 & n430 ) | ( n16 & ~n432 ) | ( n430 & ~n432 ) ;
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  assign n434 = n5 & n12 ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n437 = n359 & n435 ;
  assign n438 = n327 & ~n437 ;
  assign n439 = ( n272 & n328 ) | ( n272 & n438 ) | ( n328 & n438 ) ;
  assign n440 = n433 & n439 ;
  assign n441 = ~n36 & n58 ;
  assign n442 = n48 | n441 ;
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  assign n445 = n39 | n443 ;
  assign n446 = ( n272 & n444 ) | ( n272 & n445 ) | ( n444 & n445 ) ;
  assign n447 = n384 | n446 ;
  assign n448 = n440 & n447 ;
  buffer buf_n449( .i (n448), .o (n449) );
  assign n452 = n334 & n449 ;
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n242( .i (n241), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  assign n456 = ~n16 & n243 ;
  assign n457 = ( n16 & ~n243 ) | ( n16 & n272 ) | ( ~n243 & n272 ) ;
  assign n458 = ( n63 & n456 ) | ( n63 & n457 ) | ( n456 & n457 ) ;
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  assign n464 = n427 | n463 ;
  assign n465 = ( n428 & n455 ) | ( n428 & n464 ) | ( n455 & n464 ) ;
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n361( .i (n360), .o (n361) );
  assign n466 = ~n72 & n361 ;
  buffer buf_n467( .i (n466), .o (n467) );
  assign n468 = n414 | n467 ;
  assign n469 = n253 | n468 ;
  buffer buf_n470( .i (n469), .o (n470) );
  assign n472 = n209 & n470 ;
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n17( .i (n16), .o (n17) );
  assign n474 = ~n17 & n73 ;
  assign n475 = ( n74 & ~n422 ) | ( n74 & n474 ) | ( ~n422 & n474 ) ;
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  assign n480 = n473 & n479 ;
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n320( .i (n319), .o (n320) );
  assign n481 = ~n298 & n320 ;
  assign n482 = n96 & n481 ;
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  assign n485 = n451 & n484 ;
  buffer buf_n486( .i (n485), .o (n486) );
  assign n487 = n480 | n486 ;
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n471( .i (n470), .o (n471) );
  assign n488 = n187 & n471 ;
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  buffer buf_n109( .i (n108), .o (n109) );
  buffer buf_n190( .i (n189), .o (n190) );
  assign n489 = n109 & ~n190 ;
  assign n490 = n67 & n115 ;
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  assign n495 = ~n322 & n492 ;
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  assign n498 = ~n489 & n497 ;
  buffer buf_n199( .i (n198), .o (n199) );
  assign n499 = n288 & ~n290 ;
  buffer buf_n500( .i (n499), .o (n500) );
  assign n501 = n199 & n500 ;
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n301( .i (n300), .o (n301) );
  assign n504 = ~n91 & n125 ;
  assign n505 = n301 | n504 ;
  assign n506 = n280 & n505 ;
  assign n507 = n503 | n506 ;
  assign n508 = n498 | n507 ;
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  assign n512 = n451 & n511 ;
  assign n513 = n488 | n512 ;
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  assign n515 = n279 & n301 ;
  assign n516 = n294 | n515 ;
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n519( .i (n518), .o (n519) );
  buffer buf_n520( .i (n519), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  assign n522 = n451 & n521 ;
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n178( .i (n177), .o (n178) );
  assign n524 = n169 & ~n178 ;
  assign n525 = n118 & ~n142 ;
  assign n526 = n189 & n525 ;
  assign n527 = n524 | n526 ;
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  assign n532 = n470 & n531 ;
  buffer buf_n533( .i (n532), .o (n533) );
  assign n534 = n100 & n533 ;
  assign n535 = n523 | n534 ;
  assign n536 = ~n106 & n283 ;
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  buffer buf_n541( .i (n540), .o (n541) );
  buffer buf_n542( .i (n541), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n545( .i (n544), .o (n545) );
  buffer buf_n546( .i (n545), .o (n546) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n200( .i (n199), .o (n200) );
  assign n547 = n82 & ~n200 ;
  assign n548 = n494 & n547 ;
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  assign n554 = n453 & ~n553 ;
  buffer buf_n555( .i (n554), .o (n555) );
  assign n556 = n533 & ~n545 ;
  assign n557 = ( ~n546 & n555 ) | ( ~n546 & n556 ) | ( n555 & n556 ) ;
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  assign n558 = n282 & ~n288 ;
  buffer buf_n559( .i (n558), .o (n559) );
  assign n560 = n500 | n559 ;
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n566( .i (n565), .o (n566) );
  buffer buf_n567( .i (n566), .o (n567) );
  assign n568 = n453 & n567 ;
  buffer buf_n569( .i (n568), .o (n569) );
  assign n570 = n134 & n473 ;
  assign n571 = ( n135 & n569 ) | ( n135 & n570 ) | ( n569 & n570 ) ;
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  assign n572 = n140 | n149 ;
  assign n573 = n215 | n572 ;
  buffer buf_n395( .i (n394), .o (n395) );
  assign n574 = n88 & ~n115 ;
  buffer buf_n575( .i (n574), .o (n575) );
  assign n576 = n395 | n575 ;
  assign n577 = n573 | n576 ;
  buffer buf_n162( .i (n161), .o (n162) );
  assign n578 = n125 & n162 ;
  assign n579 = ( n285 & n577 ) | ( n285 & ~n578 ) | ( n577 & ~n578 ) ;
  buffer buf_n580( .i (n579), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  assign n583 = ~n4 & n11 ;
  assign n584 = n324 & n583 ;
  buffer buf_n585( .i (n584), .o (n585) );
  buffer buf_n586( .i (n585), .o (n586) );
  assign n587 = n23 & n491 ;
  assign n588 = n322 & n587 ;
  assign n589 = n586 & n588 ;
  assign n590 = n176 | n310 ;
  buffer buf_n591( .i (n590), .o (n591) );
  assign n594 = ~n21 & n46 ;
  assign n595 = n123 & n594 ;
  assign n596 = n66 & ~n138 ;
  buffer buf_n597( .i (n596), .o (n597) );
  assign n600 = n343 & n597 ;
  assign n601 = n595 & n600 ;
  buffer buf_n602( .i (n601), .o (n602) );
  assign n603 = n591 & n602 ;
  assign n604 = n589 | n603 ;
  buffer buf_n605( .i (n604), .o (n605) );
  assign n606 = n581 & ~n605 ;
  assign n607 = n221 | n606 ;
  buffer buf_n608( .i (n607), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n26( .i (n25), .o (n26) );
  buffer buf_n27( .i (n26), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  assign n610 = ~n31 & n608 ;
  assign n611 = ( ~n453 & n609 ) | ( ~n453 & n610 ) | ( n609 & n610 ) ;
  buffer buf_n612( .i (n611), .o (n612) );
  buffer buf_n613( .i (n612), .o (n613) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  assign n614 = n38 & n257 ;
  assign n615 = n378 | n435 ;
  assign n616 = ( n379 & ~n614 ) | ( n379 & n615 ) | ( ~n614 & n615 ) ;
  buffer buf_n617( .i (n616), .o (n617) );
  buffer buf_n618( .i (n617), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  assign n621 = n334 & n620 ;
  assign n622 = n450 & n621 ;
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n598( .i (n597), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  assign n623 = ~n397 & n599 ;
  assign n624 = ~n403 & n623 ;
  buffer buf_n625( .i (n624), .o (n625) );
  assign n626 = n314 & n625 ;
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n351( .i (n350), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  assign n628 = n353 & n591 ;
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n124), .o (n631) );
  assign n632 = n216 & n631 ;
  assign n633 = n37 | n124 ;
  buffer buf_n634( .i (n47), .o (n634) );
  assign n635 = n117 & n634 ;
  assign n636 = ( n49 & ~n633 ) | ( n49 & n635 ) | ( ~n633 & n635 ) ;
  assign n637 = n632 | n636 ;
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n640( .i (n57), .o (n640) );
  assign n641 = n227 | n640 ;
  assign n642 = n598 & ~n641 ;
  buffer buf_n643( .i (n642), .o (n643) );
  buffer buf_n644( .i (n643), .o (n644) );
  buffer buf_n645( .i (n644), .o (n645) );
  assign n646 = n638 & ~n645 ;
  assign n647 = ( ~n630 & n639 ) | ( ~n630 & n646 ) | ( n639 & n646 ) ;
  assign n648 = ~n627 & n647 ;
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  assign n649 = n300 & ~n308 ;
  assign n650 = n359 & n599 ;
  assign n651 = n649 & n650 ;
  assign n652 = n36 & n123 ;
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  assign n657 = n651 | n655 ;
  assign n658 = n580 & ~n657 ;
  assign n659 = ~n605 & n658 ;
  buffer buf_n660( .i (n659), .o (n660) );
  assign n663 = n648 | n660 ;
  assign n664 = n417 | n663 ;
  assign n665 = ~n622 & n664 ;
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  assign n666 = n42 & n155 ;
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  assign n669 = n209 & n668 ;
  assign n670 = n471 & n669 ;
  assign n671 = n665 & ~n670 ;
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n83( .i (n82), .o (n83) );
  assign n673 = ~n51 & n83 ;
  buffer buf_n674( .i (n673), .o (n674) );
  assign n675 = n111 & ~n674 ;
  assign n676 = n582 | n675 ;
  assign n677 = n311 | n653 ;
  assign n678 = ( n602 & n654 ) | ( n602 & n677 ) | ( n654 & n677 ) ;
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  assign n683 = n676 & ~n682 ;
  buffer buf_n179( .i (n178), .o (n179) );
  assign n684 = n189 & n301 ;
  assign n685 = n179 | n684 ;
  assign n686 = n625 & n685 ;
  buffer buf_n687( .i (n686), .o (n687) );
  assign n688 = n67 | n104 ;
  buffer buf_n689( .i (n688), .o (n689) );
  assign n692 = n59 & n689 ;
  assign n693 = n585 & n692 ;
  assign n694 = n643 | n693 ;
  assign n695 = n351 & n575 ;
  assign n696 = n559 & n695 ;
  buffer buf_n697( .i (n696), .o (n697) );
  assign n698 = n694 & n697 ;
  buffer buf_n699( .i (n698), .o (n699) );
  assign n702 = n40 & ~n644 ;
  assign n703 = ( n41 & ~n629 ) | ( n41 & n702 ) | ( ~n629 & n702 ) ;
  assign n704 = ~n699 & n703 ;
  assign n705 = ~n687 & n704 ;
  buffer buf_n706( .i (n705), .o (n706) );
  assign n707 = n683 | n706 ;
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n710( .i (n709), .o (n710) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  assign n711 = n593 & n625 ;
  buffer buf_n712( .i (n711), .o (n712) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n235( .i (n234), .o (n235) );
  assign n713 = ~n235 & n353 ;
  assign n714 = n655 & ~n713 ;
  buffer buf_n690( .i (n689), .o (n690) );
  buffer buf_n691( .i (n690), .o (n691) );
  buffer buf_n167( .i (n166), .o (n167) );
  assign n715 = n167 & ~n171 ;
  assign n716 = ~n691 & n715 ;
  buffer buf_n717( .i (n716), .o (n717) );
  assign n718 = ( n656 & n714 ) | ( n656 & ~n717 ) | ( n714 & ~n717 ) ;
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  assign n719 = n49 & ~n229 ;
  assign n720 = n360 & n719 ;
  buffer buf_n721( .i (n720), .o (n721) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n436( .i (n435), .o (n436) );
  assign n722 = n141 & n150 ;
  buffer buf_n723( .i (n722), .o (n723) );
  assign n730 = ( n143 & ~n436 ) | ( n143 & n723 ) | ( ~n436 & n723 ) ;
  assign n731 = n164 & ~n730 ;
  assign n732 = n721 & n731 ;
  assign n733 = n718 & ~n732 ;
  assign n734 = ~n712 & n733 ;
  buffer buf_n735( .i (n734), .o (n735) );
  assign n736 = n73 & n679 ;
  buffer buf_n84( .i (n83), .o (n84) );
  assign n737 = ( n52 & ~n84 ) | ( n52 & n580 ) | ( ~n84 & n580 ) ;
  assign n738 = ( n674 & ~n736 ) | ( n674 & n737 ) | ( ~n736 & n737 ) ;
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  buffer buf_n700( .i (n699), .o (n700) );
  buffer buf_n701( .i (n700), .o (n701) );
  assign n741 = n701 & ~n739 ;
  assign n742 = ( n735 & n740 ) | ( n735 & ~n741 ) | ( n740 & ~n741 ) ;
  buffer buf_n743( .i (n742), .o (n743) );
  buffer buf_n744( .i (n743), .o (n744) );
  buffer buf_n745( .i (n744), .o (n745) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  assign n746 = n470 | n735 ;
  assign n747 = ~n706 & n735 ;
  assign n748 = ( n662 & n746 ) | ( n662 & ~n747 ) | ( n746 & ~n747 ) ;
  buffer buf_n749( .i (n748), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n728( .i (n727), .o (n728) );
  buffer buf_n729( .i (n728), .o (n729) );
  assign n751 = n334 | n728 ;
  assign n752 = ( n450 & n729 ) | ( n450 & n751 ) | ( n729 & n751 ) ;
  buffer buf_n753( .i (n752), .o (n753) );
  assign n754 = n473 | n753 ;
  assign n755 = n749 & ~n754 ;
  assign y0 = n339 ;
  assign y1 = n392 ;
  assign y2 = n465 ;
  assign y3 = n487 ;
  assign y4 = n514 ;
  assign y5 = n535 ;
  assign y6 = n557 ;
  assign y7 = n571 ;
  assign y8 = ~n613 ;
  assign y9 = ~n672 ;
  assign y10 = ~n710 ;
  assign y11 = ~n745 ;
  assign y12 = ~n750 ;
  assign y13 = n755 ;
endmodule
