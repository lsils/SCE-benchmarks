module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G4 , G5 , G6 , G7 , G8 , G9 , G1884 , G1885 , G1886 , G1887 , G1888 , G1889 , G1890 , G1891 , G1892 , G1893 , G1894 , G1895 , G1896 , G1897 , G1898 , G1899 , G1900 , G1901 , G1902 , G1903 , G1904 , G1905 , G1906 , G1907 , G1908 );
  input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G4 , G5 , G6 , G7 , G8 , G9 ;
  output G1884 , G1885 , G1886 , G1887 , G1888 , G1889 , G1890 , G1891 , G1892 , G1893 , G1894 , G1895 , G1896 , G1897 , G1898 , G1899 , G1900 , G1901 , G1902 , G1903 , G1904 , G1905 , G1906 , G1907 , G1908 ;
  wire n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 ;
  assign n34 = G24 | G31 ;
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n38( .i (n37), .o (n38) );
  assign n39 = G18 & n38 ;
  buffer buf_n40( .i (n39), .o (n40) );
  assign n45 = G6 | G7 ;
  assign n46 = G6 & G7 ;
  assign n47 = n45 & ~n46 ;
  buffer buf_n48( .i (n47), .o (n48) );
  assign n49 = G5 & n48 ;
  assign n50 = G5 | n48 ;
  assign n51 = ~n49 & n50 ;
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  assign n55 = G4 | G8 ;
  assign n56 = G4 & G8 ;
  assign n57 = n55 & ~n56 ;
  buffer buf_n58( .i (n57), .o (n58) );
  assign n59 = G2 | G3 ;
  assign n60 = G2 & G3 ;
  assign n61 = n59 & ~n60 ;
  buffer buf_n62( .i (n61), .o (n62) );
  assign n63 = G1 & n62 ;
  assign n64 = G1 | n62 ;
  assign n65 = ~n63 & n64 ;
  buffer buf_n66( .i (n65), .o (n66) );
  assign n69 = ~n58 & n66 ;
  assign n70 = n58 & ~n66 ;
  assign n71 = n69 | n70 ;
  buffer buf_n72( .i (n71), .o (n72) );
  assign n73 = n54 | n72 ;
  assign n74 = n54 & n72 ;
  assign n75 = n73 & ~n74 ;
  buffer buf_n76( .i (n75), .o (n76) );
  assign n93 = G21 & ~G33 ;
  buffer buf_n94( .i (n93), .o (n94) );
  assign n95 = ~G9 & n94 ;
  assign n96 = G9 & ~n94 ;
  assign n97 = n95 | n96 ;
  buffer buf_n98( .i (n97), .o (n98) );
  assign n99 = G10 & ~G15 ;
  assign n100 = ~G10 & G15 ;
  assign n101 = n99 | n100 ;
  buffer buf_n102( .i (n101), .o (n102) );
  assign n103 = ~G16 & n102 ;
  assign n104 = G16 & ~n102 ;
  assign n105 = n103 | n104 ;
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  assign n109 = ~n98 & n108 ;
  assign n110 = n98 & ~n108 ;
  assign n111 = n109 | n110 ;
  buffer buf_n112( .i (n111), .o (n112) );
  assign n113 = n76 & ~n112 ;
  assign n114 = ~n76 & n112 ;
  assign n115 = n113 | n114 ;
  buffer buf_n116( .i (n115), .o (n116) );
  assign n133 = G31 | n116 ;
  buffer buf_n134( .i (n133), .o (n134) );
  assign n148 = G17 & n35 ;
  buffer buf_n149( .i (n148), .o (n149) );
  assign n161 = n134 & ~n149 ;
  assign n162 = ~n134 & n149 ;
  assign n163 = n161 | n162 ;
  buffer buf_n164( .i (n163), .o (n164) );
  assign n171 = n40 & ~n164 ;
  buffer buf_n172( .i (n171), .o (n172) );
  assign n173 = ~G11 & G13 ;
  assign n174 = G11 & ~G13 ;
  assign n175 = n173 | n174 ;
  buffer buf_n176( .i (n175), .o (n176) );
  assign n177 = G12 & ~n176 ;
  assign n178 = ~G12 & n176 ;
  assign n179 = n177 | n178 ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = ~n106 & n180 ;
  assign n182 = n106 & ~n180 ;
  assign n183 = n181 | n182 ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n202 = G24 | G33 ;
  buffer buf_n203( .i (n202), .o (n203) );
  assign n204 = G17 & ~n203 ;
  buffer buf_n205( .i (n204), .o (n205) );
  assign n206 = ~G1 & n205 ;
  assign n207 = G1 & ~n205 ;
  assign n208 = n206 | n207 ;
  buffer buf_n209( .i (n208), .o (n209) );
  assign n210 = n52 | n209 ;
  assign n211 = n52 & n209 ;
  assign n212 = n210 & ~n211 ;
  buffer buf_n213( .i (n212), .o (n213) );
  assign n214 = n184 | n213 ;
  assign n215 = n184 & n213 ;
  assign n216 = n214 & ~n215 ;
  buffer buf_n217( .i (n216), .o (n217) );
  assign n238 = G31 | n217 ;
  buffer buf_n239( .i (n238), .o (n239) );
  assign n240 = G26 | n239 ;
  assign n241 = G26 & n239 ;
  assign n242 = n240 & ~n241 ;
  assign n243 = ~G14 & G9 ;
  assign n244 = G14 & ~G9 ;
  assign n245 = n243 | n244 ;
  buffer buf_n246( .i (n245), .o (n246) );
  assign n270 = ~G16 & n246 ;
  assign n271 = G16 & ~n246 ;
  assign n272 = n270 | n271 ;
  buffer buf_n273( .i (n272), .o (n273) );
  assign n274 = G23 | G33 ;
  buffer buf_n275( .i (n274), .o (n275) );
  assign n279 = G20 & ~n275 ;
  buffer buf_n280( .i (n279), .o (n280) );
  assign n281 = ~G13 & n280 ;
  assign n282 = G13 & ~n280 ;
  assign n283 = n281 | n282 ;
  buffer buf_n284( .i (n283), .o (n284) );
  assign n285 = ~n273 & n284 ;
  assign n286 = n273 & ~n284 ;
  assign n287 = n285 | n286 ;
  buffer buf_n288( .i (n287), .o (n288) );
  assign n289 = G4 & ~G7 ;
  assign n290 = ~G4 & G7 ;
  assign n291 = n289 | n290 ;
  buffer buf_n292( .i (n291), .o (n292) );
  assign n293 = G10 & ~n292 ;
  assign n294 = ~G10 & n292 ;
  assign n295 = n293 | n294 ;
  buffer buf_n296( .i (n295), .o (n296) );
  assign n297 = n288 & n296 ;
  assign n298 = n288 | n296 ;
  assign n299 = ~n297 & n298 ;
  buffer buf_n300( .i (n299), .o (n300) );
  assign n321 = G31 | n300 ;
  buffer buf_n322( .i (n321), .o (n322) );
  assign n323 = G23 | G31 ;
  buffer buf_n324( .i (n323), .o (n324) );
  assign n329 = G19 & n324 ;
  buffer buf_n330( .i (n329), .o (n330) );
  assign n347 = n322 & n330 ;
  assign n348 = n322 | n330 ;
  assign n349 = ~n347 & n348 ;
  assign n350 = n242 & n349 ;
  assign n351 = G18 & ~n203 ;
  buffer buf_n352( .i (n351), .o (n352) );
  assign n353 = G11 | G15 ;
  assign n354 = G11 & G15 ;
  assign n355 = n353 & ~n354 ;
  buffer buf_n356( .i (n355), .o (n356) );
  assign n357 = n352 | n356 ;
  assign n358 = n352 & n356 ;
  assign n359 = n357 & ~n358 ;
  buffer buf_n360( .i (n359), .o (n360) );
  assign n361 = n273 & n360 ;
  assign n362 = n273 | n360 ;
  assign n363 = ~n361 & n362 ;
  buffer buf_n364( .i (n363), .o (n364) );
  assign n365 = G5 & ~G8 ;
  assign n366 = ~G5 & G8 ;
  assign n367 = n365 | n366 ;
  buffer buf_n368( .i (n367), .o (n368) );
  assign n369 = G2 & ~n368 ;
  assign n370 = ~G2 & n368 ;
  assign n371 = n369 | n370 ;
  buffer buf_n372( .i (n371), .o (n372) );
  assign n373 = ~n364 & n372 ;
  assign n374 = n364 & ~n372 ;
  assign n375 = n373 | n374 ;
  buffer buf_n376( .i (n375), .o (n376) );
  assign n397 = ~G31 & n376 ;
  buffer buf_n398( .i (n397), .o (n398) );
  assign n399 = G27 & n398 ;
  assign n400 = G27 | n398 ;
  assign n401 = ~n399 & n400 ;
  assign n402 = G3 | G6 ;
  assign n403 = G3 & G6 ;
  assign n404 = n402 & ~n403 ;
  buffer buf_n405( .i (n404), .o (n405) );
  assign n406 = G8 & n405 ;
  assign n407 = G8 | n405 ;
  assign n408 = ~n406 & n407 ;
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n276( .i (n275), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  assign n410 = G19 & ~n278 ;
  buffer buf_n411( .i (n410), .o (n411) );
  assign n412 = G12 & n102 ;
  assign n413 = G12 | n102 ;
  assign n414 = ~n412 & n413 ;
  buffer buf_n415( .i (n414), .o (n415) );
  assign n416 = n411 & ~n415 ;
  assign n417 = ~n411 & n415 ;
  assign n418 = n416 | n417 ;
  buffer buf_n419( .i (n418), .o (n419) );
  assign n420 = n409 | n419 ;
  assign n421 = n409 & n419 ;
  assign n422 = n420 & ~n421 ;
  buffer buf_n423( .i (n422), .o (n423) );
  assign n444 = ~G31 & n423 ;
  buffer buf_n445( .i (n444), .o (n445) );
  assign n446 = G28 & n445 ;
  assign n447 = G28 | n445 ;
  assign n448 = ~n446 & n447 ;
  assign n449 = n401 | n448 ;
  assign n450 = n350 & ~n449 ;
  buffer buf_n451( .i (n450), .o (n451) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  buffer buf_n327( .i (n326), .o (n327) );
  buffer buf_n328( .i (n327), .o (n328) );
  assign n459 = G20 & n328 ;
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  assign n466 = G22 & ~G33 ;
  buffer buf_n467( .i (n466), .o (n467) );
  assign n468 = ~G14 & G4 ;
  assign n469 = G14 & ~G4 ;
  assign n470 = n468 | n469 ;
  buffer buf_n471( .i (n470), .o (n471) );
  assign n472 = n467 & ~n471 ;
  assign n473 = ~n467 & n471 ;
  assign n474 = n472 | n473 ;
  buffer buf_n475( .i (n474), .o (n475) );
  assign n476 = n68 | n475 ;
  assign n477 = n68 & n475 ;
  assign n478 = n476 & ~n477 ;
  buffer buf_n479( .i (n478), .o (n479) );
  assign n480 = n185 | n479 ;
  assign n481 = n185 & n479 ;
  assign n482 = n480 & ~n481 ;
  buffer buf_n483( .i (n482), .o (n483) );
  assign n501 = ~G31 & n483 ;
  buffer buf_n502( .i (n501), .o (n502) );
  assign n517 = G25 | n502 ;
  assign n518 = G25 & n502 ;
  assign n519 = n517 & ~n518 ;
  buffer buf_n520( .i (n519), .o (n520) );
  assign n527 = n460 & n520 ;
  assign n528 = n451 & ~n527 ;
  buffer buf_n529( .i (n528), .o (n529) );
  assign n530 = ~n172 & n529 ;
  buffer buf_n531( .i (n530), .o (n531) );
  assign n532 = G29 | G33 ;
  buffer buf_n533( .i (n532), .o (n533) );
  assign n541 = ~G23 & G24 ;
  buffer buf_n542( .i (n541), .o (n542) );
  assign n544 = G31 | n542 ;
  buffer buf_n545( .i (n544), .o (n545) );
  assign n546 = n533 | n545 ;
  buffer buf_n543( .i (n542), .o (n543) );
  assign n547 = G32 | G33 ;
  buffer buf_n548( .i (n547), .o (n548) );
  assign n563 = n543 | n548 ;
  buffer buf_n564( .i (n563), .o (n564) );
  assign n565 = n546 & n564 ;
  buffer buf_n566( .i (n565), .o (n566) );
  assign n567 = n531 & ~n566 ;
  buffer buf_n568( .i (n567), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  buffer buf_n573( .i (n572), .o (n573) );
  buffer buf_n574( .i (n573), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  assign n576 = G1 | n575 ;
  assign n577 = G1 & n575 ;
  assign n578 = ~n576 | n577 ;
  assign n579 = G2 | n575 ;
  assign n580 = G2 & n575 ;
  assign n581 = ~n579 | n580 ;
  buffer buf_n582( .i (n574), .o (n582) );
  assign n583 = G3 | n582 ;
  assign n584 = G3 & n582 ;
  assign n585 = ~n583 | n584 ;
  assign n586 = G4 | n582 ;
  assign n587 = G4 & n582 ;
  assign n588 = ~n586 | n587 ;
  assign n589 = G30 | G33 ;
  buffer buf_n590( .i (n589), .o (n590) );
  assign n597 = n545 | n590 ;
  assign n598 = n564 & n597 ;
  buffer buf_n599( .i (n598), .o (n599) );
  assign n600 = n531 & ~n599 ;
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  buffer buf_n603( .i (n602), .o (n603) );
  buffer buf_n604( .i (n603), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  buffer buf_n607( .i (n606), .o (n607) );
  buffer buf_n608( .i (n607), .o (n608) );
  assign n609 = G10 | n608 ;
  assign n610 = G10 & n608 ;
  assign n611 = ~n609 | n610 ;
  assign n612 = G15 | n608 ;
  assign n613 = G15 & n608 ;
  assign n614 = ~n612 | n613 ;
  buffer buf_n615( .i (n607), .o (n615) );
  assign n616 = G16 | n615 ;
  assign n617 = G16 & n615 ;
  assign n618 = ~n616 | n617 ;
  buffer buf_n452( .i (n451), .o (n452) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n521( .i (n520), .o (n521) );
  assign n619 = n461 & ~n521 ;
  assign n620 = n452 & n619 ;
  assign n621 = ~n172 & n620 ;
  buffer buf_n622( .i (n621), .o (n622) );
  assign n623 = ~n566 & n622 ;
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  buffer buf_n626( .i (n625), .o (n626) );
  buffer buf_n627( .i (n626), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n631( .i (n630), .o (n631) );
  assign n632 = G5 | n631 ;
  assign n633 = G5 & n631 ;
  assign n634 = ~n632 | n633 ;
  assign n635 = G6 | n631 ;
  assign n636 = G6 & n631 ;
  assign n637 = ~n635 | n636 ;
  buffer buf_n638( .i (n630), .o (n638) );
  assign n639 = G7 | n638 ;
  assign n640 = G7 & n638 ;
  assign n641 = ~n639 | n640 ;
  assign n642 = G8 | n638 ;
  assign n643 = G8 & n638 ;
  assign n644 = ~n642 | n643 ;
  assign n645 = ~n599 & n622 ;
  buffer buf_n646( .i (n645), .o (n646) );
  assign n647 = G9 & ~n646 ;
  assign n648 = ~G9 & n646 ;
  assign n649 = n647 | n648 ;
  buffer buf_n650( .i (n649), .o (n650) );
  buffer buf_n651( .i (n650), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  buffer buf_n653( .i (n652), .o (n653) );
  buffer buf_n654( .i (n653), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  inverter inv_n656( .i (n655), .o (n656) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  assign n657 = n42 & n529 ;
  assign n658 = n167 & n657 ;
  assign n659 = ~n599 & n658 ;
  buffer buf_n660( .i (n659), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  assign n668 = G11 | n667 ;
  assign n669 = G11 & n667 ;
  assign n670 = ~n668 | n669 ;
  assign n671 = G12 | n667 ;
  assign n672 = G12 & n667 ;
  assign n673 = ~n671 | n672 ;
  buffer buf_n674( .i (n666), .o (n674) );
  assign n675 = G13 | n674 ;
  assign n676 = G13 & n674 ;
  assign n677 = ~n675 | n676 ;
  assign n678 = G14 | n674 ;
  assign n679 = G14 & n674 ;
  assign n680 = ~n678 | n679 ;
  assign n681 = n568 | n601 ;
  buffer buf_n682( .i (n681), .o (n682) );
  assign n688 = G32 & n682 ;
  buffer buf_n453( .i (n452), .o (n453) );
  buffer buf_n454( .i (n453), .o (n454) );
  buffer buf_n455( .i (n454), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  buffer buf_n525( .i (n524), .o (n525) );
  buffer buf_n526( .i (n525), .o (n526) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  assign n689 = n44 | n465 ;
  assign n690 = n526 | n689 ;
  assign n691 = n170 & ~n690 ;
  assign n692 = n458 & n691 ;
  assign n693 = G33 | n692 ;
  assign n694 = n688 | n693 ;
  buffer buf_n695( .i (n694), .o (n695) );
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n697( .i (n696), .o (n697) );
  buffer buf_n698( .i (n697), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n117( .i (n116), .o (n117) );
  buffer buf_n118( .i (n117), .o (n118) );
  buffer buf_n119( .i (n118), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n130( .i (n129), .o (n130) );
  buffer buf_n131( .i (n130), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n153( .i (n152), .o (n153) );
  buffer buf_n154( .i (n153), .o (n154) );
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  assign n700 = n160 & n682 ;
  buffer buf_n701( .i (n700), .o (n701) );
  assign n702 = ~G31 & n701 ;
  assign n703 = n132 & ~n702 ;
  buffer buf_n549( .i (n548), .o (n549) );
  buffer buf_n550( .i (n549), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n553( .i (n552), .o (n553) );
  buffer buf_n554( .i (n553), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  buffer buf_n138( .i (n137), .o (n138) );
  buffer buf_n139( .i (n138), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  buffer buf_n146( .i (n145), .o (n146) );
  buffer buf_n147( .i (n146), .o (n147) );
  assign n704 = ~n147 & n701 ;
  assign n705 = n559 & ~n704 ;
  assign n706 = ~n703 & n705 ;
  buffer buf_n707( .i (n706), .o (n707) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  assign n709 = G25 & n682 ;
  buffer buf_n710( .i (n709), .o (n710) );
  assign n711 = ~G31 & n710 ;
  assign n712 = n500 | n711 ;
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n510( .i (n509), .o (n510) );
  buffer buf_n511( .i (n510), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  buffer buf_n513( .i (n512), .o (n513) );
  buffer buf_n514( .i (n513), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  assign n713 = n516 & n710 ;
  assign n714 = n559 & ~n713 ;
  assign n715 = n712 & n714 ;
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  buffer buf_n393( .i (n392), .o (n393) );
  buffer buf_n394( .i (n393), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n684( .i (n683), .o (n684) );
  buffer buf_n685( .i (n684), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  assign n718 = G27 & ~G31 ;
  assign n719 = n686 & n718 ;
  assign n720 = n396 & ~n719 ;
  assign n721 = n562 & ~n720 ;
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  assign n722 = G28 & ~G31 ;
  assign n723 = n686 & n722 ;
  assign n724 = n443 & ~n723 ;
  assign n725 = n562 & ~n724 ;
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n335( .i (n334), .o (n335) );
  buffer buf_n336( .i (n335), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  buffer buf_n342( .i (n341), .o (n342) );
  buffer buf_n343( .i (n342), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  assign n726 = ~G31 & n346 ;
  assign n727 = n686 & n726 ;
  assign n728 = n320 | n727 ;
  assign n729 = n562 & n728 ;
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n85( .i (n84), .o (n85) );
  buffer buf_n86( .i (n85), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n91( .i (n90), .o (n91) );
  buffer buf_n92( .i (n91), .o (n92) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  buffer buf_n536( .i (n535), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  assign n730 = n92 & n540 ;
  buffer buf_n731( .i (n730), .o (n731) );
  assign n732 = G21 & G29 ;
  buffer buf_n733( .i (n732), .o (n733) );
  assign n734 = n568 | n733 ;
  assign n735 = n568 & n733 ;
  assign n736 = n734 & ~n735 ;
  assign n737 = G33 | n736 ;
  buffer buf_n738( .i (n737), .o (n738) );
  assign n739 = n731 & n738 ;
  assign n740 = n731 | n738 ;
  assign n741 = ~n739 & n740 ;
  buffer buf_n742( .i (n741), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  inverter inv_n744( .i (n743), .o (n744) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  buffer buf_n192( .i (n191), .o (n192) );
  buffer buf_n193( .i (n192), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n249( .i (n248), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  buffer buf_n252( .i (n251), .o (n252) );
  buffer buf_n253( .i (n252), .o (n253) );
  buffer buf_n254( .i (n253), .o (n254) );
  buffer buf_n255( .i (n254), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  assign n745 = n201 | n269 ;
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  buffer buf_n593( .i (n592), .o (n593) );
  buffer buf_n594( .i (n593), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  assign n746 = n200 & n268 ;
  assign n747 = n596 & ~n746 ;
  assign n748 = n745 & n747 ;
  buffer buf_n749( .i (n748), .o (n749) );
  assign n750 = G22 & G30 ;
  buffer buf_n751( .i (n750), .o (n751) );
  assign n752 = n601 | n751 ;
  assign n753 = n601 & n751 ;
  assign n754 = n752 & ~n753 ;
  assign n755 = G33 | n754 ;
  buffer buf_n756( .i (n755), .o (n756) );
  assign n757 = n749 & ~n756 ;
  assign n758 = ~n749 & n756 ;
  assign n759 = n757 | n758 ;
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  inverter inv_n762( .i (n761), .o (n762) );
  buffer buf_n687( .i (n686), .o (n687) );
  assign n763 = G26 & n687 ;
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  assign n764 = ~n237 & n561 ;
  assign n765 = ~n763 & n764 ;
  assign G1884 = n578 ;
  assign G1885 = n581 ;
  assign G1886 = n585 ;
  assign G1887 = n588 ;
  assign G1888 = n611 ;
  assign G1889 = n614 ;
  assign G1890 = n618 ;
  assign G1891 = n634 ;
  assign G1892 = n637 ;
  assign G1893 = n641 ;
  assign G1894 = n644 ;
  assign G1895 = n656 ;
  assign G1896 = n670 ;
  assign G1897 = n673 ;
  assign G1898 = n677 ;
  assign G1899 = n680 ;
  assign G1900 = n699 ;
  assign G1901 = n708 ;
  assign G1902 = n717 ;
  assign G1903 = n721 ;
  assign G1904 = n725 ;
  assign G1905 = n729 ;
  assign G1906 = n744 ;
  assign G1907 = n762 ;
  assign G1908 = n765 ;
endmodule
