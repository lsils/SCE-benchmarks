module apc128bits(in_18_,in_1_,in_7_,in_109_,in_13_,in_106_,in_54_,in_118_,in_101_,in_3_,in_0_,in_113_,in_56_,in_30_,in_89_,in_35_,in_70_,in_38_,in_100_,in_105_,in_28_,in_10_,in_9_,in_78_,in_29_,in_60_,in_94_,in_108_,in_117_,in_103_,in_67_,in_44_,in_57_,in_76_,in_47_,in_20_,in_84_,in_17_,in_72_,in_116_,in_16_,in_120_,in_104_,in_64_,in_125_,in_58_,in_42_,in_40_,in_81_,in_115_,in_88_,in_24_,in_33_,in_123_,in_61_,in_79_,in_31_,in_36_,in_82_,in_111_,in_68_,in_2_,in_87_,in_74_,in_114_,in_53_,in_83_,in_86_,in_65_,in_102_,in_6_,in_75_,in_4_,in_93_,in_45_,in_90_,in_80_,in_73_,in_46_,in_25_,in_107_,in_37_,in_85_,in_49_,in_39_,in_63_,in_12_,in_112_,in_32_,in_119_,in_77_,in_34_,in_41_,in_122_,in_124_,in_48_,in_92_,in_15_,in_55_,in_50_,in_5_,in_127_,in_96_,in_22_,in_43_,in_52_,in_51_,in_21_,in_95_,in_59_,in_69_,in_121_,in_97_,in_11_,in_98_,in_126_,in_14_,in_91_,in_26_,in_99_,in_27_,in_71_,in_8_,in_23_,in_110_,in_62_,in_66_,in_19_,out_3_,out_2_,out_5_,out_1_,out_0_,out_7_,out_4_,out_6_);
    wire jinkela_wire_0;
    wire jinkela_wire_1;
    wire jinkela_wire_2;
    wire jinkela_wire_3;
    wire jinkela_wire_4;
    wire jinkela_wire_5;
    wire jinkela_wire_6;
    wire jinkela_wire_7;
    wire jinkela_wire_8;
    wire jinkela_wire_9;
    wire jinkela_wire_10;
    wire jinkela_wire_11;
    wire jinkela_wire_12;
    wire jinkela_wire_13;
    wire jinkela_wire_14;
    wire jinkela_wire_15;
    wire jinkela_wire_16;
    wire jinkela_wire_17;
    wire jinkela_wire_18;
    wire jinkela_wire_19;
    wire jinkela_wire_20;
    wire jinkela_wire_21;
    wire jinkela_wire_22;
    wire jinkela_wire_23;
    wire jinkela_wire_24;
    wire jinkela_wire_25;
    wire jinkela_wire_26;
    wire jinkela_wire_27;
    wire jinkela_wire_28;
    wire jinkela_wire_29;
    wire jinkela_wire_30;
    wire jinkela_wire_31;
    wire jinkela_wire_32;
    wire jinkela_wire_33;
    wire jinkela_wire_34;
    wire jinkela_wire_35;
    wire jinkela_wire_36;
    wire jinkela_wire_37;
    wire jinkela_wire_38;
    wire jinkela_wire_39;
    wire jinkela_wire_40;
    wire jinkela_wire_41;
    wire jinkela_wire_42;
    wire jinkela_wire_43;
    wire jinkela_wire_44;
    wire jinkela_wire_45;
    wire jinkela_wire_46;
    wire jinkela_wire_47;
    wire jinkela_wire_48;
    wire jinkela_wire_49;
    wire jinkela_wire_50;
    wire jinkela_wire_51;
    wire jinkela_wire_52;
    wire jinkela_wire_53;
    wire jinkela_wire_54;
    wire jinkela_wire_55;
    wire jinkela_wire_56;
    wire jinkela_wire_57;
    wire jinkela_wire_58;
    wire jinkela_wire_59;
    wire jinkela_wire_60;
    wire jinkela_wire_61;
    wire jinkela_wire_62;
    wire jinkela_wire_63;
    wire jinkela_wire_64;
    wire jinkela_wire_65;
    wire jinkela_wire_66;
    wire jinkela_wire_67;
    wire jinkela_wire_68;
    wire jinkela_wire_69;
    wire jinkela_wire_70;
    wire jinkela_wire_71;
    wire jinkela_wire_72;
    wire jinkela_wire_73;
    wire jinkela_wire_74;
    wire jinkela_wire_75;
    wire jinkela_wire_76;
    wire jinkela_wire_77;
    wire jinkela_wire_78;
    wire jinkela_wire_79;
    wire jinkela_wire_80;
    wire jinkela_wire_81;
    wire jinkela_wire_82;
    wire jinkela_wire_83;
    wire jinkela_wire_84;
    wire jinkela_wire_85;
    wire jinkela_wire_86;
    wire jinkela_wire_87;
    wire jinkela_wire_88;
    wire jinkela_wire_89;
    wire jinkela_wire_90;
    wire jinkela_wire_91;
    wire jinkela_wire_92;
    wire jinkela_wire_93;
    wire jinkela_wire_94;
    wire jinkela_wire_95;
    wire jinkela_wire_96;
    wire jinkela_wire_97;
    wire jinkela_wire_98;
    wire jinkela_wire_99;
    wire jinkela_wire_100;
    wire jinkela_wire_101;
    wire jinkela_wire_102;
    wire jinkela_wire_103;
    wire jinkela_wire_104;
    wire jinkela_wire_105;
    wire jinkela_wire_106;
    wire jinkela_wire_107;
    wire jinkela_wire_108;
    wire jinkela_wire_109;
    wire jinkela_wire_110;
    wire jinkela_wire_111;
    wire jinkela_wire_112;
    wire jinkela_wire_113;
    wire jinkela_wire_114;
    wire jinkela_wire_115;
    wire jinkela_wire_116;
    wire jinkela_wire_117;
    wire jinkela_wire_118;
    wire jinkela_wire_119;
    wire jinkela_wire_120;
    wire jinkela_wire_121;
    wire jinkela_wire_122;
    wire jinkela_wire_123;
    wire jinkela_wire_124;
    wire jinkela_wire_125;
    wire jinkela_wire_126;
    wire jinkela_wire_127;
    wire jinkela_wire_128;
    wire jinkela_wire_129;
    wire jinkela_wire_130;
    wire jinkela_wire_131;
    wire jinkela_wire_132;
    wire jinkela_wire_133;
    wire jinkela_wire_134;
    wire jinkela_wire_135;
    wire jinkela_wire_136;
    wire jinkela_wire_137;
    wire jinkela_wire_138;
    wire jinkela_wire_139;
    wire jinkela_wire_140;
    wire jinkela_wire_141;
    wire jinkela_wire_142;
    wire jinkela_wire_143;
    wire jinkela_wire_144;
    wire jinkela_wire_145;
    wire jinkela_wire_146;
    wire jinkela_wire_147;
    wire jinkela_wire_148;
    wire jinkela_wire_149;
    wire jinkela_wire_150;
    wire jinkela_wire_151;
    wire jinkela_wire_152;
    wire jinkela_wire_153;
    wire jinkela_wire_154;
    wire jinkela_wire_155;
    wire jinkela_wire_156;
    wire jinkela_wire_157;
    wire jinkela_wire_158;
    wire jinkela_wire_159;
    wire jinkela_wire_160;
    wire jinkela_wire_161;
    wire jinkela_wire_162;
    wire jinkela_wire_163;
    wire jinkela_wire_164;
    wire jinkela_wire_165;
    wire jinkela_wire_166;
    wire jinkela_wire_167;
    wire jinkela_wire_168;
    wire jinkela_wire_169;
    wire jinkela_wire_170;
    wire jinkela_wire_171;
    wire jinkela_wire_172;
    wire jinkela_wire_173;
    wire jinkela_wire_174;
    wire jinkela_wire_175;
    wire jinkela_wire_176;
    wire jinkela_wire_177;
    wire jinkela_wire_178;
    wire jinkela_wire_179;
    wire jinkela_wire_180;
    wire jinkela_wire_181;
    wire jinkela_wire_182;
    wire jinkela_wire_183;
    wire jinkela_wire_184;
    wire jinkela_wire_185;
    wire jinkela_wire_186;
    wire jinkela_wire_187;
    wire jinkela_wire_188;
    wire jinkela_wire_189;
    wire jinkela_wire_190;
    wire jinkela_wire_191;
    wire jinkela_wire_192;
    wire jinkela_wire_193;
    wire jinkela_wire_194;
    wire jinkela_wire_195;
    wire jinkela_wire_196;
    wire jinkela_wire_197;
    wire jinkela_wire_198;
    wire jinkela_wire_199;
    wire jinkela_wire_200;
    wire jinkela_wire_201;
    wire jinkela_wire_202;
    wire jinkela_wire_203;
    wire jinkela_wire_204;
    wire jinkela_wire_205;
    wire jinkela_wire_206;
    wire jinkela_wire_207;
    wire jinkela_wire_208;
    wire jinkela_wire_209;
    wire jinkela_wire_210;
    wire jinkela_wire_211;
    wire jinkela_wire_212;
    wire jinkela_wire_213;
    wire jinkela_wire_214;
    wire jinkela_wire_215;
    wire jinkela_wire_216;
    wire jinkela_wire_217;
    wire jinkela_wire_218;
    wire jinkela_wire_219;
    wire jinkela_wire_220;
    wire jinkela_wire_221;
    wire jinkela_wire_222;
    wire jinkela_wire_223;
    wire jinkela_wire_224;
    wire jinkela_wire_225;
    wire jinkela_wire_226;
    wire jinkela_wire_227;
    wire jinkela_wire_228;
    wire jinkela_wire_229;
    wire jinkela_wire_230;
    wire jinkela_wire_231;
    wire jinkela_wire_232;
    wire jinkela_wire_233;
    wire jinkela_wire_234;
    wire jinkela_wire_235;
    wire jinkela_wire_236;
    wire jinkela_wire_237;
    wire jinkela_wire_238;
    wire jinkela_wire_239;
    wire jinkela_wire_240;
    wire jinkela_wire_241;
    wire jinkela_wire_242;
    wire jinkela_wire_243;
    wire jinkela_wire_244;
    wire jinkela_wire_245;
    wire jinkela_wire_246;
    wire jinkela_wire_247;
    wire jinkela_wire_248;
    wire jinkela_wire_249;
    wire jinkela_wire_250;
    wire jinkela_wire_251;
    wire jinkela_wire_252;
    wire jinkela_wire_253;
    wire jinkela_wire_254;
    wire jinkela_wire_255;
    wire jinkela_wire_256;
    wire jinkela_wire_257;
    wire jinkela_wire_258;
    wire jinkela_wire_259;
    wire jinkela_wire_260;
    wire jinkela_wire_261;
    wire jinkela_wire_262;
    wire jinkela_wire_263;
    wire jinkela_wire_264;
    wire jinkela_wire_265;
    wire jinkela_wire_266;
    wire jinkela_wire_267;
    wire jinkela_wire_268;
    wire jinkela_wire_269;
    wire jinkela_wire_270;
    wire jinkela_wire_271;
    wire jinkela_wire_272;
    wire jinkela_wire_273;
    wire jinkela_wire_274;
    wire jinkela_wire_275;
    wire jinkela_wire_276;
    wire jinkela_wire_277;
    wire jinkela_wire_278;
    wire jinkela_wire_279;
    wire jinkela_wire_280;
    wire jinkela_wire_281;
    wire jinkela_wire_282;
    wire jinkela_wire_283;
    wire jinkela_wire_284;
    wire jinkela_wire_285;
    wire jinkela_wire_286;
    wire jinkela_wire_287;
    wire jinkela_wire_288;
    wire jinkela_wire_289;
    wire jinkela_wire_290;
    wire jinkela_wire_291;
    wire jinkela_wire_292;
    wire jinkela_wire_293;
    wire jinkela_wire_294;
    wire jinkela_wire_295;
    wire jinkela_wire_296;
    wire jinkela_wire_297;
    wire jinkela_wire_298;
    wire jinkela_wire_299;
    wire jinkela_wire_300;
    wire jinkela_wire_301;
    wire jinkela_wire_302;
    wire jinkela_wire_303;
    wire jinkela_wire_304;
    wire jinkela_wire_305;
    wire jinkela_wire_306;
    wire jinkela_wire_307;
    wire jinkela_wire_308;
    wire jinkela_wire_309;
    wire jinkela_wire_310;
    wire jinkela_wire_311;
    wire jinkela_wire_312;
    wire jinkela_wire_313;
    wire jinkela_wire_314;
    wire jinkela_wire_315;
    wire jinkela_wire_316;
    wire jinkela_wire_317;
    wire jinkela_wire_318;
    wire jinkela_wire_319;
    wire jinkela_wire_320;
    wire jinkela_wire_321;
    wire jinkela_wire_322;
    wire jinkela_wire_323;
    wire jinkela_wire_324;
    wire jinkela_wire_325;
    wire jinkela_wire_326;
    wire jinkela_wire_327;
    wire jinkela_wire_328;
    wire jinkela_wire_329;
    wire jinkela_wire_330;
    wire jinkela_wire_331;
    wire jinkela_wire_332;
    wire jinkela_wire_333;
    wire jinkela_wire_334;
    wire jinkela_wire_335;
    wire jinkela_wire_336;
    wire jinkela_wire_337;
    wire jinkela_wire_338;
    wire jinkela_wire_339;
    wire jinkela_wire_340;
    wire jinkela_wire_341;
    wire jinkela_wire_342;
    wire jinkela_wire_343;
    wire jinkela_wire_344;
    wire jinkela_wire_345;
    wire jinkela_wire_346;
    wire jinkela_wire_347;
    wire jinkela_wire_348;
    wire jinkela_wire_349;
    wire jinkela_wire_350;
    wire jinkela_wire_351;
    wire jinkela_wire_352;
    wire jinkela_wire_353;
    wire jinkela_wire_354;
    wire jinkela_wire_355;
    wire jinkela_wire_356;
    wire jinkela_wire_357;
    wire jinkela_wire_358;
    wire jinkela_wire_359;
    wire jinkela_wire_360;
    wire jinkela_wire_361;
    wire jinkela_wire_362;
    wire jinkela_wire_363;
    wire jinkela_wire_364;
    wire jinkela_wire_365;
    wire jinkela_wire_366;
    wire jinkela_wire_367;
    wire jinkela_wire_368;
    wire jinkela_wire_369;
    wire jinkela_wire_370;
    wire jinkela_wire_371;
    wire jinkela_wire_372;
    wire jinkela_wire_373;
    wire jinkela_wire_374;
    wire jinkela_wire_375;
    wire jinkela_wire_376;
    wire jinkela_wire_377;
    wire jinkela_wire_378;
    wire jinkela_wire_379;
    wire jinkela_wire_380;
    wire jinkela_wire_381;
    wire jinkela_wire_382;
    wire jinkela_wire_383;
    wire jinkela_wire_384;
    wire jinkela_wire_385;
    wire jinkela_wire_386;
    wire jinkela_wire_387;
    wire jinkela_wire_388;
    wire jinkela_wire_389;
    wire jinkela_wire_390;
    wire jinkela_wire_391;
    wire jinkela_wire_392;
    wire jinkela_wire_393;
    wire jinkela_wire_394;
    wire jinkela_wire_395;
    wire jinkela_wire_396;
    wire jinkela_wire_397;
    wire jinkela_wire_398;
    wire jinkela_wire_399;
    wire jinkela_wire_400;
    wire jinkela_wire_401;
    wire jinkela_wire_402;
    wire jinkela_wire_403;
    wire jinkela_wire_404;
    wire jinkela_wire_405;
    wire jinkela_wire_406;
    wire jinkela_wire_407;
    wire jinkela_wire_408;
    wire jinkela_wire_409;
    wire jinkela_wire_410;
    wire jinkela_wire_411;
    wire jinkela_wire_412;
    wire jinkela_wire_413;
    wire jinkela_wire_414;
    wire jinkela_wire_415;
    wire jinkela_wire_416;
    wire jinkela_wire_417;
    wire jinkela_wire_418;
    wire jinkela_wire_419;
    wire jinkela_wire_420;
    wire jinkela_wire_421;
    wire jinkela_wire_422;
    wire jinkela_wire_423;
    wire jinkela_wire_424;
    wire jinkela_wire_425;
    wire jinkela_wire_426;
    wire jinkela_wire_427;
    wire jinkela_wire_428;
    wire jinkela_wire_429;
    wire jinkela_wire_430;
    wire jinkela_wire_431;
    wire jinkela_wire_432;
    wire jinkela_wire_433;
    wire jinkela_wire_434;
    wire jinkela_wire_435;
    wire jinkela_wire_436;
    wire jinkela_wire_437;
    wire jinkela_wire_438;
    wire jinkela_wire_439;
    wire jinkela_wire_440;
    wire jinkela_wire_441;
    wire jinkela_wire_442;
    wire jinkela_wire_443;
    wire jinkela_wire_444;
    wire jinkela_wire_445;
    wire jinkela_wire_446;
    wire jinkela_wire_447;
    wire jinkela_wire_448;
    wire jinkela_wire_449;
    wire jinkela_wire_450;
    wire jinkela_wire_451;
    wire jinkela_wire_452;
    wire jinkela_wire_453;
    wire jinkela_wire_454;
    wire jinkela_wire_455;
    wire jinkela_wire_456;
    wire jinkela_wire_457;
    wire jinkela_wire_458;
    wire jinkela_wire_459;
    wire jinkela_wire_460;
    wire jinkela_wire_461;
    wire jinkela_wire_462;
    wire jinkela_wire_463;
    wire jinkela_wire_464;
    wire jinkela_wire_465;
    wire jinkela_wire_466;
    wire jinkela_wire_467;
    wire jinkela_wire_468;
    input in_18_;
    input in_1_;
    input in_7_;
    input in_109_;
    input in_13_;
    input in_106_;
    input in_54_;
    input in_118_;
    input in_101_;
    input in_3_;
    input in_0_;
    input in_113_;
    input in_56_;
    input in_30_;
    input in_89_;
    input in_35_;
    input in_70_;
    input in_38_;
    input in_100_;
    input in_105_;
    input in_28_;
    input in_10_;
    input in_9_;
    input in_78_;
    input in_29_;
    input in_60_;
    input in_94_;
    input in_108_;
    input in_117_;
    input in_103_;
    input in_67_;
    input in_44_;
    input in_57_;
    input in_76_;
    input in_47_;
    input in_20_;
    input in_84_;
    input in_17_;
    input in_72_;
    input in_116_;
    input in_16_;
    input in_120_;
    input in_104_;
    input in_64_;
    input in_125_;
    input in_58_;
    input in_42_;
    input in_40_;
    input in_81_;
    input in_115_;
    input in_88_;
    input in_24_;
    input in_33_;
    input in_123_;
    input in_61_;
    input in_79_;
    input in_31_;
    input in_36_;
    input in_82_;
    input in_111_;
    input in_68_;
    input in_2_;
    input in_87_;
    input in_74_;
    input in_114_;
    input in_53_;
    input in_83_;
    input in_86_;
    input in_65_;
    input in_102_;
    input in_6_;
    input in_75_;
    input in_4_;
    input in_93_;
    input in_45_;
    input in_90_;
    input in_80_;
    input in_73_;
    input in_46_;
    input in_25_;
    input in_107_;
    input in_37_;
    input in_85_;
    input in_49_;
    input in_39_;
    input in_63_;
    input in_12_;
    input in_112_;
    input in_32_;
    input in_119_;
    input in_77_;
    input in_34_;
    input in_41_;
    input in_122_;
    input in_124_;
    input in_48_;
    input in_92_;
    input in_15_;
    input in_55_;
    input in_50_;
    input in_5_;
    input in_127_;
    input in_96_;
    input in_22_;
    input in_43_;
    input in_52_;
    input in_51_;
    input in_21_;
    input in_95_;
    input in_59_;
    input in_69_;
    input in_121_;
    input in_97_;
    input in_11_;
    input in_98_;
    input in_126_;
    input in_14_;
    input in_91_;
    input in_26_;
    input in_99_;
    input in_27_;
    input in_71_;
    input in_8_;
    input in_23_;
    input in_110_;
    input in_62_;
    input in_66_;
    input in_19_;
    output out_3_;
    output out_2_;
    output out_5_;
    output out_1_;
    output out_0_;
    output out_7_;
    output out_4_;
    output out_6_;

    and_bi _400_ (
        .a(jinkela_wire_145),
        .b(jinkela_wire_177),
        .c(jinkela_wire_303)
    );

    and_bi _401_ (
        .a(jinkela_wire_447),
        .b(jinkela_wire_303),
        .c(jinkela_wire_215)
    );

    maj_bii _402_ (
        .c(jinkela_wire_126),
        .a(jinkela_wire_145),
        .b(jinkela_wire_233),
        .d(jinkela_wire_263)
    );

    or_ii _403_ (
        .a(jinkela_wire_86),
        .b(jinkela_wire_462),
        .c(jinkela_wire_182)
    );

    and_ii _404_ (
        .a(jinkela_wire_86),
        .b(jinkela_wire_462),
        .c(jinkela_wire_253)
    );

    and_bi _405_ (
        .a(jinkela_wire_182),
        .b(jinkela_wire_253),
        .c(jinkela_wire_385)
    );

    or_bi _406_ (
        .a(jinkela_wire_263),
        .b(jinkela_wire_385),
        .c(jinkela_wire_373)
    );

    and_bi _407_ (
        .a(jinkela_wire_263),
        .b(jinkela_wire_385),
        .c(jinkela_wire_72)
    );

    and_bi _408_ (
        .a(jinkela_wire_373),
        .b(jinkela_wire_72),
        .c(jinkela_wire_141)
    );

    maj_bii _409_ (
        .c(jinkela_wire_462),
        .a(jinkela_wire_263),
        .b(jinkela_wire_86),
        .d(jinkela_wire_321)
    );

    or_ii _410_ (
        .a(jinkela_wire_455),
        .b(jinkela_wire_39),
        .c(jinkela_wire_289)
    );

    and_ii _411_ (
        .a(jinkela_wire_455),
        .b(jinkela_wire_39),
        .c(jinkela_wire_71)
    );

    and_bi _412_ (
        .a(jinkela_wire_289),
        .b(jinkela_wire_71),
        .c(jinkela_wire_167)
    );

    and_ii _524_ (
        .a(jinkela_wire_315),
        .b(jinkela_wire_433),
        .c(jinkela_wire_425)
    );

    or_bi _413_ (
        .a(jinkela_wire_321),
        .b(jinkela_wire_167),
        .c(jinkela_wire_382)
    );

    and_bi _414_ (
        .a(jinkela_wire_321),
        .b(jinkela_wire_167),
        .c(jinkela_wire_32)
    );

    and_bi _415_ (
        .a(jinkela_wire_382),
        .b(jinkela_wire_32),
        .c(jinkela_wire_394)
    );

    maj_bii _416_ (
        .c(jinkela_wire_39),
        .a(jinkela_wire_321),
        .b(jinkela_wire_455),
        .d(jinkela_wire_174)
    );

    or_ii _417_ (
        .a(jinkela_wire_193),
        .b(jinkela_wire_47),
        .c(jinkela_wire_434)
    );

    and_bi _525_ (
        .a(jinkela_wire_411),
        .b(jinkela_wire_425),
        .c(jinkela_wire_277)
    );

    and_ii _418_ (
        .a(jinkela_wire_193),
        .b(jinkela_wire_47),
        .c(jinkela_wire_374)
    );

    and_bi _419_ (
        .a(jinkela_wire_434),
        .b(jinkela_wire_374),
        .c(jinkela_wire_222)
    );

    or_bi _420_ (
        .a(jinkela_wire_174),
        .b(jinkela_wire_222),
        .c(jinkela_wire_235)
    );

    and_bi _421_ (
        .a(jinkela_wire_174),
        .b(jinkela_wire_222),
        .c(jinkela_wire_389)
    );

    and_bi _422_ (
        .a(jinkela_wire_235),
        .b(jinkela_wire_389),
        .c(jinkela_wire_232)
    );

    and_ii _423_ (
        .a(1'b0),
        .b(1'b0),
        .c(jinkela_wire_77)
    );

    maj_bbi _566_ (
        .c(jinkela_wire_260),
        .a(jinkela_wire_375),
        .b(jinkela_wire_250),
        .d(jinkela_wire_135)
    );

    and_bi _424_ (
        .a(jinkela_wire_145),
        .b(jinkela_wire_77),
        .c(jinkela_wire_34)
    );

    maj_bbi _425_ (
        .c(jinkela_wire_174),
        .a(jinkela_wire_193),
        .b(jinkela_wire_47),
        .d(jinkela_wire_310)
    );

    or_bb _426_ (
        .a(in_81_),
        .b(in_80_),
        .c(jinkela_wire_379)
    );

    and_bb _427_ (
        .a(in_83_),
        .b(in_82_),
        .c(jinkela_wire_249)
    );

    or_bb _428_ (
        .a(in_85_),
        .b(in_84_),
        .c(jinkela_wire_224)
    );

    maj_bbb _567_ (
        .c(jinkela_wire_28),
        .a(jinkela_wire_400),
        .b(jinkela_wire_44),
        .d(jinkela_wire_198)
    );

    and_bb _429_ (
        .a(in_87_),
        .b(in_86_),
        .c(jinkela_wire_305)
    );

    or_bb _430_ (
        .a(in_89_),
        .b(in_88_),
        .c(jinkela_wire_270)
    );

    and_bb _431_ (
        .a(in_91_),
        .b(in_90_),
        .c(jinkela_wire_275)
    );

    or_bb _432_ (
        .a(in_93_),
        .b(in_92_),
        .c(jinkela_wire_146)
    );

    and_bb _433_ (
        .a(in_95_),
        .b(in_94_),
        .c(jinkela_wire_84)
    );

    maj_bbb _434_ (
        .c(jinkela_wire_379),
        .a(jinkela_wire_224),
        .b(jinkela_wire_249),
        .d(jinkela_wire_138)
    );

    and_bb _608_ (
        .a(jinkela_wire_364),
        .b(jinkela_wire_156),
        .c(jinkela_wire_318)
    );

    maj_bbi _435_ (
        .c(jinkela_wire_224),
        .a(jinkela_wire_249),
        .b(jinkela_wire_379),
        .d(jinkela_wire_380)
    );

    maj_bbi _436_ (
        .c(jinkela_wire_138),
        .a(jinkela_wire_380),
        .b(jinkela_wire_224),
        .d(jinkela_wire_73)
    );

    maj_bbb _437_ (
        .c(jinkela_wire_138),
        .a(jinkela_wire_457),
        .b(jinkela_wire_360),
        .d(jinkela_wire_259)
    );

    maj_bbi _438_ (
        .c(jinkela_wire_457),
        .a(jinkela_wire_360),
        .b(jinkela_wire_138),
        .d(jinkela_wire_13)
    );

    maj_bbi _439_ (
        .c(jinkela_wire_259),
        .a(jinkela_wire_13),
        .b(jinkela_wire_457),
        .d(jinkela_wire_240)
    );

    or_bb _609_ (
        .a(jinkela_wire_364),
        .b(jinkela_wire_156),
        .c(jinkela_wire_208)
    );

    maj_bbb _440_ (
        .c(jinkela_wire_305),
        .a(jinkela_wire_275),
        .b(jinkela_wire_270),
        .d(jinkela_wire_360)
    );

    maj_bbi _441_ (
        .c(jinkela_wire_275),
        .a(jinkela_wire_270),
        .b(jinkela_wire_305),
        .d(jinkela_wire_294)
    );

    and_bi _610_ (
        .a(jinkela_wire_208),
        .b(jinkela_wire_318),
        .c(jinkela_wire_251)
    );

    maj_bbi _652_ (
        .c(jinkela_wire_185),
        .a(jinkela_wire_221),
        .b(jinkela_wire_75),
        .d(jinkela_wire_281)
    );

    or_ii _611_ (
        .a(1'b0),
        .b(1'b0),
        .c(jinkela_wire_350)
    );

    maj_bbb _653_ (
        .c(jinkela_wire_185),
        .a(jinkela_wire_202),
        .b(jinkela_wire_441),
        .d(jinkela_wire_288)
    );

    or_ii _612_ (
        .a(jinkela_wire_340),
        .b(jinkela_wire_438),
        .c(jinkela_wire_330)
    );

    maj_bbi _654_ (
        .c(jinkela_wire_202),
        .a(jinkela_wire_441),
        .b(jinkela_wire_185),
        .d(jinkela_wire_180)
    );

    and_ii _613_ (
        .a(jinkela_wire_340),
        .b(jinkela_wire_438),
        .c(jinkela_wire_409)
    );

    maj_bbi _655_ (
        .c(jinkela_wire_288),
        .a(jinkela_wire_180),
        .b(jinkela_wire_202),
        .d(jinkela_wire_406)
    );

    and_bi _614_ (
        .a(jinkela_wire_330),
        .b(jinkela_wire_409),
        .c(jinkela_wire_313)
    );

    maj_bbb _656_ (
        .c(jinkela_wire_20),
        .a(jinkela_wire_329),
        .b(jinkela_wire_31),
        .d(jinkela_wire_441)
    );

    or_bi _615_ (
        .a(jinkela_wire_350),
        .b(jinkela_wire_313),
        .c(jinkela_wire_296)
    );

    maj_bbi _657_ (
        .c(jinkela_wire_329),
        .a(jinkela_wire_31),
        .b(jinkela_wire_20),
        .d(jinkela_wire_468)
    );

    and_bi _616_ (
        .a(jinkela_wire_350),
        .b(jinkela_wire_313),
        .c(jinkela_wire_320)
    );

    maj_bbi _658_ (
        .c(jinkela_wire_441),
        .a(jinkela_wire_468),
        .b(jinkela_wire_329),
        .d(jinkela_wire_361)
    );

    and_bi _617_ (
        .a(jinkela_wire_296),
        .b(jinkela_wire_320),
        .c(jinkela_wire_426)
    );

    maj_bbb _659_ (
        .c(jinkela_wire_281),
        .a(jinkela_wire_386),
        .b(jinkela_wire_361),
        .d(jinkela_wire_202)
    );

    maj_bii _618_ (
        .c(jinkela_wire_438),
        .a(jinkela_wire_350),
        .b(jinkela_wire_340),
        .d(jinkela_wire_371)
    );

    maj_bbi _660_ (
        .c(jinkela_wire_386),
        .a(jinkela_wire_361),
        .b(jinkela_wire_281),
        .d(jinkela_wire_98)
    );

    or_ii _619_ (
        .a(jinkela_wire_186),
        .b(jinkela_wire_442),
        .c(jinkela_wire_399)
    );

    maj_bbi _661_ (
        .c(jinkela_wire_202),
        .a(jinkela_wire_98),
        .b(jinkela_wire_386),
        .d(jinkela_wire_207)
    );

    and_ii _620_ (
        .a(jinkela_wire_186),
        .b(jinkela_wire_442),
        .c(jinkela_wire_134)
    );

    and_bb _662_ (
        .a(jinkela_wire_207),
        .b(jinkela_wire_381),
        .c(jinkela_wire_159)
    );

    and_bi _621_ (
        .a(jinkela_wire_399),
        .b(jinkela_wire_134),
        .c(jinkela_wire_319)
    );

    or_bb _663_ (
        .a(jinkela_wire_207),
        .b(jinkela_wire_381),
        .c(jinkela_wire_56)
    );

    or_bi _622_ (
        .a(jinkela_wire_371),
        .b(jinkela_wire_319),
        .c(jinkela_wire_82)
    );

    and_bi _664_ (
        .a(jinkela_wire_56),
        .b(jinkela_wire_159),
        .c(jinkela_wire_438)
    );

    and_bi _623_ (
        .a(jinkela_wire_371),
        .b(jinkela_wire_319),
        .c(jinkela_wire_324)
    );

    and_bb _665_ (
        .a(jinkela_wire_159),
        .b(jinkela_wire_406),
        .c(jinkela_wire_391)
    );

    and_bi _624_ (
        .a(jinkela_wire_82),
        .b(jinkela_wire_324),
        .c(jinkela_wire_62)
    );

    or_bb _666_ (
        .a(jinkela_wire_159),
        .b(jinkela_wire_406),
        .c(jinkela_wire_439)
    );

    maj_bii _625_ (
        .c(jinkela_wire_442),
        .a(jinkela_wire_371),
        .b(jinkela_wire_186),
        .d(jinkela_wire_335)
    );

    and_bi _667_ (
        .a(jinkela_wire_439),
        .b(jinkela_wire_391),
        .c(jinkela_wire_442)
    );

    or_ii _626_ (
        .a(jinkela_wire_334),
        .b(jinkela_wire_403),
        .c(jinkela_wire_464)
    );

    and_bb _668_ (
        .a(jinkela_wire_391),
        .b(jinkela_wire_288),
        .c(jinkela_wire_217)
    );

    and_ii _627_ (
        .a(jinkela_wire_334),
        .b(jinkela_wire_403),
        .c(jinkela_wire_119)
    );

    or_bb _669_ (
        .a(jinkela_wire_391),
        .b(jinkela_wire_288),
        .c(jinkela_wire_173)
    );

    and_bi _628_ (
        .a(jinkela_wire_464),
        .b(jinkela_wire_119),
        .c(jinkela_wire_341)
    );

    and_bi _670_ (
        .a(jinkela_wire_173),
        .b(jinkela_wire_217),
        .c(jinkela_wire_403)
    );

    or_bi _629_ (
        .a(jinkela_wire_335),
        .b(jinkela_wire_341),
        .c(jinkela_wire_17)
    );

    or_bb _671_ (
        .a(in_1_),
        .b(in_0_),
        .c(jinkela_wire_239)
    );

    and_bi _630_ (
        .a(jinkela_wire_335),
        .b(jinkela_wire_341),
        .c(jinkela_wire_83)
    );

    and_bb _672_ (
        .a(in_3_),
        .b(in_2_),
        .c(jinkela_wire_333)
    );

    and_bi _631_ (
        .a(jinkela_wire_17),
        .b(jinkela_wire_83),
        .c(jinkela_wire_351)
    );

    or_bb _673_ (
        .a(in_5_),
        .b(in_4_),
        .c(jinkela_wire_465)
    );

    maj_bii _632_ (
        .c(jinkela_wire_403),
        .a(jinkela_wire_335),
        .b(jinkela_wire_334),
        .d(jinkela_wire_68)
    );

    and_bb _674_ (
        .a(in_7_),
        .b(in_6_),
        .c(jinkela_wire_191)
    );

    or_ii _633_ (
        .a(jinkela_wire_422),
        .b(jinkela_wire_217),
        .c(jinkela_wire_397)
    );

    or_bb _675_ (
        .a(in_9_),
        .b(in_8_),
        .c(jinkela_wire_266)
    );

    and_ii _634_ (
        .a(jinkela_wire_422),
        .b(jinkela_wire_217),
        .c(jinkela_wire_61)
    );

    and_bb _676_ (
        .a(in_11_),
        .b(in_10_),
        .c(jinkela_wire_440)
    );

    and_bi _635_ (
        .a(jinkela_wire_397),
        .b(jinkela_wire_61),
        .c(jinkela_wire_316)
    );

    or_bb _677_ (
        .a(in_13_),
        .b(in_12_),
        .c(jinkela_wire_161)
    );

    or_bi _636_ (
        .a(jinkela_wire_68),
        .b(jinkela_wire_316),
        .c(jinkela_wire_461)
    );

    and_bb _678_ (
        .a(in_15_),
        .b(in_14_),
        .c(jinkela_wire_19)
    );

    and_bi _637_ (
        .a(jinkela_wire_68),
        .b(jinkela_wire_316),
        .c(jinkela_wire_420)
    );

    maj_bbb _679_ (
        .c(jinkela_wire_239),
        .a(jinkela_wire_465),
        .b(jinkela_wire_333),
        .d(jinkela_wire_219)
    );

    and_bi _638_ (
        .a(jinkela_wire_461),
        .b(jinkela_wire_420),
        .c(jinkela_wire_314)
    );

    maj_bbi _680_ (
        .c(jinkela_wire_465),
        .a(jinkela_wire_333),
        .b(jinkela_wire_239),
        .d(jinkela_wire_183)
    );

    and_ii _639_ (
        .a(1'b0),
        .b(1'b0),
        .c(jinkela_wire_436)
    );

    maj_bbi _681_ (
        .c(jinkela_wire_219),
        .a(jinkela_wire_183),
        .b(jinkela_wire_465),
        .d(jinkela_wire_45)
    );

    and_bi _640_ (
        .a(jinkela_wire_350),
        .b(jinkela_wire_436),
        .c(jinkela_wire_225)
    );

    maj_bbb _682_ (
        .c(jinkela_wire_219),
        .a(jinkela_wire_206),
        .b(jinkela_wire_136),
        .d(jinkela_wire_78)
    );

    maj_bbi _641_ (
        .c(jinkela_wire_68),
        .a(jinkela_wire_422),
        .b(jinkela_wire_217),
        .d(jinkela_wire_254)
    );

    maj_bbi _683_ (
        .c(jinkela_wire_206),
        .a(jinkela_wire_136),
        .b(jinkela_wire_219),
        .d(jinkela_wire_355)
    );

    or_bb _642_ (
        .a(in_17_),
        .b(in_16_),
        .c(jinkela_wire_353)
    );

    maj_bbi _684_ (
        .c(jinkela_wire_78),
        .a(jinkela_wire_355),
        .b(jinkela_wire_206),
        .d(jinkela_wire_287)
    );

    and_bb _643_ (
        .a(in_19_),
        .b(in_18_),
        .c(jinkela_wire_92)
    );

    maj_bbb _685_ (
        .c(jinkela_wire_191),
        .a(jinkela_wire_440),
        .b(jinkela_wire_266),
        .d(jinkela_wire_136)
    );

    or_bb _644_ (
        .a(in_21_),
        .b(in_20_),
        .c(jinkela_wire_75)
    );

    maj_bbi _686_ (
        .c(jinkela_wire_440),
        .a(jinkela_wire_266),
        .b(jinkela_wire_191),
        .d(jinkela_wire_14)
    );

    and_bb _645_ (
        .a(in_23_),
        .b(in_22_),
        .c(jinkela_wire_20)
    );

    maj_bbi _687_ (
        .c(jinkela_wire_136),
        .a(jinkela_wire_14),
        .b(jinkela_wire_440),
        .d(jinkela_wire_446)
    );

    or_bb _646_ (
        .a(in_25_),
        .b(in_24_),
        .c(jinkela_wire_31)
    );

    maj_bbb _688_ (
        .c(jinkela_wire_45),
        .a(jinkela_wire_161),
        .b(jinkela_wire_446),
        .d(jinkela_wire_206)
    );

    and_bb _647_ (
        .a(in_27_),
        .b(in_26_),
        .c(jinkela_wire_329)
    );

    maj_bbi _689_ (
        .c(jinkela_wire_161),
        .a(jinkela_wire_446),
        .b(jinkela_wire_45),
        .d(jinkela_wire_269)
    );

    or_bb _648_ (
        .a(in_29_),
        .b(in_28_),
        .c(jinkela_wire_386)
    );

    maj_bbi _690_ (
        .c(jinkela_wire_206),
        .a(jinkela_wire_269),
        .b(jinkela_wire_161),
        .d(jinkela_wire_6)
    );

    and_bb _649_ (
        .a(in_31_),
        .b(in_30_),
        .c(jinkela_wire_381)
    );

    and_bb _691_ (
        .a(jinkela_wire_6),
        .b(jinkela_wire_19),
        .c(jinkela_wire_212)
    );

    maj_bbb _650_ (
        .c(jinkela_wire_353),
        .a(jinkela_wire_75),
        .b(jinkela_wire_92),
        .d(jinkela_wire_185)
    );

    or_bb _692_ (
        .a(jinkela_wire_6),
        .b(jinkela_wire_19),
        .c(jinkela_wire_448)
    );

    maj_bbi _651_ (
        .c(jinkela_wire_75),
        .a(jinkela_wire_92),
        .b(jinkela_wire_353),
        .d(jinkela_wire_221)
    );

    and_bi _693_ (
        .a(jinkela_wire_448),
        .b(jinkela_wire_212),
        .c(jinkela_wire_340)
    );

    and_bb _694_ (
        .a(jinkela_wire_212),
        .b(jinkela_wire_287),
        .c(jinkela_wire_2)
    );

    or_bb _695_ (
        .a(jinkela_wire_212),
        .b(jinkela_wire_287),
        .c(jinkela_wire_323)
    );

    and_bi _696_ (
        .a(jinkela_wire_323),
        .b(jinkela_wire_2),
        .c(jinkela_wire_186)
    );

    and_bb _697_ (
        .a(jinkela_wire_2),
        .b(jinkela_wire_78),
        .c(jinkela_wire_422)
    );

    or_bb _698_ (
        .a(jinkela_wire_2),
        .b(jinkela_wire_78),
        .c(jinkela_wire_30)
    );

    and_bi _699_ (
        .a(jinkela_wire_30),
        .b(jinkela_wire_422),
        .c(jinkela_wire_334)
    );

    maj_bbi _375_ (
        .c(jinkela_wire_122),
        .a(jinkela_wire_60),
        .b(jinkela_wire_166),
        .d(jinkela_wire_178)
    );

    maj_bbi _376_ (
        .c(jinkela_wire_279),
        .a(jinkela_wire_178),
        .b(jinkela_wire_122),
        .d(jinkela_wire_12)
    );

    maj_bbb _374_ (
        .c(jinkela_wire_166),
        .a(jinkela_wire_122),
        .b(jinkela_wire_60),
        .d(jinkela_wire_279)
    );

    or_ii _269_ (
        .a(jinkela_wire_215),
        .b(jinkela_wire_8),
        .c(jinkela_wire_450)
    );

    and_ii _270_ (
        .a(jinkela_wire_215),
        .b(jinkela_wire_8),
        .c(jinkela_wire_419)
    );

    maj_bii _313_ (
        .c(jinkela_wire_176),
        .a(jinkela_wire_114),
        .b(jinkela_wire_52),
        .d(jinkela_wire_377)
    );

    or_ii _314_ (
        .a(jinkela_wire_94),
        .b(jinkela_wire_171),
        .c(jinkela_wire_205)
    );

    and_ii _315_ (
        .a(jinkela_wire_94),
        .b(jinkela_wire_171),
        .c(jinkela_wire_273)
    );

    and_bi _316_ (
        .a(jinkela_wire_205),
        .b(jinkela_wire_273),
        .c(jinkela_wire_123)
    );

    or_bi _317_ (
        .a(jinkela_wire_377),
        .b(jinkela_wire_123),
        .c(jinkela_wire_408)
    );

    and_bi _318_ (
        .a(jinkela_wire_377),
        .b(jinkela_wire_123),
        .c(jinkela_wire_325)
    );

    and_bi _319_ (
        .a(jinkela_wire_408),
        .b(jinkela_wire_325),
        .c(jinkela_wire_268)
    );

    maj_bii _320_ (
        .c(jinkela_wire_171),
        .a(jinkela_wire_377),
        .b(jinkela_wire_94),
        .d(jinkela_wire_116)
    );

    or_ii _321_ (
        .a(jinkela_wire_190),
        .b(jinkela_wire_132),
        .c(jinkela_wire_149)
    );

    and_ii _322_ (
        .a(jinkela_wire_190),
        .b(jinkela_wire_132),
        .c(jinkela_wire_354)
    );

    and_bi _323_ (
        .a(jinkela_wire_149),
        .b(jinkela_wire_354),
        .c(jinkela_wire_358)
    );

    or_bi _324_ (
        .a(jinkela_wire_116),
        .b(jinkela_wire_358),
        .c(jinkela_wire_113)
    );

    and_bi _325_ (
        .a(jinkela_wire_116),
        .b(jinkela_wire_358),
        .c(jinkela_wire_21)
    );

    and_bi _326_ (
        .a(jinkela_wire_113),
        .b(jinkela_wire_21),
        .c(jinkela_wire_147)
    );

    maj_bii _327_ (
        .c(jinkela_wire_132),
        .a(jinkela_wire_116),
        .b(jinkela_wire_190),
        .d(jinkela_wire_337)
    );

    or_ii _328_ (
        .a(jinkela_wire_148),
        .b(jinkela_wire_36),
        .c(jinkela_wire_392)
    );

    and_ii _329_ (
        .a(jinkela_wire_148),
        .b(jinkela_wire_36),
        .c(jinkela_wire_421)
    );

    and_bi _330_ (
        .a(jinkela_wire_392),
        .b(jinkela_wire_421),
        .c(jinkela_wire_151)
    );

    or_bi _331_ (
        .a(jinkela_wire_337),
        .b(jinkela_wire_151),
        .c(jinkela_wire_264)
    );

    and_bi _332_ (
        .a(jinkela_wire_337),
        .b(jinkela_wire_151),
        .c(jinkela_wire_181)
    );

    and_bi _333_ (
        .a(jinkela_wire_264),
        .b(jinkela_wire_181),
        .c(jinkela_wire_452)
    );

    and_ii _334_ (
        .a(1'b0),
        .b(1'b0),
        .c(jinkela_wire_131)
    );

    and_bi _335_ (
        .a(jinkela_wire_114),
        .b(jinkela_wire_131),
        .c(jinkela_wire_199)
    );

    maj_bbi _336_ (
        .c(jinkela_wire_337),
        .a(jinkela_wire_148),
        .b(jinkela_wire_36),
        .d(jinkela_wire_204)
    );

    or_bb _337_ (
        .a(in_113_),
        .b(in_112_),
        .c(jinkela_wire_35)
    );

    and_bb _338_ (
        .a(in_115_),
        .b(in_114_),
        .c(jinkela_wire_396)
    );

    or_bb _339_ (
        .a(in_117_),
        .b(in_116_),
        .c(jinkela_wire_40)
    );

    and_bb _340_ (
        .a(in_119_),
        .b(in_118_),
        .c(jinkela_wire_295)
    );

    or_bb _341_ (
        .a(in_121_),
        .b(in_120_),
        .c(jinkela_wire_37)
    );

    and_bb _342_ (
        .a(in_123_),
        .b(in_122_),
        .c(jinkela_wire_144)
    );

    or_bb _343_ (
        .a(in_125_),
        .b(in_124_),
        .c(jinkela_wire_192)
    );

    and_bb _344_ (
        .a(in_127_),
        .b(in_126_),
        .c(jinkela_wire_103)
    );

    maj_bbb _345_ (
        .c(jinkela_wire_35),
        .a(jinkela_wire_40),
        .b(jinkela_wire_396),
        .d(jinkela_wire_456)
    );

    maj_bbi _346_ (
        .c(jinkela_wire_40),
        .a(jinkela_wire_396),
        .b(jinkela_wire_35),
        .d(jinkela_wire_284)
    );

    maj_bbi _347_ (
        .c(jinkela_wire_456),
        .a(jinkela_wire_284),
        .b(jinkela_wire_40),
        .d(jinkela_wire_88)
    );

    maj_bbb _348_ (
        .c(jinkela_wire_456),
        .a(jinkela_wire_104),
        .b(jinkela_wire_213),
        .d(jinkela_wire_51)
    );

    maj_bbi _349_ (
        .c(jinkela_wire_104),
        .a(jinkela_wire_213),
        .b(jinkela_wire_456),
        .d(jinkela_wire_424)
    );

    maj_bbi _350_ (
        .c(jinkela_wire_51),
        .a(jinkela_wire_424),
        .b(jinkela_wire_104),
        .d(jinkela_wire_255)
    );

    and_bi _226_ (
        .a(jinkela_wire_229),
        .b(jinkela_wire_46),
        .c(jinkela_wire_378)
    );

    or_ii _224_ (
        .a(jinkela_wire_449),
        .b(jinkela_wire_29),
        .c(jinkela_wire_229)
    );

    maj_bbb _351_ (
        .c(jinkela_wire_295),
        .a(jinkela_wire_144),
        .b(jinkela_wire_37),
        .d(jinkela_wire_213)
    );

    and_ii _225_ (
        .a(jinkela_wire_449),
        .b(jinkela_wire_29),
        .c(jinkela_wire_46)
    );

    maj_bbi _352_ (
        .c(jinkela_wire_144),
        .a(jinkela_wire_37),
        .b(jinkela_wire_295),
        .d(jinkela_wire_3)
    );

    or_ii _223_ (
        .a(jinkela_wire_168),
        .b(jinkela_wire_307),
        .c(jinkela_wire_42)
    );

    maj_bbi _353_ (
        .c(jinkela_wire_213),
        .a(jinkela_wire_3),
        .b(jinkela_wire_144),
        .d(jinkela_wire_274)
    );

    or_bi _227_ (
        .a(jinkela_wire_42),
        .b(jinkela_wire_378),
        .c(jinkela_wire_189)
    );

    and_bi _228_ (
        .a(jinkela_wire_42),
        .b(jinkela_wire_378),
        .c(jinkela_wire_293)
    );

    maj_bbb _354_ (
        .c(jinkela_wire_88),
        .a(jinkela_wire_192),
        .b(jinkela_wire_274),
        .d(jinkela_wire_104)
    );

    and_bi _271_ (
        .a(jinkela_wire_450),
        .b(jinkela_wire_419),
        .c(jinkela_wire_102)
    );

    maj_bbi _355_ (
        .c(jinkela_wire_192),
        .a(jinkela_wire_274),
        .b(jinkela_wire_88),
        .d(jinkela_wire_444)
    );

    or_bi _272_ (
        .a(jinkela_wire_344),
        .b(jinkela_wire_102),
        .c(jinkela_wire_203)
    );

    maj_bbi _356_ (
        .c(jinkela_wire_104),
        .a(jinkela_wire_444),
        .b(jinkela_wire_192),
        .d(jinkela_wire_22)
    );

    and_bi _273_ (
        .a(jinkela_wire_344),
        .b(jinkela_wire_102),
        .c(jinkela_wire_297)
    );

    and_bb _357_ (
        .a(jinkela_wire_22),
        .b(jinkela_wire_103),
        .c(jinkela_wire_317)
    );

    and_bi _274_ (
        .a(jinkela_wire_203),
        .b(jinkela_wire_297),
        .c(jinkela_wire_29)
    );

    or_bb _358_ (
        .a(jinkela_wire_22),
        .b(jinkela_wire_103),
        .c(jinkela_wire_50)
    );

    maj_bii _275_ (
        .c(jinkela_wire_8),
        .a(jinkela_wire_344),
        .b(jinkela_wire_215),
        .d(jinkela_wire_398)
    );

    and_bi _359_ (
        .a(jinkela_wire_50),
        .b(jinkela_wire_317),
        .c(jinkela_wire_176)
    );

    or_ii _276_ (
        .a(jinkela_wire_141),
        .b(jinkela_wire_268),
        .c(jinkela_wire_367)
    );

    and_bb _360_ (
        .a(jinkela_wire_317),
        .b(jinkela_wire_255),
        .c(jinkela_wire_26)
    );

    and_ii _277_ (
        .a(jinkela_wire_141),
        .b(jinkela_wire_268),
        .c(jinkela_wire_262)
    );

    or_bb _361_ (
        .a(jinkela_wire_317),
        .b(jinkela_wire_255),
        .c(jinkela_wire_276)
    );

    and_bi _278_ (
        .a(jinkela_wire_367),
        .b(jinkela_wire_262),
        .c(jinkela_wire_64)
    );

    and_bi _362_ (
        .a(jinkela_wire_276),
        .b(jinkela_wire_26),
        .c(jinkela_wire_171)
    );

    or_bi _279_ (
        .a(jinkela_wire_398),
        .b(jinkela_wire_64),
        .c(jinkela_wire_16)
    );

    and_bb _363_ (
        .a(jinkela_wire_26),
        .b(jinkela_wire_51),
        .c(jinkela_wire_36)
    );

    and_bi _280_ (
        .a(jinkela_wire_398),
        .b(jinkela_wire_64),
        .c(jinkela_wire_348)
    );

    or_bb _364_ (
        .a(jinkela_wire_26),
        .b(jinkela_wire_51),
        .c(jinkela_wire_195)
    );

    and_bi _281_ (
        .a(jinkela_wire_16),
        .b(jinkela_wire_348),
        .c(jinkela_wire_435)
    );

    and_bi _365_ (
        .a(jinkela_wire_195),
        .b(jinkela_wire_36),
        .c(jinkela_wire_132)
    );

    maj_bii _282_ (
        .c(jinkela_wire_268),
        .a(jinkela_wire_398),
        .b(jinkela_wire_141),
        .d(jinkela_wire_187)
    );

    or_bb _366_ (
        .a(in_97_),
        .b(in_96_),
        .c(jinkela_wire_166)
    );

    or_ii _283_ (
        .a(jinkela_wire_394),
        .b(jinkela_wire_147),
        .c(jinkela_wire_412)
    );

    and_bb _367_ (
        .a(in_99_),
        .b(in_98_),
        .c(jinkela_wire_60)
    );

    and_ii _284_ (
        .a(jinkela_wire_394),
        .b(jinkela_wire_147),
        .c(jinkela_wire_121)
    );

    or_bb _368_ (
        .a(in_101_),
        .b(in_100_),
        .c(jinkela_wire_122)
    );

    and_bi _285_ (
        .a(jinkela_wire_412),
        .b(jinkela_wire_121),
        .c(jinkela_wire_376)
    );

    and_bb _369_ (
        .a(in_103_),
        .b(in_102_),
        .c(jinkela_wire_388)
    );

    or_bi _286_ (
        .a(jinkela_wire_187),
        .b(jinkela_wire_376),
        .c(jinkela_wire_107)
    );

    or_bb _370_ (
        .a(in_105_),
        .b(in_104_),
        .c(jinkela_wire_69)
    );

    and_bi _287_ (
        .a(jinkela_wire_187),
        .b(jinkela_wire_376),
        .c(jinkela_wire_245)
    );

    and_bb _371_ (
        .a(in_107_),
        .b(in_106_),
        .c(jinkela_wire_194)
    );

    and_bi _288_ (
        .a(jinkela_wire_107),
        .b(jinkela_wire_245),
        .c(jinkela_wire_230)
    );

    or_bb _372_ (
        .a(in_109_),
        .b(in_108_),
        .c(jinkela_wire_223)
    );

    maj_bii _289_ (
        .c(jinkela_wire_147),
        .a(jinkela_wire_187),
        .b(jinkela_wire_394),
        .d(jinkela_wire_302)
    );

    and_bb _373_ (
        .a(in_111_),
        .b(in_110_),
        .c(jinkela_wire_164)
    );

    or_ii _290_ (
        .a(jinkela_wire_232),
        .b(jinkela_wire_452),
        .c(jinkela_wire_242)
    );

    maj_bbb _377_ (
        .c(jinkela_wire_279),
        .a(jinkela_wire_292),
        .b(jinkela_wire_445),
        .d(jinkela_wire_467)
    );

    and_ii _291_ (
        .a(jinkela_wire_232),
        .b(jinkela_wire_452),
        .c(jinkela_wire_359)
    );

    maj_bbi _378_ (
        .c(jinkela_wire_292),
        .a(jinkela_wire_445),
        .b(jinkela_wire_279),
        .d(jinkela_wire_188)
    );

    and_bi _292_ (
        .a(jinkela_wire_242),
        .b(jinkela_wire_359),
        .c(jinkela_wire_298)
    );

    maj_bbi _379_ (
        .c(jinkela_wire_467),
        .a(jinkela_wire_188),
        .b(jinkela_wire_292),
        .d(jinkela_wire_454)
    );

    or_bi _293_ (
        .a(jinkela_wire_302),
        .b(jinkela_wire_298),
        .c(jinkela_wire_286)
    );

    maj_bbb _380_ (
        .c(jinkela_wire_388),
        .a(jinkela_wire_194),
        .b(jinkela_wire_69),
        .d(jinkela_wire_445)
    );

    and_bi _294_ (
        .a(jinkela_wire_302),
        .b(jinkela_wire_298),
        .c(jinkela_wire_41)
    );

    maj_bbi _381_ (
        .c(jinkela_wire_194),
        .a(jinkela_wire_69),
        .b(jinkela_wire_388),
        .d(jinkela_wire_57)
    );

    and_bi _295_ (
        .a(jinkela_wire_286),
        .b(jinkela_wire_41),
        .c(jinkela_wire_267)
    );

    maj_bbi _382_ (
        .c(jinkela_wire_445),
        .a(jinkela_wire_57),
        .b(jinkela_wire_194),
        .d(jinkela_wire_299)
    );

    maj_bii _296_ (
        .c(jinkela_wire_452),
        .a(jinkela_wire_302),
        .b(jinkela_wire_232),
        .d(jinkela_wire_453)
    );

    maj_bbb _383_ (
        .c(jinkela_wire_12),
        .a(jinkela_wire_223),
        .b(jinkela_wire_299),
        .d(jinkela_wire_292)
    );

    or_ii _297_ (
        .a(jinkela_wire_310),
        .b(jinkela_wire_204),
        .c(jinkela_wire_67)
    );

    maj_bbi _384_ (
        .c(jinkela_wire_223),
        .a(jinkela_wire_299),
        .b(jinkela_wire_12),
        .d(jinkela_wire_216)
    );

    and_ii _298_ (
        .a(jinkela_wire_310),
        .b(jinkela_wire_204),
        .c(jinkela_wire_402)
    );

    maj_bbi _385_ (
        .c(jinkela_wire_292),
        .a(jinkela_wire_216),
        .b(jinkela_wire_223),
        .d(jinkela_wire_38)
    );

    and_bi _299_ (
        .a(jinkela_wire_67),
        .b(jinkela_wire_402),
        .c(jinkela_wire_368)
    );

    and_bb _386_ (
        .a(jinkela_wire_38),
        .b(jinkela_wire_164),
        .c(jinkela_wire_23)
    );

    or_bi _300_ (
        .a(jinkela_wire_453),
        .b(jinkela_wire_368),
        .c(jinkela_wire_97)
    );

    or_bb _387_ (
        .a(jinkela_wire_38),
        .b(jinkela_wire_164),
        .c(jinkela_wire_459)
    );

    and_bi _301_ (
        .a(jinkela_wire_453),
        .b(jinkela_wire_368),
        .c(jinkela_wire_127)
    );

    and_bi _388_ (
        .a(jinkela_wire_459),
        .b(jinkela_wire_23),
        .c(jinkela_wire_52)
    );

    and_bi _302_ (
        .a(jinkela_wire_97),
        .b(jinkela_wire_127),
        .c(jinkela_wire_140)
    );

    and_bb _389_ (
        .a(jinkela_wire_23),
        .b(jinkela_wire_454),
        .c(jinkela_wire_154)
    );

    and_ii _303_ (
        .a(jinkela_wire_34),
        .b(jinkela_wire_199),
        .c(jinkela_wire_5)
    );

    or_bb _390_ (
        .a(jinkela_wire_23),
        .b(jinkela_wire_454),
        .c(jinkela_wire_142)
    );

    and_bi _304_ (
        .a(jinkela_wire_344),
        .b(jinkela_wire_5),
        .c(jinkela_wire_307)
    );

    and_bi _391_ (
        .a(jinkela_wire_142),
        .b(jinkela_wire_154),
        .c(jinkela_wire_94)
    );

    maj_bbi _305_ (
        .c(jinkela_wire_453),
        .a(jinkela_wire_310),
        .b(jinkela_wire_204),
        .d(jinkela_wire_342)
    );

    and_bb _392_ (
        .a(jinkela_wire_154),
        .b(jinkela_wire_467),
        .c(jinkela_wire_148)
    );

    or_ii _306_ (
        .a(1'b0),
        .b(1'b0),
        .c(jinkela_wire_114)
    );

    or_bb _393_ (
        .a(jinkela_wire_154),
        .b(jinkela_wire_467),
        .c(jinkela_wire_336)
    );

    or_ii _307_ (
        .a(jinkela_wire_52),
        .b(jinkela_wire_176),
        .c(jinkela_wire_390)
    );

    and_bi _394_ (
        .a(jinkela_wire_336),
        .b(jinkela_wire_148),
        .c(jinkela_wire_190)
    );

    and_ii _308_ (
        .a(jinkela_wire_52),
        .b(jinkela_wire_176),
        .c(jinkela_wire_369)
    );

    or_ii _395_ (
        .a(1'b0),
        .b(1'b0),
        .c(jinkela_wire_145)
    );

    and_bi _309_ (
        .a(jinkela_wire_390),
        .b(jinkela_wire_369),
        .c(jinkela_wire_416)
    );

    or_ii _396_ (
        .a(jinkela_wire_233),
        .b(jinkela_wire_126),
        .c(jinkela_wire_163)
    );

    or_bi _310_ (
        .a(jinkela_wire_114),
        .b(jinkela_wire_416),
        .c(jinkela_wire_200)
    );

    and_ii _397_ (
        .a(jinkela_wire_233),
        .b(jinkela_wire_126),
        .c(jinkela_wire_110)
    );

    and_bi _311_ (
        .a(jinkela_wire_114),
        .b(jinkela_wire_416),
        .c(jinkela_wire_160)
    );

    and_bi _398_ (
        .a(jinkela_wire_163),
        .b(jinkela_wire_110),
        .c(jinkela_wire_177)
    );

    and_bi _312_ (
        .a(jinkela_wire_200),
        .b(jinkela_wire_160),
        .c(jinkela_wire_8)
    );

    or_bi _399_ (
        .a(jinkela_wire_145),
        .b(jinkela_wire_177),
        .c(jinkela_wire_447)
    );

    and_bi _229_ (
        .a(jinkela_wire_189),
        .b(jinkela_wire_293),
        .c(out_1_)
    );

    maj_bbi _442_ (
        .c(jinkela_wire_360),
        .a(jinkela_wire_294),
        .b(jinkela_wire_275),
        .d(jinkela_wire_226)
    );

    or_ii _484_ (
        .a(jinkela_wire_225),
        .b(jinkela_wire_231),
        .c(jinkela_wire_79)
    );

    or_bi _526_ (
        .a(jinkela_wire_443),
        .b(jinkela_wire_277),
        .c(jinkela_wire_363)
    );

    maj_bbi _568_ (
        .c(jinkela_wire_400),
        .a(jinkela_wire_44),
        .b(jinkela_wire_28),
        .d(jinkela_wire_328)
    );

    maj_bii _230_ (
        .c(jinkela_wire_29),
        .a(jinkela_wire_42),
        .b(jinkela_wire_449),
        .d(jinkela_wire_413)
    );

    maj_bbb _443_ (
        .c(jinkela_wire_73),
        .a(jinkela_wire_146),
        .b(jinkela_wire_226),
        .d(jinkela_wire_457)
    );

    or_ii _485_ (
        .a(jinkela_wire_426),
        .b(jinkela_wire_290),
        .c(jinkela_wire_105)
    );

    and_bi _527_ (
        .a(jinkela_wire_443),
        .b(jinkela_wire_277),
        .c(jinkela_wire_169)
    );

    maj_bbi _569_ (
        .c(jinkela_wire_198),
        .a(jinkela_wire_328),
        .b(jinkela_wire_400),
        .d(jinkela_wire_352)
    );

    or_ii _231_ (
        .a(jinkela_wire_383),
        .b(jinkela_wire_435),
        .c(jinkela_wire_306)
    );

    maj_bbi _444_ (
        .c(jinkela_wire_146),
        .a(jinkela_wire_226),
        .b(jinkela_wire_73),
        .d(jinkela_wire_430)
    );

    and_ii _486_ (
        .a(jinkela_wire_426),
        .b(jinkela_wire_290),
        .c(jinkela_wire_112)
    );

    and_bi _528_ (
        .a(jinkela_wire_363),
        .b(jinkela_wire_169),
        .c(jinkela_wire_290)
    );

    maj_bbb _570_ (
        .c(jinkela_wire_228),
        .a(jinkela_wire_129),
        .b(jinkela_wire_352),
        .d(jinkela_wire_250)
    );

    and_ii _232_ (
        .a(jinkela_wire_383),
        .b(jinkela_wire_435),
        .c(jinkela_wire_58)
    );

    maj_bbi _445_ (
        .c(jinkela_wire_457),
        .a(jinkela_wire_430),
        .b(jinkela_wire_146),
        .d(jinkela_wire_1)
    );

    and_bi _487_ (
        .a(jinkela_wire_105),
        .b(jinkela_wire_112),
        .c(jinkela_wire_55)
    );

    maj_bii _529_ (
        .c(jinkela_wire_433),
        .a(jinkela_wire_443),
        .b(jinkela_wire_315),
        .d(jinkela_wire_196)
    );

    maj_bbi _571_ (
        .c(jinkela_wire_129),
        .a(jinkela_wire_352),
        .b(jinkela_wire_228),
        .d(jinkela_wire_15)
    );

    and_bi _233_ (
        .a(jinkela_wire_306),
        .b(jinkela_wire_58),
        .c(jinkela_wire_414)
    );

    and_bb _446_ (
        .a(jinkela_wire_1),
        .b(jinkela_wire_84),
        .c(jinkela_wire_33)
    );

    or_bi _488_ (
        .a(jinkela_wire_79),
        .b(jinkela_wire_55),
        .c(jinkela_wire_405)
    );

    or_ii _530_ (
        .a(jinkela_wire_76),
        .b(jinkela_wire_133),
        .c(jinkela_wire_238)
    );

    maj_bbi _572_ (
        .c(jinkela_wire_250),
        .a(jinkela_wire_15),
        .b(jinkela_wire_129),
        .d(jinkela_wire_261)
    );

    or_bi _234_ (
        .a(jinkela_wire_413),
        .b(jinkela_wire_414),
        .c(jinkela_wire_417)
    );

    or_bb _447_ (
        .a(jinkela_wire_1),
        .b(jinkela_wire_84),
        .c(jinkela_wire_130)
    );

    and_bi _489_ (
        .a(jinkela_wire_79),
        .b(jinkela_wire_55),
        .c(jinkela_wire_308)
    );

    and_ii _531_ (
        .a(jinkela_wire_76),
        .b(jinkela_wire_133),
        .c(jinkela_wire_282)
    );

    and_bb _573_ (
        .a(jinkela_wire_261),
        .b(jinkela_wire_108),
        .c(jinkela_wire_211)
    );

    and_bi _235_ (
        .a(jinkela_wire_413),
        .b(jinkela_wire_414),
        .c(jinkela_wire_309)
    );

    and_bi _448_ (
        .a(jinkela_wire_130),
        .b(jinkela_wire_33),
        .c(jinkela_wire_126)
    );

    and_bi _490_ (
        .a(jinkela_wire_405),
        .b(jinkela_wire_308),
        .c(jinkela_wire_449)
    );

    and_bi _532_ (
        .a(jinkela_wire_238),
        .b(jinkela_wire_282),
        .c(jinkela_wire_152)
    );

    or_bb _574_ (
        .a(jinkela_wire_261),
        .b(jinkela_wire_108),
        .c(jinkela_wire_53)
    );

    and_bi _236_ (
        .a(jinkela_wire_417),
        .b(jinkela_wire_309),
        .c(out_2_)
    );

    and_bb _449_ (
        .a(jinkela_wire_33),
        .b(jinkela_wire_240),
        .c(jinkela_wire_304)
    );

    maj_bii _491_ (
        .c(jinkela_wire_290),
        .a(jinkela_wire_79),
        .b(jinkela_wire_426),
        .d(jinkela_wire_87)
    );

    or_bi _533_ (
        .a(jinkela_wire_196),
        .b(jinkela_wire_152),
        .c(jinkela_wire_395)
    );

    and_bi _575_ (
        .a(jinkela_wire_53),
        .b(jinkela_wire_211),
        .c(jinkela_wire_433)
    );

    maj_bii _237_ (
        .c(jinkela_wire_435),
        .a(jinkela_wire_413),
        .b(jinkela_wire_383),
        .d(jinkela_wire_311)
    );

    or_bb _450_ (
        .a(jinkela_wire_33),
        .b(jinkela_wire_240),
        .c(jinkela_wire_124)
    );

    or_ii _492_ (
        .a(jinkela_wire_62),
        .b(jinkela_wire_407),
        .c(jinkela_wire_248)
    );

    and_bi _534_ (
        .a(jinkela_wire_196),
        .b(jinkela_wire_152),
        .c(jinkela_wire_85)
    );

    and_bb _576_ (
        .a(jinkela_wire_211),
        .b(jinkela_wire_135),
        .c(jinkela_wire_372)
    );

    or_ii _238_ (
        .a(jinkela_wire_393),
        .b(jinkela_wire_230),
        .c(jinkela_wire_7)
    );

    and_bi _451_ (
        .a(jinkela_wire_124),
        .b(jinkela_wire_304),
        .c(jinkela_wire_462)
    );

    and_ii _493_ (
        .a(jinkela_wire_62),
        .b(jinkela_wire_407),
        .c(jinkela_wire_25)
    );

    and_bi _535_ (
        .a(jinkela_wire_395),
        .b(jinkela_wire_85),
        .c(jinkela_wire_407)
    );

    or_bb _577_ (
        .a(jinkela_wire_211),
        .b(jinkela_wire_135),
        .c(jinkela_wire_91)
    );

    and_ii _239_ (
        .a(jinkela_wire_393),
        .b(jinkela_wire_230),
        .c(jinkela_wire_285)
    );

    and_bb _452_ (
        .a(jinkela_wire_304),
        .b(jinkela_wire_259),
        .c(jinkela_wire_47)
    );

    and_bi _494_ (
        .a(jinkela_wire_248),
        .b(jinkela_wire_25),
        .c(jinkela_wire_70)
    );

    maj_bii _536_ (
        .c(jinkela_wire_133),
        .a(jinkela_wire_196),
        .b(jinkela_wire_76),
        .d(jinkela_wire_283)
    );

    and_bi _578_ (
        .a(jinkela_wire_91),
        .b(jinkela_wire_372),
        .c(jinkela_wire_133)
    );

    and_bi _240_ (
        .a(jinkela_wire_7),
        .b(jinkela_wire_285),
        .c(jinkela_wire_118)
    );

    or_bb _453_ (
        .a(jinkela_wire_304),
        .b(jinkela_wire_259),
        .c(jinkela_wire_175)
    );

    or_bi _495_ (
        .a(jinkela_wire_87),
        .b(jinkela_wire_70),
        .c(jinkela_wire_301)
    );

    or_ii _537_ (
        .a(jinkela_wire_251),
        .b(jinkela_wire_89),
        .c(jinkela_wire_278)
    );

    and_bb _579_ (
        .a(jinkela_wire_372),
        .b(jinkela_wire_260),
        .c(jinkela_wire_63)
    );

    or_bi _241_ (
        .a(jinkela_wire_311),
        .b(jinkela_wire_118),
        .c(jinkela_wire_65)
    );

    and_bi _454_ (
        .a(jinkela_wire_175),
        .b(jinkela_wire_47),
        .c(jinkela_wire_39)
    );

    and_bi _496_ (
        .a(jinkela_wire_87),
        .b(jinkela_wire_70),
        .c(jinkela_wire_257)
    );

    and_ii _538_ (
        .a(jinkela_wire_251),
        .b(jinkela_wire_89),
        .c(jinkela_wire_214)
    );

    or_bb _580_ (
        .a(jinkela_wire_372),
        .b(jinkela_wire_260),
        .c(jinkela_wire_384)
    );

    and_bi _242_ (
        .a(jinkela_wire_311),
        .b(jinkela_wire_118),
        .c(jinkela_wire_93)
    );

    or_bb _455_ (
        .a(in_65_),
        .b(in_64_),
        .c(jinkela_wire_179)
    );

    and_bi _497_ (
        .a(jinkela_wire_301),
        .b(jinkela_wire_257),
        .c(jinkela_wire_383)
    );

    and_bi _539_ (
        .a(jinkela_wire_278),
        .b(jinkela_wire_214),
        .c(jinkela_wire_210)
    );

    and_bi _581_ (
        .a(jinkela_wire_384),
        .b(jinkela_wire_63),
        .c(jinkela_wire_89)
    );

    and_bi _243_ (
        .a(jinkela_wire_65),
        .b(jinkela_wire_93),
        .c(out_3_)
    );

    and_bb _456_ (
        .a(in_67_),
        .b(in_66_),
        .c(jinkela_wire_150)
    );

    maj_bii _498_ (
        .c(jinkela_wire_407),
        .a(jinkela_wire_87),
        .b(jinkela_wire_62),
        .d(jinkela_wire_49)
    );

    or_bi _540_ (
        .a(jinkela_wire_283),
        .b(jinkela_wire_210),
        .c(jinkela_wire_59)
    );

    or_bb _582_ (
        .a(in_33_),
        .b(in_32_),
        .c(jinkela_wire_0)
    );

    maj_bii _244_ (
        .c(jinkela_wire_230),
        .a(jinkela_wire_311),
        .b(jinkela_wire_393),
        .d(jinkela_wire_271)
    );

    or_bb _457_ (
        .a(in_69_),
        .b(in_68_),
        .c(jinkela_wire_415)
    );

    or_ii _499_ (
        .a(jinkela_wire_351),
        .b(jinkela_wire_256),
        .c(jinkela_wire_209)
    );

    and_bi _541_ (
        .a(jinkela_wire_283),
        .b(jinkela_wire_210),
        .c(jinkela_wire_345)
    );

    and_bb _583_ (
        .a(in_35_),
        .b(in_34_),
        .c(jinkela_wire_370)
    );

    or_ii _245_ (
        .a(jinkela_wire_280),
        .b(jinkela_wire_267),
        .c(jinkela_wire_427)
    );

    and_bb _458_ (
        .a(in_71_),
        .b(in_70_),
        .c(jinkela_wire_197)
    );

    and_ii _500_ (
        .a(jinkela_wire_351),
        .b(jinkela_wire_256),
        .c(jinkela_wire_153)
    );

    and_bi _542_ (
        .a(jinkela_wire_59),
        .b(jinkela_wire_345),
        .c(jinkela_wire_256)
    );

    or_bb _584_ (
        .a(in_37_),
        .b(in_36_),
        .c(jinkela_wire_404)
    );

    and_ii _246_ (
        .a(jinkela_wire_280),
        .b(jinkela_wire_267),
        .c(jinkela_wire_258)
    );

    or_bb _459_ (
        .a(in_73_),
        .b(in_72_),
        .c(jinkela_wire_80)
    );

    and_bi _501_ (
        .a(jinkela_wire_209),
        .b(jinkela_wire_153),
        .c(jinkela_wire_109)
    );

    maj_bii _543_ (
        .c(jinkela_wire_89),
        .a(jinkela_wire_283),
        .b(jinkela_wire_251),
        .d(jinkela_wire_432)
    );

    and_bb _585_ (
        .a(in_39_),
        .b(in_38_),
        .c(jinkela_wire_227)
    );

    and_bi _247_ (
        .a(jinkela_wire_427),
        .b(jinkela_wire_258),
        .c(jinkela_wire_111)
    );

    and_bb _460_ (
        .a(in_75_),
        .b(in_74_),
        .c(jinkela_wire_66)
    );

    or_bi _502_ (
        .a(jinkela_wire_49),
        .b(jinkela_wire_109),
        .c(jinkela_wire_162)
    );

    or_ii _544_ (
        .a(jinkela_wire_318),
        .b(jinkela_wire_63),
        .c(jinkela_wire_410)
    );

    or_bb _586_ (
        .a(in_41_),
        .b(in_40_),
        .c(jinkela_wire_172)
    );

    or_bi _248_ (
        .a(jinkela_wire_271),
        .b(jinkela_wire_111),
        .c(jinkela_wire_401)
    );

    or_bb _461_ (
        .a(in_77_),
        .b(in_76_),
        .c(jinkela_wire_365)
    );

    and_bi _503_ (
        .a(jinkela_wire_49),
        .b(jinkela_wire_109),
        .c(jinkela_wire_143)
    );

    and_ii _545_ (
        .a(jinkela_wire_318),
        .b(jinkela_wire_63),
        .c(jinkela_wire_458)
    );

    and_bb _587_ (
        .a(in_43_),
        .b(in_42_),
        .c(jinkela_wire_106)
    );

    and_bi _249_ (
        .a(jinkela_wire_271),
        .b(jinkela_wire_111),
        .c(jinkela_wire_265)
    );

    and_bb _462_ (
        .a(in_79_),
        .b(in_78_),
        .c(jinkela_wire_234)
    );

    and_bi _504_ (
        .a(jinkela_wire_162),
        .b(jinkela_wire_143),
        .c(jinkela_wire_393)
    );

    and_bi _546_ (
        .a(jinkela_wire_410),
        .b(jinkela_wire_458),
        .c(jinkela_wire_139)
    );

    or_bb _588_ (
        .a(in_45_),
        .b(in_44_),
        .c(jinkela_wire_366)
    );

    and_bi _250_ (
        .a(jinkela_wire_401),
        .b(jinkela_wire_265),
        .c(out_4_)
    );

    maj_bbb _463_ (
        .c(jinkela_wire_179),
        .a(jinkela_wire_415),
        .b(jinkela_wire_150),
        .d(jinkela_wire_247)
    );

    maj_bii _505_ (
        .c(jinkela_wire_256),
        .a(jinkela_wire_49),
        .b(jinkela_wire_351),
        .d(jinkela_wire_100)
    );

    or_bi _547_ (
        .a(jinkela_wire_432),
        .b(jinkela_wire_139),
        .c(jinkela_wire_96)
    );

    and_bb _589_ (
        .a(in_47_),
        .b(in_46_),
        .c(jinkela_wire_4)
    );

    maj_bii _251_ (
        .c(jinkela_wire_267),
        .a(jinkela_wire_271),
        .b(jinkela_wire_280),
        .d(jinkela_wire_338)
    );

    maj_bbi _464_ (
        .c(jinkela_wire_415),
        .a(jinkela_wire_150),
        .b(jinkela_wire_179),
        .d(jinkela_wire_18)
    );

    or_ii _506_ (
        .a(jinkela_wire_314),
        .b(jinkela_wire_252),
        .c(jinkela_wire_244)
    );

    and_bi _548_ (
        .a(jinkela_wire_432),
        .b(jinkela_wire_139),
        .c(jinkela_wire_347)
    );

    maj_bbb _590_ (
        .c(jinkela_wire_0),
        .a(jinkela_wire_404),
        .b(jinkela_wire_370),
        .d(jinkela_wire_165)
    );

    or_ii _252_ (
        .a(jinkela_wire_158),
        .b(jinkela_wire_140),
        .c(jinkela_wire_429)
    );

    maj_bbi _465_ (
        .c(jinkela_wire_247),
        .a(jinkela_wire_18),
        .b(jinkela_wire_415),
        .d(jinkela_wire_331)
    );

    and_ii _507_ (
        .a(jinkela_wire_314),
        .b(jinkela_wire_252),
        .c(jinkela_wire_101)
    );

    and_bi _549_ (
        .a(jinkela_wire_96),
        .b(jinkela_wire_347),
        .c(jinkela_wire_252)
    );

    maj_bbi _591_ (
        .c(jinkela_wire_404),
        .a(jinkela_wire_370),
        .b(jinkela_wire_0),
        .d(jinkela_wire_99)
    );

    and_ii _253_ (
        .a(jinkela_wire_158),
        .b(jinkela_wire_140),
        .c(jinkela_wire_246)
    );

    maj_bbb _466_ (
        .c(jinkela_wire_247),
        .a(jinkela_wire_437),
        .b(jinkela_wire_332),
        .d(jinkela_wire_362)
    );

    and_bi _508_ (
        .a(jinkela_wire_244),
        .b(jinkela_wire_101),
        .c(jinkela_wire_339)
    );

    and_ii _550_ (
        .a(1'b0),
        .b(1'b0),
        .c(jinkela_wire_463)
    );

    maj_bbi _592_ (
        .c(jinkela_wire_165),
        .a(jinkela_wire_99),
        .b(jinkela_wire_404),
        .d(jinkela_wire_243)
    );

    and_bi _254_ (
        .a(jinkela_wire_429),
        .b(jinkela_wire_246),
        .c(jinkela_wire_466)
    );

    maj_bbi _467_ (
        .c(jinkela_wire_437),
        .a(jinkela_wire_332),
        .b(jinkela_wire_247),
        .d(jinkela_wire_300)
    );

    or_bi _509_ (
        .a(jinkela_wire_100),
        .b(jinkela_wire_339),
        .c(jinkela_wire_11)
    );

    and_bi _551_ (
        .a(jinkela_wire_443),
        .b(jinkela_wire_463),
        .c(jinkela_wire_231)
    );

    maj_bbb _593_ (
        .c(jinkela_wire_165),
        .a(jinkela_wire_237),
        .b(jinkela_wire_125),
        .d(jinkela_wire_156)
    );

    or_bi _255_ (
        .a(jinkela_wire_338),
        .b(jinkela_wire_466),
        .c(jinkela_wire_272)
    );

    maj_bbi _468_ (
        .c(jinkela_wire_362),
        .a(jinkela_wire_300),
        .b(jinkela_wire_437),
        .d(jinkela_wire_291)
    );

    and_bi _510_ (
        .a(jinkela_wire_100),
        .b(jinkela_wire_339),
        .c(jinkela_wire_418)
    );

    maj_bbi _552_ (
        .c(jinkela_wire_432),
        .a(jinkela_wire_318),
        .b(jinkela_wire_63),
        .d(jinkela_wire_220)
    );

    maj_bbi _594_ (
        .c(jinkela_wire_237),
        .a(jinkela_wire_125),
        .b(jinkela_wire_165),
        .d(jinkela_wire_95)
    );

    and_bi _256_ (
        .a(jinkela_wire_338),
        .b(jinkela_wire_466),
        .c(jinkela_wire_322)
    );

    maj_bbb _469_ (
        .c(jinkela_wire_197),
        .a(jinkela_wire_66),
        .b(jinkela_wire_80),
        .d(jinkela_wire_332)
    );

    and_bi _511_ (
        .a(jinkela_wire_11),
        .b(jinkela_wire_418),
        .c(jinkela_wire_280)
    );

    or_bb _553_ (
        .a(in_49_),
        .b(in_48_),
        .c(jinkela_wire_349)
    );

    maj_bbi _595_ (
        .c(jinkela_wire_156),
        .a(jinkela_wire_95),
        .b(jinkela_wire_237),
        .d(jinkela_wire_24)
    );

    and_bi _257_ (
        .a(jinkela_wire_272),
        .b(jinkela_wire_322),
        .c(out_5_)
    );

    maj_bbi _470_ (
        .c(jinkela_wire_66),
        .a(jinkela_wire_80),
        .b(jinkela_wire_197),
        .d(jinkela_wire_218)
    );

    maj_bii _512_ (
        .c(jinkela_wire_252),
        .a(jinkela_wire_100),
        .b(jinkela_wire_314),
        .d(jinkela_wire_343)
    );

    and_bb _554_ (
        .a(in_51_),
        .b(in_50_),
        .c(jinkela_wire_157)
    );

    maj_bbb _596_ (
        .c(jinkela_wire_227),
        .a(jinkela_wire_106),
        .b(jinkela_wire_172),
        .d(jinkela_wire_125)
    );

    maj_bii _258_ (
        .c(jinkela_wire_140),
        .a(jinkela_wire_338),
        .b(jinkela_wire_158),
        .d(jinkela_wire_460)
    );

    maj_bbi _471_ (
        .c(jinkela_wire_332),
        .a(jinkela_wire_218),
        .b(jinkela_wire_66),
        .d(jinkela_wire_120)
    );

    or_ii _513_ (
        .a(jinkela_wire_254),
        .b(jinkela_wire_220),
        .c(jinkela_wire_10)
    );

    or_bb _555_ (
        .a(in_53_),
        .b(in_52_),
        .c(jinkela_wire_74)
    );

    maj_bbi _597_ (
        .c(jinkela_wire_106),
        .a(jinkela_wire_172),
        .b(jinkela_wire_227),
        .d(jinkela_wire_326)
    );

    or_ii _259_ (
        .a(jinkela_wire_117),
        .b(jinkela_wire_342),
        .c(jinkela_wire_327)
    );

    maj_bbb _472_ (
        .c(jinkela_wire_331),
        .a(jinkela_wire_365),
        .b(jinkela_wire_120),
        .d(jinkela_wire_437)
    );

    and_ii _514_ (
        .a(jinkela_wire_254),
        .b(jinkela_wire_220),
        .c(jinkela_wire_27)
    );

    and_bb _556_ (
        .a(in_55_),
        .b(in_54_),
        .c(jinkela_wire_28)
    );

    maj_bbi _598_ (
        .c(jinkela_wire_125),
        .a(jinkela_wire_326),
        .b(jinkela_wire_106),
        .d(jinkela_wire_115)
    );

    and_ii _260_ (
        .a(jinkela_wire_117),
        .b(jinkela_wire_342),
        .c(jinkela_wire_387)
    );

    maj_bbi _473_ (
        .c(jinkela_wire_365),
        .a(jinkela_wire_120),
        .b(jinkela_wire_331),
        .d(jinkela_wire_431)
    );

    and_bi _515_ (
        .a(jinkela_wire_10),
        .b(jinkela_wire_27),
        .c(jinkela_wire_236)
    );

    or_bb _557_ (
        .a(in_57_),
        .b(in_56_),
        .c(jinkela_wire_44)
    );

    maj_bbb _599_ (
        .c(jinkela_wire_243),
        .a(jinkela_wire_366),
        .b(jinkela_wire_115),
        .d(jinkela_wire_237)
    );

    and_bi _261_ (
        .a(jinkela_wire_327),
        .b(jinkela_wire_387),
        .c(jinkela_wire_312)
    );

    maj_bbi _474_ (
        .c(jinkela_wire_437),
        .a(jinkela_wire_431),
        .b(jinkela_wire_365),
        .d(jinkela_wire_357)
    );

    or_bi _516_ (
        .a(jinkela_wire_343),
        .b(jinkela_wire_236),
        .c(jinkela_wire_48)
    );

    and_bb _558_ (
        .a(in_59_),
        .b(in_58_),
        .c(jinkela_wire_400)
    );

    maj_bbi _600_ (
        .c(jinkela_wire_366),
        .a(jinkela_wire_115),
        .b(jinkela_wire_243),
        .d(jinkela_wire_346)
    );

    or_bi _262_ (
        .a(jinkela_wire_460),
        .b(jinkela_wire_312),
        .c(jinkela_wire_155)
    );

    and_bb _475_ (
        .a(jinkela_wire_357),
        .b(jinkela_wire_234),
        .c(jinkela_wire_170)
    );

    and_bi _517_ (
        .a(jinkela_wire_343),
        .b(jinkela_wire_236),
        .c(jinkela_wire_423)
    );

    or_bb _559_ (
        .a(in_61_),
        .b(in_60_),
        .c(jinkela_wire_129)
    );

    maj_bbi _601_ (
        .c(jinkela_wire_237),
        .a(jinkela_wire_346),
        .b(jinkela_wire_366),
        .d(jinkela_wire_43)
    );

    and_bi _263_ (
        .a(jinkela_wire_460),
        .b(jinkela_wire_312),
        .c(jinkela_wire_128)
    );

    or_bb _476_ (
        .a(jinkela_wire_357),
        .b(jinkela_wire_234),
        .c(jinkela_wire_137)
    );

    and_bi _518_ (
        .a(jinkela_wire_48),
        .b(jinkela_wire_423),
        .c(jinkela_wire_158)
    );

    and_bb _560_ (
        .a(in_63_),
        .b(in_62_),
        .c(jinkela_wire_108)
    );

    and_bb _602_ (
        .a(jinkela_wire_43),
        .b(jinkela_wire_4),
        .c(jinkela_wire_9)
    );

    and_bi _264_ (
        .a(jinkela_wire_155),
        .b(jinkela_wire_128),
        .c(out_6_)
    );

    and_bi _477_ (
        .a(jinkela_wire_137),
        .b(jinkela_wire_170),
        .c(jinkela_wire_233)
    );

    and_ii _519_ (
        .a(jinkela_wire_225),
        .b(jinkela_wire_231),
        .c(jinkela_wire_81)
    );

    maj_bbb _561_ (
        .c(jinkela_wire_349),
        .a(jinkela_wire_74),
        .b(jinkela_wire_157),
        .d(jinkela_wire_428)
    );

    or_bb _603_ (
        .a(jinkela_wire_43),
        .b(jinkela_wire_4),
        .c(jinkela_wire_184)
    );

    maj_bbi _265_ (
        .c(jinkela_wire_460),
        .a(jinkela_wire_117),
        .b(jinkela_wire_342),
        .d(out_7_)
    );

    and_bb _478_ (
        .a(jinkela_wire_170),
        .b(jinkela_wire_291),
        .c(jinkela_wire_90)
    );

    and_bi _520_ (
        .a(jinkela_wire_79),
        .b(jinkela_wire_81),
        .c(jinkela_wire_168)
    );

    maj_bbi _562_ (
        .c(jinkela_wire_74),
        .a(jinkela_wire_157),
        .b(jinkela_wire_349),
        .d(jinkela_wire_201)
    );

    and_bi _604_ (
        .a(jinkela_wire_184),
        .b(jinkela_wire_9),
        .c(jinkela_wire_315)
    );

    and_ii _266_ (
        .a(jinkela_wire_168),
        .b(jinkela_wire_307),
        .c(jinkela_wire_54)
    );

    or_bb _479_ (
        .a(jinkela_wire_170),
        .b(jinkela_wire_291),
        .c(jinkela_wire_241)
    );

    maj_bbi _521_ (
        .c(jinkela_wire_343),
        .a(jinkela_wire_254),
        .b(jinkela_wire_220),
        .d(jinkela_wire_117)
    );

    maj_bbi _563_ (
        .c(jinkela_wire_428),
        .a(jinkela_wire_201),
        .b(jinkela_wire_74),
        .d(jinkela_wire_228)
    );

    and_bb _605_ (
        .a(jinkela_wire_9),
        .b(jinkela_wire_24),
        .c(jinkela_wire_364)
    );

    and_bi _267_ (
        .a(jinkela_wire_42),
        .b(jinkela_wire_54),
        .c(out_0_)
    );

    and_bi _480_ (
        .a(jinkela_wire_241),
        .b(jinkela_wire_90),
        .c(jinkela_wire_86)
    );

    or_ii _522_ (
        .a(1'b0),
        .b(1'b0),
        .c(jinkela_wire_443)
    );

    maj_bbb _564_ (
        .c(jinkela_wire_428),
        .a(jinkela_wire_250),
        .b(jinkela_wire_198),
        .d(jinkela_wire_260)
    );

    or_bb _606_ (
        .a(jinkela_wire_9),
        .b(jinkela_wire_24),
        .c(jinkela_wire_356)
    );

    or_ii _268_ (
        .a(jinkela_wire_34),
        .b(jinkela_wire_199),
        .c(jinkela_wire_344)
    );

    and_bb _481_ (
        .a(jinkela_wire_90),
        .b(jinkela_wire_362),
        .c(jinkela_wire_193)
    );

    or_ii _523_ (
        .a(jinkela_wire_315),
        .b(jinkela_wire_433),
        .c(jinkela_wire_411)
    );

    maj_bbi _565_ (
        .c(jinkela_wire_250),
        .a(jinkela_wire_198),
        .b(jinkela_wire_428),
        .d(jinkela_wire_375)
    );

    and_bi _607_ (
        .a(jinkela_wire_356),
        .b(jinkela_wire_364),
        .c(jinkela_wire_76)
    );

    or_bb _482_ (
        .a(jinkela_wire_90),
        .b(jinkela_wire_362),
        .c(jinkela_wire_451)
    );

    and_bi _483_ (
        .a(jinkela_wire_451),
        .b(jinkela_wire_193),
        .c(jinkela_wire_455)
    );

endmodule
