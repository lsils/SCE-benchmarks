module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n40 , n41 , n42 , n43 , n44 , n45 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n86 , n87 , n89 , n90 , n92 , n93 , n95 , n96 , n98 , n100 , n102 , n103 , n105 , n106 , n107 , n109 , n111 , n112 , n113 , n115 , n116 , n117 , n119 , n120 , n121 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n148 , n149 , n150 , n151 , n152 , n153 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n224 , n225 , n227 , n228 , n230 , n231 , n233 , n234 , n236 , n237 , n238 , n239 , n240 , n242 , n243 , n244 , n246 , n247 , n248 , n250 , n251 , n253 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n266 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n300 , n301 , n302 , n303 , n304 , n305 , n307 , n308 , n309 , n310 , n311 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n322 , n323 , n324 , n325 , n326 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n336 , n337 , n338 , n339 , n340 , n341 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n351 , n352 , n353 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n363 , n364 , n365 , n366 , n367 , n368 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n402 , n403 , n404 , n405 , n406 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n417 , n418 , n419 , n420 , n421 , n422 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n453 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n480 , n481 , n482 , n483 , n484 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n511 , n512 , n514 , n515 , n516 , n517 , n518 , n520 , n521 , n522 , n523 , n524 , n526 , n527 , n528 , n529 , n531 , n532 , n533 , n534 , n536 , n537 , n538 , n539 , n540 , n542 , n543 , n544 , n546 , n547 , n548 , n550 , n551 , n552 , n554 , n555 , n556 , n557 , n558 , n560 , n561 , n562 , n564 , n566 , n568 , n569 , n570 , n571 , n572 , n574 , n575 , n576 , n577 , n578 , n580 , n581 , n582 , n583 , n584 , n586 , n587 , n588 , n590 , n591 , n592 , n594 , n595 , n596 , n598 , n599 , n600 , n601 , n602 , n604 , n605 , n606 , n608 , n609 , n610 , n611 , n613 , n614 , n615 , n616 , n618 , n619 , n620 , n621 , n623 , n624 , n625 , n627 , n628 , n629 , n630 , n631 , n633 , n634 , n635 , n637 , n638 , n639 , n640 , n642 , n643 , n645 , n646 , n647 , n648 , n649 , n651 , n652 , n654 , n655 , n656 , n657 , n658 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n685 , n686 , n687 , n688 , n689 , n690 , n692 , n693 , n694 , n695 , n696 , n698 , n699 , n700 , n701 , n702 , n704 , n705 , n706 , n707 , n708 , n709 , n711 , n712 , n714 , n715 , n716 , n717 , n719 , n720 , n722 , n723 , n724 , n725 , n726 , n727 , n729 , n730 , n731 , n733 , n734 , n735 , n736 , n738 , n739 , n740 , n742 , n743 , n744 , n746 , n747 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n799 , n800 , n801 , n802 , n803 , n805 , n806 , n807 , n808 , n809 , n811 , n812 , n813 , n814 , n816 , n817 , n818 , n819 , n820 , n821 , n823 , n824 , n825 , n826 , n828 , n829 , n830 , n831 , n832 , n834 , n835 , n836 , n837 , n838 , n840 , n841 , n842 , n843 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n856 , n857 , n858 , n859 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n886 , n887 , n888 , n889 , n890 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n917 , n918 , n919 , n920 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n947 , n948 , n949 , n950 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n986 , n987 , n988 , n989 , n990 , n992 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1314 , n1315 , n1316 , n1317 , n1318 , n1320 , n1321 , n1322 , n1324 , n1325 , n1326 , n1327 , n1328 , n1330 , n1331 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1343 , n1344 , n1345 , n1347 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1374 , n1375 , n1376 , n1377 , n1378 , n1380 , n1381 , n1382 , n1383 , n1384 , n1386 , n1387 , n1388 , n1389 , n1390 , n1392 , n1393 , n1394 , n1395 , n1396 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 ;
  buffer buf_n486( .i (x65), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  buffer buf_n489( .i (n488), .o (n489) );
  buffer buf_n490( .i (n489), .o (n490) );
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  buffer buf_n496( .i (n495), .o (n496) );
  buffer buf_n497( .i (n496), .o (n497) );
  buffer buf_n498( .i (n497), .o (n498) );
  buffer buf_n499( .i (n498), .o (n499) );
  buffer buf_n500( .i (n499), .o (n500) );
  buffer buf_n501( .i (n500), .o (n501) );
  buffer buf_n502( .i (n501), .o (n502) );
  buffer buf_n503( .i (n502), .o (n503) );
  buffer buf_n504( .i (n503), .o (n504) );
  buffer buf_n505( .i (n504), .o (n505) );
  buffer buf_n506( .i (n505), .o (n506) );
  buffer buf_n507( .i (n506), .o (n507) );
  buffer buf_n508( .i (n507), .o (n508) );
  buffer buf_n509( .i (n508), .o (n509) );
  buffer buf_n749( .i (x112), .o (n749) );
  buffer buf_n750( .i (n749), .o (n750) );
  buffer buf_n751( .i (n750), .o (n751) );
  buffer buf_n752( .i (n751), .o (n752) );
  buffer buf_n753( .i (n752), .o (n753) );
  buffer buf_n754( .i (n753), .o (n754) );
  buffer buf_n755( .i (n754), .o (n755) );
  buffer buf_n756( .i (n755), .o (n756) );
  buffer buf_n757( .i (n756), .o (n757) );
  buffer buf_n758( .i (n757), .o (n758) );
  buffer buf_n759( .i (n758), .o (n759) );
  buffer buf_n760( .i (n759), .o (n760) );
  buffer buf_n761( .i (n760), .o (n761) );
  buffer buf_n762( .i (n761), .o (n762) );
  buffer buf_n763( .i (n762), .o (n763) );
  buffer buf_n764( .i (n763), .o (n764) );
  buffer buf_n765( .i (n764), .o (n765) );
  buffer buf_n766( .i (n765), .o (n766) );
  buffer buf_n767( .i (n766), .o (n767) );
  buffer buf_n768( .i (n767), .o (n768) );
  buffer buf_n769( .i (n768), .o (n769) );
  buffer buf_n770( .i (n769), .o (n770) );
  buffer buf_n771( .i (n770), .o (n771) );
  buffer buf_n772( .i (n771), .o (n772) );
  buffer buf_n1349( .i (x164), .o (n1349) );
  buffer buf_n1350( .i (n1349), .o (n1350) );
  buffer buf_n1351( .i (n1350), .o (n1351) );
  buffer buf_n1352( .i (n1351), .o (n1352) );
  buffer buf_n1353( .i (n1352), .o (n1353) );
  buffer buf_n1354( .i (n1353), .o (n1354) );
  buffer buf_n1355( .i (n1354), .o (n1355) );
  buffer buf_n1356( .i (n1355), .o (n1356) );
  buffer buf_n1357( .i (n1356), .o (n1357) );
  buffer buf_n1358( .i (n1357), .o (n1358) );
  buffer buf_n1359( .i (n1358), .o (n1359) );
  buffer buf_n1360( .i (n1359), .o (n1360) );
  buffer buf_n1361( .i (n1360), .o (n1361) );
  buffer buf_n1362( .i (n1361), .o (n1362) );
  buffer buf_n1363( .i (n1362), .o (n1363) );
  buffer buf_n1364( .i (n1363), .o (n1364) );
  buffer buf_n1365( .i (n1364), .o (n1365) );
  buffer buf_n1366( .i (n1365), .o (n1366) );
  buffer buf_n1367( .i (n1366), .o (n1367) );
  buffer buf_n1368( .i (n1367), .o (n1368) );
  buffer buf_n1369( .i (n1368), .o (n1369) );
  buffer buf_n1370( .i (n1369), .o (n1370) );
  buffer buf_n1371( .i (n1370), .o (n1371) );
  buffer buf_n1372( .i (n1371), .o (n1372) );
  buffer buf_n1179( .i (x150), .o (n1179) );
  buffer buf_n1180( .i (n1179), .o (n1180) );
  buffer buf_n1181( .i (n1180), .o (n1181) );
  buffer buf_n1182( .i (n1181), .o (n1182) );
  buffer buf_n1183( .i (n1182), .o (n1183) );
  buffer buf_n1184( .i (n1183), .o (n1184) );
  buffer buf_n1185( .i (n1184), .o (n1185) );
  buffer buf_n1186( .i (n1185), .o (n1186) );
  buffer buf_n1187( .i (n1186), .o (n1187) );
  buffer buf_n1188( .i (n1187), .o (n1188) );
  buffer buf_n1189( .i (n1188), .o (n1189) );
  buffer buf_n1190( .i (n1189), .o (n1190) );
  buffer buf_n1191( .i (n1190), .o (n1191) );
  buffer buf_n1192( .i (n1191), .o (n1192) );
  buffer buf_n1193( .i (n1192), .o (n1193) );
  buffer buf_n1194( .i (n1193), .o (n1194) );
  buffer buf_n1195( .i (n1194), .o (n1195) );
  buffer buf_n1196( .i (n1195), .o (n1196) );
  buffer buf_n1197( .i (n1196), .o (n1197) );
  buffer buf_n1198( .i (n1197), .o (n1198) );
  buffer buf_n1199( .i (n1198), .o (n1199) );
  buffer buf_n1200( .i (n1199), .o (n1200) );
  buffer buf_n1201( .i (n1200), .o (n1201) );
  buffer buf_n1202( .i (n1201), .o (n1202) );
  buffer buf_n892( .i (x126), .o (n892) );
  buffer buf_n893( .i (n892), .o (n893) );
  buffer buf_n894( .i (n893), .o (n894) );
  buffer buf_n895( .i (n894), .o (n895) );
  buffer buf_n896( .i (n895), .o (n896) );
  buffer buf_n897( .i (n896), .o (n897) );
  buffer buf_n898( .i (n897), .o (n898) );
  buffer buf_n899( .i (n898), .o (n899) );
  buffer buf_n900( .i (n899), .o (n900) );
  buffer buf_n901( .i (n900), .o (n901) );
  buffer buf_n902( .i (n901), .o (n902) );
  buffer buf_n903( .i (n902), .o (n903) );
  buffer buf_n904( .i (n903), .o (n904) );
  buffer buf_n905( .i (n904), .o (n905) );
  buffer buf_n906( .i (n905), .o (n906) );
  buffer buf_n907( .i (n906), .o (n907) );
  buffer buf_n908( .i (n907), .o (n908) );
  buffer buf_n909( .i (n908), .o (n909) );
  buffer buf_n910( .i (n909), .o (n910) );
  buffer buf_n911( .i (n910), .o (n911) );
  buffer buf_n912( .i (n911), .o (n912) );
  buffer buf_n913( .i (n912), .o (n913) );
  buffer buf_n914( .i (n913), .o (n914) );
  buffer buf_n915( .i (n914), .o (n915) );
  buffer buf_n952( .i (x130), .o (n952) );
  buffer buf_n953( .i (n952), .o (n953) );
  buffer buf_n954( .i (n953), .o (n954) );
  buffer buf_n955( .i (n954), .o (n955) );
  buffer buf_n956( .i (n955), .o (n956) );
  buffer buf_n957( .i (n956), .o (n957) );
  buffer buf_n958( .i (n957), .o (n958) );
  buffer buf_n959( .i (n958), .o (n959) );
  buffer buf_n960( .i (n959), .o (n960) );
  buffer buf_n961( .i (n960), .o (n961) );
  buffer buf_n962( .i (n961), .o (n962) );
  buffer buf_n963( .i (n962), .o (n963) );
  buffer buf_n964( .i (n963), .o (n964) );
  buffer buf_n965( .i (n964), .o (n965) );
  buffer buf_n966( .i (n965), .o (n966) );
  buffer buf_n967( .i (n966), .o (n967) );
  buffer buf_n968( .i (n967), .o (n968) );
  buffer buf_n969( .i (n968), .o (n969) );
  buffer buf_n970( .i (n969), .o (n970) );
  buffer buf_n971( .i (n970), .o (n971) );
  buffer buf_n972( .i (n971), .o (n972) );
  buffer buf_n973( .i (n972), .o (n973) );
  buffer buf_n974( .i (n973), .o (n974) );
  buffer buf_n975( .i (n974), .o (n975) );
  buffer buf_n1229( .i (x152), .o (n1229) );
  buffer buf_n1230( .i (n1229), .o (n1230) );
  buffer buf_n1231( .i (n1230), .o (n1231) );
  buffer buf_n1232( .i (n1231), .o (n1232) );
  buffer buf_n1233( .i (n1232), .o (n1233) );
  buffer buf_n1234( .i (n1233), .o (n1234) );
  buffer buf_n1280( .i (x155), .o (n1280) );
  buffer buf_n1281( .i (n1280), .o (n1281) );
  buffer buf_n1282( .i (n1281), .o (n1282) );
  buffer buf_n1283( .i (n1282), .o (n1283) );
  buffer buf_n1284( .i (n1283), .o (n1284) );
  buffer buf_n1285( .i (n1284), .o (n1285) );
  assign n1535 = n1234 & n1285 ;
  buffer buf_n1536( .i (n1535), .o (n1536) );
  buffer buf_n1537( .i (n1536), .o (n1537) );
  buffer buf_n1538( .i (n1537), .o (n1538) );
  buffer buf_n1539( .i (n1538), .o (n1539) );
  buffer buf_n1540( .i (n1539), .o (n1540) );
  buffer buf_n1541( .i (n1540), .o (n1541) );
  buffer buf_n1542( .i (n1541), .o (n1542) );
  buffer buf_n1543( .i (n1542), .o (n1543) );
  buffer buf_n1544( .i (n1543), .o (n1544) );
  buffer buf_n1545( .i (n1544), .o (n1545) );
  buffer buf_n1546( .i (n1545), .o (n1546) );
  buffer buf_n1547( .i (n1546), .o (n1547) );
  buffer buf_n1548( .i (n1547), .o (n1548) );
  buffer buf_n1549( .i (n1548), .o (n1549) );
  buffer buf_n1550( .i (n1549), .o (n1550) );
  buffer buf_n1551( .i (n1550), .o (n1551) );
  buffer buf_n1552( .i (n1551), .o (n1552) );
  buffer buf_n1204( .i (x151), .o (n1204) );
  buffer buf_n1205( .i (n1204), .o (n1205) );
  buffer buf_n1206( .i (n1205), .o (n1206) );
  buffer buf_n1207( .i (n1206), .o (n1207) );
  buffer buf_n1208( .i (n1207), .o (n1208) );
  buffer buf_n1209( .i (n1208), .o (n1209) );
  buffer buf_n1210( .i (n1209), .o (n1210) );
  buffer buf_n1211( .i (n1210), .o (n1211) );
  buffer buf_n1212( .i (n1211), .o (n1212) );
  buffer buf_n1213( .i (n1212), .o (n1213) );
  buffer buf_n1214( .i (n1213), .o (n1214) );
  buffer buf_n1215( .i (n1214), .o (n1215) );
  buffer buf_n1216( .i (n1215), .o (n1216) );
  buffer buf_n1217( .i (n1216), .o (n1217) );
  buffer buf_n1218( .i (n1217), .o (n1218) );
  buffer buf_n1219( .i (n1218), .o (n1219) );
  buffer buf_n1220( .i (n1219), .o (n1220) );
  buffer buf_n1221( .i (n1220), .o (n1221) );
  buffer buf_n1222( .i (n1221), .o (n1222) );
  buffer buf_n1223( .i (n1222), .o (n1223) );
  buffer buf_n1224( .i (n1223), .o (n1224) );
  buffer buf_n1225( .i (n1224), .o (n1225) );
  buffer buf_n1226( .i (n1225), .o (n1226) );
  buffer buf_n1227( .i (n1226), .o (n1227) );
  buffer buf_n861( .i (x124), .o (n861) );
  buffer buf_n862( .i (n861), .o (n862) );
  buffer buf_n863( .i (n862), .o (n863) );
  buffer buf_n864( .i (n863), .o (n864) );
  buffer buf_n865( .i (n864), .o (n865) );
  buffer buf_n866( .i (n865), .o (n866) );
  buffer buf_n867( .i (n866), .o (n867) );
  buffer buf_n868( .i (n867), .o (n868) );
  buffer buf_n869( .i (n868), .o (n869) );
  buffer buf_n870( .i (n869), .o (n870) );
  buffer buf_n871( .i (n870), .o (n871) );
  buffer buf_n872( .i (n871), .o (n872) );
  buffer buf_n873( .i (n872), .o (n873) );
  buffer buf_n874( .i (n873), .o (n874) );
  buffer buf_n875( .i (n874), .o (n875) );
  buffer buf_n876( .i (n875), .o (n876) );
  buffer buf_n877( .i (n876), .o (n877) );
  buffer buf_n878( .i (n877), .o (n878) );
  buffer buf_n879( .i (n878), .o (n879) );
  buffer buf_n880( .i (n879), .o (n880) );
  buffer buf_n881( .i (n880), .o (n881) );
  buffer buf_n882( .i (n881), .o (n882) );
  buffer buf_n883( .i (n882), .o (n883) );
  buffer buf_n884( .i (n883), .o (n884) );
  buffer buf_n922( .i (x128), .o (n922) );
  buffer buf_n923( .i (n922), .o (n923) );
  buffer buf_n924( .i (n923), .o (n924) );
  buffer buf_n925( .i (n924), .o (n925) );
  buffer buf_n926( .i (n925), .o (n926) );
  buffer buf_n927( .i (n926), .o (n927) );
  buffer buf_n928( .i (n927), .o (n928) );
  buffer buf_n929( .i (n928), .o (n929) );
  buffer buf_n930( .i (n929), .o (n930) );
  buffer buf_n931( .i (n930), .o (n931) );
  buffer buf_n932( .i (n931), .o (n932) );
  buffer buf_n933( .i (n932), .o (n933) );
  buffer buf_n934( .i (n933), .o (n934) );
  buffer buf_n935( .i (n934), .o (n935) );
  buffer buf_n936( .i (n935), .o (n936) );
  buffer buf_n937( .i (n936), .o (n937) );
  buffer buf_n938( .i (n937), .o (n938) );
  buffer buf_n939( .i (n938), .o (n939) );
  buffer buf_n940( .i (n939), .o (n940) );
  buffer buf_n941( .i (n940), .o (n941) );
  buffer buf_n942( .i (n941), .o (n942) );
  buffer buf_n943( .i (n942), .o (n943) );
  buffer buf_n944( .i (n943), .o (n944) );
  buffer buf_n945( .i (n944), .o (n945) );
  buffer buf_n511( .i (x66), .o (n511) );
  buffer buf_n512( .i (n511), .o (n512) );
  assign n1553 = n487 & n512 ;
  buffer buf_n1554( .i (n1553), .o (n1554) );
  buffer buf_n1555( .i (n1554), .o (n1555) );
  buffer buf_n1556( .i (n1555), .o (n1556) );
  buffer buf_n1557( .i (n1556), .o (n1557) );
  buffer buf_n1558( .i (n1557), .o (n1558) );
  buffer buf_n1559( .i (n1558), .o (n1559) );
  buffer buf_n1560( .i (n1559), .o (n1560) );
  buffer buf_n1561( .i (n1560), .o (n1561) );
  buffer buf_n1562( .i (n1561), .o (n1562) );
  buffer buf_n1563( .i (n1562), .o (n1563) );
  buffer buf_n1564( .i (n1563), .o (n1564) );
  buffer buf_n1565( .i (n1564), .o (n1565) );
  buffer buf_n1566( .i (n1565), .o (n1566) );
  buffer buf_n1567( .i (n1566), .o (n1567) );
  buffer buf_n1568( .i (n1567), .o (n1568) );
  buffer buf_n1569( .i (n1568), .o (n1569) );
  buffer buf_n1570( .i (n1569), .o (n1570) );
  buffer buf_n1571( .i (n1570), .o (n1571) );
  buffer buf_n1572( .i (n1571), .o (n1572) );
  buffer buf_n1573( .i (n1572), .o (n1573) );
  buffer buf_n1574( .i (n1573), .o (n1574) );
  buffer buf_n660( .i (x98), .o (n660) );
  buffer buf_n661( .i (n660), .o (n661) );
  buffer buf_n662( .i (n661), .o (n662) );
  buffer buf_n663( .i (n662), .o (n663) );
  buffer buf_n664( .i (n663), .o (n664) );
  buffer buf_n665( .i (n664), .o (n665) );
  buffer buf_n666( .i (n665), .o (n666) );
  buffer buf_n667( .i (n666), .o (n667) );
  buffer buf_n668( .i (n667), .o (n668) );
  buffer buf_n669( .i (n668), .o (n669) );
  buffer buf_n670( .i (n669), .o (n670) );
  buffer buf_n671( .i (n670), .o (n671) );
  buffer buf_n672( .i (n671), .o (n672) );
  buffer buf_n673( .i (n672), .o (n673) );
  buffer buf_n674( .i (n673), .o (n674) );
  buffer buf_n675( .i (n674), .o (n675) );
  buffer buf_n676( .i (n675), .o (n676) );
  buffer buf_n677( .i (n676), .o (n677) );
  buffer buf_n678( .i (n677), .o (n678) );
  buffer buf_n679( .i (n678), .o (n679) );
  buffer buf_n680( .i (n679), .o (n680) );
  buffer buf_n681( .i (n680), .o (n681) );
  buffer buf_n682( .i (n681), .o (n682) );
  buffer buf_n683( .i (n682), .o (n683) );
  buffer buf_n1235( .i (n1234), .o (n1235) );
  buffer buf_n1236( .i (n1235), .o (n1236) );
  buffer buf_n1237( .i (n1236), .o (n1237) );
  buffer buf_n1238( .i (n1237), .o (n1238) );
  buffer buf_n1239( .i (n1238), .o (n1239) );
  buffer buf_n1240( .i (n1239), .o (n1240) );
  buffer buf_n1241( .i (n1240), .o (n1241) );
  buffer buf_n1242( .i (n1241), .o (n1242) );
  buffer buf_n1243( .i (n1242), .o (n1243) );
  buffer buf_n1244( .i (n1243), .o (n1244) );
  buffer buf_n1245( .i (n1244), .o (n1245) );
  buffer buf_n1246( .i (n1245), .o (n1246) );
  buffer buf_n1247( .i (n1246), .o (n1247) );
  buffer buf_n1248( .i (n1247), .o (n1248) );
  buffer buf_n1249( .i (n1248), .o (n1249) );
  buffer buf_n1250( .i (n1249), .o (n1250) );
  buffer buf_n1251( .i (n1250), .o (n1251) );
  buffer buf_n1252( .i (n1251), .o (n1252) );
  buffer buf_n1286( .i (n1285), .o (n1286) );
  buffer buf_n1287( .i (n1286), .o (n1287) );
  buffer buf_n1288( .i (n1287), .o (n1288) );
  buffer buf_n1289( .i (n1288), .o (n1289) );
  buffer buf_n1290( .i (n1289), .o (n1290) );
  buffer buf_n1291( .i (n1290), .o (n1291) );
  buffer buf_n1292( .i (n1291), .o (n1292) );
  buffer buf_n1293( .i (n1292), .o (n1293) );
  buffer buf_n1294( .i (n1293), .o (n1294) );
  buffer buf_n1295( .i (n1294), .o (n1295) );
  buffer buf_n1296( .i (n1295), .o (n1296) );
  buffer buf_n1297( .i (n1296), .o (n1297) );
  buffer buf_n1298( .i (n1297), .o (n1298) );
  buffer buf_n1299( .i (n1298), .o (n1299) );
  buffer buf_n1300( .i (n1299), .o (n1300) );
  buffer buf_n1301( .i (n1300), .o (n1301) );
  buffer buf_n1302( .i (n1301), .o (n1302) );
  buffer buf_n1303( .i (n1302), .o (n1303) );
  buffer buf_n1255( .i (x154), .o (n1255) );
  buffer buf_n1256( .i (n1255), .o (n1256) );
  buffer buf_n1257( .i (n1256), .o (n1257) );
  buffer buf_n1258( .i (n1257), .o (n1258) );
  buffer buf_n1259( .i (n1258), .o (n1259) );
  buffer buf_n1260( .i (n1259), .o (n1260) );
  buffer buf_n1261( .i (n1260), .o (n1261) );
  buffer buf_n1262( .i (n1261), .o (n1262) );
  buffer buf_n1263( .i (n1262), .o (n1263) );
  buffer buf_n1264( .i (n1263), .o (n1264) );
  buffer buf_n1265( .i (n1264), .o (n1265) );
  buffer buf_n1266( .i (n1265), .o (n1266) );
  buffer buf_n1267( .i (n1266), .o (n1267) );
  buffer buf_n1268( .i (n1267), .o (n1268) );
  buffer buf_n1269( .i (n1268), .o (n1269) );
  buffer buf_n1270( .i (n1269), .o (n1270) );
  buffer buf_n1271( .i (n1270), .o (n1271) );
  buffer buf_n1272( .i (n1271), .o (n1272) );
  buffer buf_n1273( .i (n1272), .o (n1273) );
  buffer buf_n1274( .i (n1273), .o (n1274) );
  buffer buf_n1275( .i (n1274), .o (n1275) );
  buffer buf_n1276( .i (n1275), .o (n1276) );
  buffer buf_n1277( .i (n1276), .o (n1277) );
  buffer buf_n1278( .i (n1277), .o (n1278) );
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n992( .i (x133), .o (n992) );
  assign n1575 = n2 & n992 ;
  buffer buf_n1576( .i (n1575), .o (n1576) );
  buffer buf_n1577( .i (n1576), .o (n1577) );
  buffer buf_n1578( .i (n1577), .o (n1578) );
  buffer buf_n1579( .i (n1578), .o (n1579) );
  buffer buf_n1580( .i (n1579), .o (n1580) );
  buffer buf_n1581( .i (n1580), .o (n1581) );
  buffer buf_n1582( .i (n1581), .o (n1582) );
  buffer buf_n1583( .i (n1582), .o (n1583) );
  buffer buf_n1584( .i (n1583), .o (n1584) );
  buffer buf_n1585( .i (n1584), .o (n1585) );
  buffer buf_n1586( .i (n1585), .o (n1586) );
  buffer buf_n1587( .i (n1586), .o (n1587) );
  buffer buf_n1588( .i (n1587), .o (n1588) );
  buffer buf_n1589( .i (n1588), .o (n1589) );
  buffer buf_n1590( .i (n1589), .o (n1590) );
  buffer buf_n1591( .i (n1590), .o (n1591) );
  buffer buf_n1592( .i (n1591), .o (n1592) );
  buffer buf_n1593( .i (n1592), .o (n1593) );
  buffer buf_n1594( .i (n1593), .o (n1594) );
  buffer buf_n1595( .i (n1594), .o (n1595) );
  buffer buf_n1596( .i (n1595), .o (n1596) );
  buffer buf_n1597( .i (n1596), .o (n1597) );
  buffer buf_n453( .i (x62), .o (n453) );
  assign n1598 = n453 & ~n1349 ;
  buffer buf_n1599( .i (n1598), .o (n1599) );
  buffer buf_n1600( .i (n1599), .o (n1600) );
  buffer buf_n1601( .i (n1600), .o (n1601) );
  buffer buf_n1602( .i (n1601), .o (n1602) );
  buffer buf_n1603( .i (n1602), .o (n1603) );
  buffer buf_n1604( .i (n1603), .o (n1604) );
  buffer buf_n1605( .i (n1604), .o (n1605) );
  buffer buf_n1606( .i (n1605), .o (n1606) );
  buffer buf_n1607( .i (n1606), .o (n1607) );
  buffer buf_n1608( .i (n1607), .o (n1608) );
  buffer buf_n1609( .i (n1608), .o (n1609) );
  buffer buf_n1610( .i (n1609), .o (n1610) );
  buffer buf_n1611( .i (n1610), .o (n1611) );
  buffer buf_n1612( .i (n1611), .o (n1612) );
  buffer buf_n1613( .i (n1612), .o (n1613) );
  buffer buf_n1614( .i (n1613), .o (n1614) );
  buffer buf_n1615( .i (n1614), .o (n1615) );
  buffer buf_n1616( .i (n1615), .o (n1616) );
  buffer buf_n1617( .i (n1616), .o (n1617) );
  buffer buf_n1618( .i (n1617), .o (n1618) );
  buffer buf_n1619( .i (n1618), .o (n1619) );
  buffer buf_n1620( .i (n1619), .o (n1620) );
  buffer buf_n98( .i (x10), .o (n98) );
  buffer buf_n1347( .i (x163), .o (n1347) );
  assign n1621 = n98 & ~n1347 ;
  buffer buf_n1622( .i (n1621), .o (n1622) );
  buffer buf_n1623( .i (n1622), .o (n1623) );
  buffer buf_n1624( .i (n1623), .o (n1624) );
  buffer buf_n1625( .i (n1624), .o (n1625) );
  buffer buf_n1626( .i (n1625), .o (n1626) );
  buffer buf_n1627( .i (n1626), .o (n1627) );
  buffer buf_n1628( .i (n1627), .o (n1628) );
  buffer buf_n1629( .i (n1628), .o (n1629) );
  buffer buf_n1630( .i (n1629), .o (n1630) );
  buffer buf_n1631( .i (n1630), .o (n1631) );
  buffer buf_n1632( .i (n1631), .o (n1632) );
  buffer buf_n1633( .i (n1632), .o (n1633) );
  buffer buf_n1634( .i (n1633), .o (n1634) );
  buffer buf_n1635( .i (n1634), .o (n1635) );
  buffer buf_n1636( .i (n1635), .o (n1636) );
  buffer buf_n1637( .i (n1636), .o (n1637) );
  buffer buf_n1638( .i (n1637), .o (n1638) );
  buffer buf_n1639( .i (n1638), .o (n1639) );
  buffer buf_n1640( .i (n1639), .o (n1640) );
  buffer buf_n1641( .i (n1640), .o (n1641) );
  buffer buf_n1642( .i (n1641), .o (n1642) );
  buffer buf_n1643( .i (n1642), .o (n1643) );
  assign n1644 = x135 & x153 ;
  buffer buf_n1645( .i (n1644), .o (n1645) );
  buffer buf_n1646( .i (n1645), .o (n1646) );
  buffer buf_n1647( .i (n1646), .o (n1647) );
  buffer buf_n1648( .i (n1647), .o (n1648) );
  buffer buf_n1649( .i (n1648), .o (n1649) );
  buffer buf_n1650( .i (n1649), .o (n1650) );
  buffer buf_n1651( .i (n1650), .o (n1651) );
  buffer buf_n1652( .i (n1651), .o (n1652) );
  buffer buf_n1653( .i (n1652), .o (n1653) );
  buffer buf_n1654( .i (n1653), .o (n1654) );
  buffer buf_n1655( .i (n1654), .o (n1655) );
  buffer buf_n1656( .i (n1655), .o (n1656) );
  buffer buf_n1657( .i (n1656), .o (n1657) );
  buffer buf_n1658( .i (n1657), .o (n1658) );
  buffer buf_n1659( .i (n1658), .o (n1659) );
  buffer buf_n1660( .i (n1659), .o (n1660) );
  buffer buf_n1661( .i (n1660), .o (n1661) );
  buffer buf_n1662( .i (n1661), .o (n1662) );
  buffer buf_n1663( .i (n1662), .o (n1663) );
  buffer buf_n1664( .i (n1663), .o (n1664) );
  buffer buf_n1665( .i (n1664), .o (n1665) );
  buffer buf_n1666( .i (n1665), .o (n1666) );
  buffer buf_n1667( .i (n1666), .o (n1667) );
  buffer buf_n455( .i (x63), .o (n455) );
  buffer buf_n456( .i (n455), .o (n456) );
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n458( .i (n457), .o (n458) );
  buffer buf_n459( .i (n458), .o (n459) );
  buffer buf_n460( .i (n459), .o (n460) );
  buffer buf_n461( .i (n460), .o (n461) );
  buffer buf_n462( .i (n461), .o (n462) );
  buffer buf_n463( .i (n462), .o (n463) );
  buffer buf_n464( .i (n463), .o (n464) );
  buffer buf_n465( .i (n464), .o (n465) );
  buffer buf_n466( .i (n465), .o (n466) );
  buffer buf_n467( .i (n466), .o (n467) );
  buffer buf_n468( .i (n467), .o (n468) );
  buffer buf_n469( .i (n468), .o (n469) );
  buffer buf_n470( .i (n469), .o (n470) );
  buffer buf_n471( .i (n470), .o (n471) );
  buffer buf_n472( .i (n471), .o (n472) );
  buffer buf_n473( .i (n472), .o (n473) );
  buffer buf_n474( .i (n473), .o (n474) );
  buffer buf_n475( .i (n474), .o (n475) );
  buffer buf_n476( .i (n475), .o (n476) );
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n10( .i (n9), .o (n10) );
  buffer buf_n11( .i (n10), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n18( .i (n17), .o (n18) );
  buffer buf_n19( .i (n18), .o (n19) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  buffer buf_n774( .i (x113), .o (n774) );
  buffer buf_n775( .i (n774), .o (n775) );
  buffer buf_n776( .i (n775), .o (n776) );
  buffer buf_n777( .i (n776), .o (n777) );
  buffer buf_n778( .i (n777), .o (n778) );
  buffer buf_n779( .i (n778), .o (n779) );
  buffer buf_n780( .i (n779), .o (n780) );
  buffer buf_n781( .i (n780), .o (n781) );
  buffer buf_n782( .i (n781), .o (n782) );
  buffer buf_n783( .i (n782), .o (n783) );
  buffer buf_n784( .i (n783), .o (n784) );
  buffer buf_n785( .i (n784), .o (n785) );
  buffer buf_n786( .i (n785), .o (n786) );
  buffer buf_n787( .i (n786), .o (n787) );
  buffer buf_n788( .i (n787), .o (n788) );
  buffer buf_n789( .i (n788), .o (n789) );
  buffer buf_n790( .i (n789), .o (n790) );
  buffer buf_n791( .i (n790), .o (n791) );
  buffer buf_n792( .i (n791), .o (n792) );
  buffer buf_n793( .i (n792), .o (n793) );
  buffer buf_n794( .i (n793), .o (n794) );
  buffer buf_n795( .i (n794), .o (n795) );
  buffer buf_n796( .i (n795), .o (n796) );
  buffer buf_n797( .i (n796), .o (n797) );
  buffer buf_n480( .i (x64), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n100( .i (x11), .o (n100) );
  assign n1668 = n98 & n100 ;
  buffer buf_n1669( .i (n1668), .o (n1669) );
  buffer buf_n1670( .i (n1669), .o (n1670) );
  buffer buf_n1671( .i (n1670), .o (n1671) );
  assign n1691 = n484 & n1671 ;
  buffer buf_n1692( .i (n1691), .o (n1692) );
  buffer buf_n1693( .i (n1692), .o (n1693) );
  buffer buf_n1694( .i (n1693), .o (n1694) );
  buffer buf_n1695( .i (n1694), .o (n1695) );
  buffer buf_n1696( .i (n1695), .o (n1696) );
  buffer buf_n1697( .i (n1696), .o (n1697) );
  buffer buf_n1698( .i (n1697), .o (n1698) );
  buffer buf_n1699( .i (n1698), .o (n1699) );
  buffer buf_n1700( .i (n1699), .o (n1700) );
  buffer buf_n1701( .i (n1700), .o (n1701) );
  buffer buf_n1702( .i (n1701), .o (n1702) );
  buffer buf_n1703( .i (n1702), .o (n1703) );
  buffer buf_n1704( .i (n1703), .o (n1704) );
  buffer buf_n1705( .i (n1704), .o (n1705) );
  buffer buf_n1706( .i (n1705), .o (n1706) );
  buffer buf_n1707( .i (n1706), .o (n1707) );
  buffer buf_n1708( .i (n1707), .o (n1708) );
  buffer buf_n1709( .i (n1708), .o (n1709) );
  buffer buf_n1672( .i (n1671), .o (n1672) );
  buffer buf_n1673( .i (n1672), .o (n1673) );
  buffer buf_n1674( .i (n1673), .o (n1674) );
  buffer buf_n1675( .i (n1674), .o (n1675) );
  buffer buf_n1676( .i (n1675), .o (n1676) );
  buffer buf_n1677( .i (n1676), .o (n1677) );
  buffer buf_n1678( .i (n1677), .o (n1678) );
  buffer buf_n1679( .i (n1678), .o (n1679) );
  buffer buf_n1680( .i (n1679), .o (n1680) );
  buffer buf_n1681( .i (n1680), .o (n1681) );
  buffer buf_n1682( .i (n1681), .o (n1682) );
  buffer buf_n1683( .i (n1682), .o (n1683) );
  buffer buf_n1684( .i (n1683), .o (n1684) );
  buffer buf_n1685( .i (n1684), .o (n1685) );
  buffer buf_n1686( .i (n1685), .o (n1686) );
  buffer buf_n1687( .i (n1686), .o (n1687) );
  buffer buf_n1688( .i (n1687), .o (n1688) );
  buffer buf_n1689( .i (n1688), .o (n1689) );
  buffer buf_n1690( .i (n1689), .o (n1690) );
  buffer buf_n4913( .i (n24), .o (n4913) );
  buffer buf_n246( .i (x33), .o (n246) );
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  buffer buf_n1343( .i (x162), .o (n1343) );
  buffer buf_n1344( .i (n1343), .o (n1344) );
  buffer buf_n1345( .i (n1344), .o (n1345) );
  assign n1710 = n248 & n1345 ;
  buffer buf_n242( .i (x32), .o (n242) );
  buffer buf_n243( .i (n242), .o (n243) );
  buffer buf_n244( .i (n243), .o (n244) );
  assign n1711 = n244 & ~n1345 ;
  assign n1712 = ( n1670 & n1710 ) | ( n1670 & n1711 ) | ( n1710 & n1711 ) ;
  buffer buf_n1713( .i (n1712), .o (n1713) );
  buffer buf_n1714( .i (n1713), .o (n1714) );
  buffer buf_n1715( .i (n1714), .o (n1715) );
  buffer buf_n1716( .i (n1715), .o (n1716) );
  buffer buf_n1717( .i (n1716), .o (n1717) );
  buffer buf_n1718( .i (n1717), .o (n1718) );
  buffer buf_n1719( .i (n1718), .o (n1719) );
  buffer buf_n1720( .i (n1719), .o (n1720) );
  buffer buf_n1721( .i (n1720), .o (n1721) );
  buffer buf_n1722( .i (n1721), .o (n1722) );
  buffer buf_n1723( .i (n1722), .o (n1723) );
  buffer buf_n1724( .i (n1723), .o (n1724) );
  buffer buf_n1725( .i (n1724), .o (n1725) );
  buffer buf_n1726( .i (n1725), .o (n1726) );
  buffer buf_n1727( .i (n1726), .o (n1727) );
  buffer buf_n1728( .i (n1727), .o (n1728) );
  buffer buf_n1729( .i (n1728), .o (n1729) );
  buffer buf_n1730( .i (n1729), .o (n1730) );
  buffer buf_n1731( .i (n1730), .o (n1731) );
  buffer buf_n102( .i (x12), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  assign n1732 = n103 & n1344 ;
  buffer buf_n1733( .i (n1732), .o (n1733) );
  buffer buf_n250( .i (x34), .o (n250) );
  buffer buf_n251( .i (n250), .o (n251) );
  assign n1734 = n251 & ~n1344 ;
  buffer buf_n1735( .i (n1734), .o (n1735) );
  assign n1736 = ( n1670 & n1733 ) | ( n1670 & n1735 ) | ( n1733 & n1735 ) ;
  buffer buf_n1737( .i (n1736), .o (n1737) );
  buffer buf_n1738( .i (n1737), .o (n1738) );
  buffer buf_n1739( .i (n1738), .o (n1739) );
  buffer buf_n1740( .i (n1739), .o (n1740) );
  buffer buf_n1741( .i (n1740), .o (n1741) );
  buffer buf_n1742( .i (n1741), .o (n1742) );
  buffer buf_n1743( .i (n1742), .o (n1743) );
  buffer buf_n1744( .i (n1743), .o (n1744) );
  buffer buf_n1745( .i (n1744), .o (n1745) );
  buffer buf_n1746( .i (n1745), .o (n1746) );
  buffer buf_n1747( .i (n1746), .o (n1747) );
  buffer buf_n1748( .i (n1747), .o (n1748) );
  buffer buf_n1749( .i (n1748), .o (n1749) );
  buffer buf_n1750( .i (n1749), .o (n1750) );
  buffer buf_n1751( .i (n1750), .o (n1751) );
  buffer buf_n1752( .i (n1751), .o (n1752) );
  buffer buf_n1753( .i (n1752), .o (n1753) );
  buffer buf_n1754( .i (n1753), .o (n1754) );
  buffer buf_n1755( .i (n1754), .o (n1755) );
  buffer buf_n236( .i (x31), .o (n236) );
  buffer buf_n237( .i (n236), .o (n237) );
  buffer buf_n238( .i (n237), .o (n238) );
  buffer buf_n239( .i (n238), .o (n239) );
  buffer buf_n240( .i (n239), .o (n240) );
  assign n1756 = n240 & n1671 ;
  buffer buf_n1757( .i (n1756), .o (n1757) );
  buffer buf_n1758( .i (n1757), .o (n1758) );
  buffer buf_n1759( .i (n1758), .o (n1759) );
  buffer buf_n1760( .i (n1759), .o (n1760) );
  buffer buf_n1761( .i (n1760), .o (n1761) );
  buffer buf_n1762( .i (n1761), .o (n1762) );
  buffer buf_n1763( .i (n1762), .o (n1763) );
  buffer buf_n1764( .i (n1763), .o (n1764) );
  buffer buf_n1765( .i (n1764), .o (n1765) );
  buffer buf_n1766( .i (n1765), .o (n1766) );
  buffer buf_n1767( .i (n1766), .o (n1767) );
  buffer buf_n1768( .i (n1767), .o (n1768) );
  buffer buf_n1769( .i (n1768), .o (n1769) );
  buffer buf_n1770( .i (n1769), .o (n1770) );
  buffer buf_n1771( .i (n1770), .o (n1771) );
  buffer buf_n1772( .i (n1771), .o (n1772) );
  buffer buf_n1773( .i (n1772), .o (n1773) );
  buffer buf_n1774( .i (n1773), .o (n1774) );
  buffer buf_n92( .i (x8), .o (n92) );
  buffer buf_n93( .i (n92), .o (n93) );
  assign n1775 = ~n93 & n1344 ;
  buffer buf_n89( .i (x7), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  buffer buf_n1776( .i (n1343), .o (n1776) );
  assign n1777 = n90 | n1776 ;
  assign n1778 = ( n1669 & n1775 ) | ( n1669 & ~n1777 ) | ( n1775 & ~n1777 ) ;
  assign n1779 = n489 & ~n1778 ;
  buffer buf_n1780( .i (n1779), .o (n1780) );
  buffer buf_n1781( .i (n1780), .o (n1781) );
  buffer buf_n1782( .i (n1781), .o (n1782) );
  buffer buf_n1783( .i (n1782), .o (n1783) );
  buffer buf_n1784( .i (n1783), .o (n1784) );
  buffer buf_n1785( .i (n1784), .o (n1785) );
  buffer buf_n1786( .i (n1785), .o (n1786) );
  buffer buf_n1787( .i (n1786), .o (n1787) );
  buffer buf_n1788( .i (n1787), .o (n1788) );
  buffer buf_n1789( .i (n1788), .o (n1789) );
  buffer buf_n1790( .i (n1789), .o (n1790) );
  buffer buf_n1791( .i (n1790), .o (n1791) );
  buffer buf_n1792( .i (n1791), .o (n1792) );
  buffer buf_n1793( .i (n1792), .o (n1793) );
  buffer buf_n1794( .i (n1793), .o (n1794) );
  buffer buf_n1795( .i (n1794), .o (n1795) );
  buffer buf_n1796( .i (n1795), .o (n1796) );
  buffer buf_n1797( .i (n1796), .o (n1797) );
  buffer buf_n1798( .i (n1797), .o (n1798) );
  buffer buf_n230( .i (x29), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  assign n1799 = ~n231 & n1776 ;
  buffer buf_n95( .i (x9), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  assign n1800 = n96 | n1776 ;
  assign n1801 = ( n1669 & n1799 ) | ( n1669 & ~n1800 ) | ( n1799 & ~n1800 ) ;
  assign n1802 = n489 & ~n1801 ;
  buffer buf_n1803( .i (n1802), .o (n1803) );
  buffer buf_n1804( .i (n1803), .o (n1804) );
  buffer buf_n1805( .i (n1804), .o (n1805) );
  buffer buf_n1806( .i (n1805), .o (n1806) );
  buffer buf_n1807( .i (n1806), .o (n1807) );
  buffer buf_n1808( .i (n1807), .o (n1808) );
  buffer buf_n1809( .i (n1808), .o (n1809) );
  buffer buf_n1810( .i (n1809), .o (n1810) );
  buffer buf_n1811( .i (n1810), .o (n1811) );
  buffer buf_n1812( .i (n1811), .o (n1812) );
  buffer buf_n1813( .i (n1812), .o (n1813) );
  buffer buf_n1814( .i (n1813), .o (n1814) );
  buffer buf_n1815( .i (n1814), .o (n1815) );
  buffer buf_n1816( .i (n1815), .o (n1816) );
  buffer buf_n1817( .i (n1816), .o (n1817) );
  buffer buf_n1818( .i (n1817), .o (n1818) );
  buffer buf_n1819( .i (n1818), .o (n1819) );
  buffer buf_n1820( .i (n1819), .o (n1820) );
  buffer buf_n1821( .i (n1820), .o (n1821) );
  buffer buf_n86( .i (x6), .o (n86) );
  buffer buf_n87( .i (n86), .o (n87) );
  assign n1822 = ~n87 & n1776 ;
  buffer buf_n1823( .i (n1822), .o (n1823) );
  buffer buf_n224( .i (x27), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n1824( .i (n1343), .o (n1824) );
  assign n1825 = n225 | n1824 ;
  buffer buf_n1826( .i (n1825), .o (n1826) );
  assign n1827 = ( n1670 & n1823 ) | ( n1670 & ~n1826 ) | ( n1823 & ~n1826 ) ;
  assign n1828 = n490 & ~n1827 ;
  buffer buf_n1829( .i (n1828), .o (n1829) );
  buffer buf_n1830( .i (n1829), .o (n1830) );
  buffer buf_n1831( .i (n1830), .o (n1831) );
  buffer buf_n1832( .i (n1831), .o (n1832) );
  buffer buf_n1833( .i (n1832), .o (n1833) );
  buffer buf_n1834( .i (n1833), .o (n1834) );
  buffer buf_n1835( .i (n1834), .o (n1835) );
  buffer buf_n1836( .i (n1835), .o (n1836) );
  buffer buf_n1837( .i (n1836), .o (n1837) );
  buffer buf_n1838( .i (n1837), .o (n1838) );
  buffer buf_n1839( .i (n1838), .o (n1839) );
  buffer buf_n1840( .i (n1839), .o (n1840) );
  buffer buf_n1841( .i (n1840), .o (n1841) );
  buffer buf_n1842( .i (n1841), .o (n1842) );
  buffer buf_n1843( .i (n1842), .o (n1843) );
  buffer buf_n1844( .i (n1843), .o (n1844) );
  buffer buf_n1845( .i (n1844), .o (n1845) );
  buffer buf_n1846( .i (n1845), .o (n1846) );
  buffer buf_n227( .i (x28), .o (n227) );
  buffer buf_n228( .i (n227), .o (n228) );
  assign n1847 = ~n228 & n1824 ;
  buffer buf_n1848( .i (n1847), .o (n1848) );
  buffer buf_n233( .i (x30), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  assign n1849 = n234 | n1824 ;
  buffer buf_n1850( .i (n1849), .o (n1850) );
  buffer buf_n1851( .i (n1669), .o (n1851) );
  assign n1852 = ( n1848 & ~n1850 ) | ( n1848 & n1851 ) | ( ~n1850 & n1851 ) ;
  assign n1853 = n490 & ~n1852 ;
  buffer buf_n1854( .i (n1853), .o (n1854) );
  buffer buf_n1855( .i (n1854), .o (n1855) );
  buffer buf_n1856( .i (n1855), .o (n1856) );
  buffer buf_n1857( .i (n1856), .o (n1857) );
  buffer buf_n1858( .i (n1857), .o (n1858) );
  buffer buf_n1859( .i (n1858), .o (n1859) );
  buffer buf_n1860( .i (n1859), .o (n1860) );
  buffer buf_n1861( .i (n1860), .o (n1861) );
  buffer buf_n1862( .i (n1861), .o (n1862) );
  buffer buf_n1863( .i (n1862), .o (n1863) );
  buffer buf_n1864( .i (n1863), .o (n1864) );
  buffer buf_n1865( .i (n1864), .o (n1865) );
  buffer buf_n1866( .i (n1865), .o (n1866) );
  buffer buf_n1867( .i (n1866), .o (n1867) );
  buffer buf_n1868( .i (n1867), .o (n1868) );
  buffer buf_n1869( .i (n1868), .o (n1869) );
  buffer buf_n1870( .i (n1869), .o (n1870) );
  buffer buf_n1871( .i (n1870), .o (n1871) );
  buffer buf_n811( .i (x116), .o (n811) );
  buffer buf_n812( .i (n811), .o (n812) );
  buffer buf_n813( .i (n812), .o (n813) );
  buffer buf_n814( .i (n813), .o (n814) );
  buffer buf_n654( .i (x97), .o (n654) );
  buffer buf_n655( .i (n654), .o (n655) );
  buffer buf_n656( .i (n655), .o (n656) );
  buffer buf_n1096( .i (x144), .o (n1096) );
  buffer buf_n1097( .i (n1096), .o (n1097) );
  buffer buf_n1098( .i (n1097), .o (n1098) );
  assign n1872 = n656 | n1098 ;
  buffer buf_n685( .i (x99), .o (n685) );
  buffer buf_n686( .i (n685), .o (n686) );
  buffer buf_n687( .i (n686), .o (n687) );
  assign n1873 = n687 & n1098 ;
  assign n1874 = ( n814 & ~n1872 ) | ( n814 & n1873 ) | ( ~n1872 & n1873 ) ;
  buffer buf_n698( .i (x101), .o (n698) );
  buffer buf_n699( .i (n698), .o (n699) );
  buffer buf_n700( .i (n699), .o (n700) );
  assign n1875 = n700 | n1098 ;
  buffer buf_n692( .i (x100), .o (n692) );
  buffer buf_n693( .i (n692), .o (n693) );
  buffer buf_n694( .i (n693), .o (n694) );
  buffer buf_n1876( .i (n1097), .o (n1876) );
  assign n1877 = n694 & n1876 ;
  assign n1878 = ( n814 & n1875 ) | ( n814 & ~n1877 ) | ( n1875 & ~n1877 ) ;
  assign n1879 = ~n1874 & n1878 ;
  buffer buf_n1880( .i (n1879), .o (n1880) );
  buffer buf_n1881( .i (n1880), .o (n1881) );
  buffer buf_n1882( .i (n1881), .o (n1882) );
  buffer buf_n823( .i (x118), .o (n823) );
  buffer buf_n824( .i (n823), .o (n824) );
  buffer buf_n825( .i (n824), .o (n825) );
  buffer buf_n826( .i (n825), .o (n826) );
  buffer buf_n1110( .i (x145), .o (n1110) );
  buffer buf_n1111( .i (n1110), .o (n1111) );
  buffer buf_n1112( .i (n1111), .o (n1112) );
  assign n1883 = n656 | n1112 ;
  assign n1884 = n687 & n1112 ;
  assign n1885 = ( n826 & ~n1883 ) | ( n826 & n1884 ) | ( ~n1883 & n1884 ) ;
  assign n1886 = n700 | n1112 ;
  buffer buf_n1887( .i (n1111), .o (n1887) );
  assign n1888 = n694 & n1887 ;
  assign n1889 = ( n826 & n1886 ) | ( n826 & ~n1888 ) | ( n1886 & ~n1888 ) ;
  assign n1890 = ~n1885 & n1889 ;
  buffer buf_n1891( .i (n1890), .o (n1891) );
  buffer buf_n1892( .i (n1891), .o (n1892) );
  buffer buf_n1893( .i (n1892), .o (n1893) );
  assign n1894 = n1882 | n1893 ;
  buffer buf_n834( .i (x120), .o (n834) );
  buffer buf_n835( .i (n834), .o (n835) );
  buffer buf_n836( .i (n835), .o (n836) );
  buffer buf_n837( .i (n836), .o (n837) );
  buffer buf_n838( .i (n837), .o (n838) );
  buffer buf_n1126( .i (x146), .o (n1126) );
  buffer buf_n1127( .i (n1126), .o (n1127) );
  buffer buf_n1128( .i (n1127), .o (n1128) );
  buffer buf_n1129( .i (n1128), .o (n1129) );
  buffer buf_n1392( .i (x168), .o (n1392) );
  buffer buf_n1393( .i (n1392), .o (n1393) );
  buffer buf_n1394( .i (n1393), .o (n1394) );
  buffer buf_n1395( .i (n1394), .o (n1395) );
  assign n1895 = n1129 & n1395 ;
  buffer buf_n1374( .i (x165), .o (n1374) );
  buffer buf_n1375( .i (n1374), .o (n1375) );
  buffer buf_n1376( .i (n1375), .o (n1376) );
  buffer buf_n1377( .i (n1376), .o (n1377) );
  assign n1896 = n1129 | n1377 ;
  assign n1897 = ( n838 & n1895 ) | ( n838 & ~n1896 ) | ( n1895 & ~n1896 ) ;
  buffer buf_n1386( .i (x167), .o (n1386) );
  buffer buf_n1387( .i (n1386), .o (n1387) );
  buffer buf_n1388( .i (n1387), .o (n1388) );
  buffer buf_n1389( .i (n1388), .o (n1389) );
  assign n1898 = n1129 & n1389 ;
  buffer buf_n1380( .i (x166), .o (n1380) );
  buffer buf_n1381( .i (n1380), .o (n1381) );
  buffer buf_n1382( .i (n1381), .o (n1382) );
  buffer buf_n1383( .i (n1382), .o (n1383) );
  buffer buf_n1899( .i (n1128), .o (n1899) );
  assign n1900 = n1383 | n1899 ;
  assign n1901 = ( n838 & ~n1898 ) | ( n838 & n1900 ) | ( ~n1898 & n1900 ) ;
  assign n1902 = ~n1897 & n1901 ;
  buffer buf_n1903( .i (n1902), .o (n1903) );
  buffer buf_n1140( .i (x147), .o (n1140) );
  buffer buf_n1141( .i (n1140), .o (n1141) );
  buffer buf_n1142( .i (n1141), .o (n1142) );
  assign n1904 = ~n1142 & n1376 ;
  assign n1905 = n1142 & ~n1394 ;
  assign n1906 = n1904 | n1905 ;
  buffer buf_n1907( .i (n1906), .o (n1907) );
  buffer buf_n799( .i (x114), .o (n799) );
  buffer buf_n800( .i (n799), .o (n800) );
  buffer buf_n801( .i (n800), .o (n801) );
  assign n1908 = ~n687 & n801 ;
  assign n1909 = n694 | n801 ;
  assign n1910 = ~n1908 & n1909 ;
  buffer buf_n1911( .i (n1910), .o (n1911) );
  assign n1912 = n1907 & n1911 ;
  buffer buf_n947( .i (x129), .o (n947) );
  buffer buf_n948( .i (n947), .o (n948) );
  buffer buf_n949( .i (n948), .o (n949) );
  buffer buf_n1913( .i (n686), .o (n1913) );
  assign n1914 = n949 & ~n1913 ;
  buffer buf_n1915( .i (n693), .o (n1915) );
  assign n1916 = n949 | n1915 ;
  assign n1917 = ~n1914 & n1916 ;
  buffer buf_n1918( .i (n1917), .o (n1918) );
  assign n1919 = n656 & n751 ;
  assign n1920 = n700 & ~n751 ;
  assign n1921 = n1919 | n1920 ;
  buffer buf_n1922( .i (n1921), .o (n1922) );
  assign n1925 = n1918 & ~n1922 ;
  assign n1926 = n1912 & n1925 ;
  assign n1927 = n1903 & n1926 ;
  buffer buf_n886( .i (x125), .o (n886) );
  buffer buf_n887( .i (n886), .o (n887) );
  buffer buf_n888( .i (n887), .o (n888) );
  buffer buf_n889( .i (n888), .o (n889) );
  buffer buf_n890( .i (n889), .o (n890) );
  buffer buf_n1152( .i (x148), .o (n1152) );
  buffer buf_n1153( .i (n1152), .o (n1153) );
  buffer buf_n1154( .i (n1153), .o (n1154) );
  buffer buf_n1155( .i (n1154), .o (n1155) );
  assign n1928 = n1155 & n1395 ;
  assign n1929 = n1155 | n1377 ;
  assign n1930 = ( n890 & n1928 ) | ( n890 & ~n1929 ) | ( n1928 & ~n1929 ) ;
  assign n1931 = n1155 & n1389 ;
  buffer buf_n1932( .i (n1154), .o (n1932) );
  assign n1933 = n1383 | n1932 ;
  assign n1934 = ( n890 & ~n1931 ) | ( n890 & n1933 ) | ( ~n1931 & n1933 ) ;
  assign n1935 = ~n1930 & n1934 ;
  buffer buf_n1936( .i (n1935), .o (n1936) );
  buffer buf_n1162( .i (x149), .o (n1162) );
  buffer buf_n1163( .i (n1162), .o (n1163) );
  buffer buf_n1164( .i (n1163), .o (n1164) );
  buffer buf_n1165( .i (n1164), .o (n1165) );
  buffer buf_n1166( .i (n1165), .o (n1166) );
  buffer buf_n917( .i (x127), .o (n917) );
  buffer buf_n918( .i (n917), .o (n918) );
  buffer buf_n919( .i (n918), .o (n919) );
  buffer buf_n920( .i (n919), .o (n920) );
  assign n1937 = n920 & ~n1395 ;
  assign n1938 = n920 | n1389 ;
  assign n1939 = ( n1166 & n1937 ) | ( n1166 & ~n1938 ) | ( n1937 & ~n1938 ) ;
  assign n1940 = ~n920 & n1383 ;
  assign n1941 = n920 & n1377 ;
  assign n1942 = ( ~n1166 & n1940 ) | ( ~n1166 & n1941 ) | ( n1940 & n1941 ) ;
  assign n1943 = n1939 | n1942 ;
  buffer buf_n1944( .i (n1943), .o (n1944) );
  assign n1945 = n1936 & n1944 ;
  assign n1946 = n1927 & n1945 ;
  assign n1947 = ~n1894 & n1946 ;
  buffer buf_n1948( .i (n1947), .o (n1948) );
  buffer buf_n1949( .i (n1948), .o (n1949) );
  buffer buf_n1950( .i (n1949), .o (n1950) );
  buffer buf_n1951( .i (n1950), .o (n1951) );
  buffer buf_n1952( .i (n1951), .o (n1952) );
  buffer buf_n1953( .i (n1952), .o (n1953) );
  buffer buf_n1954( .i (n1953), .o (n1954) );
  buffer buf_n1955( .i (n1954), .o (n1955) );
  buffer buf_n1956( .i (n1955), .o (n1956) );
  buffer buf_n1957( .i (n1956), .o (n1957) );
  buffer buf_n1958( .i (n1957), .o (n1958) );
  buffer buf_n1959( .i (n1958), .o (n1959) );
  buffer buf_n1960( .i (n1959), .o (n1960) );
  buffer buf_n722( .i (x106), .o (n722) );
  buffer buf_n723( .i (n722), .o (n723) );
  buffer buf_n724( .i (n723), .o (n724) );
  buffer buf_n725( .i (n724), .o (n725) );
  buffer buf_n726( .i (n725), .o (n726) );
  buffer buf_n727( .i (n726), .o (n727) );
  buffer buf_n1028( .i (x138), .o (n1028) );
  buffer buf_n1029( .i (n1028), .o (n1029) );
  buffer buf_n1030( .i (n1029), .o (n1030) );
  buffer buf_n1031( .i (n1030), .o (n1031) );
  buffer buf_n1032( .i (n1031), .o (n1032) );
  buffer buf_n1396( .i (n1395), .o (n1396) );
  assign n1961 = n1032 & n1396 ;
  buffer buf_n1378( .i (n1377), .o (n1378) );
  assign n1962 = n1032 | n1378 ;
  assign n1963 = ( n727 & n1961 ) | ( n727 & ~n1962 ) | ( n1961 & ~n1962 ) ;
  buffer buf_n1390( .i (n1389), .o (n1390) );
  assign n1964 = n1032 & n1390 ;
  buffer buf_n1384( .i (n1383), .o (n1384) );
  buffer buf_n1965( .i (n1031), .o (n1965) );
  assign n1966 = n1384 | n1965 ;
  assign n1967 = ( n727 & ~n1964 ) | ( n727 & n1966 ) | ( ~n1964 & n1966 ) ;
  assign n1968 = ~n1963 & n1967 ;
  buffer buf_n1969( .i (n1968), .o (n1969) );
  buffer buf_n1088( .i (x143), .o (n1088) );
  buffer buf_n1089( .i (n1088), .o (n1089) );
  buffer buf_n1090( .i (n1089), .o (n1090) );
  buffer buf_n1091( .i (n1090), .o (n1091) );
  buffer buf_n1092( .i (n1091), .o (n1092) );
  buffer buf_n627( .i (x91), .o (n627) );
  buffer buf_n628( .i (n627), .o (n628) );
  buffer buf_n629( .i (n628), .o (n629) );
  buffer buf_n630( .i (n629), .o (n630) );
  buffer buf_n1970( .i (n1394), .o (n1970) );
  assign n1971 = n630 & n1970 ;
  buffer buf_n1972( .i (n1388), .o (n1972) );
  assign n1973 = ~n630 & n1972 ;
  assign n1974 = ( n1092 & n1971 ) | ( n1092 & n1973 ) | ( n1971 & n1973 ) ;
  buffer buf_n1975( .i (n1382), .o (n1975) );
  assign n1976 = n630 | n1975 ;
  buffer buf_n1977( .i (n629), .o (n1977) );
  buffer buf_n1978( .i (n1376), .o (n1978) );
  assign n1979 = n1977 & ~n1978 ;
  assign n1980 = ( n1092 & n1976 ) | ( n1092 & ~n1979 ) | ( n1976 & ~n1979 ) ;
  assign n1981 = ~n1974 & n1980 ;
  buffer buf_n1982( .i (n1981), .o (n1982) );
  buffer buf_n1018( .i (x137), .o (n1018) );
  buffer buf_n1019( .i (n1018), .o (n1019) );
  buffer buf_n1020( .i (n1019), .o (n1020) );
  buffer buf_n1021( .i (n1020), .o (n1021) );
  buffer buf_n1022( .i (n1021), .o (n1022) );
  buffer buf_n714( .i (x104), .o (n714) );
  buffer buf_n715( .i (n714), .o (n715) );
  buffer buf_n716( .i (n715), .o (n716) );
  buffer buf_n717( .i (n716), .o (n717) );
  assign n1983 = n717 & ~n1970 ;
  assign n1984 = n717 | n1972 ;
  assign n1985 = ( n1022 & n1983 ) | ( n1022 & ~n1984 ) | ( n1983 & ~n1984 ) ;
  assign n1986 = ~n717 & n1975 ;
  assign n1987 = n717 & n1978 ;
  assign n1988 = ( ~n1022 & n1986 ) | ( ~n1022 & n1987 ) | ( n1986 & n1987 ) ;
  assign n1989 = n1985 | n1988 ;
  buffer buf_n1990( .i (n1989), .o (n1990) );
  assign n1991 = n1982 & n1990 ;
  assign n1992 = n1969 & n1991 ;
  buffer buf_n1993( .i (n1992), .o (n1993) );
  buffer buf_n1054( .i (x140), .o (n1054) );
  buffer buf_n1055( .i (n1054), .o (n1055) );
  buffer buf_n1056( .i (n1055), .o (n1056) );
  buffer buf_n1057( .i (n1056), .o (n1057) );
  buffer buf_n1058( .i (n1057), .o (n1058) );
  buffer buf_n645( .i (x95), .o (n645) );
  buffer buf_n646( .i (n645), .o (n646) );
  buffer buf_n647( .i (n646), .o (n647) );
  buffer buf_n648( .i (n647), .o (n648) );
  assign n1994 = n648 & ~n1970 ;
  assign n1995 = n648 | n1972 ;
  assign n1996 = ( n1058 & n1994 ) | ( n1058 & ~n1995 ) | ( n1994 & ~n1995 ) ;
  assign n1997 = ~n648 & n1975 ;
  buffer buf_n1998( .i (n647), .o (n1998) );
  assign n1999 = n1978 & n1998 ;
  assign n2000 = ( ~n1058 & n1997 ) | ( ~n1058 & n1999 ) | ( n1997 & n1999 ) ;
  assign n2001 = n1996 | n2000 ;
  buffer buf_n2002( .i (n2001), .o (n2002) );
  buffer buf_n1080( .i (x142), .o (n1080) );
  buffer buf_n1081( .i (n1080), .o (n1081) );
  buffer buf_n1082( .i (n1081), .o (n1082) );
  buffer buf_n1083( .i (n1082), .o (n1083) );
  buffer buf_n1084( .i (n1083), .o (n1084) );
  buffer buf_n618( .i (x89), .o (n618) );
  buffer buf_n619( .i (n618), .o (n619) );
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  assign n2003 = n621 & ~n1970 ;
  assign n2004 = n621 | n1972 ;
  assign n2005 = ( n1084 & n2003 ) | ( n1084 & ~n2004 ) | ( n2003 & ~n2004 ) ;
  assign n2006 = ~n621 & n1975 ;
  assign n2007 = n621 & n1978 ;
  assign n2008 = ( ~n1084 & n2006 ) | ( ~n1084 & n2007 ) | ( n2006 & n2007 ) ;
  assign n2009 = n2005 | n2008 ;
  buffer buf_n2010( .i (n2009), .o (n2010) );
  assign n2011 = n2002 & n2010 ;
  buffer buf_n2012( .i (n2011), .o (n2012) );
  buffer buf_n1062( .i (x141), .o (n1062) );
  buffer buf_n1063( .i (n1062), .o (n1063) );
  buffer buf_n1064( .i (n1063), .o (n1064) );
  buffer buf_n1065( .i (n1064), .o (n1065) );
  buffer buf_n1066( .i (n1065), .o (n1066) );
  buffer buf_n608( .i (x87), .o (n608) );
  buffer buf_n609( .i (n608), .o (n609) );
  buffer buf_n610( .i (n609), .o (n610) );
  buffer buf_n611( .i (n610), .o (n611) );
  buffer buf_n688( .i (n687), .o (n688) );
  assign n2013 = n611 & n688 ;
  buffer buf_n695( .i (n694), .o (n695) );
  assign n2014 = ~n611 & n695 ;
  assign n2015 = ( n1066 & n2013 ) | ( n1066 & n2014 ) | ( n2013 & n2014 ) ;
  buffer buf_n701( .i (n700), .o (n701) );
  assign n2016 = n611 | n701 ;
  buffer buf_n657( .i (n656), .o (n657) );
  assign n2017 = n611 & ~n657 ;
  assign n2018 = ( n1066 & n2016 ) | ( n1066 & ~n2017 ) | ( n2016 & ~n2017 ) ;
  assign n2019 = ~n2015 & n2018 ;
  buffer buf_n2020( .i (n2019), .o (n2020) );
  buffer buf_n994( .i (x134), .o (n994) );
  buffer buf_n995( .i (n994), .o (n995) );
  buffer buf_n996( .i (n995), .o (n996) );
  buffer buf_n997( .i (n996), .o (n997) );
  buffer buf_n998( .i (n997), .o (n998) );
  buffer buf_n733( .i (x108), .o (n733) );
  buffer buf_n734( .i (n733), .o (n734) );
  buffer buf_n735( .i (n734), .o (n735) );
  buffer buf_n736( .i (n735), .o (n736) );
  buffer buf_n2024( .i (n1394), .o (n2024) );
  assign n2025 = n736 & n2024 ;
  buffer buf_n2026( .i (n1388), .o (n2026) );
  assign n2027 = ~n736 & n2026 ;
  assign n2028 = ( n998 & n2025 ) | ( n998 & n2027 ) | ( n2025 & n2027 ) ;
  buffer buf_n2029( .i (n1382), .o (n2029) );
  assign n2030 = n736 | n2029 ;
  buffer buf_n2031( .i (n1376), .o (n2031) );
  assign n2032 = n736 & ~n2031 ;
  assign n2033 = ( n998 & n2030 ) | ( n998 & ~n2032 ) | ( n2030 & ~n2032 ) ;
  assign n2034 = ~n2028 & n2033 ;
  buffer buf_n2035( .i (n2034), .o (n2035) );
  assign n2036 = ~n2020 & n2035 ;
  buffer buf_n1005( .i (x136), .o (n1005) );
  buffer buf_n1006( .i (n1005), .o (n1006) );
  buffer buf_n1007( .i (n1006), .o (n1007) );
  buffer buf_n1008( .i (n1007), .o (n1008) );
  buffer buf_n1009( .i (n1008), .o (n1009) );
  buffer buf_n704( .i (x102), .o (n704) );
  buffer buf_n705( .i (n704), .o (n705) );
  buffer buf_n706( .i (n705), .o (n706) );
  buffer buf_n707( .i (n706), .o (n707) );
  assign n2037 = n707 & n2024 ;
  assign n2038 = ~n707 & n2026 ;
  assign n2039 = ( n1009 & n2037 ) | ( n1009 & n2038 ) | ( n2037 & n2038 ) ;
  assign n2040 = n707 | n2029 ;
  buffer buf_n2041( .i (n706), .o (n2041) );
  assign n2042 = ~n2031 & n2041 ;
  assign n2043 = ( n1009 & n2040 ) | ( n1009 & ~n2042 ) | ( n2040 & ~n2042 ) ;
  assign n2044 = ~n2039 & n2043 ;
  buffer buf_n2045( .i (n2044), .o (n2045) );
  buffer buf_n1039( .i (x139), .o (n1039) );
  buffer buf_n1040( .i (n1039), .o (n1040) );
  buffer buf_n1041( .i (n1040), .o (n1041) );
  buffer buf_n1042( .i (n1041), .o (n1042) );
  buffer buf_n1043( .i (n1042), .o (n1043) );
  buffer buf_n637( .i (x93), .o (n637) );
  buffer buf_n638( .i (n637), .o (n638) );
  buffer buf_n639( .i (n638), .o (n639) );
  buffer buf_n640( .i (n639), .o (n640) );
  assign n2046 = n640 & n2024 ;
  assign n2047 = ~n640 & n2026 ;
  assign n2048 = ( n1043 & n2046 ) | ( n1043 & n2047 ) | ( n2046 & n2047 ) ;
  assign n2049 = n640 | n2029 ;
  assign n2050 = n640 & ~n2031 ;
  assign n2051 = ( n1043 & n2049 ) | ( n1043 & ~n2050 ) | ( n2049 & ~n2050 ) ;
  assign n2052 = ~n2048 & n2051 ;
  buffer buf_n2053( .i (n2052), .o (n2053) );
  assign n2054 = n2045 & n2053 ;
  assign n2055 = n2036 & n2054 ;
  assign n2056 = n2012 & n2055 ;
  assign n2057 = n1993 & n2056 ;
  buffer buf_n2058( .i (n2057), .o (n2058) );
  buffer buf_n2059( .i (n2058), .o (n2059) );
  buffer buf_n2060( .i (n2059), .o (n2060) );
  buffer buf_n2061( .i (n2060), .o (n2061) );
  buffer buf_n2062( .i (n2061), .o (n2062) );
  buffer buf_n2063( .i (n2062), .o (n2063) );
  buffer buf_n2064( .i (n2063), .o (n2064) );
  buffer buf_n2065( .i (n2064), .o (n2065) );
  buffer buf_n2066( .i (n2065), .o (n2066) );
  buffer buf_n2067( .i (n2066), .o (n2067) );
  buffer buf_n2068( .i (n2067), .o (n2068) );
  buffer buf_n2069( .i (n2068), .o (n2069) );
  buffer buf_n1033( .i (n1032), .o (n1033) );
  buffer buf_n729( .i (x107), .o (n729) );
  buffer buf_n730( .i (n729), .o (n730) );
  buffer buf_n731( .i (n730), .o (n731) );
  buffer buf_n856( .i (x123), .o (n856) );
  buffer buf_n857( .i (n856), .o (n857) );
  buffer buf_n858( .i (n857), .o (n858) );
  assign n2070 = n731 & n858 ;
  assign n2071 = n724 & ~n858 ;
  assign n2072 = n2070 | n2071 ;
  buffer buf_n2073( .i (n2072), .o (n2073) );
  assign n2079 = n1033 | n2073 ;
  buffer buf_n2080( .i (n2079), .o (n2080) );
  assign n2081 = n1033 & n2073 ;
  buffer buf_n2082( .i (n2081), .o (n2082) );
  assign n2085 = n2080 & ~n2082 ;
  buffer buf_n2086( .i (n2085), .o (n2086) );
  buffer buf_n711( .i (x103), .o (n711) );
  buffer buf_n712( .i (n711), .o (n712) );
  assign n2089 = ~n712 & n857 ;
  assign n2090 = n705 | n857 ;
  assign n2091 = ~n2089 & n2090 ;
  buffer buf_n2092( .i (n2091), .o (n2092) );
  assign n2100 = n1009 | n2092 ;
  buffer buf_n2101( .i (n2100), .o (n2101) );
  buffer buf_n2106( .i (n1008), .o (n2106) );
  assign n2107 = n2092 & n2106 ;
  buffer buf_n2108( .i (n2107), .o (n2108) );
  assign n2111 = n2101 & ~n2108 ;
  buffer buf_n2112( .i (n2111), .o (n2112) );
  buffer buf_n2113( .i (n2112), .o (n2113) );
  assign n2117 = n2086 & n2113 ;
  buffer buf_n999( .i (n998), .o (n999) );
  buffer buf_n1000( .i (n999), .o (n1000) );
  buffer buf_n738( .i (x109), .o (n738) );
  buffer buf_n739( .i (n738), .o (n739) );
  buffer buf_n740( .i (n739), .o (n740) );
  assign n2118 = n740 & n858 ;
  buffer buf_n2119( .i (n857), .o (n2119) );
  assign n2120 = n735 & ~n2119 ;
  assign n2121 = n2118 | n2120 ;
  buffer buf_n2122( .i (n2121), .o (n2122) );
  buffer buf_n2123( .i (n2122), .o (n2123) );
  assign n2128 = n1000 | n2123 ;
  assign n2129 = n999 & n2122 ;
  buffer buf_n2130( .i (n2129), .o (n2130) );
  assign n2131 = n2128 & ~n2130 ;
  buffer buf_n2132( .i (n2131), .o (n2132) );
  buffer buf_n719( .i (x105), .o (n719) );
  buffer buf_n720( .i (n719), .o (n720) );
  buffer buf_n2135( .i (n856), .o (n2135) );
  assign n2136 = ~n720 & n2135 ;
  assign n2137 = n715 | n2135 ;
  assign n2138 = ~n2136 & n2137 ;
  buffer buf_n2139( .i (n2138), .o (n2139) );
  assign n2147 = n1022 | n2139 ;
  buffer buf_n2148( .i (n2147), .o (n2148) );
  buffer buf_n2151( .i (n1021), .o (n2151) );
  assign n2152 = n2139 & n2151 ;
  buffer buf_n2153( .i (n2152), .o (n2153) );
  assign n2154 = n2148 & ~n2153 ;
  buffer buf_n2155( .i (n2154), .o (n2155) );
  buffer buf_n2156( .i (n2155), .o (n2156) );
  assign n2159 = n2132 & n2156 ;
  assign n2160 = n2117 & n2159 ;
  buffer buf_n2161( .i (n2160), .o (n2161) );
  buffer buf_n2162( .i (n2161), .o (n2162) );
  buffer buf_n2163( .i (n2162), .o (n2163) );
  buffer buf_n2164( .i (n2163), .o (n2164) );
  buffer buf_n651( .i (x96), .o (n651) );
  buffer buf_n652( .i (n651), .o (n652) );
  assign n2165 = ~n652 & n2135 ;
  assign n2166 = n646 | n2135 ;
  assign n2167 = ~n2165 & n2166 ;
  buffer buf_n2168( .i (n2167), .o (n2168) );
  assign n2173 = n1058 | n2168 ;
  buffer buf_n2174( .i (n2173), .o (n2174) );
  buffer buf_n2175( .i (n2174), .o (n2175) );
  buffer buf_n2176( .i (n2175), .o (n2176) );
  buffer buf_n2177( .i (n2176), .o (n2177) );
  buffer buf_n2178( .i (n2177), .o (n2178) );
  buffer buf_n2179( .i (n2178), .o (n2179) );
  buffer buf_n1093( .i (n1092), .o (n1093) );
  buffer buf_n633( .i (x92), .o (n633) );
  buffer buf_n634( .i (n633), .o (n634) );
  buffer buf_n635( .i (n634), .o (n635) );
  assign n2182 = ~n635 & n2119 ;
  assign n2183 = n629 | n2119 ;
  assign n2184 = ~n2182 & n2183 ;
  buffer buf_n2185( .i (n2184), .o (n2185) );
  assign n2187 = n1093 & n2185 ;
  buffer buf_n2188( .i (n2187), .o (n2188) );
  assign n2189 = n1093 | n2185 ;
  buffer buf_n2190( .i (n2189), .o (n2190) );
  assign n2192 = ~n2188 & n2190 ;
  buffer buf_n2193( .i (n2192), .o (n2193) );
  buffer buf_n1085( .i (n1084), .o (n1085) );
  buffer buf_n623( .i (x90), .o (n623) );
  buffer buf_n624( .i (n623), .o (n624) );
  buffer buf_n625( .i (n624), .o (n625) );
  assign n2200 = ~n625 & n2119 ;
  buffer buf_n2201( .i (n856), .o (n2201) );
  buffer buf_n2202( .i (n2201), .o (n2202) );
  assign n2203 = n620 | n2202 ;
  assign n2204 = ~n2200 & n2203 ;
  buffer buf_n2205( .i (n2204), .o (n2205) );
  assign n2215 = n1085 | n2205 ;
  buffer buf_n2216( .i (n2215), .o (n2216) );
  assign n2224 = n1085 & n2205 ;
  buffer buf_n2225( .i (n2224), .o (n2225) );
  assign n2234 = n2216 & ~n2225 ;
  buffer buf_n2235( .i (n2234), .o (n2235) );
  assign n2242 = n2193 & ~n2235 ;
  buffer buf_n2243( .i (n2242), .o (n2243) );
  buffer buf_n642( .i (x94), .o (n642) );
  buffer buf_n643( .i (n642), .o (n643) );
  assign n2244 = ~n643 & n2201 ;
  assign n2245 = n638 | n2201 ;
  assign n2246 = ~n2244 & n2245 ;
  buffer buf_n2247( .i (n2246), .o (n2247) );
  assign n2257 = n1043 | n2247 ;
  buffer buf_n2258( .i (n2257), .o (n2258) );
  buffer buf_n2263( .i (n1042), .o (n2263) );
  assign n2264 = n2247 & n2263 ;
  buffer buf_n2265( .i (n2264), .o (n2265) );
  assign n2267 = n2258 & ~n2265 ;
  buffer buf_n2268( .i (n2267), .o (n2268) );
  buffer buf_n2269( .i (n2268), .o (n2269) );
  buffer buf_n2270( .i (n2269), .o (n2270) );
  assign n2277 = n2178 & ~n2270 ;
  assign n2278 = ( n2179 & n2243 ) | ( n2179 & n2277 ) | ( n2243 & n2277 ) ;
  buffer buf_n2279( .i (n2278), .o (n2279) );
  buffer buf_n2087( .i (n2086), .o (n2087) );
  buffer buf_n2124( .i (n2123), .o (n2124) );
  buffer buf_n2125( .i (n2124), .o (n2125) );
  buffer buf_n2126( .i (n2125), .o (n2126) );
  buffer buf_n2127( .i (n2126), .o (n2127) );
  assign n2280 = ~n2087 & n2127 ;
  buffer buf_n2102( .i (n2101), .o (n2102) );
  buffer buf_n2103( .i (n2102), .o (n2103) );
  buffer buf_n2104( .i (n2103), .o (n2104) );
  buffer buf_n2105( .i (n2104), .o (n2105) );
  buffer buf_n1059( .i (n1058), .o (n1059) );
  buffer buf_n2169( .i (n2168), .o (n2169) );
  assign n2281 = n1059 & n2169 ;
  assign n2282 = n2174 & ~n2281 ;
  buffer buf_n2283( .i (n2282), .o (n2283) );
  buffer buf_n2284( .i (n2283), .o (n2284) );
  buffer buf_n2285( .i (n2284), .o (n2285) );
  assign n2289 = n2105 & ~n2285 ;
  assign n2290 = n2280 | n2289 ;
  buffer buf_n2217( .i (n2216), .o (n2217) );
  buffer buf_n2218( .i (n2217), .o (n2218) );
  buffer buf_n2219( .i (n2218), .o (n2219) );
  buffer buf_n1067( .i (n1066), .o (n1067) );
  buffer buf_n1068( .i (n1067), .o (n1068) );
  buffer buf_n613( .i (x88), .o (n613) );
  buffer buf_n614( .i (n613), .o (n614) );
  buffer buf_n615( .i (n614), .o (n615) );
  buffer buf_n616( .i (n615), .o (n616) );
  buffer buf_n859( .i (n858), .o (n859) );
  assign n2291 = ~n616 & n859 ;
  buffer buf_n2292( .i (n610), .o (n2292) );
  assign n2293 = n859 | n2292 ;
  assign n2294 = ~n2291 & n2293 ;
  buffer buf_n2295( .i (n2294), .o (n2295) );
  assign n2306 = n1068 & n2295 ;
  assign n2307 = n1068 | n2295 ;
  assign n2308 = ~n2306 & n2307 ;
  buffer buf_n2309( .i (n2308), .o (n2309) );
  buffer buf_n2310( .i (n2309), .o (n2310) );
  assign n2315 = n2219 & ~n2310 ;
  buffer buf_n2194( .i (n2193), .o (n2194) );
  buffer buf_n2259( .i (n2258), .o (n2259) );
  buffer buf_n2260( .i (n2259), .o (n2260) );
  buffer buf_n2261( .i (n2260), .o (n2261) );
  buffer buf_n2262( .i (n2261), .o (n2262) );
  assign n2316 = ~n2194 & n2262 ;
  assign n2317 = n2315 | n2316 ;
  assign n2318 = n2290 | n2317 ;
  assign n2319 = n2279 | n2318 ;
  buffer buf_n2320( .i (n2319), .o (n2320) );
  assign n2322 = n2164 & ~n2320 ;
  buffer buf_n2323( .i (n2322), .o (n2323) );
  buffer buf_n2324( .i (n2323), .o (n2324) );
  buffer buf_n2325( .i (n2324), .o (n2325) );
  buffer buf_n2326( .i (n2325), .o (n2326) );
  buffer buf_n2327( .i (n2326), .o (n2327) );
  buffer buf_n2328( .i (n2327), .o (n2328) );
  buffer buf_n2329( .i (n2328), .o (n2329) );
  buffer buf_n845( .i (x122), .o (n845) );
  buffer buf_n846( .i (n845), .o (n846) );
  buffer buf_n847( .i (n846), .o (n847) );
  buffer buf_n848( .i (n847), .o (n848) );
  buffer buf_n950( .i (n949), .o (n950) );
  assign n2330 = n848 | n950 ;
  assign n2331 = n848 & ~n955 ;
  assign n2332 = n2330 & ~n2331 ;
  buffer buf_n2333( .i (n2332), .o (n2333) );
  buffer buf_n2334( .i (n2333), .o (n2334) );
  buffer buf_n2335( .i (n2334), .o (n2335) );
  buffer buf_n2336( .i (n2335), .o (n2336) );
  buffer buf_n2337( .i (n2336), .o (n2337) );
  buffer buf_n2338( .i (n2337), .o (n2338) );
  buffer buf_n2339( .i (n2338), .o (n2339) );
  buffer buf_n2340( .i (n2339), .o (n2340) );
  buffer buf_n2341( .i (n2340), .o (n2341) );
  buffer buf_n2342( .i (n2341), .o (n2342) );
  buffer buf_n2343( .i (n2342), .o (n2343) );
  buffer buf_n2344( .i (n2343), .o (n2344) );
  buffer buf_n2345( .i (n2344), .o (n2345) );
  buffer buf_n1130( .i (n1129), .o (n1130) );
  buffer buf_n1131( .i (n1130), .o (n1131) );
  buffer buf_n1132( .i (n1131), .o (n1132) );
  buffer buf_n840( .i (x121), .o (n840) );
  buffer buf_n841( .i (n840), .o (n841) );
  buffer buf_n842( .i (n841), .o (n842) );
  buffer buf_n843( .i (n842), .o (n843) );
  assign n2346 = n843 & n848 ;
  buffer buf_n2347( .i (n847), .o (n2347) );
  assign n2348 = n837 & ~n2347 ;
  assign n2349 = n2346 | n2348 ;
  buffer buf_n2350( .i (n2349), .o (n2350) );
  assign n2357 = n1132 & n2350 ;
  assign n2358 = n1132 | n2350 ;
  assign n2359 = ~n2357 & n2358 ;
  buffer buf_n2360( .i (n2359), .o (n2360) );
  buffer buf_n1143( .i (n1142), .o (n1143) );
  assign n2364 = n846 & ~n862 ;
  buffer buf_n2365( .i (n2364), .o (n2365) );
  assign n2373 = n1143 & ~n2365 ;
  buffer buf_n2374( .i (n2373), .o (n2374) );
  assign n2380 = ~n1143 & n2365 ;
  buffer buf_n2381( .i (n2380), .o (n2381) );
  assign n2385 = n2374 | n2381 ;
  buffer buf_n2386( .i (n2385), .o (n2386) );
  assign n2391 = n845 & n892 ;
  assign n2392 = ~n845 & n886 ;
  assign n2393 = n2391 | n2392 ;
  buffer buf_n2394( .i (n2393), .o (n2394) );
  assign n2399 = n1932 & n2394 ;
  buffer buf_n2400( .i (n2399), .o (n2400) );
  buffer buf_n1156( .i (n1155), .o (n1156) );
  buffer buf_n2395( .i (n2394), .o (n2395) );
  assign n2404 = n1156 | n2395 ;
  assign n2405 = ~n2400 & n2404 ;
  buffer buf_n2406( .i (n2405), .o (n2406) );
  assign n2410 = ~n2386 & n2406 ;
  buffer buf_n2411( .i (n2410), .o (n2411) );
  assign n2414 = n2360 & n2411 ;
  buffer buf_n2415( .i (n2414), .o (n2415) );
  buffer buf_n1099( .i (n1098), .o (n1099) );
  buffer buf_n1100( .i (n1099), .o (n1100) );
  buffer buf_n816( .i (x117), .o (n816) );
  buffer buf_n817( .i (n816), .o (n817) );
  assign n2416 = ~n817 & n846 ;
  assign n2417 = n812 | n846 ;
  assign n2418 = ~n2416 & n2417 ;
  buffer buf_n2419( .i (n2418), .o (n2419) );
  assign n2428 = n1100 & n2419 ;
  buffer buf_n2429( .i (n2428), .o (n2429) );
  assign n2436 = n1100 | n2419 ;
  buffer buf_n2437( .i (n2436), .o (n2437) );
  assign n2443 = ~n2429 & n2437 ;
  buffer buf_n2444( .i (n2443), .o (n2444) );
  buffer buf_n1113( .i (n1112), .o (n1113) );
  buffer buf_n1114( .i (n1113), .o (n1114) );
  buffer buf_n1115( .i (n1114), .o (n1115) );
  buffer buf_n1116( .i (n1115), .o (n1116) );
  buffer buf_n828( .i (x119), .o (n828) );
  buffer buf_n829( .i (n828), .o (n829) );
  buffer buf_n830( .i (n829), .o (n830) );
  buffer buf_n831( .i (n830), .o (n831) );
  assign n2453 = ~n831 & n2347 ;
  assign n2454 = n826 | n2347 ;
  assign n2455 = ~n2453 & n2454 ;
  buffer buf_n2456( .i (n2455), .o (n2456) );
  assign n2465 = n1116 | n2456 ;
  buffer buf_n2466( .i (n2465), .o (n2466) );
  assign n2471 = n2444 & n2466 ;
  buffer buf_n2472( .i (n2471), .o (n2472) );
  buffer buf_n2473( .i (n2472), .o (n2473) );
  assign n2474 = n2415 & n2473 ;
  buffer buf_n2475( .i (n2474), .o (n2475) );
  buffer buf_n2476( .i (n2475), .o (n2476) );
  buffer buf_n2477( .i (n2476), .o (n2477) );
  buffer buf_n2478( .i (n2477), .o (n2478) );
  buffer buf_n1167( .i (n1166), .o (n1167) );
  buffer buf_n1168( .i (n1167), .o (n1168) );
  buffer buf_n1169( .i (n1168), .o (n1169) );
  buffer buf_n2479( .i (n919), .o (n2479) );
  assign n2480 = n2347 | n2479 ;
  buffer buf_n2481( .i (n847), .o (n2481) );
  assign n2482 = ~n925 & n2481 ;
  assign n2483 = n2480 & ~n2482 ;
  buffer buf_n2484( .i (n2483), .o (n2484) );
  buffer buf_n2485( .i (n2484), .o (n2485) );
  assign n2487 = n1169 & n2485 ;
  assign n2488 = n1168 | n2484 ;
  buffer buf_n2489( .i (n2488), .o (n2489) );
  assign n2490 = ~n2487 & n2489 ;
  buffer buf_n2491( .i (n2490), .o (n2491) );
  buffer buf_n2492( .i (n2491), .o (n2492) );
  buffer buf_n2493( .i (n2492), .o (n2493) );
  buffer buf_n2494( .i (n2493), .o (n2494) );
  buffer buf_n2495( .i (n2494), .o (n2495) );
  buffer buf_n2496( .i (n2495), .o (n2496) );
  buffer buf_n849( .i (n848), .o (n849) );
  buffer buf_n850( .i (n849), .o (n850) );
  buffer buf_n851( .i (n850), .o (n851) );
  buffer buf_n852( .i (n851), .o (n852) );
  buffer buf_n853( .i (n852), .o (n853) );
  buffer buf_n854( .i (n853), .o (n854) );
  assign n2497 = ~n783 & n854 ;
  assign n2498 = n758 | n854 ;
  assign n2499 = ~n2497 & n2498 ;
  buffer buf_n2500( .i (n2499), .o (n2500) );
  buffer buf_n805( .i (x115), .o (n805) );
  buffer buf_n806( .i (n805), .o (n806) );
  buffer buf_n807( .i (n806), .o (n807) );
  buffer buf_n808( .i (n807), .o (n808) );
  buffer buf_n809( .i (n808), .o (n809) );
  assign n2507 = n809 & n849 ;
  buffer buf_n802( .i (n801), .o (n802) );
  buffer buf_n803( .i (n802), .o (n803) );
  assign n2508 = n803 & ~n849 ;
  assign n2509 = n2507 | n2508 ;
  buffer buf_n2510( .i (n2509), .o (n2510) );
  buffer buf_n2511( .i (n2510), .o (n2511) );
  buffer buf_n2512( .i (n2511), .o (n2512) );
  buffer buf_n2513( .i (n2512), .o (n2513) );
  buffer buf_n2514( .i (n2513), .o (n2514) );
  buffer buf_n2515( .i (n2514), .o (n2515) );
  assign n2520 = n2500 | n2515 ;
  buffer buf_n2521( .i (n2520), .o (n2521) );
  buffer buf_n1117( .i (n1116), .o (n1117) );
  buffer buf_n1118( .i (n1117), .o (n1118) );
  buffer buf_n1119( .i (n1118), .o (n1119) );
  buffer buf_n1120( .i (n1119), .o (n1120) );
  buffer buf_n2457( .i (n2456), .o (n2457) );
  buffer buf_n2458( .i (n2457), .o (n2458) );
  buffer buf_n2459( .i (n2458), .o (n2459) );
  buffer buf_n2460( .i (n2459), .o (n2460) );
  assign n2523 = n1120 & n2460 ;
  buffer buf_n2524( .i (n2523), .o (n2524) );
  buffer buf_n2525( .i (n2524), .o (n2525) );
  buffer buf_n2526( .i (n2525), .o (n2526) );
  assign n2527 = n2521 | n2526 ;
  assign n2528 = n2496 & ~n2527 ;
  assign n2529 = n2478 & n2528 ;
  buffer buf_n2530( .i (n2529), .o (n2530) );
  assign n2531 = ~n2345 & n2530 ;
  buffer buf_n2532( .i (n2531), .o (n2532) );
  buffer buf_n2533( .i (n2532), .o (n2533) );
  buffer buf_n2534( .i (n2533), .o (n2534) );
  buffer buf_n2535( .i (n2534), .o (n2535) );
  buffer buf_n977( .i (x131), .o (n977) );
  buffer buf_n978( .i (n977), .o (n978) );
  buffer buf_n979( .i (n978), .o (n979) );
  buffer buf_n980( .i (n979), .o (n980) );
  buffer buf_n981( .i (n980), .o (n981) );
  buffer buf_n982( .i (n981), .o (n982) );
  buffer buf_n983( .i (n982), .o (n983) );
  buffer buf_n984( .i (n983), .o (n984) );
  assign n2536 = ( ~n799 & n811 ) | ( ~n799 & n823 ) | ( n811 & n823 ) ;
  assign n2537 = ( n799 & n811 ) | ( n799 & n823 ) | ( n811 & n823 ) ;
  assign n2538 = ( n800 & n2536 ) | ( n800 & ~n2537 ) | ( n2536 & ~n2537 ) ;
  buffer buf_n2539( .i (n2538), .o (n2539) );
  assign n2540 = ( ~n889 & n950 ) | ( ~n889 & n2539 ) | ( n950 & n2539 ) ;
  assign n2541 = ( n889 & n950 ) | ( n889 & n2539 ) | ( n950 & n2539 ) ;
  assign n2542 = ( n890 & n2540 ) | ( n890 & ~n2541 ) | ( n2540 & ~n2541 ) ;
  buffer buf_n2543( .i (n2542), .o (n2543) );
  assign n2544 = ( ~n750 & n835 ) | ( ~n750 & n918 ) | ( n835 & n918 ) ;
  assign n2545 = ( n750 & n835 ) | ( n750 & n918 ) | ( n835 & n918 ) ;
  assign n2546 = ( n751 & n2544 ) | ( n751 & ~n2545 ) | ( n2544 & ~n2545 ) ;
  buffer buf_n2547( .i (n2546), .o (n2547) );
  buffer buf_n2548( .i (n2547), .o (n2548) );
  buffer buf_n2549( .i (n2548), .o (n2549) );
  assign n2550 = ( n983 & n2543 ) | ( n983 & ~n2549 ) | ( n2543 & ~n2549 ) ;
  assign n2551 = ( n983 & ~n2543 ) | ( n983 & n2549 ) | ( ~n2543 & n2549 ) ;
  assign n2552 = ( ~n984 & n2550 ) | ( ~n984 & n2551 ) | ( n2550 & n2551 ) ;
  buffer buf_n2553( .i (n2552), .o (n2553) );
  buffer buf_n2554( .i (n2553), .o (n2554) );
  buffer buf_n2555( .i (n2554), .o (n2555) );
  buffer buf_n2556( .i (n2555), .o (n2556) );
  buffer buf_n2557( .i (n2556), .o (n2557) );
  buffer buf_n2558( .i (n2557), .o (n2558) );
  buffer buf_n2559( .i (n2558), .o (n2559) );
  buffer buf_n2560( .i (n2559), .o (n2560) );
  buffer buf_n2561( .i (n2560), .o (n2561) );
  buffer buf_n2562( .i (n2561), .o (n2562) );
  buffer buf_n2563( .i (n2562), .o (n2563) );
  buffer buf_n2564( .i (n2563), .o (n2564) );
  buffer buf_n2565( .i (n2564), .o (n2565) );
  buffer buf_n2566( .i (n2565), .o (n2566) );
  buffer buf_n2567( .i (n2566), .o (n2567) );
  buffer buf_n649( .i (n648), .o (n649) );
  assign n2568 = ( ~n618 & n627 ) | ( ~n618 & n637 ) | ( n627 & n637 ) ;
  assign n2569 = ( n618 & n627 ) | ( n618 & n637 ) | ( n627 & n637 ) ;
  assign n2570 = ( n619 & n2568 ) | ( n619 & ~n2569 ) | ( n2568 & ~n2569 ) ;
  buffer buf_n2571( .i (n2570), .o (n2571) );
  buffer buf_n2572( .i (n716), .o (n2572) );
  assign n2573 = ( ~n1998 & n2571 ) | ( ~n1998 & n2572 ) | ( n2571 & n2572 ) ;
  assign n2574 = ( n1998 & n2571 ) | ( n1998 & n2572 ) | ( n2571 & n2572 ) ;
  assign n2575 = ( n649 & n2573 ) | ( n649 & ~n2574 ) | ( n2573 & ~n2574 ) ;
  buffer buf_n2576( .i (n2575), .o (n2576) );
  buffer buf_n2577( .i (n2576), .o (n2577) );
  buffer buf_n708( .i (n707), .o (n708) );
  buffer buf_n709( .i (n708), .o (n709) );
  buffer buf_n742( .i (x110), .o (n742) );
  buffer buf_n743( .i (n742), .o (n743) );
  assign n2578 = ( ~n609 & n734 ) | ( ~n609 & n743 ) | ( n734 & n743 ) ;
  assign n2579 = ( n609 & n734 ) | ( n609 & n743 ) | ( n734 & n743 ) ;
  assign n2580 = ( n610 & n2578 ) | ( n610 & ~n2579 ) | ( n2578 & ~n2579 ) ;
  buffer buf_n2581( .i (n2580), .o (n2581) );
  assign n2582 = ( n708 & ~n726 ) | ( n708 & n2581 ) | ( ~n726 & n2581 ) ;
  assign n2583 = ( n708 & n726 ) | ( n708 & ~n2581 ) | ( n726 & ~n2581 ) ;
  assign n2584 = ( ~n709 & n2582 ) | ( ~n709 & n2583 ) | ( n2582 & n2583 ) ;
  buffer buf_n2585( .i (n2584), .o (n2585) );
  assign n2586 = ~n2577 & n2585 ;
  assign n2587 = n2577 & ~n2585 ;
  assign n2588 = n2586 | n2587 ;
  buffer buf_n2589( .i (n2588), .o (n2589) );
  buffer buf_n2590( .i (n2589), .o (n2590) );
  buffer buf_n2591( .i (n2590), .o (n2591) );
  buffer buf_n2592( .i (n2591), .o (n2592) );
  buffer buf_n2593( .i (n2592), .o (n2593) );
  buffer buf_n2594( .i (n2593), .o (n2594) );
  buffer buf_n2595( .i (n2594), .o (n2595) );
  buffer buf_n2596( .i (n2595), .o (n2596) );
  buffer buf_n2597( .i (n2596), .o (n2597) );
  buffer buf_n2598( .i (n2597), .o (n2598) );
  buffer buf_n2599( .i (n2598), .o (n2599) );
  buffer buf_n2600( .i (n2599), .o (n2600) );
  buffer buf_n2601( .i (n2600), .o (n2601) );
  buffer buf_n2602( .i (n2601), .o (n2602) );
  buffer buf_n1069( .i (n1068), .o (n1069) );
  buffer buf_n1070( .i (n1069), .o (n1070) );
  buffer buf_n1071( .i (n1070), .o (n1071) );
  buffer buf_n1072( .i (n1071), .o (n1072) );
  buffer buf_n1073( .i (n1072), .o (n1073) );
  buffer buf_n1074( .i (n1073), .o (n1074) );
  buffer buf_n1075( .i (n1074), .o (n1075) );
  buffer buf_n1076( .i (n1075), .o (n1076) );
  buffer buf_n1077( .i (n1076), .o (n1077) );
  buffer buf_n1078( .i (n1077), .o (n1078) );
  buffer buf_n2296( .i (n2295), .o (n2296) );
  buffer buf_n2297( .i (n2296), .o (n2297) );
  buffer buf_n2298( .i (n2297), .o (n2298) );
  buffer buf_n2299( .i (n2298), .o (n2299) );
  buffer buf_n2300( .i (n2299), .o (n2300) );
  buffer buf_n2301( .i (n2300), .o (n2301) );
  buffer buf_n2302( .i (n2301), .o (n2302) );
  buffer buf_n2303( .i (n2302), .o (n2303) );
  buffer buf_n2304( .i (n2303), .o (n2304) );
  buffer buf_n2305( .i (n2304), .o (n2305) );
  buffer buf_n2226( .i (n2225), .o (n2226) );
  buffer buf_n2227( .i (n2226), .o (n2227) );
  buffer buf_n2228( .i (n2227), .o (n2228) );
  buffer buf_n2229( .i (n2228), .o (n2229) );
  buffer buf_n2230( .i (n2229), .o (n2230) );
  buffer buf_n2231( .i (n2230), .o (n2231) );
  buffer buf_n2232( .i (n2231), .o (n2232) );
  buffer buf_n2233( .i (n2232), .o (n2233) );
  buffer buf_n2220( .i (n2219), .o (n2220) );
  buffer buf_n2221( .i (n2220), .o (n2221) );
  buffer buf_n2222( .i (n2221), .o (n2222) );
  buffer buf_n2223( .i (n2222), .o (n2223) );
  buffer buf_n2180( .i (n2179), .o (n2180) );
  buffer buf_n2181( .i (n2180), .o (n2181) );
  buffer buf_n1094( .i (n1093), .o (n1094) );
  buffer buf_n2186( .i (n2185), .o (n2186) );
  assign n2603 = ( n1094 & n2186 ) | ( n1094 & n2265 ) | ( n2186 & n2265 ) ;
  buffer buf_n2604( .i (n2603), .o (n2604) );
  buffer buf_n2605( .i (n2604), .o (n2605) );
  buffer buf_n2606( .i (n2605), .o (n2606) );
  buffer buf_n2607( .i (n2606), .o (n2607) );
  buffer buf_n2608( .i (n2607), .o (n2608) );
  buffer buf_n2609( .i (n2608), .o (n2609) );
  buffer buf_n1034( .i (n1033), .o (n1034) );
  buffer buf_n1035( .i (n1034), .o (n1035) );
  buffer buf_n2074( .i (n2073), .o (n2074) );
  buffer buf_n2075( .i (n2074), .o (n2075) );
  assign n2610 = ( n1035 & n2075 ) | ( n1035 & n2130 ) | ( n2075 & n2130 ) ;
  buffer buf_n2611( .i (n2610), .o (n2611) );
  buffer buf_n2149( .i (n2148), .o (n2149) );
  assign n2612 = n2102 & n2149 ;
  buffer buf_n2613( .i (n2612), .o (n2613) );
  assign n2616 = n2611 & n2613 ;
  buffer buf_n1010( .i (n1009), .o (n1010) );
  buffer buf_n1011( .i (n1010), .o (n1011) );
  buffer buf_n2093( .i (n2092), .o (n2093) );
  buffer buf_n2094( .i (n2093), .o (n2094) );
  assign n2617 = ( n1011 & n2094 ) | ( n1011 & n2153 ) | ( n2094 & n2153 ) ;
  buffer buf_n2618( .i (n2617), .o (n2618) );
  buffer buf_n2619( .i (n2618), .o (n2619) );
  assign n2621 = n2284 & ~n2619 ;
  assign n2622 = ~n2616 & n2621 ;
  buffer buf_n2623( .i (n2622), .o (n2623) );
  assign n2625 = n2190 & n2259 ;
  buffer buf_n2626( .i (n2625), .o (n2626) );
  buffer buf_n2627( .i (n2626), .o (n2627) );
  buffer buf_n2628( .i (n2627), .o (n2628) );
  buffer buf_n2629( .i (n2628), .o (n2629) );
  assign n2631 = ( n2608 & ~n2623 ) | ( n2608 & n2629 ) | ( ~n2623 & n2629 ) ;
  assign n2632 = ( n2181 & n2609 ) | ( n2181 & n2631 ) | ( n2609 & n2631 ) ;
  assign n2633 = n2223 & n2632 ;
  assign n2634 = n2233 | n2633 ;
  assign n2635 = ( n1078 & n2305 ) | ( n1078 & n2634 ) | ( n2305 & n2634 ) ;
  buffer buf_n2636( .i (n2635), .o (n2636) );
  buffer buf_n2637( .i (n2636), .o (n2637) );
  buffer buf_n2638( .i (n2637), .o (n2638) );
  buffer buf_n2639( .i (n2638), .o (n2639) );
  buffer buf_n2640( .i (n2639), .o (n2640) );
  buffer buf_n2641( .i (n2640), .o (n2641) );
  buffer buf_n2522( .i (n2521), .o (n2522) );
  buffer buf_n1101( .i (n1100), .o (n1101) );
  buffer buf_n1102( .i (n1101), .o (n1102) );
  buffer buf_n1103( .i (n1102), .o (n1103) );
  buffer buf_n1104( .i (n1103), .o (n1104) );
  buffer buf_n1105( .i (n1104), .o (n1105) );
  buffer buf_n1106( .i (n1105), .o (n1106) );
  buffer buf_n1107( .i (n1106), .o (n1107) );
  buffer buf_n1108( .i (n1107), .o (n1108) );
  buffer buf_n2420( .i (n2419), .o (n2420) );
  buffer buf_n2421( .i (n2420), .o (n2421) );
  buffer buf_n2422( .i (n2421), .o (n2422) );
  buffer buf_n2423( .i (n2422), .o (n2423) );
  buffer buf_n2424( .i (n2423), .o (n2424) );
  buffer buf_n2425( .i (n2424), .o (n2425) );
  buffer buf_n2426( .i (n2425), .o (n2426) );
  buffer buf_n2427( .i (n2426), .o (n2427) );
  buffer buf_n2467( .i (n2466), .o (n2467) );
  buffer buf_n2468( .i (n2467), .o (n2468) );
  buffer buf_n2469( .i (n2468), .o (n2469) );
  buffer buf_n2412( .i (n2411), .o (n2412) );
  assign n2642 = ( n1168 & n2333 ) | ( n1168 & n2484 ) | ( n2333 & n2484 ) ;
  buffer buf_n2643( .i (n2642), .o (n2643) );
  buffer buf_n2644( .i (n2643), .o (n2644) );
  assign n2645 = n2360 & n2644 ;
  assign n2646 = n2412 & n2645 ;
  buffer buf_n1133( .i (n1132), .o (n1133) );
  buffer buf_n1134( .i (n1133), .o (n1134) );
  buffer buf_n2351( .i (n2350), .o (n2351) );
  buffer buf_n2352( .i (n2351), .o (n2352) );
  buffer buf_n2375( .i (n2374), .o (n2375) );
  buffer buf_n2376( .i (n2375), .o (n2376) );
  buffer buf_n2401( .i (n2400), .o (n2401) );
  buffer buf_n2402( .i (n2401), .o (n2402) );
  buffer buf_n2382( .i (n2381), .o (n2382) );
  assign n2647 = ~n2375 & n2382 ;
  assign n2648 = ( n2376 & n2402 ) | ( n2376 & ~n2647 ) | ( n2402 & ~n2647 ) ;
  assign n2649 = ( n1134 & n2352 ) | ( n1134 & n2648 ) | ( n2352 & n2648 ) ;
  buffer buf_n2650( .i (n2649), .o (n2650) );
  assign n2653 = ( n1120 & n2460 ) | ( n1120 & n2650 ) | ( n2460 & n2650 ) ;
  assign n2654 = ( n2469 & n2646 ) | ( n2469 & n2653 ) | ( n2646 & n2653 ) ;
  assign n2655 = ( n1108 & n2427 ) | ( n1108 & n2654 ) | ( n2427 & n2654 ) ;
  buffer buf_n2656( .i (n2655), .o (n2656) );
  buffer buf_n2657( .i (n2656), .o (n2657) );
  assign n2658 = n2522 | n2657 ;
  buffer buf_n2659( .i (n2658), .o (n2659) );
  buffer buf_n2660( .i (n2659), .o (n2660) );
  buffer buf_n2661( .i (n2660), .o (n2661) );
  buffer buf_n2662( .i (n2661), .o (n2662) );
  buffer buf_n2663( .i (n2662), .o (n2663) );
  buffer buf_n2664( .i (n2663), .o (n2664) );
  buffer buf_n2665( .i (n2664), .o (n2665) );
  buffer buf_n1506( .i (x175), .o (n1506) );
  buffer buf_n1507( .i (n1506), .o (n1507) );
  buffer buf_n1508( .i (n1507), .o (n1508) );
  buffer buf_n1523( .i (x176), .o (n1523) );
  buffer buf_n1524( .i (n1523), .o (n1524) );
  buffer buf_n1525( .i (n1524), .o (n1525) );
  assign n2666 = n1508 | n1525 ;
  buffer buf_n2667( .i (n2666), .o (n2667) );
  buffer buf_n2668( .i (n2667), .o (n2668) );
  assign n2679 = n1918 & ~n2668 ;
  buffer buf_n2680( .i (n2679), .o (n2680) );
  buffer buf_n2681( .i (n2680), .o (n2681) );
  buffer buf_n2682( .i (n2681), .o (n2682) );
  buffer buf_n2683( .i (n2682), .o (n2683) );
  buffer buf_n2684( .i (n2683), .o (n2684) );
  buffer buf_n2685( .i (n2684), .o (n2685) );
  buffer buf_n1509( .i (n1508), .o (n1509) );
  buffer buf_n1510( .i (n1509), .o (n1510) );
  buffer buf_n1511( .i (n1510), .o (n1511) );
  buffer buf_n1512( .i (n1511), .o (n1512) );
  buffer buf_n1513( .i (n1512), .o (n1513) );
  buffer buf_n1514( .i (n1513), .o (n1514) );
  buffer buf_n1515( .i (n1514), .o (n1515) );
  buffer buf_n1516( .i (n1515), .o (n1516) );
  buffer buf_n1517( .i (n1516), .o (n1517) );
  buffer buf_n1526( .i (n1525), .o (n1526) );
  buffer buf_n1527( .i (n1526), .o (n1527) );
  buffer buf_n1528( .i (n1527), .o (n1528) );
  buffer buf_n1529( .i (n1528), .o (n1529) );
  buffer buf_n1530( .i (n1529), .o (n1530) );
  buffer buf_n1531( .i (n1530), .o (n1531) );
  buffer buf_n1532( .i (n1531), .o (n1532) );
  buffer buf_n1533( .i (n1532), .o (n1533) );
  buffer buf_n139( .i (x20), .o (n139) );
  buffer buf_n140( .i (n139), .o (n140) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  buffer buf_n143( .i (n142), .o (n143) );
  buffer buf_n144( .i (n143), .o (n144) );
  buffer buf_n145( .i (n144), .o (n145) );
  assign n2686 = n145 | n2333 ;
  buffer buf_n2687( .i (n2686), .o (n2687) );
  buffer buf_n146( .i (n145), .o (n146) );
  assign n2690 = n146 & n2334 ;
  assign n2691 = n2687 & ~n2690 ;
  buffer buf_n2692( .i (n2691), .o (n2692) );
  assign n2701 = n1533 | n2692 ;
  buffer buf_n424( .i (x59), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  buffer buf_n427( .i (n426), .o (n427) );
  buffer buf_n428( .i (n427), .o (n428) );
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  assign n2702 = ~n431 & n1530 ;
  buffer buf_n2703( .i (n2702), .o (n2703) );
  buffer buf_n2704( .i (n2703), .o (n2704) );
  buffer buf_n2705( .i (n2704), .o (n2705) );
  assign n2706 = ( n1517 & n2701 ) | ( n1517 & n2705 ) | ( n2701 & n2705 ) ;
  assign n2707 = n2685 | n2706 ;
  buffer buf_n2708( .i (n2707), .o (n2708) );
  buffer buf_n2709( .i (n2708), .o (n2709) );
  buffer buf_n2710( .i (n2709), .o (n2710) );
  buffer buf_n2711( .i (n2710), .o (n2711) );
  buffer buf_n2712( .i (n2711), .o (n2712) );
  buffer buf_n2713( .i (n2712), .o (n2713) );
  buffer buf_n2714( .i (n2713), .o (n2714) );
  buffer buf_n2715( .i (n2714), .o (n2715) );
  buffer buf_n2716( .i (n2715), .o (n2716) );
  buffer buf_n2717( .i (n2716), .o (n2717) );
  buffer buf_n2669( .i (n2668), .o (n2669) );
  buffer buf_n2670( .i (n2669), .o (n2670) );
  assign n2718 = n1944 & ~n2670 ;
  buffer buf_n2719( .i (n2718), .o (n2719) );
  buffer buf_n2720( .i (n2719), .o (n2720) );
  buffer buf_n2721( .i (n2720), .o (n2721) );
  buffer buf_n2722( .i (n2721), .o (n2722) );
  buffer buf_n2688( .i (n2687), .o (n2688) );
  buffer buf_n2689( .i (n2688), .o (n2689) );
  assign n2723 = n2491 & n2689 ;
  assign n2724 = ( ~n1533 & n2491 ) | ( ~n1533 & n2689 ) | ( n2491 & n2689 ) ;
  buffer buf_n408( .i (x57), .o (n408) );
  buffer buf_n409( .i (n408), .o (n409) );
  buffer buf_n410( .i (n409), .o (n410) );
  buffer buf_n411( .i (n410), .o (n411) );
  buffer buf_n412( .i (n411), .o (n412) );
  buffer buf_n413( .i (n412), .o (n413) );
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  assign n2725 = ( ~n415 & n1513 ) | ( ~n415 & n2670 ) | ( n1513 & n2670 ) ;
  buffer buf_n2726( .i (n2725), .o (n2726) );
  buffer buf_n2727( .i (n2726), .o (n2727) );
  buffer buf_n2728( .i (n2727), .o (n2728) );
  assign n2729 = ( n2723 & ~n2724 ) | ( n2723 & n2728 ) | ( ~n2724 & n2728 ) ;
  assign n2730 = n2722 | n2729 ;
  buffer buf_n2731( .i (n2730), .o (n2731) );
  buffer buf_n2732( .i (n2731), .o (n2732) );
  buffer buf_n2733( .i (n2732), .o (n2733) );
  buffer buf_n2734( .i (n2733), .o (n2734) );
  buffer buf_n2735( .i (n2734), .o (n2735) );
  buffer buf_n2736( .i (n2735), .o (n2736) );
  buffer buf_n2737( .i (n2736), .o (n2737) );
  buffer buf_n2738( .i (n2737), .o (n2738) );
  buffer buf_n2739( .i (n2738), .o (n2739) );
  buffer buf_n2740( .i (n2739), .o (n2740) );
  buffer buf_n336( .i (x47), .o (n336) );
  buffer buf_n337( .i (n336), .o (n337) );
  buffer buf_n338( .i (n337), .o (n338) );
  buffer buf_n339( .i (n338), .o (n339) );
  buffer buf_n340( .i (n339), .o (n340) );
  buffer buf_n341( .i (n340), .o (n341) );
  assign n2741 = ~n1508 & n1525 ;
  buffer buf_n2742( .i (n2741), .o (n2742) );
  buffer buf_n2743( .i (n2742), .o (n2743) );
  assign n2745 = n341 & n2743 ;
  buffer buf_n2746( .i (n2745), .o (n2746) );
  buffer buf_n2747( .i (n2746), .o (n2747) );
  assign n2748 = n2035 | n2670 ;
  assign n2749 = ~n2747 & n2748 ;
  buffer buf_n2750( .i (n2749), .o (n2750) );
  buffer buf_n2751( .i (n2750), .o (n2751) );
  buffer buf_n27( .i (x1), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  buffer buf_n32( .i (n31), .o (n32) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n37( .i (n36), .o (n37) );
  buffer buf_n2133( .i (n2132), .o (n2133) );
  assign n2752 = n37 | n2133 ;
  assign n2753 = n1510 & ~n1527 ;
  buffer buf_n2754( .i (n2753), .o (n2754) );
  buffer buf_n2755( .i (n2754), .o (n2755) );
  buffer buf_n2756( .i (n2755), .o (n2756) );
  buffer buf_n2757( .i (n2756), .o (n2757) );
  buffer buf_n2758( .i (n2757), .o (n2758) );
  assign n2769 = ( n37 & n2133 ) | ( n37 & ~n2758 ) | ( n2133 & ~n2758 ) ;
  assign n2770 = ( n2751 & ~n2752 ) | ( n2751 & n2769 ) | ( ~n2752 & n2769 ) ;
  buffer buf_n2771( .i (n2770), .o (n2771) );
  buffer buf_n2772( .i (n2771), .o (n2772) );
  buffer buf_n2773( .i (n2772), .o (n2773) );
  buffer buf_n2774( .i (n2773), .o (n2774) );
  buffer buf_n2775( .i (n2774), .o (n2775) );
  buffer buf_n2776( .i (n2775), .o (n2776) );
  buffer buf_n2777( .i (n2776), .o (n2777) );
  buffer buf_n2778( .i (n2777), .o (n2778) );
  buffer buf_n2779( .i (n2778), .o (n2779) );
  buffer buf_n2780( .i (n2779), .o (n2780) );
  buffer buf_n2781( .i (n2780), .o (n2781) );
  buffer buf_n2501( .i (n2500), .o (n2501) );
  buffer buf_n2502( .i (n2501), .o (n2502) );
  buffer buf_n2503( .i (n2502), .o (n2503) );
  buffer buf_n2504( .i (n2503), .o (n2504) );
  buffer buf_n2516( .i (n2515), .o (n2516) );
  buffer buf_n1157( .i (n1156), .o (n1157) );
  buffer buf_n1158( .i (n1157), .o (n1158) );
  buffer buf_n1159( .i (n1158), .o (n1159) );
  buffer buf_n2396( .i (n2395), .o (n2396) );
  buffer buf_n2397( .i (n2396), .o (n2397) );
  buffer buf_n2398( .i (n2397), .o (n2398) );
  assign n2782 = ( n1159 & n1169 ) | ( n1159 & n2398 ) | ( n1169 & n2398 ) ;
  assign n2783 = ( n1159 & n2398 ) | ( n1159 & n2485 ) | ( n2398 & n2485 ) ;
  assign n2784 = ( n2687 & n2782 ) | ( n2687 & n2783 ) | ( n2782 & n2783 ) ;
  buffer buf_n2785( .i (n2784), .o (n2785) );
  assign n2787 = n2472 & n2785 ;
  assign n2788 = n2415 & n2787 ;
  buffer buf_n2789( .i (n2788), .o (n2789) );
  assign n2791 = n2516 | n2789 ;
  assign n2792 = n2656 | n2791 ;
  buffer buf_n2793( .i (n2792), .o (n2793) );
  assign n2795 = ~n2504 & n2793 ;
  assign n2796 = n2504 & ~n2793 ;
  assign n2797 = n2795 | n2796 ;
  buffer buf_n2798( .i (n2797), .o (n2798) );
  buffer buf_n2799( .i (n2798), .o (n2799) );
  buffer buf_n2800( .i (n2799), .o (n2800) );
  buffer buf_n2801( .i (n2800), .o (n2801) );
  buffer buf_n2802( .i (n2801), .o (n2802) );
  buffer buf_n1435( .i (x171), .o (n1435) );
  buffer buf_n1436( .i (n1435), .o (n1436) );
  buffer buf_n1449( .i (x172), .o (n1449) );
  buffer buf_n1450( .i (n1449), .o (n1450) );
  assign n2803 = n1436 | n1450 ;
  buffer buf_n2804( .i (n2803), .o (n2804) );
  buffer buf_n2805( .i (n2804), .o (n2805) );
  buffer buf_n2806( .i (n2805), .o (n2806) );
  buffer buf_n2807( .i (n2806), .o (n2807) );
  buffer buf_n2808( .i (n2807), .o (n2808) );
  buffer buf_n2809( .i (n2808), .o (n2809) );
  buffer buf_n2810( .i (n2809), .o (n2810) );
  buffer buf_n2811( .i (n2810), .o (n2811) );
  buffer buf_n2812( .i (n2811), .o (n2812) );
  buffer buf_n2813( .i (n2812), .o (n2813) );
  buffer buf_n2814( .i (n2813), .o (n2814) );
  buffer buf_n2815( .i (n2814), .o (n2815) );
  assign n2822 = n2708 | n2815 ;
  buffer buf_n1437( .i (n1436), .o (n1437) );
  buffer buf_n1438( .i (n1437), .o (n1438) );
  buffer buf_n1439( .i (n1438), .o (n1439) );
  buffer buf_n1440( .i (n1439), .o (n1440) );
  buffer buf_n1441( .i (n1440), .o (n1441) );
  buffer buf_n1442( .i (n1441), .o (n1442) );
  buffer buf_n1443( .i (n1442), .o (n1443) );
  buffer buf_n1444( .i (n1443), .o (n1444) );
  buffer buf_n1445( .i (n1444), .o (n1445) );
  buffer buf_n1446( .i (n1445), .o (n1446) );
  buffer buf_n1451( .i (n1450), .o (n1451) );
  buffer buf_n1452( .i (n1451), .o (n1452) );
  buffer buf_n1453( .i (n1452), .o (n1453) );
  buffer buf_n1454( .i (n1453), .o (n1454) );
  buffer buf_n1455( .i (n1454), .o (n1455) );
  buffer buf_n1456( .i (n1455), .o (n1456) );
  buffer buf_n1457( .i (n1456), .o (n1457) );
  buffer buf_n1458( .i (n1457), .o (n1458) );
  buffer buf_n1459( .i (n1458), .o (n1459) );
  buffer buf_n1460( .i (n1459), .o (n1460) );
  assign n2823 = ~n1446 & n1460 ;
  buffer buf_n2824( .i (n2823), .o (n2824) );
  assign n2833 = ~n2771 & n2824 ;
  buffer buf_n40( .i (x2), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  buffer buf_n44( .i (n43), .o (n44) );
  assign n2834 = n44 & ~n1453 ;
  buffer buf_n148( .i (x21), .o (n148) );
  buffer buf_n149( .i (n148), .o (n149) );
  buffer buf_n150( .i (n149), .o (n150) );
  buffer buf_n151( .i (n150), .o (n151) );
  buffer buf_n152( .i (n151), .o (n152) );
  assign n2835 = n152 & n1453 ;
  assign n2836 = ( n1440 & n2834 ) | ( n1440 & n2835 ) | ( n2834 & n2835 ) ;
  buffer buf_n2837( .i (n2836), .o (n2837) );
  buffer buf_n2838( .i (n2837), .o (n2838) );
  buffer buf_n2839( .i (n2838), .o (n2839) );
  buffer buf_n2840( .i (n2839), .o (n2840) );
  buffer buf_n2841( .i (n2840), .o (n2841) );
  buffer buf_n2842( .i (n2841), .o (n2842) );
  buffer buf_n2843( .i (n2842), .o (n2843) );
  buffer buf_n2844( .i (n2843), .o (n2844) );
  assign n2845 = n2833 | n2844 ;
  assign n2846 = n2822 & ~n2845 ;
  buffer buf_n2847( .i (n2846), .o (n2847) );
  buffer buf_n2848( .i (n2847), .o (n2848) );
  buffer buf_n2849( .i (n2848), .o (n2849) );
  buffer buf_n2850( .i (n2849), .o (n2850) );
  buffer buf_n2851( .i (n2850), .o (n2851) );
  buffer buf_n2852( .i (n2851), .o (n2852) );
  buffer buf_n2853( .i (n2852), .o (n2853) );
  buffer buf_n123( .i (x18), .o (n123) );
  buffer buf_n124( .i (n123), .o (n124) );
  buffer buf_n125( .i (n124), .o (n125) );
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  buffer buf_n129( .i (n128), .o (n129) );
  buffer buf_n2744( .i (n2743), .o (n2744) );
  assign n2854 = n129 & n2744 ;
  buffer buf_n2855( .i (n2854), .o (n2855) );
  buffer buf_n2856( .i (n2669), .o (n2856) );
  assign n2857 = n1903 | n2856 ;
  assign n2858 = ~n2855 & n2857 ;
  buffer buf_n2859( .i (n2858), .o (n2859) );
  buffer buf_n2860( .i (n2859), .o (n2860) );
  buffer buf_n2861( .i (n2860), .o (n2861) );
  buffer buf_n2862( .i (n2861), .o (n2862) );
  buffer buf_n2361( .i (n2360), .o (n2361) );
  buffer buf_n2362( .i (n2361), .o (n2362) );
  buffer buf_n2363( .i (n2362), .o (n2363) );
  buffer buf_n1144( .i (n1143), .o (n1144) );
  buffer buf_n1145( .i (n1144), .o (n1145) );
  buffer buf_n1146( .i (n1145), .o (n1146) );
  buffer buf_n1147( .i (n1146), .o (n1147) );
  buffer buf_n1148( .i (n1147), .o (n1148) );
  buffer buf_n1149( .i (n1148), .o (n1149) );
  buffer buf_n1150( .i (n1149), .o (n1150) );
  buffer buf_n2366( .i (n2365), .o (n2366) );
  buffer buf_n2367( .i (n2366), .o (n2367) );
  buffer buf_n2368( .i (n2367), .o (n2368) );
  buffer buf_n2369( .i (n2368), .o (n2369) );
  buffer buf_n2370( .i (n2369), .o (n2370) );
  buffer buf_n2371( .i (n2370), .o (n2371) );
  buffer buf_n2372( .i (n2371), .o (n2372) );
  assign n2863 = ( n1150 & ~n2372 ) | ( n1150 & n2785 ) | ( ~n2372 & n2785 ) ;
  buffer buf_n2864( .i (n2863), .o (n2864) );
  assign n2865 = n2363 & n2864 ;
  buffer buf_n2759( .i (n2758), .o (n2759) );
  buffer buf_n2760( .i (n2759), .o (n2760) );
  assign n2866 = ( n2363 & n2760 ) | ( n2363 & n2864 ) | ( n2760 & n2864 ) ;
  assign n2867 = ( n2862 & n2865 ) | ( n2862 & ~n2866 ) | ( n2865 & ~n2866 ) ;
  buffer buf_n2868( .i (n2867), .o (n2868) );
  buffer buf_n2869( .i (n2868), .o (n2869) );
  buffer buf_n2870( .i (n2869), .o (n2870) );
  buffer buf_n2871( .i (n2870), .o (n2871) );
  buffer buf_n2872( .i (n2871), .o (n2872) );
  buffer buf_n2873( .i (n2872), .o (n2873) );
  buffer buf_n2874( .i (n2873), .o (n2874) );
  buffer buf_n2875( .i (n2874), .o (n2875) );
  buffer buf_n2876( .i (n2875), .o (n2876) );
  assign n2877 = n1907 | n2668 ;
  buffer buf_n417( .i (x58), .o (n417) );
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  assign n2878 = n422 & n2743 ;
  assign n2879 = n2877 & ~n2878 ;
  buffer buf_n2880( .i (n2879), .o (n2880) );
  buffer buf_n2881( .i (n2880), .o (n2881) );
  buffer buf_n2882( .i (n2881), .o (n2882) );
  buffer buf_n2883( .i (n2882), .o (n2883) );
  buffer buf_n2884( .i (n2883), .o (n2884) );
  buffer buf_n2387( .i (n2386), .o (n2387) );
  buffer buf_n2388( .i (n2387), .o (n2388) );
  buffer buf_n2389( .i (n2388), .o (n2389) );
  buffer buf_n2390( .i (n2389), .o (n2390) );
  buffer buf_n2786( .i (n2785), .o (n2786) );
  assign n2885 = n2390 & ~n2786 ;
  assign n2886 = ( n2390 & n2759 ) | ( n2390 & ~n2786 ) | ( n2759 & ~n2786 ) ;
  assign n2887 = ( n2884 & n2885 ) | ( n2884 & ~n2886 ) | ( n2885 & ~n2886 ) ;
  buffer buf_n2888( .i (n2887), .o (n2888) );
  buffer buf_n2889( .i (n2888), .o (n2889) );
  buffer buf_n2890( .i (n2889), .o (n2890) );
  buffer buf_n2891( .i (n2890), .o (n2891) );
  buffer buf_n2892( .i (n2891), .o (n2892) );
  buffer buf_n2893( .i (n2892), .o (n2893) );
  buffer buf_n2894( .i (n2893), .o (n2894) );
  buffer buf_n2895( .i (n2894), .o (n2895) );
  buffer buf_n2896( .i (n2895), .o (n2896) );
  buffer buf_n2897( .i (n2896), .o (n2897) );
  buffer buf_n351( .i (x49), .o (n351) );
  buffer buf_n352( .i (n351), .o (n352) );
  buffer buf_n353( .i (n352), .o (n353) );
  assign n2898 = n353 & n1525 ;
  assign n2899 = ~n1509 & n2898 ;
  buffer buf_n2900( .i (n2899), .o (n2900) );
  assign n2905 = n1528 & ~n2900 ;
  buffer buf_n2906( .i (n2905), .o (n2906) );
  buffer buf_n2907( .i (n2906), .o (n2907) );
  buffer buf_n2908( .i (n2907), .o (n2908) );
  buffer buf_n2901( .i (n2900), .o (n2901) );
  buffer buf_n2902( .i (n2901), .o (n2902) );
  assign n2909 = ( n1936 & ~n2902 ) | ( n1936 & n2906 ) | ( ~n2902 & n2906 ) ;
  buffer buf_n2910( .i (n2909), .o (n2910) );
  assign n2911 = ( ~n1515 & n2908 ) | ( ~n1515 & n2910 ) | ( n2908 & n2910 ) ;
  buffer buf_n2912( .i (n2911), .o (n2912) );
  buffer buf_n2913( .i (n2912), .o (n2913) );
  buffer buf_n2914( .i (n2913), .o (n2914) );
  buffer buf_n2407( .i (n2406), .o (n2407) );
  buffer buf_n2408( .i (n2407), .o (n2408) );
  buffer buf_n2409( .i (n2408), .o (n2409) );
  buffer buf_n1170( .i (n1169), .o (n1170) );
  buffer buf_n2486( .i (n2485), .o (n2486) );
  assign n2915 = ( n1170 & n2486 ) | ( n1170 & n2687 ) | ( n2486 & n2687 ) ;
  buffer buf_n2916( .i (n2915), .o (n2916) );
  assign n2917 = n2409 & n2916 ;
  buffer buf_n2918( .i (n2917), .o (n2918) );
  assign n2919 = n2409 | n2916 ;
  buffer buf_n2920( .i (n2919), .o (n2920) );
  assign n2921 = ~n2918 & n2920 ;
  buffer buf_n2903( .i (n2902), .o (n2903) );
  buffer buf_n2904( .i (n2903), .o (n2904) );
  assign n2922 = ( n1515 & ~n2904 ) | ( n1515 & n2910 ) | ( ~n2904 & n2910 ) ;
  buffer buf_n2923( .i (n2922), .o (n2923) );
  buffer buf_n2924( .i (n2923), .o (n2924) );
  buffer buf_n2925( .i (n2924), .o (n2925) );
  assign n2926 = ( n2914 & ~n2921 ) | ( n2914 & n2925 ) | ( ~n2921 & n2925 ) ;
  buffer buf_n2927( .i (n2926), .o (n2927) );
  buffer buf_n2928( .i (n2927), .o (n2928) );
  buffer buf_n2929( .i (n2928), .o (n2929) );
  buffer buf_n2930( .i (n2929), .o (n2930) );
  buffer buf_n2931( .i (n2930), .o (n2931) );
  buffer buf_n2932( .i (n2931), .o (n2932) );
  buffer buf_n2933( .i (n2932), .o (n2933) );
  buffer buf_n2934( .i (n2933), .o (n2934) );
  buffer buf_n2935( .i (n2934), .o (n2935) );
  buffer buf_n1462( .i (x173), .o (n1462) );
  buffer buf_n1463( .i (n1462), .o (n1463) );
  buffer buf_n1464( .i (n1463), .o (n1464) );
  buffer buf_n1465( .i (n1464), .o (n1465) );
  buffer buf_n1466( .i (n1465), .o (n1466) );
  buffer buf_n1467( .i (n1466), .o (n1467) );
  buffer buf_n1468( .i (n1467), .o (n1468) );
  buffer buf_n1469( .i (n1468), .o (n1469) );
  buffer buf_n1485( .i (x174), .o (n1485) );
  buffer buf_n1486( .i (n1485), .o (n1486) );
  buffer buf_n1487( .i (n1486), .o (n1487) );
  buffer buf_n1488( .i (n1487), .o (n1488) );
  buffer buf_n1489( .i (n1488), .o (n1489) );
  buffer buf_n1490( .i (n1489), .o (n1490) );
  buffer buf_n1491( .i (n1490), .o (n1491) );
  buffer buf_n1492( .i (n1491), .o (n1492) );
  assign n2936 = n1469 | n1492 ;
  buffer buf_n2937( .i (n2936), .o (n2937) );
  buffer buf_n2938( .i (n2937), .o (n2938) );
  buffer buf_n2939( .i (n2938), .o (n2939) );
  buffer buf_n2940( .i (n2939), .o (n2940) );
  buffer buf_n2941( .i (n2940), .o (n2941) );
  buffer buf_n2942( .i (n2941), .o (n2942) );
  buffer buf_n2943( .i (n2942), .o (n2943) );
  assign n2947 = n2709 & ~n2943 ;
  assign n2948 = n1463 & ~n1486 ;
  buffer buf_n2949( .i (n2948), .o (n2949) );
  buffer buf_n2950( .i (n2949), .o (n2950) );
  buffer buf_n2951( .i (n2950), .o (n2951) );
  buffer buf_n2952( .i (n2951), .o (n2952) );
  buffer buf_n2953( .i (n2952), .o (n2953) );
  buffer buf_n2954( .i (n2953), .o (n2954) );
  buffer buf_n2955( .i (n2954), .o (n2955) );
  buffer buf_n2956( .i (n2955), .o (n2956) );
  buffer buf_n2957( .i (n2956), .o (n2957) );
  buffer buf_n2958( .i (n2957), .o (n2958) );
  buffer buf_n2959( .i (n2958), .o (n2959) );
  buffer buf_n2960( .i (n2959), .o (n2960) );
  assign n2966 = n2772 & n2960 ;
  buffer buf_n153( .i (n152), .o (n153) );
  assign n2967 = ~n153 & n1467 ;
  buffer buf_n45( .i (n44), .o (n45) );
  assign n2968 = n45 | n1467 ;
  assign n2969 = ( n1491 & n2967 ) | ( n1491 & ~n2968 ) | ( n2967 & ~n2968 ) ;
  buffer buf_n2970( .i (n2969), .o (n2970) );
  buffer buf_n2971( .i (n2970), .o (n2971) );
  buffer buf_n2972( .i (n2971), .o (n2972) );
  buffer buf_n2973( .i (n2972), .o (n2973) );
  buffer buf_n2974( .i (n2973), .o (n2974) );
  buffer buf_n2975( .i (n2974), .o (n2975) );
  buffer buf_n2976( .i (n2975), .o (n2976) );
  buffer buf_n2977( .i (n2976), .o (n2977) );
  assign n2978 = n2966 | n2977 ;
  assign n2979 = n2947 | n2978 ;
  buffer buf_n2980( .i (n2979), .o (n2980) );
  buffer buf_n2981( .i (n2980), .o (n2981) );
  buffer buf_n2982( .i (n2981), .o (n2982) );
  buffer buf_n2983( .i (n2982), .o (n2983) );
  buffer buf_n2984( .i (n2983), .o (n2984) );
  buffer buf_n2985( .i (n2984), .o (n2985) );
  buffer buf_n370( .i (x52), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  assign n2986 = n376 & n2744 ;
  buffer buf_n2987( .i (n2986), .o (n2987) );
  assign n2988 = n2002 | n2856 ;
  assign n2989 = ~n2987 & n2988 ;
  buffer buf_n2990( .i (n2989), .o (n2990) );
  buffer buf_n2991( .i (n2990), .o (n2991) );
  buffer buf_n2992( .i (n2991), .o (n2992) );
  buffer buf_n2993( .i (n2992), .o (n2993) );
  buffer buf_n2994( .i (n2993), .o (n2994) );
  buffer buf_n2286( .i (n2285), .o (n2286) );
  buffer buf_n2287( .i (n2286), .o (n2287) );
  buffer buf_n2288( .i (n2287), .o (n2288) );
  buffer buf_n1012( .i (n1011), .o (n1012) );
  buffer buf_n1013( .i (n1012), .o (n1013) );
  buffer buf_n1014( .i (n1013), .o (n1014) );
  buffer buf_n1015( .i (n1014), .o (n1015) );
  buffer buf_n1016( .i (n1015), .o (n1016) );
  buffer buf_n2095( .i (n2094), .o (n2095) );
  buffer buf_n2096( .i (n2095), .o (n2096) );
  buffer buf_n2097( .i (n2096), .o (n2097) );
  buffer buf_n2098( .i (n2097), .o (n2098) );
  buffer buf_n2099( .i (n2098), .o (n2099) );
  buffer buf_n1001( .i (n1000), .o (n1001) );
  assign n2995 = ( n34 & n1001 ) | ( n34 & n2124 ) | ( n1001 & n2124 ) ;
  buffer buf_n2996( .i (n2995), .o (n2996) );
  buffer buf_n1023( .i (n1022), .o (n1023) );
  buffer buf_n1024( .i (n1023), .o (n1024) );
  buffer buf_n1025( .i (n1024), .o (n1025) );
  buffer buf_n1026( .i (n1025), .o (n1026) );
  buffer buf_n1036( .i (n1035), .o (n1036) );
  buffer buf_n2140( .i (n2139), .o (n2140) );
  buffer buf_n2141( .i (n2140), .o (n2141) );
  buffer buf_n2142( .i (n2141), .o (n2142) );
  buffer buf_n2143( .i (n2142), .o (n2143) );
  assign n2999 = ( n1026 & n1036 ) | ( n1026 & n2143 ) | ( n1036 & n2143 ) ;
  buffer buf_n2076( .i (n2075), .o (n2076) );
  assign n3000 = ( n1026 & n2076 ) | ( n1026 & n2143 ) | ( n2076 & n2143 ) ;
  assign n3001 = ( n2996 & n2999 ) | ( n2996 & n3000 ) | ( n2999 & n3000 ) ;
  buffer buf_n3002( .i (n3001), .o (n3002) );
  assign n3004 = ( n1016 & n2099 ) | ( n1016 & n3002 ) | ( n2099 & n3002 ) ;
  buffer buf_n3005( .i (n3004), .o (n3005) );
  assign n3006 = n2288 & n3005 ;
  buffer buf_n2761( .i (n2760), .o (n2761) );
  assign n3007 = ( n2288 & n2761 ) | ( n2288 & n3005 ) | ( n2761 & n3005 ) ;
  assign n3008 = ( n2994 & n3006 ) | ( n2994 & ~n3007 ) | ( n3006 & ~n3007 ) ;
  buffer buf_n3009( .i (n3008), .o (n3009) );
  buffer buf_n3010( .i (n3009), .o (n3010) );
  buffer buf_n3011( .i (n3010), .o (n3011) );
  buffer buf_n3012( .i (n3011), .o (n3012) );
  buffer buf_n3013( .i (n3012), .o (n3013) );
  buffer buf_n3014( .i (n3013), .o (n3014) );
  buffer buf_n3015( .i (n3014), .o (n3015) );
  buffer buf_n3016( .i (n3015), .o (n3016) );
  buffer buf_n402( .i (x56), .o (n402) );
  buffer buf_n403( .i (n402), .o (n403) );
  buffer buf_n404( .i (n403), .o (n404) );
  buffer buf_n405( .i (n404), .o (n405) );
  buffer buf_n406( .i (n405), .o (n406) );
  assign n3017 = n406 & ~n1510 ;
  buffer buf_n3018( .i (n3017), .o (n3018) );
  buffer buf_n3019( .i (n3018), .o (n3019) );
  assign n3020 = n1530 & ~n3019 ;
  assign n3021 = n2045 & ~n2856 ;
  assign n3022 = n3020 | n3021 ;
  buffer buf_n3023( .i (n3022), .o (n3023) );
  buffer buf_n3024( .i (n3023), .o (n3024) );
  buffer buf_n3025( .i (n3024), .o (n3025) );
  buffer buf_n3026( .i (n3025), .o (n3026) );
  buffer buf_n2114( .i (n2113), .o (n2114) );
  buffer buf_n2115( .i (n2114), .o (n2115) );
  buffer buf_n2116( .i (n2115), .o (n2116) );
  buffer buf_n3003( .i (n3002), .o (n3003) );
  assign n3027 = n2116 & ~n3003 ;
  buffer buf_n1518( .i (n1517), .o (n1518) );
  assign n3028 = ( n1518 & n2116 ) | ( n1518 & ~n3003 ) | ( n2116 & ~n3003 ) ;
  assign n3029 = ( n3026 & ~n3027 ) | ( n3026 & n3028 ) | ( ~n3027 & n3028 ) ;
  buffer buf_n3030( .i (n3029), .o (n3030) );
  buffer buf_n3031( .i (n3030), .o (n3031) );
  buffer buf_n3032( .i (n3031), .o (n3032) );
  buffer buf_n3033( .i (n3032), .o (n3033) );
  buffer buf_n3034( .i (n3033), .o (n3034) );
  buffer buf_n3035( .i (n3034), .o (n3035) );
  buffer buf_n3036( .i (n3035), .o (n3036) );
  buffer buf_n3037( .i (n3036), .o (n3037) );
  buffer buf_n3038( .i (n3037), .o (n3038) );
  assign n3039 = n1990 | n2856 ;
  buffer buf_n394( .i (x55), .o (n394) );
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n396( .i (n395), .o (n396) );
  buffer buf_n397( .i (n396), .o (n397) );
  buffer buf_n398( .i (n397), .o (n398) );
  buffer buf_n399( .i (n398), .o (n399) );
  buffer buf_n400( .i (n399), .o (n400) );
  assign n3040 = n400 & n2744 ;
  buffer buf_n3041( .i (n3040), .o (n3041) );
  assign n3042 = n3039 & ~n3041 ;
  buffer buf_n3043( .i (n3042), .o (n3043) );
  buffer buf_n3044( .i (n3043), .o (n3044) );
  buffer buf_n3045( .i (n3044), .o (n3045) );
  buffer buf_n2157( .i (n2156), .o (n2157) );
  buffer buf_n2158( .i (n2157), .o (n2158) );
  buffer buf_n1037( .i (n1036), .o (n1037) );
  buffer buf_n2077( .i (n2076), .o (n2077) );
  assign n3046 = ( n1037 & n2077 ) | ( n1037 & n2996 ) | ( n2077 & n2996 ) ;
  buffer buf_n3047( .i (n3046), .o (n3047) );
  assign n3048 = n2158 & n3047 ;
  assign n3049 = ( n2158 & n2759 ) | ( n2158 & n3047 ) | ( n2759 & n3047 ) ;
  assign n3050 = ( n3045 & n3048 ) | ( n3045 & ~n3049 ) | ( n3048 & ~n3049 ) ;
  buffer buf_n3051( .i (n3050), .o (n3051) );
  buffer buf_n3052( .i (n3051), .o (n3052) );
  buffer buf_n3053( .i (n3052), .o (n3053) );
  buffer buf_n3054( .i (n3053), .o (n3054) );
  buffer buf_n3055( .i (n3054), .o (n3055) );
  buffer buf_n3056( .i (n3055), .o (n3056) );
  buffer buf_n3057( .i (n3056), .o (n3057) );
  buffer buf_n3058( .i (n3057), .o (n3058) );
  buffer buf_n3059( .i (n3058), .o (n3059) );
  buffer buf_n3060( .i (n3059), .o (n3060) );
  assign n3061 = ( n1531 & n1969 ) | ( n1531 & ~n2756 ) | ( n1969 & ~n2756 ) ;
  buffer buf_n386( .i (x54), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  buffer buf_n390( .i (n389), .o (n390) );
  buffer buf_n391( .i (n390), .o (n391) );
  buffer buf_n392( .i (n391), .o (n392) );
  assign n3062 = n392 & n2744 ;
  buffer buf_n3063( .i (n3062), .o (n3063) );
  buffer buf_n3064( .i (n3063), .o (n3064) );
  assign n3065 = n3061 & ~n3064 ;
  buffer buf_n3066( .i (n3065), .o (n3066) );
  buffer buf_n3067( .i (n3066), .o (n3067) );
  buffer buf_n2088( .i (n2087), .o (n2088) );
  buffer buf_n2997( .i (n2996), .o (n2997) );
  buffer buf_n2998( .i (n2997), .o (n2998) );
  assign n3068 = n2088 & ~n2998 ;
  assign n3069 = ( n1517 & n2088 ) | ( n1517 & ~n2998 ) | ( n2088 & ~n2998 ) ;
  assign n3070 = ( n3067 & ~n3068 ) | ( n3067 & n3069 ) | ( ~n3068 & n3069 ) ;
  buffer buf_n3071( .i (n3070), .o (n3071) );
  buffer buf_n3072( .i (n3071), .o (n3072) );
  buffer buf_n3073( .i (n3072), .o (n3073) );
  buffer buf_n3074( .i (n3073), .o (n3074) );
  buffer buf_n3075( .i (n3074), .o (n3075) );
  buffer buf_n3076( .i (n3075), .o (n3076) );
  buffer buf_n3077( .i (n3076), .o (n3077) );
  buffer buf_n3078( .i (n3077), .o (n3078) );
  buffer buf_n3079( .i (n3078), .o (n3079) );
  buffer buf_n3080( .i (n3079), .o (n3080) );
  buffer buf_n986( .i (x132), .o (n986) );
  buffer buf_n987( .i (n986), .o (n987) );
  buffer buf_n988( .i (n987), .o (n988) );
  buffer buf_n989( .i (n988), .o (n989) );
  buffer buf_n990( .i (n989), .o (n990) );
  assign n3081 = ( ~n806 & n862 ) | ( ~n806 & n893 ) | ( n862 & n893 ) ;
  assign n3082 = ( n806 & n862 ) | ( n806 & n893 ) | ( n862 & n893 ) ;
  assign n3083 = ( n807 & n3081 ) | ( n807 & ~n3082 ) | ( n3081 & ~n3082 ) ;
  buffer buf_n3084( .i (n3083), .o (n3084) );
  assign n3085 = ( ~n956 & n990 ) | ( ~n956 & n3084 ) | ( n990 & n3084 ) ;
  assign n3086 = ( n956 & n990 ) | ( n956 & n3084 ) | ( n990 & n3084 ) ;
  assign n3087 = ( n957 & n3085 ) | ( n957 & ~n3086 ) | ( n3085 & ~n3086 ) ;
  buffer buf_n3088( .i (n3087), .o (n3088) );
  buffer buf_n818( .i (n817), .o (n818) );
  buffer buf_n819( .i (n818), .o (n819) );
  buffer buf_n820( .i (n819), .o (n820) );
  buffer buf_n821( .i (n820), .o (n821) );
  buffer buf_n832( .i (n831), .o (n832) );
  assign n3089 = ( ~n775 & n841 ) | ( ~n775 & n923 ) | ( n841 & n923 ) ;
  assign n3090 = ( n775 & n841 ) | ( n775 & n923 ) | ( n841 & n923 ) ;
  assign n3091 = ( n776 & n3089 ) | ( n776 & ~n3090 ) | ( n3089 & ~n3090 ) ;
  buffer buf_n3092( .i (n3091), .o (n3092) );
  assign n3094 = ( ~n820 & n832 ) | ( ~n820 & n3092 ) | ( n832 & n3092 ) ;
  assign n3095 = ( n820 & n832 ) | ( n820 & n3092 ) | ( n832 & n3092 ) ;
  assign n3096 = ( n821 & n3094 ) | ( n821 & ~n3095 ) | ( n3094 & ~n3095 ) ;
  buffer buf_n3097( .i (n3096), .o (n3097) );
  assign n3098 = ( ~n852 & n3088 ) | ( ~n852 & n3097 ) | ( n3088 & n3097 ) ;
  assign n3099 = ( n852 & n3088 ) | ( n852 & n3097 ) | ( n3088 & n3097 ) ;
  assign n3100 = ~n3098 & n3099 ;
  buffer buf_n3101( .i (n3100), .o (n3101) );
  assign n3102 = n854 | n2553 ;
  assign n3103 = ~n3101 & n3102 ;
  buffer buf_n3104( .i (n3103), .o (n3104) );
  buffer buf_n3105( .i (n3104), .o (n3105) );
  buffer buf_n3106( .i (n3105), .o (n3106) );
  buffer buf_n3107( .i (n3106), .o (n3107) );
  buffer buf_n3108( .i (n3107), .o (n3108) );
  buffer buf_n3109( .i (n3108), .o (n3109) );
  buffer buf_n3110( .i (n3109), .o (n3110) );
  buffer buf_n3111( .i (n3110), .o (n3111) );
  buffer buf_n3112( .i (n3111), .o (n3112) );
  buffer buf_n3113( .i (n3112), .o (n3113) );
  buffer buf_n3114( .i (n3113), .o (n3114) );
  buffer buf_n3115( .i (n3114), .o (n3115) );
  buffer buf_n2078( .i (n2077), .o (n2078) );
  assign n3116 = ( n2077 & n2097 ) | ( n2077 & ~n2126 ) | ( n2097 & ~n2126 ) ;
  assign n3117 = ( n2077 & ~n2097 ) | ( n2077 & n2126 ) | ( ~n2097 & n2126 ) ;
  assign n3118 = ( ~n2078 & n3116 ) | ( ~n2078 & n3117 ) | ( n3116 & n3117 ) ;
  buffer buf_n3119( .i (n3118), .o (n3119) );
  buffer buf_n3120( .i (n3119), .o (n3120) );
  buffer buf_n3121( .i (n3120), .o (n3121) );
  buffer buf_n746( .i (x111), .o (n746) );
  buffer buf_n747( .i (n746), .o (n747) );
  assign n3122 = ( n634 & n747 ) | ( n634 & n2201 ) | ( n747 & n2201 ) ;
  buffer buf_n3123( .i (n856), .o (n3123) );
  assign n3124 = ( n634 & n747 ) | ( n634 & ~n3123 ) | ( n747 & ~n3123 ) ;
  assign n3125 = n3122 & ~n3124 ;
  buffer buf_n744( .i (n743), .o (n744) );
  assign n3126 = n629 | n744 ;
  buffer buf_n3127( .i (n628), .o (n3127) );
  assign n3128 = ( n744 & n2202 ) | ( n744 & n3127 ) | ( n2202 & n3127 ) ;
  assign n3129 = ( n3125 & n3126 ) | ( n3125 & ~n3128 ) | ( n3126 & ~n3128 ) ;
  buffer buf_n3130( .i (n3129), .o (n3130) );
  buffer buf_n3131( .i (n3130), .o (n3131) );
  buffer buf_n3132( .i (n3131), .o (n3132) );
  buffer buf_n3133( .i (n3132), .o (n3133) );
  buffer buf_n3134( .i (n3133), .o (n3134) );
  buffer buf_n3135( .i (n3134), .o (n3135) );
  buffer buf_n3136( .i (n3135), .o (n3136) );
  buffer buf_n3137( .i (n3136), .o (n3137) );
  buffer buf_n3138( .i (n3137), .o (n3138) );
  buffer buf_n2144( .i (n2143), .o (n2144) );
  buffer buf_n2145( .i (n2144), .o (n2145) );
  buffer buf_n2146( .i (n2145), .o (n2146) );
  buffer buf_n2206( .i (n2205), .o (n2206) );
  buffer buf_n2207( .i (n2206), .o (n2207) );
  buffer buf_n2208( .i (n2207), .o (n2208) );
  buffer buf_n2209( .i (n2208), .o (n2209) );
  buffer buf_n2210( .i (n2209), .o (n2210) );
  buffer buf_n2170( .i (n2169), .o (n2170) );
  buffer buf_n2171( .i (n2170), .o (n2171) );
  buffer buf_n2172( .i (n2171), .o (n2172) );
  buffer buf_n2248( .i (n2247), .o (n2248) );
  buffer buf_n2249( .i (n2248), .o (n2249) );
  buffer buf_n2250( .i (n2249), .o (n2250) );
  assign n3139 = ( ~n2171 & n2250 ) | ( ~n2171 & n2296 ) | ( n2250 & n2296 ) ;
  assign n3140 = ( n2171 & n2250 ) | ( n2171 & n2296 ) | ( n2250 & n2296 ) ;
  assign n3141 = ( n2172 & n3139 ) | ( n2172 & ~n3140 ) | ( n3139 & ~n3140 ) ;
  buffer buf_n3142( .i (n3141), .o (n3142) );
  assign n3143 = ( ~n2145 & n2210 ) | ( ~n2145 & n3142 ) | ( n2210 & n3142 ) ;
  assign n3144 = ( n2145 & n2210 ) | ( n2145 & n3142 ) | ( n2210 & n3142 ) ;
  assign n3145 = ( n2146 & n3143 ) | ( n2146 & ~n3144 ) | ( n3143 & ~n3144 ) ;
  buffer buf_n3146( .i (n3145), .o (n3146) );
  assign n3147 = ( ~n3120 & n3138 ) | ( ~n3120 & n3146 ) | ( n3138 & n3146 ) ;
  assign n3148 = ( n3120 & n3138 ) | ( n3120 & n3146 ) | ( n3138 & n3146 ) ;
  assign n3149 = ( n3121 & n3147 ) | ( n3121 & ~n3148 ) | ( n3147 & ~n3148 ) ;
  buffer buf_n3150( .i (n3149), .o (n3150) );
  buffer buf_n3151( .i (n3150), .o (n3151) );
  buffer buf_n3152( .i (n3151), .o (n3152) );
  buffer buf_n3153( .i (n3152), .o (n3153) );
  buffer buf_n3154( .i (n3153), .o (n3154) );
  buffer buf_n3155( .i (n3154), .o (n3155) );
  buffer buf_n3156( .i (n3155), .o (n3156) );
  buffer buf_n3157( .i (n3156), .o (n3157) );
  buffer buf_n2150( .i (n2149), .o (n2150) );
  assign n3158 = ~n2112 & n2150 ;
  assign n3159 = n1001 | n2080 ;
  assign n3160 = ~n2155 & n3159 ;
  assign n3161 = n3158 | n3160 ;
  assign n3162 = ( ~n37 & n2133 ) | ( ~n37 & n3161 ) | ( n2133 & n3161 ) ;
  buffer buf_n3163( .i (n3162), .o (n3163) );
  buffer buf_n38( .i (n37), .o (n38) );
  buffer buf_n2134( .i (n2133), .o (n2134) );
  assign n3164 = ~n2218 & n2309 ;
  buffer buf_n1002( .i (n1001), .o (n1002) );
  buffer buf_n2083( .i (n2082), .o (n2083) );
  assign n3165 = n1002 & n2083 ;
  buffer buf_n3166( .i (n3165), .o (n3166) );
  assign n3167 = n3164 | n3166 ;
  assign n3168 = ( n38 & ~n2134 ) | ( n38 & n3167 ) | ( ~n2134 & n3167 ) ;
  assign n3169 = n3163 | n3168 ;
  buffer buf_n2236( .i (n2235), .o (n2236) );
  buffer buf_n2237( .i (n2236), .o (n2237) );
  buffer buf_n2238( .i (n2237), .o (n2238) );
  assign n3170 = ~n2158 & n2243 ;
  assign n3171 = ( ~n2238 & n2608 ) | ( ~n2238 & n3170 ) | ( n2608 & n3170 ) ;
  assign n3172 = n3169 | n3171 ;
  buffer buf_n3173( .i (n3172), .o (n3173) );
  buffer buf_n3174( .i (n3173), .o (n3174) );
  buffer buf_n3175( .i (n3174), .o (n3175) );
  buffer buf_n2321( .i (n2320), .o (n2321) );
  buffer buf_n2239( .i (n2238), .o (n2239) );
  assign n3176 = n2239 & ~n2609 ;
  buffer buf_n3177( .i (n3176), .o (n3177) );
  buffer buf_n2211( .i (n2210), .o (n2211) );
  buffer buf_n2212( .i (n2211), .o (n2212) );
  buffer buf_n2213( .i (n2212), .o (n2213) );
  buffer buf_n2214( .i (n2213), .o (n2214) );
  buffer buf_n1060( .i (n1059), .o (n1060) );
  assign n3178 = ( n1011 & n1060 ) | ( n1011 & n2170 ) | ( n1060 & n2170 ) ;
  buffer buf_n3179( .i (n3178), .o (n3179) );
  buffer buf_n3180( .i (n3179), .o (n3180) );
  buffer buf_n3181( .i (n3180), .o (n3181) );
  buffer buf_n3182( .i (n3181), .o (n3182) );
  assign n3183 = ( n1060 & n2094 ) | ( n1060 & n2170 ) | ( n2094 & n2170 ) ;
  buffer buf_n3184( .i (n3183), .o (n3184) );
  buffer buf_n3185( .i (n3184), .o (n3185) );
  buffer buf_n3186( .i (n3185), .o (n3186) );
  buffer buf_n3187( .i (n3186), .o (n3187) );
  assign n3188 = ( n3002 & n3182 ) | ( n3002 & n3187 ) | ( n3182 & n3187 ) ;
  buffer buf_n3189( .i (n3188), .o (n3189) );
  buffer buf_n3190( .i (n3189), .o (n3190) );
  buffer buf_n2630( .i (n2629), .o (n2630) );
  assign n3192 = n2630 & n3189 ;
  assign n3193 = ( ~n2214 & n3190 ) | ( ~n2214 & n3192 ) | ( n3190 & n3192 ) ;
  assign n3194 = n3177 & ~n3193 ;
  assign n3195 = n2321 | n3194 ;
  assign n3196 = n3175 | n3195 ;
  buffer buf_n3197( .i (n3196), .o (n3197) );
  buffer buf_n3198( .i (n3197), .o (n3198) );
  buffer buf_n3199( .i (n3198), .o (n3199) );
  buffer buf_n3200( .i (n3199), .o (n3200) );
  buffer buf_n3201( .i (n3200), .o (n3201) );
  buffer buf_n2693( .i (n2692), .o (n2693) );
  buffer buf_n2694( .i (n2693), .o (n2694) );
  buffer buf_n2695( .i (n2694), .o (n2695) );
  buffer buf_n2696( .i (n2695), .o (n2696) );
  buffer buf_n2697( .i (n2696), .o (n2697) );
  buffer buf_n2698( .i (n2697), .o (n2698) );
  buffer buf_n2699( .i (n2698), .o (n2699) );
  buffer buf_n2700( .i (n2699), .o (n2700) );
  assign n3202 = n2530 & n2700 ;
  buffer buf_n3203( .i (n3202), .o (n3203) );
  buffer buf_n3204( .i (n3203), .o (n3204) );
  buffer buf_n3205( .i (n3204), .o (n3205) );
  buffer buf_n3206( .i (n3205), .o (n3206) );
  buffer buf_n1314( .i (x157), .o (n1314) );
  buffer buf_n1315( .i (n1314), .o (n1315) );
  buffer buf_n1316( .i (n1315), .o (n1316) );
  buffer buf_n1317( .i (n1316), .o (n1317) );
  buffer buf_n1318( .i (n1317), .o (n1318) );
  buffer buf_n1320( .i (x158), .o (n1320) );
  buffer buf_n1321( .i (n1320), .o (n1321) );
  buffer buf_n1322( .i (n1321), .o (n1322) );
  assign n3207 = n457 & ~n1322 ;
  buffer buf_n3208( .i (n3207), .o (n3208) );
  assign n3209 = ~n1318 & n3208 ;
  buffer buf_n3210( .i (n3209), .o (n3210) );
  buffer buf_n3211( .i (n3210), .o (n3211) );
  buffer buf_n3212( .i (n3211), .o (n3212) );
  buffer buf_n3213( .i (n3212), .o (n3213) );
  buffer buf_n3214( .i (n3213), .o (n3214) );
  buffer buf_n3215( .i (n3214), .o (n3215) );
  buffer buf_n3216( .i (n3215), .o (n3216) );
  buffer buf_n3217( .i (n3216), .o (n3217) );
  buffer buf_n3218( .i (n3217), .o (n3218) );
  buffer buf_n3219( .i (n3218), .o (n3219) );
  assign n3225 = ~n2709 & n3219 ;
  assign n3226 = n1318 & n3208 ;
  buffer buf_n3227( .i (n3226), .o (n3227) );
  buffer buf_n3228( .i (n3227), .o (n3228) );
  buffer buf_n3229( .i (n3228), .o (n3229) );
  buffer buf_n3230( .i (n3229), .o (n3230) );
  buffer buf_n3231( .i (n3230), .o (n3231) );
  buffer buf_n3232( .i (n3231), .o (n3232) );
  buffer buf_n3233( .i (n3232), .o (n3233) );
  buffer buf_n3234( .i (n3233), .o (n3234) );
  buffer buf_n3235( .i (n3234), .o (n3235) );
  assign n3243 = ~n2772 & n3235 ;
  assign n3244 = n457 & n1322 ;
  buffer buf_n3245( .i (n3244), .o (n3245) );
  buffer buf_n3246( .i (n3245), .o (n3246) );
  buffer buf_n574( .i (x80), .o (n574) );
  buffer buf_n575( .i (n574), .o (n575) );
  buffer buf_n576( .i (n575), .o (n576) );
  buffer buf_n577( .i (n576), .o (n577) );
  buffer buf_n578( .i (n577), .o (n578) );
  assign n3247 = n578 & n1318 ;
  buffer buf_n568( .i (x79), .o (n568) );
  buffer buf_n569( .i (n568), .o (n569) );
  buffer buf_n570( .i (n569), .o (n570) );
  buffer buf_n571( .i (n570), .o (n571) );
  buffer buf_n572( .i (n571), .o (n572) );
  assign n3248 = n572 & ~n1318 ;
  assign n3249 = ( n3246 & n3247 ) | ( n3246 & n3248 ) | ( n3247 & n3248 ) ;
  buffer buf_n3250( .i (n3249), .o (n3250) );
  buffer buf_n3251( .i (n3250), .o (n3251) );
  buffer buf_n3252( .i (n3251), .o (n3252) );
  buffer buf_n3253( .i (n3252), .o (n3253) );
  buffer buf_n3254( .i (n3253), .o (n3254) );
  buffer buf_n3255( .i (n3254), .o (n3255) );
  buffer buf_n3256( .i (n3255), .o (n3256) );
  buffer buf_n3257( .i (n3256), .o (n3257) );
  buffer buf_n3258( .i (n3257), .o (n3258) );
  assign n3259 = n3243 | n3258 ;
  assign n3260 = n3225 | n3259 ;
  buffer buf_n3261( .i (n3260), .o (n3261) );
  buffer buf_n3262( .i (n3261), .o (n3262) );
  buffer buf_n3263( .i (n3262), .o (n3263) );
  buffer buf_n3264( .i (n3263), .o (n3264) );
  buffer buf_n3265( .i (n3264), .o (n3265) );
  buffer buf_n3266( .i (n3265), .o (n3266) );
  buffer buf_n1324( .i (x159), .o (n1324) );
  buffer buf_n1325( .i (n1324), .o (n1325) );
  buffer buf_n1326( .i (n1325), .o (n1326) );
  buffer buf_n1327( .i (n1326), .o (n1327) );
  buffer buf_n1330( .i (x160), .o (n1330) );
  buffer buf_n1331( .i (n1330), .o (n1331) );
  assign n3267 = n456 & ~n1331 ;
  buffer buf_n3268( .i (n3267), .o (n3268) );
  assign n3269 = ~n1327 & n3268 ;
  buffer buf_n3270( .i (n3269), .o (n3270) );
  buffer buf_n3271( .i (n3270), .o (n3271) );
  buffer buf_n3272( .i (n3271), .o (n3272) );
  buffer buf_n3273( .i (n3272), .o (n3273) );
  buffer buf_n3274( .i (n3273), .o (n3274) );
  buffer buf_n3275( .i (n3274), .o (n3275) );
  buffer buf_n3276( .i (n3275), .o (n3276) );
  buffer buf_n3277( .i (n3276), .o (n3277) );
  buffer buf_n3278( .i (n3277), .o (n3278) );
  buffer buf_n3279( .i (n3278), .o (n3279) );
  buffer buf_n3280( .i (n3279), .o (n3280) );
  assign n3286 = ~n2709 & n3280 ;
  assign n3287 = n1327 & n3268 ;
  buffer buf_n3288( .i (n3287), .o (n3288) );
  buffer buf_n3289( .i (n3288), .o (n3289) );
  buffer buf_n3290( .i (n3289), .o (n3290) );
  buffer buf_n3291( .i (n3290), .o (n3291) );
  buffer buf_n3292( .i (n3291), .o (n3292) );
  buffer buf_n3293( .i (n3292), .o (n3293) );
  buffer buf_n3294( .i (n3293), .o (n3294) );
  buffer buf_n3295( .i (n3294), .o (n3295) );
  buffer buf_n3296( .i (n3295), .o (n3296) );
  buffer buf_n3297( .i (n3296), .o (n3297) );
  assign n3305 = ~n2772 & n3297 ;
  assign n3306 = n456 & n1331 ;
  buffer buf_n3307( .i (n3306), .o (n3307) );
  buffer buf_n3308( .i (n3307), .o (n3308) );
  buffer buf_n3309( .i (n3308), .o (n3309) );
  buffer buf_n1328( .i (n1327), .o (n1328) );
  assign n3310 = n578 & n1328 ;
  assign n3311 = n572 & ~n1328 ;
  assign n3312 = ( n3309 & n3310 ) | ( n3309 & n3311 ) | ( n3310 & n3311 ) ;
  buffer buf_n3313( .i (n3312), .o (n3313) );
  buffer buf_n3314( .i (n3313), .o (n3314) );
  buffer buf_n3315( .i (n3314), .o (n3315) );
  buffer buf_n3316( .i (n3315), .o (n3316) );
  buffer buf_n3317( .i (n3316), .o (n3317) );
  buffer buf_n3318( .i (n3317), .o (n3318) );
  buffer buf_n3319( .i (n3318), .o (n3319) );
  buffer buf_n3320( .i (n3319), .o (n3320) );
  buffer buf_n3321( .i (n3320), .o (n3321) );
  assign n3322 = n3305 | n3321 ;
  assign n3323 = n3286 | n3322 ;
  buffer buf_n3324( .i (n3323), .o (n3324) );
  buffer buf_n3325( .i (n3324), .o (n3325) );
  buffer buf_n3326( .i (n3325), .o (n3326) );
  buffer buf_n3327( .i (n3326), .o (n3327) );
  buffer buf_n3328( .i (n3327), .o (n3328) );
  buffer buf_n3329( .i (n3328), .o (n3329) );
  buffer buf_n2825( .i (n2824), .o (n2825) );
  buffer buf_n2826( .i (n2825), .o (n2826) );
  buffer buf_n2827( .i (n2826), .o (n2827) );
  buffer buf_n2828( .i (n2827), .o (n2828) );
  buffer buf_n2829( .i (n2828), .o (n2829) );
  buffer buf_n2830( .i (n2829), .o (n2830) );
  assign n3330 = n2830 & ~n3012 ;
  buffer buf_n111( .i (x15), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  buffer buf_n113( .i (n112), .o (n113) );
  assign n3331 = n113 & ~n1451 ;
  buffer buf_n105( .i (x13), .o (n105) );
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  assign n3332 = n107 & n1451 ;
  assign n3333 = ( n1438 & n3331 ) | ( n1438 & n3332 ) | ( n3331 & n3332 ) ;
  buffer buf_n3334( .i (n3333), .o (n3334) );
  buffer buf_n3335( .i (n3334), .o (n3335) );
  buffer buf_n3336( .i (n3335), .o (n3336) );
  buffer buf_n3337( .i (n3336), .o (n3337) );
  buffer buf_n3338( .i (n3337), .o (n3338) );
  buffer buf_n3339( .i (n3338), .o (n3339) );
  buffer buf_n3340( .i (n3339), .o (n3340) );
  buffer buf_n3341( .i (n3340), .o (n3341) );
  buffer buf_n3342( .i (n3341), .o (n3342) );
  buffer buf_n3343( .i (n3342), .o (n3343) );
  buffer buf_n3344( .i (n3343), .o (n3344) );
  buffer buf_n3345( .i (n3344), .o (n3345) );
  buffer buf_n2816( .i (n2815), .o (n2816) );
  assign n3346 = n2816 & ~n3344 ;
  assign n3347 = ( n2869 & ~n3345 ) | ( n2869 & n3346 ) | ( ~n3345 & n3346 ) ;
  buffer buf_n3348( .i (n3347), .o (n3348) );
  buffer buf_n3349( .i (n3348), .o (n3349) );
  buffer buf_n3350( .i (n3349), .o (n3350) );
  assign n3351 = ~n3330 & n3350 ;
  buffer buf_n3352( .i (n3351), .o (n3352) );
  buffer buf_n3353( .i (n3352), .o (n3353) );
  assign n3354 = n2828 & n3032 ;
  buffer buf_n209( .i (x26), .o (n209) );
  buffer buf_n210( .i (n209), .o (n210) );
  buffer buf_n211( .i (n210), .o (n211) );
  buffer buf_n212( .i (n211), .o (n212) );
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n215( .i (n214), .o (n215) );
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  assign n3355 = n219 | n1459 ;
  buffer buf_n71( .i (x5), .o (n71) );
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  buffer buf_n75( .i (n74), .o (n75) );
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  buffer buf_n79( .i (n78), .o (n79) );
  buffer buf_n80( .i (n79), .o (n80) );
  buffer buf_n81( .i (n80), .o (n81) );
  assign n3356 = ~n81 & n1459 ;
  assign n3357 = ( n1446 & ~n3355 ) | ( n1446 & n3356 ) | ( ~n3355 & n3356 ) ;
  buffer buf_n3358( .i (n3357), .o (n3358) );
  buffer buf_n3359( .i (n3358), .o (n3359) );
  assign n3360 = n2814 & ~n3358 ;
  assign n3361 = ( n2888 & n3359 ) | ( n2888 & ~n3360 ) | ( n3359 & ~n3360 ) ;
  buffer buf_n3362( .i (n3361), .o (n3362) );
  buffer buf_n3363( .i (n3362), .o (n3363) );
  buffer buf_n3364( .i (n3363), .o (n3364) );
  assign n3365 = n3354 | n3364 ;
  buffer buf_n3366( .i (n3365), .o (n3366) );
  buffer buf_n3367( .i (n3366), .o (n3367) );
  buffer buf_n3368( .i (n3367), .o (n3368) );
  buffer buf_n3369( .i (n3368), .o (n3369) );
  assign n3370 = n2826 & ~n3052 ;
  buffer buf_n1447( .i (n1446), .o (n1447) );
  buffer buf_n193( .i (x25), .o (n193) );
  buffer buf_n194( .i (n193), .o (n194) );
  buffer buf_n195( .i (n194), .o (n195) );
  buffer buf_n196( .i (n195), .o (n196) );
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  buffer buf_n199( .i (n198), .o (n199) );
  buffer buf_n200( .i (n199), .o (n200) );
  buffer buf_n201( .i (n200), .o (n201) );
  buffer buf_n202( .i (n201), .o (n202) );
  buffer buf_n203( .i (n202), .o (n203) );
  buffer buf_n204( .i (n203), .o (n204) );
  assign n3371 = n204 & ~n1460 ;
  buffer buf_n55( .i (x4), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  buffer buf_n59( .i (n58), .o (n59) );
  buffer buf_n60( .i (n59), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  buffer buf_n64( .i (n63), .o (n64) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  assign n3372 = n66 & n1460 ;
  assign n3373 = ( n1447 & n3371 ) | ( n1447 & n3372 ) | ( n3371 & n3372 ) ;
  buffer buf_n3374( .i (n3373), .o (n3374) );
  buffer buf_n3375( .i (n3374), .o (n3375) );
  assign n3376 = n2815 & ~n3374 ;
  assign n3377 = ( n2927 & ~n3375 ) | ( n2927 & n3376 ) | ( ~n3375 & n3376 ) ;
  assign n3378 = ~n3370 & n3377 ;
  buffer buf_n3379( .i (n3378), .o (n3379) );
  buffer buf_n3380( .i (n3379), .o (n3380) );
  buffer buf_n3381( .i (n3380), .o (n3381) );
  buffer buf_n3382( .i (n3381), .o (n3382) );
  buffer buf_n3383( .i (n3382), .o (n3383) );
  buffer buf_n3384( .i (n3383), .o (n3384) );
  assign n3385 = n2732 | n2816 ;
  buffer buf_n163( .i (x23), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  buffer buf_n167( .i (n166), .o (n167) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  assign n3386 = n173 & ~n1459 ;
  buffer buf_n178( .i (x24), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n185( .i (n184), .o (n185) );
  buffer buf_n186( .i (n185), .o (n186) );
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  buffer buf_n3387( .i (n1458), .o (n3387) );
  assign n3388 = n188 & n3387 ;
  assign n3389 = ( n1446 & n3386 ) | ( n1446 & n3388 ) | ( n3386 & n3388 ) ;
  buffer buf_n3390( .i (n3389), .o (n3390) );
  buffer buf_n3391( .i (n3390), .o (n3391) );
  buffer buf_n3392( .i (n3391), .o (n3392) );
  assign n3393 = n2825 | n3391 ;
  assign n3394 = ( ~n3072 & n3392 ) | ( ~n3072 & n3393 ) | ( n3392 & n3393 ) ;
  assign n3395 = n3385 & ~n3394 ;
  buffer buf_n3396( .i (n3395), .o (n3396) );
  buffer buf_n3397( .i (n3396), .o (n3397) );
  buffer buf_n3398( .i (n3397), .o (n3398) );
  buffer buf_n3399( .i (n3398), .o (n3399) );
  buffer buf_n3400( .i (n3399), .o (n3400) );
  buffer buf_n3401( .i (n3400), .o (n3401) );
  buffer buf_n2961( .i (n2960), .o (n2961) );
  buffer buf_n2962( .i (n2961), .o (n2962) );
  buffer buf_n2963( .i (n2962), .o (n2963) );
  buffer buf_n2964( .i (n2963), .o (n2964) );
  buffer buf_n2965( .i (n2964), .o (n2965) );
  assign n3402 = n2965 & n3012 ;
  assign n3403 = n2868 & ~n2943 ;
  assign n3404 = ~n107 & n1464 ;
  assign n3405 = n113 | n1464 ;
  assign n3406 = ( n1488 & n3404 ) | ( n1488 & ~n3405 ) | ( n3404 & ~n3405 ) ;
  buffer buf_n3407( .i (n3406), .o (n3407) );
  buffer buf_n3408( .i (n3407), .o (n3408) );
  buffer buf_n3409( .i (n3408), .o (n3409) );
  buffer buf_n3410( .i (n3409), .o (n3410) );
  buffer buf_n3411( .i (n3410), .o (n3411) );
  buffer buf_n3412( .i (n3411), .o (n3412) );
  buffer buf_n3413( .i (n3412), .o (n3413) );
  buffer buf_n3414( .i (n3413), .o (n3414) );
  buffer buf_n3415( .i (n3414), .o (n3415) );
  buffer buf_n3416( .i (n3415), .o (n3416) );
  buffer buf_n3417( .i (n3416), .o (n3417) );
  buffer buf_n3418( .i (n3417), .o (n3418) );
  assign n3419 = n3403 | n3418 ;
  buffer buf_n3420( .i (n3419), .o (n3420) );
  buffer buf_n3421( .i (n3420), .o (n3421) );
  buffer buf_n3422( .i (n3421), .o (n3422) );
  assign n3423 = n3402 | n3422 ;
  buffer buf_n3424( .i (n3423), .o (n3424) );
  buffer buf_n3425( .i (n3424), .o (n3425) );
  assign n3426 = n2963 & ~n3032 ;
  assign n3427 = n2888 | n2942 ;
  buffer buf_n1493( .i (n1492), .o (n1493) );
  buffer buf_n1494( .i (n1493), .o (n1494) );
  buffer buf_n1495( .i (n1494), .o (n1495) );
  buffer buf_n1496( .i (n1495), .o (n1496) );
  buffer buf_n1497( .i (n1496), .o (n1497) );
  buffer buf_n1498( .i (n1497), .o (n1498) );
  buffer buf_n1499( .i (n1498), .o (n1499) );
  buffer buf_n82( .i (n81), .o (n82) );
  buffer buf_n83( .i (n82), .o (n83) );
  buffer buf_n84( .i (n83), .o (n84) );
  buffer buf_n1470( .i (n1469), .o (n1470) );
  buffer buf_n1471( .i (n1470), .o (n1471) );
  buffer buf_n1472( .i (n1471), .o (n1472) );
  buffer buf_n1473( .i (n1472), .o (n1473) );
  buffer buf_n1474( .i (n1473), .o (n1474) );
  buffer buf_n1475( .i (n1474), .o (n1475) );
  assign n3428 = n84 & n1475 ;
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  assign n3429 = n222 & ~n1475 ;
  assign n3430 = ( n1499 & n3428 ) | ( n1499 & n3429 ) | ( n3428 & n3429 ) ;
  assign n3431 = n3427 & ~n3430 ;
  buffer buf_n3432( .i (n3431), .o (n3432) );
  buffer buf_n3433( .i (n3432), .o (n3433) );
  assign n3434 = ~n3426 & n3433 ;
  buffer buf_n3435( .i (n3434), .o (n3435) );
  buffer buf_n3436( .i (n3435), .o (n3436) );
  buffer buf_n3437( .i (n3436), .o (n3437) );
  buffer buf_n3438( .i (n3437), .o (n3438) );
  assign n3439 = n2962 & ~n3053 ;
  assign n3440 = n2927 | n2943 ;
  buffer buf_n1500( .i (n1499), .o (n1500) );
  buffer buf_n67( .i (n66), .o (n67) );
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n1476( .i (n1475), .o (n1476) );
  assign n3441 = n69 & n1476 ;
  buffer buf_n205( .i (n204), .o (n205) );
  buffer buf_n206( .i (n205), .o (n206) );
  buffer buf_n207( .i (n206), .o (n207) );
  assign n3442 = n207 & ~n1476 ;
  assign n3443 = ( n1500 & n3441 ) | ( n1500 & n3442 ) | ( n3441 & n3442 ) ;
  assign n3444 = n3440 & ~n3443 ;
  assign n3445 = ~n3439 & n3444 ;
  buffer buf_n3446( .i (n3445), .o (n3446) );
  buffer buf_n3447( .i (n3446), .o (n3447) );
  buffer buf_n3448( .i (n3447), .o (n3448) );
  buffer buf_n3449( .i (n3448), .o (n3449) );
  buffer buf_n3450( .i (n3449), .o (n3450) );
  buffer buf_n3451( .i (n2942), .o (n3451) );
  assign n3452 = n2732 | n3451 ;
  assign n3453 = n2960 & ~n3071 ;
  buffer buf_n189( .i (n188), .o (n189) );
  buffer buf_n190( .i (n189), .o (n190) );
  buffer buf_n191( .i (n190), .o (n191) );
  assign n3454 = n191 & n1475 ;
  buffer buf_n174( .i (n173), .o (n174) );
  buffer buf_n175( .i (n174), .o (n175) );
  buffer buf_n176( .i (n175), .o (n176) );
  buffer buf_n3455( .i (n1474), .o (n3455) );
  assign n3456 = n176 & ~n3455 ;
  assign n3457 = ( n1499 & n3454 ) | ( n1499 & n3456 ) | ( n3454 & n3456 ) ;
  assign n3458 = n3453 | n3457 ;
  assign n3459 = n3452 & ~n3458 ;
  buffer buf_n3460( .i (n3459), .o (n3460) );
  buffer buf_n3461( .i (n3460), .o (n3461) );
  buffer buf_n3462( .i (n3461), .o (n3462) );
  buffer buf_n3463( .i (n3462), .o (n3463) );
  buffer buf_n3464( .i (n3463), .o (n3464) );
  buffer buf_n3465( .i (n3464), .o (n3465) );
  buffer buf_n3236( .i (n3235), .o (n3236) );
  buffer buf_n3237( .i (n3236), .o (n3237) );
  buffer buf_n3238( .i (n3237), .o (n3238) );
  buffer buf_n3239( .i (n3238), .o (n3239) );
  buffer buf_n3240( .i (n3239), .o (n3240) );
  assign n3466 = ~n3012 & n3240 ;
  buffer buf_n554( .i (x75), .o (n554) );
  buffer buf_n555( .i (n554), .o (n555) );
  buffer buf_n556( .i (n555), .o (n556) );
  buffer buf_n557( .i (n556), .o (n557) );
  buffer buf_n558( .i (n557), .o (n558) );
  buffer buf_n3467( .i (n1317), .o (n3467) );
  assign n3468 = n558 & n3467 ;
  buffer buf_n598( .i (x85), .o (n598) );
  buffer buf_n599( .i (n598), .o (n599) );
  buffer buf_n600( .i (n599), .o (n600) );
  buffer buf_n601( .i (n600), .o (n601) );
  buffer buf_n602( .i (n601), .o (n602) );
  assign n3469 = n602 & ~n3467 ;
  assign n3470 = ( n3246 & n3468 ) | ( n3246 & n3469 ) | ( n3468 & n3469 ) ;
  buffer buf_n3471( .i (n3470), .o (n3471) );
  buffer buf_n3472( .i (n3471), .o (n3472) );
  buffer buf_n3473( .i (n3472), .o (n3473) );
  buffer buf_n3474( .i (n3473), .o (n3474) );
  buffer buf_n3475( .i (n3474), .o (n3475) );
  buffer buf_n3476( .i (n3475), .o (n3476) );
  buffer buf_n3477( .i (n3476), .o (n3477) );
  buffer buf_n3478( .i (n3477), .o (n3478) );
  buffer buf_n3479( .i (n3478), .o (n3479) );
  buffer buf_n3480( .i (n3479), .o (n3480) );
  assign n3481 = ~n2868 & n3219 ;
  assign n3482 = n3480 | n3481 ;
  buffer buf_n3483( .i (n3482), .o (n3483) );
  buffer buf_n3484( .i (n3483), .o (n3484) );
  buffer buf_n3485( .i (n3484), .o (n3485) );
  assign n3486 = n3466 | n3485 ;
  buffer buf_n3487( .i (n3486), .o (n3487) );
  buffer buf_n3488( .i (n3487), .o (n3488) );
  assign n3489 = ~n2732 & n3219 ;
  buffer buf_n536( .i (x71), .o (n536) );
  buffer buf_n537( .i (n536), .o (n537) );
  buffer buf_n538( .i (n537), .o (n538) );
  buffer buf_n539( .i (n538), .o (n539) );
  buffer buf_n540( .i (n539), .o (n540) );
  assign n3490 = n540 & n3467 ;
  buffer buf_n580( .i (x81), .o (n580) );
  buffer buf_n581( .i (n580), .o (n581) );
  buffer buf_n582( .i (n581), .o (n582) );
  buffer buf_n583( .i (n582), .o (n583) );
  buffer buf_n584( .i (n583), .o (n584) );
  assign n3491 = n584 & ~n3467 ;
  assign n3492 = ( n3246 & n3490 ) | ( n3246 & n3491 ) | ( n3490 & n3491 ) ;
  buffer buf_n3493( .i (n3492), .o (n3493) );
  buffer buf_n3494( .i (n3493), .o (n3494) );
  buffer buf_n3495( .i (n3494), .o (n3495) );
  buffer buf_n3496( .i (n3495), .o (n3496) );
  buffer buf_n3497( .i (n3496), .o (n3497) );
  buffer buf_n3498( .i (n3497), .o (n3498) );
  buffer buf_n3499( .i (n3498), .o (n3499) );
  buffer buf_n3500( .i (n3499), .o (n3500) );
  buffer buf_n3501( .i (n3500), .o (n3501) );
  assign n3502 = ~n3071 & n3235 ;
  assign n3503 = n3501 | n3502 ;
  assign n3504 = n3489 | n3503 ;
  buffer buf_n3505( .i (n3504), .o (n3505) );
  buffer buf_n3506( .i (n3505), .o (n3506) );
  buffer buf_n3507( .i (n3506), .o (n3507) );
  buffer buf_n3508( .i (n3507), .o (n3508) );
  buffer buf_n3509( .i (n3508), .o (n3509) );
  buffer buf_n3510( .i (n3509), .o (n3510) );
  assign n3511 = ~n3051 & n3235 ;
  assign n3512 = n2759 & n3215 ;
  assign n3513 = ~n2918 & n3512 ;
  buffer buf_n526( .i (x69), .o (n526) );
  buffer buf_n527( .i (n526), .o (n527) );
  buffer buf_n528( .i (n527), .o (n528) );
  buffer buf_n529( .i (n528), .o (n529) );
  assign n3514 = n529 & n1317 ;
  buffer buf_n531( .i (x70), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  assign n3515 = n534 & ~n1317 ;
  assign n3516 = ( n3245 & n3514 ) | ( n3245 & n3515 ) | ( n3514 & n3515 ) ;
  buffer buf_n3517( .i (n3516), .o (n3517) );
  buffer buf_n3518( .i (n3517), .o (n3518) );
  buffer buf_n3519( .i (n3518), .o (n3519) );
  buffer buf_n3520( .i (n3519), .o (n3520) );
  buffer buf_n3521( .i (n3520), .o (n3521) );
  buffer buf_n3522( .i (n3521), .o (n3522) );
  buffer buf_n3523( .i (n3522), .o (n3523) );
  buffer buf_n3524( .i (n3523), .o (n3524) );
  assign n3525 = n3513 | n3524 ;
  assign n3526 = ~n2923 & n3215 ;
  buffer buf_n3527( .i (n3526), .o (n3527) );
  buffer buf_n3528( .i (n3527), .o (n3528) );
  assign n3529 = ~n2920 & n3216 ;
  assign n3530 = ~n3527 & n3529 ;
  assign n3531 = ( n3525 & n3528 ) | ( n3525 & ~n3530 ) | ( n3528 & ~n3530 ) ;
  assign n3532 = n3511 | n3531 ;
  buffer buf_n3533( .i (n3532), .o (n3533) );
  buffer buf_n3534( .i (n3533), .o (n3534) );
  buffer buf_n3535( .i (n3534), .o (n3535) );
  buffer buf_n3536( .i (n3535), .o (n3536) );
  buffer buf_n3537( .i (n3536), .o (n3537) );
  buffer buf_n3538( .i (n3537), .o (n3538) );
  buffer buf_n3539( .i (n3538), .o (n3539) );
  assign n3540 = ~n3030 & n3236 ;
  buffer buf_n514( .i (x67), .o (n514) );
  buffer buf_n515( .i (n514), .o (n515) );
  buffer buf_n516( .i (n515), .o (n516) );
  buffer buf_n517( .i (n516), .o (n517) );
  buffer buf_n518( .i (n517), .o (n518) );
  buffer buf_n3541( .i (n1316), .o (n3541) );
  buffer buf_n3542( .i (n3541), .o (n3542) );
  assign n3543 = n518 & n3542 ;
  buffer buf_n520( .i (x68), .o (n520) );
  buffer buf_n521( .i (n520), .o (n521) );
  buffer buf_n522( .i (n521), .o (n522) );
  buffer buf_n523( .i (n522), .o (n523) );
  buffer buf_n524( .i (n523), .o (n524) );
  assign n3544 = n524 & ~n3542 ;
  assign n3545 = ( n3246 & n3543 ) | ( n3246 & n3544 ) | ( n3543 & n3544 ) ;
  assign n3546 = n3210 | n3545 ;
  buffer buf_n3547( .i (n3546), .o (n3547) );
  buffer buf_n3548( .i (n3547), .o (n3548) );
  buffer buf_n3549( .i (n3548), .o (n3549) );
  buffer buf_n3550( .i (n3549), .o (n3550) );
  buffer buf_n3551( .i (n3550), .o (n3551) );
  buffer buf_n3552( .i (n3551), .o (n3552) );
  buffer buf_n3553( .i (n3552), .o (n3553) );
  buffer buf_n3554( .i (n3553), .o (n3554) );
  buffer buf_n3555( .i (n3554), .o (n3555) );
  buffer buf_n3556( .i (n3218), .o (n3556) );
  assign n3557 = n2889 & n3556 ;
  assign n3558 = ( n3540 & n3555 ) | ( n3540 & ~n3557 ) | ( n3555 & ~n3557 ) ;
  buffer buf_n3559( .i (n3558), .o (n3559) );
  buffer buf_n3560( .i (n3559), .o (n3560) );
  buffer buf_n3561( .i (n3560), .o (n3561) );
  buffer buf_n3562( .i (n3561), .o (n3562) );
  buffer buf_n3563( .i (n3562), .o (n3563) );
  buffer buf_n3564( .i (n3563), .o (n3564) );
  buffer buf_n3298( .i (n3297), .o (n3298) );
  buffer buf_n3299( .i (n3298), .o (n3299) );
  buffer buf_n3300( .i (n3299), .o (n3300) );
  buffer buf_n3301( .i (n3300), .o (n3301) );
  buffer buf_n3302( .i (n3301), .o (n3302) );
  buffer buf_n3565( .i (n3011), .o (n3565) );
  assign n3566 = n3302 & ~n3565 ;
  assign n3567 = n558 & n1328 ;
  assign n3568 = n602 & ~n1328 ;
  assign n3569 = ( n3309 & n3567 ) | ( n3309 & n3568 ) | ( n3567 & n3568 ) ;
  buffer buf_n3570( .i (n3569), .o (n3570) );
  buffer buf_n3571( .i (n3570), .o (n3571) );
  buffer buf_n3572( .i (n3571), .o (n3572) );
  buffer buf_n3573( .i (n3572), .o (n3573) );
  buffer buf_n3574( .i (n3573), .o (n3574) );
  buffer buf_n3575( .i (n3574), .o (n3575) );
  buffer buf_n3576( .i (n3575), .o (n3576) );
  buffer buf_n3577( .i (n3576), .o (n3577) );
  buffer buf_n3578( .i (n3577), .o (n3578) );
  buffer buf_n3579( .i (n3578), .o (n3579) );
  assign n3580 = ~n2868 & n3280 ;
  assign n3581 = n3579 | n3580 ;
  buffer buf_n3582( .i (n3581), .o (n3582) );
  buffer buf_n3583( .i (n3582), .o (n3583) );
  buffer buf_n3584( .i (n3583), .o (n3584) );
  assign n3585 = n3566 | n3584 ;
  buffer buf_n3586( .i (n3585), .o (n3586) );
  buffer buf_n3587( .i (n3586), .o (n3587) );
  buffer buf_n3588( .i (n2731), .o (n3588) );
  assign n3589 = n3280 & ~n3588 ;
  buffer buf_n3590( .i (n1327), .o (n3590) );
  assign n3591 = n540 & n3590 ;
  assign n3592 = n584 & ~n3590 ;
  assign n3593 = ( n3309 & n3591 ) | ( n3309 & n3592 ) | ( n3591 & n3592 ) ;
  buffer buf_n3594( .i (n3593), .o (n3594) );
  buffer buf_n3595( .i (n3594), .o (n3595) );
  buffer buf_n3596( .i (n3595), .o (n3596) );
  buffer buf_n3597( .i (n3596), .o (n3597) );
  buffer buf_n3598( .i (n3597), .o (n3598) );
  buffer buf_n3599( .i (n3598), .o (n3599) );
  buffer buf_n3600( .i (n3599), .o (n3600) );
  buffer buf_n3601( .i (n3600), .o (n3601) );
  buffer buf_n3602( .i (n3601), .o (n3602) );
  assign n3603 = ~n3071 & n3297 ;
  assign n3604 = n3602 | n3603 ;
  assign n3605 = n3589 | n3604 ;
  buffer buf_n3606( .i (n3605), .o (n3606) );
  buffer buf_n3607( .i (n3606), .o (n3607) );
  buffer buf_n3608( .i (n3607), .o (n3608) );
  buffer buf_n3609( .i (n3608), .o (n3609) );
  buffer buf_n3610( .i (n3609), .o (n3610) );
  buffer buf_n3611( .i (n3610), .o (n3611) );
  assign n3612 = ~n3051 & n3297 ;
  buffer buf_n3613( .i (n2758), .o (n3613) );
  assign n3614 = n3276 & n3613 ;
  assign n3615 = ~n2918 & n3614 ;
  buffer buf_n3616( .i (n1326), .o (n3616) );
  assign n3617 = n529 & n3616 ;
  assign n3618 = n534 & ~n3616 ;
  assign n3619 = ( n3308 & n3617 ) | ( n3308 & n3618 ) | ( n3617 & n3618 ) ;
  buffer buf_n3620( .i (n3619), .o (n3620) );
  buffer buf_n3621( .i (n3620), .o (n3621) );
  buffer buf_n3622( .i (n3621), .o (n3622) );
  buffer buf_n3623( .i (n3622), .o (n3623) );
  buffer buf_n3624( .i (n3623), .o (n3624) );
  buffer buf_n3625( .i (n3624), .o (n3625) );
  buffer buf_n3626( .i (n3625), .o (n3626) );
  buffer buf_n3627( .i (n3626), .o (n3627) );
  assign n3628 = n3615 | n3627 ;
  assign n3629 = ~n2923 & n3276 ;
  buffer buf_n3630( .i (n3629), .o (n3630) );
  buffer buf_n3631( .i (n3630), .o (n3631) );
  assign n3632 = ~n2920 & n3277 ;
  assign n3633 = ~n3630 & n3632 ;
  assign n3634 = ( n3628 & n3631 ) | ( n3628 & ~n3633 ) | ( n3631 & ~n3633 ) ;
  assign n3635 = n3612 | n3634 ;
  buffer buf_n3636( .i (n3635), .o (n3636) );
  buffer buf_n3637( .i (n3636), .o (n3637) );
  buffer buf_n3638( .i (n3637), .o (n3638) );
  buffer buf_n3639( .i (n3638), .o (n3639) );
  buffer buf_n3640( .i (n3639), .o (n3640) );
  buffer buf_n3641( .i (n3640), .o (n3641) );
  buffer buf_n3642( .i (n3641), .o (n3642) );
  assign n3643 = ~n3030 & n3298 ;
  assign n3644 = n518 & n3590 ;
  assign n3645 = n524 & ~n3590 ;
  assign n3646 = ( n3309 & n3644 ) | ( n3309 & n3645 ) | ( n3644 & n3645 ) ;
  assign n3647 = n3271 | n3646 ;
  buffer buf_n3648( .i (n3647), .o (n3648) );
  buffer buf_n3649( .i (n3648), .o (n3649) );
  buffer buf_n3650( .i (n3649), .o (n3650) );
  buffer buf_n3651( .i (n3650), .o (n3651) );
  buffer buf_n3652( .i (n3651), .o (n3652) );
  buffer buf_n3653( .i (n3652), .o (n3653) );
  buffer buf_n3654( .i (n3653), .o (n3654) );
  buffer buf_n3655( .i (n3654), .o (n3655) );
  buffer buf_n3656( .i (n3655), .o (n3656) );
  buffer buf_n3657( .i (n3279), .o (n3657) );
  assign n3658 = n2889 & n3657 ;
  assign n3659 = ( n3643 & n3656 ) | ( n3643 & ~n3658 ) | ( n3656 & ~n3658 ) ;
  buffer buf_n3660( .i (n3659), .o (n3660) );
  buffer buf_n3661( .i (n3660), .o (n3661) );
  buffer buf_n3662( .i (n3661), .o (n3662) );
  buffer buf_n3663( .i (n3662), .o (n3663) );
  buffer buf_n3664( .i (n3663), .o (n3664) );
  buffer buf_n3665( .i (n3664), .o (n3665) );
  assign n3666 = x61 & x177 ;
  buffer buf_n3667( .i (n3666), .o (n3667) );
  buffer buf_n3668( .i (n3667), .o (n3668) );
  buffer buf_n3669( .i (n3668), .o (n3669) );
  buffer buf_n3670( .i (n3669), .o (n3670) );
  buffer buf_n3671( .i (n3670), .o (n3671) );
  buffer buf_n3672( .i (n3671), .o (n3672) );
  buffer buf_n3673( .i (n3672), .o (n3673) );
  buffer buf_n3674( .i (n3673), .o (n3674) );
  buffer buf_n1415( .i (x170), .o (n1415) );
  buffer buf_n1416( .i (n1415), .o (n1416) );
  buffer buf_n1417( .i (n1416), .o (n1417) );
  buffer buf_n1418( .i (n1417), .o (n1418) );
  buffer buf_n1419( .i (n1418), .o (n1419) );
  buffer buf_n1420( .i (n1419), .o (n1420) );
  buffer buf_n1421( .i (n1420), .o (n1421) );
  buffer buf_n1422( .i (n1421), .o (n1422) );
  buffer buf_n378( .i (x53), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  buffer buf_n380( .i (n379), .o (n380) );
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n1398( .i (x169), .o (n1398) );
  buffer buf_n1399( .i (n1398), .o (n1399) );
  buffer buf_n1400( .i (n1399), .o (n1400) );
  buffer buf_n1401( .i (n1400), .o (n1401) );
  buffer buf_n1402( .i (n1401), .o (n1402) );
  buffer buf_n1403( .i (n1402), .o (n1403) );
  buffer buf_n1404( .i (n1403), .o (n1404) );
  assign n3675 = ~n384 & n1404 ;
  buffer buf_n1923( .i (n1922), .o (n1923) );
  assign n3676 = n1404 | n1923 ;
  assign n3677 = ( n1422 & ~n3675 ) | ( n1422 & n3676 ) | ( ~n3675 & n3676 ) ;
  assign n3678 = ~n3674 & n3677 ;
  buffer buf_n3679( .i (n3678), .o (n3679) );
  buffer buf_n3680( .i (n3679), .o (n3680) );
  buffer buf_n3681( .i (n3680), .o (n3681) );
  buffer buf_n3682( .i (n3681), .o (n3682) );
  buffer buf_n3683( .i (n3682), .o (n3683) );
  buffer buf_n3684( .i (n3683), .o (n3684) );
  buffer buf_n3685( .i (n3684), .o (n3685) );
  buffer buf_n3686( .i (n3685), .o (n3686) );
  buffer buf_n3687( .i (n3686), .o (n3687) );
  buffer buf_n3688( .i (n3687), .o (n3688) );
  buffer buf_n2505( .i (n2504), .o (n2505) );
  buffer buf_n2506( .i (n2505), .o (n2506) );
  buffer buf_n433( .i (x60), .o (n433) );
  buffer buf_n434( .i (n433), .o (n434) );
  buffer buf_n435( .i (n434), .o (n435) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n444( .i (n443), .o (n444) );
  buffer buf_n445( .i (n444), .o (n445) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n1405( .i (n1404), .o (n1405) );
  buffer buf_n1406( .i (n1405), .o (n1406) );
  buffer buf_n1407( .i (n1406), .o (n1407) );
  buffer buf_n1408( .i (n1407), .o (n1408) );
  buffer buf_n1409( .i (n1408), .o (n1409) );
  buffer buf_n1410( .i (n1409), .o (n1410) );
  buffer buf_n1411( .i (n1410), .o (n1411) );
  assign n3689 = n446 & ~n1411 ;
  buffer buf_n3690( .i (n3689), .o (n3690) );
  buffer buf_n3691( .i (n3690), .o (n3691) );
  buffer buf_n1412( .i (n1411), .o (n1412) );
  buffer buf_n1413( .i (n1412), .o (n1413) );
  assign n3692 = n1413 | n3690 ;
  assign n3693 = ( n2793 & n3691 ) | ( n2793 & n3692 ) | ( n3691 & n3692 ) ;
  buffer buf_n3694( .i (n3693), .o (n3694) );
  assign n3695 = n2506 | n3694 ;
  buffer buf_n1423( .i (n1422), .o (n1423) );
  buffer buf_n1424( .i (n1423), .o (n1424) );
  buffer buf_n1425( .i (n1424), .o (n1425) );
  buffer buf_n1426( .i (n1425), .o (n1426) );
  buffer buf_n1427( .i (n1426), .o (n1427) );
  buffer buf_n1428( .i (n1427), .o (n1428) );
  buffer buf_n1429( .i (n1428), .o (n1429) );
  buffer buf_n1430( .i (n1429), .o (n1430) );
  buffer buf_n1431( .i (n1430), .o (n1431) );
  buffer buf_n1432( .i (n1431), .o (n1432) );
  buffer buf_n1433( .i (n1432), .o (n1433) );
  assign n3696 = ( ~n1433 & n2506 ) | ( ~n1433 & n3694 ) | ( n2506 & n3694 ) ;
  assign n3697 = ( n3688 & ~n3695 ) | ( n3688 & n3696 ) | ( ~n3695 & n3696 ) ;
  buffer buf_n3698( .i (n3697), .o (n3698) );
  buffer buf_n3699( .i (n3698), .o (n3699) );
  buffer buf_n3700( .i (n3699), .o (n3700) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  buffer buf_n2794( .i (n2793), .o (n2794) );
  assign n3701 = ~n450 & n2794 ;
  assign n3702 = n450 & ~n2794 ;
  assign n3703 = n3701 | n3702 ;
  buffer buf_n3704( .i (n3703), .o (n3704) );
  buffer buf_n3705( .i (n3704), .o (n3705) );
  buffer buf_n3706( .i (n3705), .o (n3706) );
  buffer buf_n3707( .i (n3706), .o (n3707) );
  buffer buf_n1924( .i (n1923), .o (n1924) );
  buffer buf_n3708( .i (n2669), .o (n3708) );
  assign n3709 = n1924 & ~n3708 ;
  buffer buf_n3710( .i (n3709), .o (n3710) );
  assign n3711 = n382 & n2742 ;
  buffer buf_n3712( .i (n3711), .o (n3712) );
  buffer buf_n3713( .i (n3712), .o (n3713) );
  buffer buf_n3714( .i (n3713), .o (n3714) );
  buffer buf_n3715( .i (n3714), .o (n3715) );
  assign n3716 = n3710 | n3715 ;
  buffer buf_n3717( .i (n3716), .o (n3717) );
  buffer buf_n3718( .i (n3717), .o (n3718) );
  buffer buf_n3719( .i (n3718), .o (n3719) );
  buffer buf_n3720( .i (n3719), .o (n3720) );
  buffer buf_n3721( .i (n3720), .o (n3721) );
  buffer buf_n3722( .i (n3721), .o (n3722) );
  buffer buf_n3723( .i (n3722), .o (n3723) );
  buffer buf_n3724( .i (n3723), .o (n3724) );
  buffer buf_n3725( .i (n3724), .o (n3725) );
  assign n3726 = n2756 | n3714 ;
  assign n3727 = n3710 | n3726 ;
  buffer buf_n3728( .i (n3727), .o (n3728) );
  buffer buf_n3729( .i (n3728), .o (n3729) );
  buffer buf_n3730( .i (n3729), .o (n3730) );
  buffer buf_n3731( .i (n3730), .o (n3731) );
  buffer buf_n3732( .i (n3731), .o (n3732) );
  buffer buf_n3733( .i (n3732), .o (n3733) );
  buffer buf_n3734( .i (n3733), .o (n3734) );
  buffer buf_n3735( .i (n3734), .o (n3735) );
  buffer buf_n3736( .i (n3735), .o (n3736) );
  assign n3737 = ( ~n2798 & n3725 ) | ( ~n2798 & n3736 ) | ( n3725 & n3736 ) ;
  buffer buf_n3738( .i (n3737), .o (n3738) );
  buffer buf_n3739( .i (n3738), .o (n3739) );
  buffer buf_n3740( .i (n3739), .o (n3740) );
  assign n3741 = n1911 | n2668 ;
  buffer buf_n363( .i (x51), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  buffer buf_n367( .i (n366), .o (n367) );
  buffer buf_n368( .i (n367), .o (n368) );
  assign n3742 = n368 & n2743 ;
  assign n3743 = n3741 & ~n3742 ;
  buffer buf_n3744( .i (n3743), .o (n3744) );
  buffer buf_n3745( .i (n3744), .o (n3745) );
  buffer buf_n3746( .i (n3745), .o (n3746) );
  buffer buf_n3747( .i (n3746), .o (n3747) );
  buffer buf_n3748( .i (n3747), .o (n3748) );
  buffer buf_n3749( .i (n3748), .o (n3749) );
  buffer buf_n3750( .i (n3749), .o (n3750) );
  buffer buf_n3751( .i (n3750), .o (n3751) );
  buffer buf_n3752( .i (n3751), .o (n3752) );
  buffer buf_n3753( .i (n3752), .o (n3753) );
  buffer buf_n2517( .i (n2516), .o (n2517) );
  buffer buf_n2518( .i (n2517), .o (n2518) );
  buffer buf_n2519( .i (n2518), .o (n2519) );
  buffer buf_n2790( .i (n2789), .o (n2790) );
  assign n3754 = n2656 | n2790 ;
  buffer buf_n3755( .i (n3754), .o (n3755) );
  assign n3756 = ~n2519 & n3755 ;
  buffer buf_n2762( .i (n2761), .o (n2762) );
  buffer buf_n2763( .i (n2762), .o (n2763) );
  buffer buf_n2764( .i (n2763), .o (n2764) );
  assign n3757 = ( ~n2519 & n2764 ) | ( ~n2519 & n3755 ) | ( n2764 & n3755 ) ;
  assign n3758 = ( n3753 & n3756 ) | ( n3753 & ~n3757 ) | ( n3756 & ~n3757 ) ;
  buffer buf_n3759( .i (n3758), .o (n3759) );
  buffer buf_n3760( .i (n3759), .o (n3760) );
  buffer buf_n3761( .i (n3760), .o (n3761) );
  buffer buf_n3762( .i (n3761), .o (n3762) );
  buffer buf_n3763( .i (n3762), .o (n3763) );
  buffer buf_n328( .i (x46), .o (n328) );
  buffer buf_n329( .i (n328), .o (n329) );
  buffer buf_n330( .i (n329), .o (n330) );
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n333( .i (n332), .o (n333) );
  buffer buf_n334( .i (n333), .o (n334) );
  buffer buf_n3764( .i (n2742), .o (n3764) );
  buffer buf_n3765( .i (n3764), .o (n3765) );
  assign n3766 = n334 & n3765 ;
  buffer buf_n3767( .i (n3766), .o (n3767) );
  buffer buf_n3768( .i (n3767), .o (n3768) );
  buffer buf_n2671( .i (n2670), .o (n2671) );
  assign n3769 = n1882 & ~n2671 ;
  assign n3770 = n3768 | n3769 ;
  buffer buf_n3771( .i (n3770), .o (n3771) );
  buffer buf_n3772( .i (n3771), .o (n3772) );
  buffer buf_n3773( .i (n3772), .o (n3773) );
  buffer buf_n3774( .i (n3773), .o (n3774) );
  buffer buf_n3775( .i (n3774), .o (n3775) );
  buffer buf_n3776( .i (n3775), .o (n3776) );
  buffer buf_n3777( .i (n3776), .o (n3777) );
  buffer buf_n2445( .i (n2444), .o (n2445) );
  buffer buf_n2446( .i (n2445), .o (n2446) );
  buffer buf_n2447( .i (n2446), .o (n2447) );
  buffer buf_n2448( .i (n2447), .o (n2448) );
  buffer buf_n2449( .i (n2448), .o (n2449) );
  buffer buf_n2450( .i (n2449), .o (n2450) );
  buffer buf_n2451( .i (n2450), .o (n2451) );
  buffer buf_n2452( .i (n2451), .o (n2452) );
  buffer buf_n1121( .i (n1120), .o (n1121) );
  buffer buf_n1122( .i (n1121), .o (n1122) );
  buffer buf_n1123( .i (n1122), .o (n1123) );
  buffer buf_n1124( .i (n1123), .o (n1124) );
  buffer buf_n2461( .i (n2460), .o (n2461) );
  buffer buf_n2462( .i (n2461), .o (n2462) );
  buffer buf_n2463( .i (n2462), .o (n2463) );
  buffer buf_n2464( .i (n2463), .o (n2464) );
  buffer buf_n1135( .i (n1134), .o (n1135) );
  buffer buf_n1136( .i (n1135), .o (n1136) );
  buffer buf_n1137( .i (n1136), .o (n1137) );
  buffer buf_n1138( .i (n1137), .o (n1138) );
  buffer buf_n2353( .i (n2352), .o (n2353) );
  buffer buf_n2354( .i (n2353), .o (n2354) );
  buffer buf_n2355( .i (n2354), .o (n2355) );
  buffer buf_n2356( .i (n2355), .o (n2356) );
  assign n3778 = ( n1138 & n2356 ) | ( n1138 & n2864 ) | ( n2356 & n2864 ) ;
  buffer buf_n3779( .i (n3778), .o (n3779) );
  assign n3780 = ( n1124 & n2464 ) | ( n1124 & n3779 ) | ( n2464 & n3779 ) ;
  buffer buf_n3781( .i (n3780), .o (n3781) );
  assign n3782 = n2452 & n3781 ;
  assign n3783 = ( n2452 & n2764 ) | ( n2452 & n3781 ) | ( n2764 & n3781 ) ;
  assign n3784 = ( n3777 & ~n3782 ) | ( n3777 & n3783 ) | ( ~n3782 & n3783 ) ;
  buffer buf_n3785( .i (n3784), .o (n3785) );
  buffer buf_n3786( .i (n3785), .o (n3786) );
  buffer buf_n3787( .i (n3786), .o (n3787) );
  buffer buf_n3788( .i (n3787), .o (n3788) );
  buffer buf_n3789( .i (n3788), .o (n3789) );
  buffer buf_n300( .i (x42), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  assign n3790 = n305 & n3764 ;
  buffer buf_n3791( .i (n3790), .o (n3791) );
  buffer buf_n3792( .i (n3791), .o (n3792) );
  assign n3793 = n1892 & ~n3708 ;
  assign n3794 = n3792 | n3793 ;
  buffer buf_n3795( .i (n3794), .o (n3795) );
  buffer buf_n3796( .i (n3795), .o (n3796) );
  buffer buf_n3797( .i (n3796), .o (n3797) );
  buffer buf_n3798( .i (n3797), .o (n3798) );
  buffer buf_n3799( .i (n3798), .o (n3799) );
  buffer buf_n3800( .i (n3799), .o (n3800) );
  buffer buf_n2470( .i (n2469), .o (n2470) );
  assign n3801 = n2470 & ~n2524 ;
  buffer buf_n3802( .i (n3801), .o (n3802) );
  assign n3803 = n3779 & n3802 ;
  assign n3804 = ( n2762 & n3779 ) | ( n2762 & n3802 ) | ( n3779 & n3802 ) ;
  assign n3805 = ( n3800 & ~n3803 ) | ( n3800 & n3804 ) | ( ~n3803 & n3804 ) ;
  buffer buf_n3806( .i (n3805), .o (n3806) );
  buffer buf_n3807( .i (n3806), .o (n3807) );
  buffer buf_n3808( .i (n3807), .o (n3808) );
  buffer buf_n3809( .i (n3808), .o (n3809) );
  buffer buf_n3810( .i (n3809), .o (n3810) );
  buffer buf_n3811( .i (n3810), .o (n3811) );
  buffer buf_n3812( .i (n3811), .o (n3812) );
  assign n3813 = n666 & n1261 ;
  assign n3814 = n1536 & n3813 ;
  assign n3815 = n1652 & n3814 ;
  assign n3816 = n2553 & n3815 ;
  buffer buf_n3817( .i (n3816), .o (n3817) );
  assign n3818 = n2589 | n3101 ;
  assign n3819 = n3817 & ~n3818 ;
  buffer buf_n3820( .i (n3819), .o (n3820) );
  buffer buf_n3821( .i (n3820), .o (n3821) );
  buffer buf_n3822( .i (n3821), .o (n3822) );
  buffer buf_n3823( .i (n3822), .o (n3823) );
  assign n3824 = ~n3150 & n3823 ;
  buffer buf_n3825( .i (n3824), .o (n3825) );
  buffer buf_n3826( .i (n3825), .o (n3826) );
  buffer buf_n3827( .i (n3826), .o (n3827) );
  buffer buf_n3828( .i (n3827), .o (n3828) );
  buffer buf_n3829( .i (n3828), .o (n3829) );
  buffer buf_n3830( .i (n3829), .o (n3830) );
  buffer buf_n2311( .i (n2310), .o (n2311) );
  assign n3831 = n2228 & n2758 ;
  assign n3832 = ~n2311 & n3831 ;
  buffer buf_n322( .i (x45), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  buffer buf_n324( .i (n323), .o (n324) );
  buffer buf_n325( .i (n324), .o (n325) );
  buffer buf_n326( .i (n325), .o (n326) );
  assign n3833 = n326 & n2742 ;
  buffer buf_n3834( .i (n3833), .o (n3834) );
  buffer buf_n3835( .i (n3834), .o (n3835) );
  assign n3836 = n2669 & ~n3834 ;
  assign n3837 = ( n2020 & n3835 ) | ( n2020 & ~n3836 ) | ( n3835 & ~n3836 ) ;
  buffer buf_n3838( .i (n3837), .o (n3838) );
  buffer buf_n3839( .i (n3838), .o (n3839) );
  buffer buf_n3840( .i (n3839), .o (n3840) );
  buffer buf_n3841( .i (n3840), .o (n3841) );
  assign n3842 = n3832 | n3841 ;
  buffer buf_n3843( .i (n3842), .o (n3843) );
  buffer buf_n3844( .i (n3843), .o (n3844) );
  buffer buf_n3845( .i (n3844), .o (n3845) );
  assign n3846 = n2608 | n2629 ;
  assign n3847 = ( n2609 & n3189 ) | ( n2609 & n3846 ) | ( n3189 & n3846 ) ;
  buffer buf_n3848( .i (n3847), .o (n3848) );
  buffer buf_n2312( .i (n2311), .o (n2312) );
  buffer buf_n2313( .i (n2312), .o (n2313) );
  assign n3849 = ~n2313 & n2761 ;
  assign n3850 = n2223 & ~n3849 ;
  assign n3851 = n3848 & n3850 ;
  buffer buf_n1086( .i (n1085), .o (n1086) );
  assign n3852 = ~n1086 & n2754 ;
  assign n3853 = ( ~n2207 & n2755 ) | ( ~n2207 & n3852 ) | ( n2755 & n3852 ) ;
  buffer buf_n3854( .i (n3853), .o (n3854) );
  assign n3855 = n2309 & n3854 ;
  buffer buf_n3856( .i (n3855), .o (n3856) );
  buffer buf_n3857( .i (n3856), .o (n3857) );
  buffer buf_n3858( .i (n3857), .o (n3858) );
  buffer buf_n3859( .i (n3858), .o (n3859) );
  buffer buf_n3860( .i (n3859), .o (n3860) );
  assign n3861 = n2223 | n3859 ;
  assign n3862 = ( n3848 & n3860 ) | ( n3848 & n3861 ) | ( n3860 & n3861 ) ;
  assign n3863 = ( n3845 & ~n3851 ) | ( n3845 & n3862 ) | ( ~n3851 & n3862 ) ;
  buffer buf_n3864( .i (n3863), .o (n3864) );
  buffer buf_n3865( .i (n3864), .o (n3865) );
  buffer buf_n3866( .i (n3865), .o (n3866) );
  buffer buf_n3867( .i (n3866), .o (n3867) );
  buffer buf_n3868( .i (n3867), .o (n3868) );
  buffer buf_n3869( .i (n3868), .o (n3869) );
  buffer buf_n1519( .i (n1518), .o (n1519) );
  buffer buf_n1520( .i (n1519), .o (n1520) );
  buffer buf_n1521( .i (n1520), .o (n1521) );
  buffer buf_n2240( .i (n2239), .o (n2240) );
  buffer buf_n2241( .i (n2240), .o (n2241) );
  assign n3870 = ( n1521 & ~n2241 ) | ( n1521 & n3848 ) | ( ~n2241 & n3848 ) ;
  assign n3871 = ( n1521 & n2241 ) | ( n1521 & ~n3848 ) | ( n2241 & ~n3848 ) ;
  assign n3872 = n3870 & n3871 ;
  buffer buf_n3873( .i (n3872), .o (n3873) );
  buffer buf_n313( .i (x44), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  buffer buf_n316( .i (n315), .o (n316) );
  buffer buf_n317( .i (n316), .o (n317) );
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n319( .i (n318), .o (n319) );
  buffer buf_n320( .i (n319), .o (n320) );
  assign n3874 = ( ~n320 & n1513 ) | ( ~n320 & n1530 ) | ( n1513 & n1530 ) ;
  buffer buf_n3875( .i (n1529), .o (n3875) );
  assign n3876 = ( n2010 & ~n2755 ) | ( n2010 & n3875 ) | ( ~n2755 & n3875 ) ;
  assign n3877 = ( ~n2671 & n3874 ) | ( ~n2671 & n3876 ) | ( n3874 & n3876 ) ;
  buffer buf_n3878( .i (n3877), .o (n3878) );
  buffer buf_n3879( .i (n3878), .o (n3879) );
  buffer buf_n3880( .i (n3879), .o (n3880) );
  buffer buf_n3881( .i (n3880), .o (n3881) );
  buffer buf_n3882( .i (n3881), .o (n3882) );
  buffer buf_n3883( .i (n3882), .o (n3883) );
  buffer buf_n3884( .i (n3883), .o (n3884) );
  buffer buf_n3885( .i (n3884), .o (n3885) );
  buffer buf_n3886( .i (n3885), .o (n3886) );
  assign n3887 = n3873 | n3886 ;
  buffer buf_n3888( .i (n3887), .o (n3888) );
  buffer buf_n3889( .i (n3888), .o (n3889) );
  buffer buf_n3890( .i (n3889), .o (n3890) );
  buffer buf_n3891( .i (n3890), .o (n3891) );
  assign n3892 = n1982 | n3708 ;
  buffer buf_n131( .i (x19), .o (n131) );
  buffer buf_n132( .i (n131), .o (n132) );
  buffer buf_n133( .i (n132), .o (n133) );
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  buffer buf_n137( .i (n136), .o (n137) );
  assign n3893 = n137 & n3765 ;
  buffer buf_n3894( .i (n3893), .o (n3894) );
  assign n3895 = n3892 & ~n3894 ;
  buffer buf_n3896( .i (n3895), .o (n3896) );
  buffer buf_n3897( .i (n3896), .o (n3897) );
  buffer buf_n3898( .i (n3897), .o (n3898) );
  buffer buf_n3899( .i (n3898), .o (n3899) );
  buffer buf_n3900( .i (n3899), .o (n3900) );
  buffer buf_n3901( .i (n3900), .o (n3901) );
  buffer buf_n3902( .i (n3901), .o (n3902) );
  buffer buf_n2195( .i (n2194), .o (n2195) );
  buffer buf_n2196( .i (n2195), .o (n2196) );
  buffer buf_n2197( .i (n2196), .o (n2197) );
  buffer buf_n2198( .i (n2197), .o (n2198) );
  buffer buf_n2199( .i (n2198), .o (n2199) );
  buffer buf_n1044( .i (n1043), .o (n1044) );
  buffer buf_n1045( .i (n1044), .o (n1045) );
  buffer buf_n1046( .i (n1045), .o (n1046) );
  buffer buf_n1047( .i (n1046), .o (n1047) );
  buffer buf_n1048( .i (n1047), .o (n1048) );
  buffer buf_n1049( .i (n1048), .o (n1049) );
  buffer buf_n1050( .i (n1049), .o (n1050) );
  buffer buf_n1051( .i (n1050), .o (n1051) );
  buffer buf_n1052( .i (n1051), .o (n1052) );
  buffer buf_n2251( .i (n2250), .o (n2251) );
  buffer buf_n2252( .i (n2251), .o (n2252) );
  buffer buf_n2253( .i (n2252), .o (n2253) );
  buffer buf_n2254( .i (n2253), .o (n2254) );
  buffer buf_n2255( .i (n2254), .o (n2255) );
  buffer buf_n2256( .i (n2255), .o (n2256) );
  assign n3903 = ( n1052 & n2256 ) | ( n1052 & n3189 ) | ( n2256 & n3189 ) ;
  buffer buf_n3904( .i (n3903), .o (n3904) );
  assign n3905 = n2199 & n3904 ;
  assign n3906 = ( n2199 & n2763 ) | ( n2199 & n3904 ) | ( n2763 & n3904 ) ;
  assign n3907 = ( n3902 & n3905 ) | ( n3902 & ~n3906 ) | ( n3905 & ~n3906 ) ;
  buffer buf_n3908( .i (n3907), .o (n3908) );
  buffer buf_n3909( .i (n3908), .o (n3909) );
  buffer buf_n3910( .i (n3909), .o (n3910) );
  buffer buf_n3911( .i (n3910), .o (n3911) );
  buffer buf_n3912( .i (n3911), .o (n3912) );
  buffer buf_n3913( .i (n3912), .o (n3913) );
  assign n3914 = n2176 | n2268 ;
  buffer buf_n307( .i (x43), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  buffer buf_n310( .i (n309), .o (n310) );
  buffer buf_n311( .i (n310), .o (n311) );
  assign n3915 = ( ~n311 & n1510 ) | ( ~n311 & n2667 ) | ( n1510 & n2667 ) ;
  buffer buf_n3916( .i (n3915), .o (n3916) );
  buffer buf_n3917( .i (n3916), .o (n3917) );
  buffer buf_n3918( .i (n3917), .o (n3918) );
  buffer buf_n3919( .i (n3918), .o (n3919) );
  assign n3920 = n1531 & n3918 ;
  assign n3921 = ( ~n3914 & n3919 ) | ( ~n3914 & n3920 ) | ( n3919 & n3920 ) ;
  buffer buf_n3922( .i (n3921), .o (n3922) );
  buffer buf_n3923( .i (n3922), .o (n3923) );
  buffer buf_n3924( .i (n3923), .o (n3924) );
  buffer buf_n3925( .i (n3924), .o (n3925) );
  buffer buf_n3926( .i (n3925), .o (n3926) );
  buffer buf_n3927( .i (n3926), .o (n3927) );
  buffer buf_n3928( .i (n3927), .o (n3928) );
  buffer buf_n3929( .i (n3928), .o (n3929) );
  assign n3930 = n1529 & ~n3916 ;
  assign n3931 = ( n2053 & n3917 ) | ( n2053 & ~n3930 ) | ( n3917 & ~n3930 ) ;
  buffer buf_n3932( .i (n3931), .o (n3932) );
  buffer buf_n3933( .i (n3932), .o (n3933) );
  buffer buf_n3934( .i (n3933), .o (n3934) );
  buffer buf_n3935( .i (n3934), .o (n3935) );
  buffer buf_n3936( .i (n3935), .o (n3936) );
  buffer buf_n3937( .i (n3936), .o (n3937) );
  buffer buf_n3938( .i (n3937), .o (n3938) );
  buffer buf_n3939( .i (n3938), .o (n3939) );
  buffer buf_n3940( .i (n3939), .o (n3940) );
  buffer buf_n2271( .i (n2270), .o (n2271) );
  buffer buf_n2272( .i (n2271), .o (n2272) );
  buffer buf_n2273( .i (n2272), .o (n2273) );
  buffer buf_n2274( .i (n2273), .o (n2274) );
  buffer buf_n2275( .i (n2274), .o (n2275) );
  buffer buf_n2276( .i (n2275), .o (n2276) );
  buffer buf_n3191( .i (n3190), .o (n3191) );
  buffer buf_n2672( .i (n2671), .o (n2672) );
  buffer buf_n2673( .i (n2672), .o (n2673) );
  buffer buf_n2674( .i (n2673), .o (n2674) );
  buffer buf_n2675( .i (n2674), .o (n2675) );
  buffer buf_n2676( .i (n2675), .o (n2676) );
  assign n3941 = ( n2273 & n2676 ) | ( n2273 & n3005 ) | ( n2676 & n3005 ) ;
  buffer buf_n3942( .i (n3941), .o (n3942) );
  assign n3943 = ~n3191 & n3942 ;
  buffer buf_n2677( .i (n2676), .o (n2677) );
  buffer buf_n2678( .i (n2677), .o (n2678) );
  assign n3944 = ( n2678 & n3191 ) | ( n2678 & n3942 ) | ( n3191 & n3942 ) ;
  assign n3945 = ( ~n2276 & n3943 ) | ( ~n2276 & n3944 ) | ( n3943 & n3944 ) ;
  assign n3946 = n3940 & ~n3945 ;
  assign n3947 = n3929 | n3946 ;
  buffer buf_n3948( .i (n3947), .o (n3948) );
  buffer buf_n3949( .i (n3948), .o (n3949) );
  buffer buf_n3950( .i (n3949), .o (n3950) );
  buffer buf_n3951( .i (n3950), .o (n3951) );
  assign n3952 = n2964 & ~n3864 ;
  buffer buf_n3953( .i (n3952), .o (n3953) );
  buffer buf_n284( .i (x40), .o (n284) );
  buffer buf_n285( .i (n284), .o (n285) );
  buffer buf_n286( .i (n285), .o (n286) );
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  buffer buf_n290( .i (n289), .o (n290) );
  assign n3954 = ~n290 & n1468 ;
  buffer buf_n292( .i (x41), .o (n292) );
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  buffer buf_n295( .i (n294), .o (n295) );
  buffer buf_n296( .i (n295), .o (n296) );
  buffer buf_n297( .i (n296), .o (n297) );
  buffer buf_n298( .i (n297), .o (n298) );
  assign n3955 = n298 | n1468 ;
  assign n3956 = ( n1492 & n3954 ) | ( n1492 & ~n3955 ) | ( n3954 & ~n3955 ) ;
  buffer buf_n3957( .i (n3956), .o (n3957) );
  buffer buf_n3958( .i (n3957), .o (n3958) );
  buffer buf_n3959( .i (n3958), .o (n3959) );
  assign n3960 = n2937 & ~n3957 ;
  buffer buf_n3961( .i (n3960), .o (n3961) );
  assign n3962 = ( n3717 & ~n3959 ) | ( n3717 & n3961 ) | ( ~n3959 & n3961 ) ;
  buffer buf_n3963( .i (n3962), .o (n3963) );
  buffer buf_n3964( .i (n3963), .o (n3964) );
  buffer buf_n3965( .i (n3964), .o (n3965) );
  buffer buf_n3966( .i (n3965), .o (n3966) );
  buffer buf_n3967( .i (n3966), .o (n3967) );
  buffer buf_n3968( .i (n3967), .o (n3968) );
  buffer buf_n3969( .i (n3968), .o (n3969) );
  buffer buf_n3970( .i (n3969), .o (n3970) );
  assign n3971 = ~n3953 & n3970 ;
  assign n3972 = ( n3728 & ~n3959 ) | ( n3728 & n3961 ) | ( ~n3959 & n3961 ) ;
  buffer buf_n3973( .i (n3972), .o (n3973) );
  buffer buf_n3974( .i (n3973), .o (n3974) );
  buffer buf_n3975( .i (n3974), .o (n3975) );
  buffer buf_n3976( .i (n3975), .o (n3976) );
  buffer buf_n3977( .i (n3976), .o (n3977) );
  buffer buf_n3978( .i (n3977), .o (n3978) );
  buffer buf_n3979( .i (n3978), .o (n3979) );
  buffer buf_n3980( .i (n3979), .o (n3980) );
  assign n3981 = ~n3953 & n3980 ;
  assign n3982 = ( ~n2800 & n3971 ) | ( ~n2800 & n3981 ) | ( n3971 & n3981 ) ;
  buffer buf_n3983( .i (n3982), .o (n3983) );
  buffer buf_n2831( .i (n2830), .o (n2831) );
  buffer buf_n2832( .i (n2831), .o (n2832) );
  assign n3984 = n2832 & ~n3867 ;
  assign n3985 = n294 | n1451 ;
  buffer buf_n3986( .i (n1450), .o (n3986) );
  assign n3987 = ~n286 & n3986 ;
  assign n3988 = ( n1438 & ~n3985 ) | ( n1438 & n3987 ) | ( ~n3985 & n3987 ) ;
  buffer buf_n3989( .i (n3988), .o (n3989) );
  buffer buf_n3990( .i (n3989), .o (n3990) );
  buffer buf_n3991( .i (n3990), .o (n3991) );
  buffer buf_n3992( .i (n3991), .o (n3992) );
  buffer buf_n3993( .i (n3992), .o (n3993) );
  buffer buf_n3994( .i (n3993), .o (n3994) );
  buffer buf_n3995( .i (n3994), .o (n3995) );
  buffer buf_n3996( .i (n3995), .o (n3996) );
  buffer buf_n3997( .i (n3996), .o (n3997) );
  buffer buf_n3998( .i (n3997), .o (n3998) );
  buffer buf_n3999( .i (n3998), .o (n3999) );
  buffer buf_n4000( .i (n3999), .o (n4000) );
  buffer buf_n4001( .i (n4000), .o (n4001) );
  buffer buf_n4002( .i (n4001), .o (n4002) );
  buffer buf_n4003( .i (n4002), .o (n4003) );
  buffer buf_n4004( .i (n4003), .o (n4004) );
  buffer buf_n4005( .i (n4004), .o (n4005) );
  buffer buf_n2817( .i (n2816), .o (n2817) );
  buffer buf_n2818( .i (n2817), .o (n2818) );
  buffer buf_n2819( .i (n2818), .o (n2819) );
  buffer buf_n2820( .i (n2819), .o (n2820) );
  buffer buf_n2821( .i (n2820), .o (n2821) );
  assign n4006 = n2821 & ~n4004 ;
  assign n4007 = ( n3738 & ~n4005 ) | ( n3738 & n4006 ) | ( ~n4005 & n4006 ) ;
  assign n4008 = ~n3984 & n4007 ;
  assign n4009 = n2831 & n3888 ;
  buffer buf_n115( .i (x16), .o (n115) );
  buffer buf_n116( .i (n115), .o (n116) );
  buffer buf_n117( .i (n116), .o (n117) );
  assign n4010 = n117 | n3986 ;
  buffer buf_n119( .i (x17), .o (n119) );
  buffer buf_n120( .i (n119), .o (n120) );
  buffer buf_n121( .i (n120), .o (n121) );
  assign n4011 = ~n121 & n3986 ;
  assign n4012 = ( n1438 & ~n4010 ) | ( n1438 & n4011 ) | ( ~n4010 & n4011 ) ;
  buffer buf_n4013( .i (n4012), .o (n4013) );
  buffer buf_n4014( .i (n4013), .o (n4014) );
  buffer buf_n4015( .i (n4014), .o (n4015) );
  buffer buf_n4016( .i (n4015), .o (n4016) );
  buffer buf_n4017( .i (n4016), .o (n4017) );
  buffer buf_n4018( .i (n4017), .o (n4018) );
  buffer buf_n4019( .i (n4018), .o (n4019) );
  buffer buf_n4020( .i (n4019), .o (n4020) );
  buffer buf_n4021( .i (n4020), .o (n4021) );
  buffer buf_n4022( .i (n4021), .o (n4022) );
  buffer buf_n4023( .i (n4022), .o (n4023) );
  buffer buf_n4024( .i (n4023), .o (n4024) );
  buffer buf_n4025( .i (n4024), .o (n4025) );
  buffer buf_n4026( .i (n4025), .o (n4026) );
  buffer buf_n4027( .i (n4026), .o (n4027) );
  buffer buf_n4028( .i (n4027), .o (n4028) );
  assign n4029 = n2820 & ~n4027 ;
  assign n4030 = ( n3760 & n4028 ) | ( n3760 & ~n4029 ) | ( n4028 & ~n4029 ) ;
  assign n4031 = n4009 | n4030 ;
  buffer buf_n4032( .i (n4031), .o (n4032) );
  assign n4033 = n2830 & ~n3909 ;
  buffer buf_n268( .i (x38), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  assign n4034 = n270 & ~n3986 ;
  buffer buf_n276( .i (x39), .o (n276) );
  buffer buf_n277( .i (n276), .o (n277) );
  buffer buf_n278( .i (n277), .o (n278) );
  buffer buf_n4035( .i (n1450), .o (n4035) );
  assign n4036 = n278 & n4035 ;
  buffer buf_n4037( .i (n1437), .o (n4037) );
  assign n4038 = ( n4034 & n4036 ) | ( n4034 & n4037 ) | ( n4036 & n4037 ) ;
  buffer buf_n4039( .i (n4038), .o (n4039) );
  buffer buf_n4040( .i (n4039), .o (n4040) );
  buffer buf_n4041( .i (n4040), .o (n4041) );
  buffer buf_n4042( .i (n4041), .o (n4042) );
  buffer buf_n4043( .i (n4042), .o (n4043) );
  buffer buf_n4044( .i (n4043), .o (n4044) );
  buffer buf_n4045( .i (n4044), .o (n4045) );
  buffer buf_n4046( .i (n4045), .o (n4046) );
  buffer buf_n4047( .i (n4046), .o (n4047) );
  buffer buf_n4048( .i (n4047), .o (n4048) );
  buffer buf_n4049( .i (n4048), .o (n4049) );
  buffer buf_n4050( .i (n4049), .o (n4050) );
  buffer buf_n4051( .i (n4050), .o (n4051) );
  buffer buf_n4052( .i (n4051), .o (n4052) );
  buffer buf_n4053( .i (n4052), .o (n4053) );
  assign n4054 = n2819 & ~n4052 ;
  assign n4055 = ( n3785 & n4053 ) | ( n3785 & ~n4054 ) | ( n4053 & ~n4054 ) ;
  assign n4056 = n4033 | n4055 ;
  buffer buf_n4057( .i (n4056), .o (n4057) );
  buffer buf_n4058( .i (n4057), .o (n4058) );
  buffer buf_n253( .i (x35), .o (n253) );
  assign n4059 = n253 | n1449 ;
  buffer buf_n109( .i (x14), .o (n109) );
  assign n4060 = ~n109 & n1449 ;
  assign n4061 = ( n1436 & ~n4059 ) | ( n1436 & n4060 ) | ( ~n4059 & n4060 ) ;
  buffer buf_n4062( .i (n4061), .o (n4062) );
  buffer buf_n4063( .i (n4062), .o (n4063) );
  buffer buf_n4064( .i (n4063), .o (n4064) );
  buffer buf_n4065( .i (n4064), .o (n4065) );
  buffer buf_n4066( .i (n4065), .o (n4066) );
  buffer buf_n4067( .i (n4066), .o (n4067) );
  buffer buf_n4068( .i (n4067), .o (n4068) );
  buffer buf_n4069( .i (n4068), .o (n4069) );
  buffer buf_n4070( .i (n4069), .o (n4070) );
  buffer buf_n4071( .i (n4070), .o (n4071) );
  buffer buf_n4072( .i (n4071), .o (n4072) );
  buffer buf_n4073( .i (n4072), .o (n4073) );
  buffer buf_n4074( .i (n4073), .o (n4074) );
  buffer buf_n4075( .i (n4074), .o (n4075) );
  buffer buf_n4076( .i (n4075), .o (n4076) );
  assign n4077 = n2817 & ~n4075 ;
  assign n4078 = ( n3806 & ~n4076 ) | ( n3806 & n4077 ) | ( ~n4076 & n4077 ) ;
  buffer buf_n4079( .i (n4078), .o (n4079) );
  buffer buf_n4080( .i (n4079), .o (n4080) );
  assign n4081 = ~n2830 & n4079 ;
  assign n4082 = ( ~n3948 & n4080 ) | ( ~n3948 & n4081 ) | ( n4080 & n4081 ) ;
  buffer buf_n4083( .i (n4082), .o (n4083) );
  buffer buf_n4084( .i (n4083), .o (n4084) );
  buffer buf_n1477( .i (n1476), .o (n1477) );
  buffer buf_n1478( .i (n1477), .o (n1478) );
  buffer buf_n1479( .i (n1478), .o (n1479) );
  buffer buf_n1480( .i (n1479), .o (n1480) );
  buffer buf_n1481( .i (n1480), .o (n1481) );
  buffer buf_n1482( .i (n1481), .o (n1482) );
  buffer buf_n1483( .i (n1482), .o (n1483) );
  assign n4085 = n120 & n1463 ;
  assign n4086 = n116 & ~n1463 ;
  assign n4087 = ( n1487 & n4085 ) | ( n1487 & n4086 ) | ( n4085 & n4086 ) ;
  buffer buf_n4088( .i (n4087), .o (n4088) );
  buffer buf_n4089( .i (n4088), .o (n4089) );
  buffer buf_n4090( .i (n4089), .o (n4090) );
  buffer buf_n4091( .i (n4090), .o (n4091) );
  buffer buf_n4092( .i (n4091), .o (n4092) );
  buffer buf_n4093( .i (n4092), .o (n4093) );
  buffer buf_n4094( .i (n4093), .o (n4094) );
  assign n4095 = n2955 | n4093 ;
  assign n4096 = ( ~n3878 & n4094 ) | ( ~n3878 & n4095 ) | ( n4094 & n4095 ) ;
  buffer buf_n4097( .i (n4096), .o (n4097) );
  buffer buf_n4098( .i (n4097), .o (n4098) );
  buffer buf_n4099( .i (n4098), .o (n4099) );
  buffer buf_n4100( .i (n4099), .o (n4100) );
  buffer buf_n4101( .i (n4100), .o (n4101) );
  buffer buf_n4102( .i (n4101), .o (n4102) );
  buffer buf_n4103( .i (n4102), .o (n4103) );
  buffer buf_n4104( .i (n4103), .o (n4104) );
  buffer buf_n4105( .i (n4104), .o (n4105) );
  buffer buf_n1501( .i (n1500), .o (n1501) );
  buffer buf_n1502( .i (n1501), .o (n1502) );
  buffer buf_n1503( .i (n1502), .o (n1503) );
  buffer buf_n1504( .i (n1503), .o (n1504) );
  assign n4106 = n1504 | n3759 ;
  assign n4107 = ~n4105 & n4106 ;
  assign n4108 = ~n1503 & n3873 ;
  assign n4109 = n4104 & ~n4108 ;
  buffer buf_n4110( .i (n4109), .o (n4110) );
  assign n4111 = ( n1483 & n4107 ) | ( n1483 & ~n4110 ) | ( n4107 & ~n4110 ) ;
  buffer buf_n4112( .i (n4111), .o (n4112) );
  assign n4113 = n2965 & n3909 ;
  buffer buf_n279( .i (n278), .o (n279) );
  buffer buf_n280( .i (n279), .o (n280) );
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n282( .i (n281), .o (n282) );
  assign n4114 = ~n282 & n1468 ;
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n273( .i (n272), .o (n273) );
  buffer buf_n274( .i (n273), .o (n274) );
  buffer buf_n4115( .i (n1467), .o (n4115) );
  assign n4116 = n274 | n4115 ;
  assign n4117 = ( n1492 & n4114 ) | ( n1492 & ~n4116 ) | ( n4114 & ~n4116 ) ;
  buffer buf_n4118( .i (n4117), .o (n4118) );
  buffer buf_n4119( .i (n4118), .o (n4119) );
  buffer buf_n4120( .i (n4119), .o (n4120) );
  buffer buf_n4121( .i (n4120), .o (n4121) );
  buffer buf_n4122( .i (n4121), .o (n4122) );
  buffer buf_n4123( .i (n4122), .o (n4123) );
  buffer buf_n4124( .i (n4123), .o (n4124) );
  buffer buf_n4125( .i (n4124), .o (n4125) );
  buffer buf_n4126( .i (n4125), .o (n4126) );
  buffer buf_n4127( .i (n4126), .o (n4127) );
  buffer buf_n4128( .i (n4127), .o (n4128) );
  buffer buf_n2944( .i (n2943), .o (n2944) );
  buffer buf_n2945( .i (n2944), .o (n2945) );
  buffer buf_n2946( .i (n2945), .o (n2946) );
  assign n4129 = n2946 & ~n4127 ;
  assign n4130 = ( n3785 & ~n4128 ) | ( n3785 & n4129 ) | ( ~n4128 & n4129 ) ;
  assign n4131 = ~n4113 & n4130 ;
  buffer buf_n4132( .i (n4131), .o (n4132) );
  buffer buf_n4133( .i (n4132), .o (n4133) );
  assign n4134 = ( n2274 & n2762 ) | ( n2274 & n3190 ) | ( n2762 & n3190 ) ;
  assign n4135 = ( n2274 & ~n2762 ) | ( n2274 & n3190 ) | ( ~n2762 & n3190 ) ;
  assign n4136 = n4134 & ~n4135 ;
  buffer buf_n4137( .i (n4136), .o (n4137) );
  assign n4138 = n2963 & n4137 ;
  assign n4139 = n109 & n1462 ;
  assign n4140 = n253 & ~n1462 ;
  assign n4141 = ( n1486 & n4139 ) | ( n1486 & n4140 ) | ( n4139 & n4140 ) ;
  buffer buf_n4142( .i (n4141), .o (n4142) );
  buffer buf_n4143( .i (n4142), .o (n4143) );
  buffer buf_n4144( .i (n4143), .o (n4144) );
  buffer buf_n4145( .i (n4144), .o (n4145) );
  buffer buf_n4146( .i (n4145), .o (n4146) );
  buffer buf_n4147( .i (n4146), .o (n4147) );
  buffer buf_n4148( .i (n4147), .o (n4148) );
  assign n4149 = n2954 | n4147 ;
  assign n4150 = ( ~n3932 & n4148 ) | ( ~n3932 & n4149 ) | ( n4148 & n4149 ) ;
  buffer buf_n4151( .i (n4150), .o (n4151) );
  buffer buf_n4152( .i (n4151), .o (n4152) );
  buffer buf_n4153( .i (n4152), .o (n4153) );
  buffer buf_n4154( .i (n4153), .o (n4154) );
  buffer buf_n4155( .i (n4154), .o (n4155) );
  buffer buf_n4156( .i (n4155), .o (n4156) );
  buffer buf_n4157( .i (n4156), .o (n4157) );
  assign n4158 = n2944 & ~n4156 ;
  assign n4159 = ( n3806 & n4157 ) | ( n3806 & ~n4158 ) | ( n4157 & ~n4158 ) ;
  assign n4160 = n4138 | n4159 ;
  buffer buf_n4161( .i (n4160), .o (n4161) );
  buffer buf_n4162( .i (n4161), .o (n4162) );
  buffer buf_n4163( .i (n4162), .o (n4163) );
  buffer buf_n4164( .i (n4163), .o (n4164) );
  assign n4165 = n3940 & ~n4137 ;
  buffer buf_n4166( .i (n4165), .o (n4166) );
  assign n4167 = n3240 & ~n4166 ;
  buffer buf_n560( .i (x76), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  assign n4168 = n562 & n1316 ;
  buffer buf_n4169( .i (n4168), .o (n4169) );
  buffer buf_n4170( .i (n4169), .o (n4170) );
  buffer buf_n604( .i (x86), .o (n604) );
  buffer buf_n605( .i (n604), .o (n605) );
  buffer buf_n606( .i (n605), .o (n606) );
  assign n4171 = n606 & ~n1316 ;
  buffer buf_n4172( .i (n4171), .o (n4172) );
  buffer buf_n4173( .i (n4172), .o (n4173) );
  buffer buf_n4174( .i (n3245), .o (n4174) );
  assign n4175 = ( n4170 & n4173 ) | ( n4170 & n4174 ) | ( n4173 & n4174 ) ;
  buffer buf_n4176( .i (n4175), .o (n4176) );
  buffer buf_n4177( .i (n4176), .o (n4177) );
  buffer buf_n4178( .i (n4177), .o (n4178) );
  buffer buf_n4179( .i (n4178), .o (n4179) );
  buffer buf_n4180( .i (n4179), .o (n4180) );
  buffer buf_n4181( .i (n4180), .o (n4181) );
  buffer buf_n4182( .i (n4181), .o (n4182) );
  buffer buf_n4183( .i (n4182), .o (n4183) );
  buffer buf_n4184( .i (n4183), .o (n4184) );
  buffer buf_n4185( .i (n4184), .o (n4185) );
  buffer buf_n4186( .i (n4185), .o (n4186) );
  buffer buf_n4187( .i (n4186), .o (n4187) );
  buffer buf_n4188( .i (n4187), .o (n4188) );
  buffer buf_n3220( .i (n3219), .o (n3220) );
  buffer buf_n3221( .i (n3220), .o (n3221) );
  buffer buf_n3222( .i (n3221), .o (n3222) );
  assign n4189 = n3222 | n4187 ;
  assign n4190 = ( n3808 & n4188 ) | ( n3808 & n4189 ) | ( n4188 & n4189 ) ;
  assign n4191 = n4167 | n4190 ;
  buffer buf_n4192( .i (n4191), .o (n4192) );
  buffer buf_n4193( .i (n4192), .o (n4193) );
  buffer buf_n3241( .i (n3240), .o (n3241) );
  assign n4194 = n3241 & ~n3910 ;
  buffer buf_n550( .i (x74), .o (n550) );
  buffer buf_n551( .i (n550), .o (n551) );
  buffer buf_n552( .i (n551), .o (n552) );
  buffer buf_n4195( .i (n1315), .o (n4195) );
  assign n4196 = n552 & n4195 ;
  buffer buf_n4197( .i (n4196), .o (n4197) );
  buffer buf_n4198( .i (n4197), .o (n4198) );
  buffer buf_n594( .i (x84), .o (n594) );
  buffer buf_n595( .i (n594), .o (n595) );
  buffer buf_n596( .i (n595), .o (n596) );
  assign n4199 = n596 & ~n4195 ;
  buffer buf_n4200( .i (n4199), .o (n4200) );
  buffer buf_n4201( .i (n4200), .o (n4201) );
  assign n4202 = ( n4174 & n4198 ) | ( n4174 & n4201 ) | ( n4198 & n4201 ) ;
  buffer buf_n4203( .i (n4202), .o (n4203) );
  buffer buf_n4204( .i (n4203), .o (n4204) );
  buffer buf_n4205( .i (n4204), .o (n4205) );
  buffer buf_n4206( .i (n4205), .o (n4206) );
  buffer buf_n4207( .i (n4206), .o (n4207) );
  buffer buf_n4208( .i (n4207), .o (n4208) );
  buffer buf_n4209( .i (n4208), .o (n4209) );
  buffer buf_n4210( .i (n4209), .o (n4210) );
  buffer buf_n4211( .i (n4210), .o (n4211) );
  buffer buf_n4212( .i (n4211), .o (n4212) );
  buffer buf_n4213( .i (n4212), .o (n4213) );
  buffer buf_n4214( .i (n4213), .o (n4214) );
  buffer buf_n4215( .i (n4214), .o (n4215) );
  buffer buf_n4216( .i (n4215), .o (n4216) );
  buffer buf_n3223( .i (n3222), .o (n3223) );
  assign n4217 = n3223 | n4215 ;
  assign n4218 = ( n3786 & n4216 ) | ( n3786 & n4217 ) | ( n4216 & n4217 ) ;
  assign n4219 = n4194 | n4218 ;
  buffer buf_n4220( .i (n4219), .o (n4220) );
  assign n4221 = n3241 & ~n3888 ;
  buffer buf_n546( .i (x73), .o (n546) );
  buffer buf_n547( .i (n546), .o (n547) );
  buffer buf_n548( .i (n547), .o (n548) );
  assign n4222 = n548 & n4195 ;
  buffer buf_n4223( .i (n4222), .o (n4223) );
  buffer buf_n4224( .i (n4223), .o (n4224) );
  buffer buf_n590( .i (x83), .o (n590) );
  buffer buf_n591( .i (n590), .o (n591) );
  buffer buf_n592( .i (n591), .o (n592) );
  assign n4225 = n592 & ~n4195 ;
  buffer buf_n4226( .i (n4225), .o (n4226) );
  buffer buf_n4227( .i (n4226), .o (n4227) );
  assign n4228 = ( n4174 & n4224 ) | ( n4174 & n4227 ) | ( n4224 & n4227 ) ;
  buffer buf_n4229( .i (n4228), .o (n4229) );
  buffer buf_n4230( .i (n4229), .o (n4230) );
  buffer buf_n4231( .i (n4230), .o (n4231) );
  buffer buf_n4232( .i (n4231), .o (n4232) );
  buffer buf_n4233( .i (n4232), .o (n4233) );
  buffer buf_n4234( .i (n4233), .o (n4234) );
  buffer buf_n4235( .i (n4234), .o (n4235) );
  buffer buf_n4236( .i (n4235), .o (n4236) );
  buffer buf_n4237( .i (n4236), .o (n4237) );
  buffer buf_n4238( .i (n4237), .o (n4238) );
  buffer buf_n4239( .i (n4238), .o (n4239) );
  buffer buf_n4240( .i (n4239), .o (n4240) );
  buffer buf_n4241( .i (n4240), .o (n4241) );
  buffer buf_n4242( .i (n4241), .o (n4242) );
  assign n4243 = n3223 | n4241 ;
  assign n4244 = ( ~n3760 & n4242 ) | ( ~n3760 & n4243 ) | ( n4242 & n4243 ) ;
  assign n4245 = n4221 | n4244 ;
  buffer buf_n4246( .i (n4245), .o (n4246) );
  buffer buf_n3242( .i (n3241), .o (n3242) );
  assign n4247 = n3242 & n3867 ;
  buffer buf_n542( .i (x72), .o (n542) );
  buffer buf_n543( .i (n542), .o (n543) );
  buffer buf_n544( .i (n543), .o (n544) );
  buffer buf_n4248( .i (n1315), .o (n4248) );
  assign n4249 = n544 & n4248 ;
  buffer buf_n4250( .i (n4249), .o (n4250) );
  buffer buf_n4251( .i (n4250), .o (n4251) );
  buffer buf_n586( .i (x82), .o (n586) );
  buffer buf_n587( .i (n586), .o (n587) );
  buffer buf_n588( .i (n587), .o (n588) );
  assign n4252 = n588 & ~n4248 ;
  buffer buf_n4253( .i (n4252), .o (n4253) );
  buffer buf_n4254( .i (n4253), .o (n4254) );
  assign n4255 = ( n4174 & n4251 ) | ( n4174 & n4254 ) | ( n4251 & n4254 ) ;
  buffer buf_n4256( .i (n4255), .o (n4256) );
  buffer buf_n4257( .i (n4256), .o (n4257) );
  buffer buf_n4258( .i (n4257), .o (n4258) );
  buffer buf_n4259( .i (n4258), .o (n4259) );
  buffer buf_n4260( .i (n4259), .o (n4260) );
  buffer buf_n4261( .i (n4260), .o (n4261) );
  buffer buf_n4262( .i (n4261), .o (n4262) );
  buffer buf_n4263( .i (n4262), .o (n4263) );
  buffer buf_n4264( .i (n4263), .o (n4264) );
  buffer buf_n4265( .i (n4264), .o (n4265) );
  buffer buf_n4266( .i (n4265), .o (n4266) );
  buffer buf_n4267( .i (n4266), .o (n4267) );
  buffer buf_n4268( .i (n4267), .o (n4268) );
  buffer buf_n4269( .i (n4268), .o (n4269) );
  buffer buf_n4270( .i (n4269), .o (n4270) );
  buffer buf_n3224( .i (n3223), .o (n3224) );
  assign n4271 = n3224 | n4269 ;
  assign n4272 = ( n3738 & n4270 ) | ( n3738 & n4271 ) | ( n4270 & n4271 ) ;
  assign n4273 = n4247 | n4272 ;
  assign n4274 = n3302 & ~n4166 ;
  assign n4275 = n562 & n1326 ;
  assign n4276 = n606 & ~n1326 ;
  assign n4277 = ( n3307 & n4275 ) | ( n3307 & n4276 ) | ( n4275 & n4276 ) ;
  buffer buf_n4278( .i (n4277), .o (n4278) );
  buffer buf_n4279( .i (n4278), .o (n4279) );
  buffer buf_n4280( .i (n4279), .o (n4280) );
  buffer buf_n4281( .i (n4280), .o (n4281) );
  buffer buf_n4282( .i (n4281), .o (n4282) );
  buffer buf_n4283( .i (n4282), .o (n4283) );
  buffer buf_n4284( .i (n4283), .o (n4284) );
  buffer buf_n4285( .i (n4284), .o (n4285) );
  buffer buf_n4286( .i (n4285), .o (n4286) );
  buffer buf_n4287( .i (n4286), .o (n4287) );
  buffer buf_n4288( .i (n4287), .o (n4288) );
  buffer buf_n4289( .i (n4288), .o (n4289) );
  buffer buf_n4290( .i (n4289), .o (n4290) );
  buffer buf_n4291( .i (n4290), .o (n4291) );
  buffer buf_n4292( .i (n4291), .o (n4292) );
  buffer buf_n3281( .i (n3280), .o (n3281) );
  buffer buf_n3282( .i (n3281), .o (n3282) );
  buffer buf_n3283( .i (n3282), .o (n3283) );
  assign n4293 = n3283 | n4291 ;
  assign n4294 = ( n3808 & n4292 ) | ( n3808 & n4293 ) | ( n4292 & n4293 ) ;
  assign n4295 = n4274 | n4294 ;
  buffer buf_n4296( .i (n4295), .o (n4296) );
  buffer buf_n4297( .i (n4296), .o (n4297) );
  buffer buf_n3303( .i (n3302), .o (n3303) );
  assign n4298 = n3303 & ~n3910 ;
  buffer buf_n4299( .i (n1325), .o (n4299) );
  assign n4300 = n552 & n4299 ;
  assign n4301 = n596 & ~n4299 ;
  assign n4302 = ( n3307 & n4300 ) | ( n3307 & n4301 ) | ( n4300 & n4301 ) ;
  buffer buf_n4303( .i (n4302), .o (n4303) );
  buffer buf_n4304( .i (n4303), .o (n4304) );
  buffer buf_n4305( .i (n4304), .o (n4305) );
  buffer buf_n4306( .i (n4305), .o (n4306) );
  buffer buf_n4307( .i (n4306), .o (n4307) );
  buffer buf_n4308( .i (n4307), .o (n4308) );
  buffer buf_n4309( .i (n4308), .o (n4309) );
  buffer buf_n4310( .i (n4309), .o (n4310) );
  buffer buf_n4311( .i (n4310), .o (n4311) );
  buffer buf_n4312( .i (n4311), .o (n4312) );
  buffer buf_n4313( .i (n4312), .o (n4313) );
  buffer buf_n4314( .i (n4313), .o (n4314) );
  buffer buf_n4315( .i (n4314), .o (n4315) );
  buffer buf_n4316( .i (n4315), .o (n4316) );
  buffer buf_n4317( .i (n4316), .o (n4317) );
  buffer buf_n4318( .i (n4317), .o (n4318) );
  buffer buf_n3284( .i (n3283), .o (n3284) );
  assign n4319 = n3284 | n4317 ;
  assign n4320 = ( n3786 & n4318 ) | ( n3786 & n4319 ) | ( n4318 & n4319 ) ;
  assign n4321 = n4298 | n4320 ;
  buffer buf_n4322( .i (n4321), .o (n4322) );
  assign n4323 = n3303 & ~n3888 ;
  assign n4324 = n548 & n4299 ;
  buffer buf_n4325( .i (n4324), .o (n4325) );
  assign n4326 = n592 & ~n4299 ;
  buffer buf_n4327( .i (n4326), .o (n4327) );
  assign n4328 = ( n3308 & n4325 ) | ( n3308 & n4327 ) | ( n4325 & n4327 ) ;
  buffer buf_n4329( .i (n4328), .o (n4329) );
  buffer buf_n4330( .i (n4329), .o (n4330) );
  buffer buf_n4331( .i (n4330), .o (n4331) );
  buffer buf_n4332( .i (n4331), .o (n4332) );
  buffer buf_n4333( .i (n4332), .o (n4333) );
  buffer buf_n4334( .i (n4333), .o (n4334) );
  buffer buf_n4335( .i (n4334), .o (n4335) );
  buffer buf_n4336( .i (n4335), .o (n4336) );
  buffer buf_n4337( .i (n4336), .o (n4337) );
  buffer buf_n4338( .i (n4337), .o (n4338) );
  buffer buf_n4339( .i (n4338), .o (n4339) );
  buffer buf_n4340( .i (n4339), .o (n4340) );
  buffer buf_n4341( .i (n4340), .o (n4341) );
  buffer buf_n4342( .i (n4341), .o (n4342) );
  buffer buf_n4343( .i (n4342), .o (n4343) );
  assign n4344 = n3284 | n4342 ;
  assign n4345 = ( ~n3760 & n4343 ) | ( ~n3760 & n4344 ) | ( n4343 & n4344 ) ;
  assign n4346 = n4323 | n4345 ;
  buffer buf_n4347( .i (n4346), .o (n4347) );
  buffer buf_n3304( .i (n3303), .o (n3304) );
  assign n4348 = n3304 & n3867 ;
  buffer buf_n4349( .i (n1325), .o (n4349) );
  assign n4350 = n544 & n4349 ;
  buffer buf_n4351( .i (n4350), .o (n4351) );
  buffer buf_n4352( .i (n4351), .o (n4352) );
  assign n4353 = n588 & ~n4349 ;
  buffer buf_n4354( .i (n4353), .o (n4354) );
  buffer buf_n4355( .i (n4354), .o (n4355) );
  buffer buf_n4356( .i (n3308), .o (n4356) );
  assign n4357 = ( n4352 & n4355 ) | ( n4352 & n4356 ) | ( n4355 & n4356 ) ;
  buffer buf_n4358( .i (n4357), .o (n4358) );
  buffer buf_n4359( .i (n4358), .o (n4359) );
  buffer buf_n4360( .i (n4359), .o (n4360) );
  buffer buf_n4361( .i (n4360), .o (n4361) );
  buffer buf_n4362( .i (n4361), .o (n4362) );
  buffer buf_n4363( .i (n4362), .o (n4363) );
  buffer buf_n4364( .i (n4363), .o (n4364) );
  buffer buf_n4365( .i (n4364), .o (n4365) );
  buffer buf_n4366( .i (n4365), .o (n4366) );
  buffer buf_n4367( .i (n4366), .o (n4367) );
  buffer buf_n4368( .i (n4367), .o (n4368) );
  buffer buf_n4369( .i (n4368), .o (n4369) );
  buffer buf_n4370( .i (n4369), .o (n4370) );
  buffer buf_n4371( .i (n4370), .o (n4371) );
  buffer buf_n4372( .i (n4371), .o (n4372) );
  buffer buf_n3285( .i (n3284), .o (n3285) );
  assign n4373 = n3285 | n4371 ;
  assign n4374 = ( n3738 & n4372 ) | ( n3738 & n4373 ) | ( n4372 & n4373 ) ;
  assign n4375 = n4348 | n4374 ;
  buffer buf_n2765( .i (n2764), .o (n2765) );
  buffer buf_n2766( .i (n2765), .o (n2766) );
  buffer buf_n2767( .i (n2766), .o (n2767) );
  buffer buf_n2768( .i (n2767), .o (n2768) );
  buffer buf_n2651( .i (n2650), .o (n2651) );
  buffer buf_n2652( .i (n2651), .o (n2652) );
  buffer buf_n2413( .i (n2412), .o (n2413) );
  buffer buf_n1333( .i (x161), .o (n1333) );
  buffer buf_n1334( .i (n1333), .o (n1334) );
  buffer buf_n1335( .i (n1334), .o (n1335) );
  buffer buf_n1336( .i (n1335), .o (n1336) );
  buffer buf_n1337( .i (n1336), .o (n1337) );
  buffer buf_n1338( .i (n1337), .o (n1338) );
  buffer buf_n1339( .i (n1338), .o (n1339) );
  buffer buf_n1340( .i (n1339), .o (n1340) );
  buffer buf_n1341( .i (n1340), .o (n1341) );
  assign n4376 = ( n1341 & n2489 ) | ( n1341 & n2643 ) | ( n2489 & n2643 ) ;
  buffer buf_n4377( .i (n4376), .o (n4377) );
  assign n4380 = n2361 & n4377 ;
  assign n4381 = n2413 & n4380 ;
  assign n4382 = n2652 | n4381 ;
  buffer buf_n4383( .i (n4382), .o (n4383) );
  buffer buf_n2430( .i (n2429), .o (n2430) );
  buffer buf_n2431( .i (n2430), .o (n2431) );
  buffer buf_n2432( .i (n2431), .o (n2432) );
  buffer buf_n2433( .i (n2432), .o (n2433) );
  buffer buf_n2438( .i (n2437), .o (n2438) );
  buffer buf_n2439( .i (n2438), .o (n2439) );
  assign n4384 = n1117 & n2510 ;
  assign n4385 = n2439 & ~n4384 ;
  buffer buf_n4386( .i (n4385), .o (n4386) );
  assign n4387 = ( n1136 & n2433 ) | ( n1136 & n4386 ) | ( n2433 & n4386 ) ;
  assign n4388 = ( n1136 & ~n2433 ) | ( n1136 & n4386 ) | ( ~n2433 & n4386 ) ;
  assign n4389 = ~n4387 & n4388 ;
  buffer buf_n4390( .i (n4389), .o (n4390) );
  assign n4391 = ~n1134 & n2511 ;
  assign n4392 = n1134 & ~n2511 ;
  assign n4393 = ( n2432 & n4391 ) | ( n2432 & n4392 ) | ( n4391 & n4392 ) ;
  buffer buf_n4394( .i (n4393), .o (n4394) );
  buffer buf_n4395( .i (n4394), .o (n4395) );
  assign n4397 = n2462 & ~n4395 ;
  assign n4398 = ~n4390 & n4397 ;
  assign n4399 = n4383 | n4398 ;
  buffer buf_n2434( .i (n2433), .o (n2434) );
  buffer buf_n2435( .i (n2434), .o (n2435) );
  buffer buf_n2440( .i (n2439), .o (n2440) );
  buffer buf_n2441( .i (n2440), .o (n2441) );
  buffer buf_n2442( .i (n2441), .o (n2442) );
  assign n4400 = ( ~n1137 & n2442 ) | ( ~n1137 & n4394 ) | ( n2442 & n4394 ) ;
  assign n4401 = ( n1137 & ~n2447 ) | ( n1137 & n4394 ) | ( ~n2447 & n4394 ) ;
  assign n4402 = ( ~n2435 & n4400 ) | ( ~n2435 & n4401 ) | ( n4400 & n4401 ) ;
  buffer buf_n4403( .i (n4402), .o (n4403) );
  assign n4404 = n1124 & n4403 ;
  assign n4405 = ( n1124 & ~n2464 ) | ( n1124 & n4403 ) | ( ~n2464 & n4403 ) ;
  assign n4406 = ( n4399 & ~n4404 ) | ( n4399 & n4405 ) | ( ~n4404 & n4405 ) ;
  buffer buf_n4407( .i (n4406), .o (n4407) );
  buffer buf_n1171( .i (n1170), .o (n1171) );
  buffer buf_n1172( .i (n1171), .o (n1172) );
  buffer buf_n1173( .i (n1172), .o (n1173) );
  buffer buf_n1174( .i (n1173), .o (n1174) );
  buffer buf_n1175( .i (n1174), .o (n1175) );
  buffer buf_n1176( .i (n1175), .o (n1176) );
  buffer buf_n1177( .i (n1176), .o (n1177) );
  buffer buf_n4378( .i (n4377), .o (n4378) );
  buffer buf_n4379( .i (n4378), .o (n4379) );
  buffer buf_n2377( .i (n2376), .o (n2377) );
  buffer buf_n2378( .i (n2377), .o (n2378) );
  buffer buf_n2379( .i (n2378), .o (n2379) );
  assign n4408 = ~n2379 & n2409 ;
  buffer buf_n4409( .i (n4408), .o (n4409) );
  buffer buf_n2383( .i (n2382), .o (n2383) );
  buffer buf_n2384( .i (n2383), .o (n2384) );
  buffer buf_n2403( .i (n2402), .o (n2403) );
  assign n4410 = ~n2384 & n2403 ;
  buffer buf_n4411( .i (n4410), .o (n4411) );
  buffer buf_n4412( .i (n4411), .o (n4412) );
  buffer buf_n1160( .i (n1159), .o (n1160) );
  assign n4413 = ( n1160 & n2377 ) | ( n1160 & ~n2384 ) | ( n2377 & ~n2384 ) ;
  assign n4414 = n1147 | n1159 ;
  assign n4415 = n2370 & ~n4414 ;
  assign n4416 = ( n2408 & ~n4413 ) | ( n2408 & n4415 ) | ( ~n4413 & n4415 ) ;
  buffer buf_n4417( .i (n4416), .o (n4417) );
  assign n4418 = ( n2390 & n4412 ) | ( n2390 & n4417 ) | ( n4412 & n4417 ) ;
  assign n4419 = ( n4379 & n4409 ) | ( n4379 & n4418 ) | ( n4409 & n4418 ) ;
  buffer buf_n4420( .i (n4419), .o (n4420) );
  assign n4421 = n949 & n1335 ;
  buffer buf_n4422( .i (n4421), .o (n4422) );
  assign n4423 = ( n849 & ~n2547 ) | ( n849 & n4422 ) | ( ~n2547 & n4422 ) ;
  buffer buf_n4424( .i (n2481), .o (n4424) );
  assign n4425 = ( n2547 & ~n4422 ) | ( n2547 & n4424 ) | ( ~n4422 & n4424 ) ;
  assign n4426 = n4423 | n4425 ;
  buffer buf_n3093( .i (n3092), .o (n3093) );
  assign n4427 = n954 & n1335 ;
  buffer buf_n4428( .i (n4427), .o (n4428) );
  buffer buf_n4429( .i (n4428), .o (n4429) );
  assign n4430 = n3093 & ~n4429 ;
  assign n4431 = ( n850 & n3093 ) | ( n850 & ~n4429 ) | ( n3093 & ~n4429 ) ;
  assign n4432 = ( n4426 & n4430 ) | ( n4426 & ~n4431 ) | ( n4430 & ~n4431 ) ;
  buffer buf_n4433( .i (n4432), .o (n4433) );
  buffer buf_n4434( .i (n4433), .o (n4434) );
  buffer buf_n4435( .i (n4434), .o (n4435) );
  buffer buf_n4436( .i (n4435), .o (n4436) );
  buffer buf_n4437( .i (n4436), .o (n4437) );
  buffer buf_n4438( .i (n4437), .o (n4438) );
  assign n4439 = ( ~n2389 & n2409 ) | ( ~n2389 & n4377 ) | ( n2409 & n4377 ) ;
  buffer buf_n4440( .i (n2408), .o (n4440) );
  assign n4441 = ( n4377 & ~n4411 ) | ( n4377 & n4440 ) | ( ~n4411 & n4440 ) ;
  assign n4442 = ( ~n4417 & n4439 ) | ( ~n4417 & n4441 ) | ( n4439 & n4441 ) ;
  buffer buf_n4443( .i (n4442), .o (n4443) );
  assign n4444 = ( ~n1175 & n4438 ) | ( ~n1175 & n4443 ) | ( n4438 & n4443 ) ;
  assign n4445 = n2389 & ~n4440 ;
  assign n4446 = n4411 & ~n4440 ;
  assign n4447 = ( n4417 & n4445 ) | ( n4417 & n4446 ) | ( n4445 & n4446 ) ;
  buffer buf_n4448( .i (n4447), .o (n4448) );
  assign n4449 = ( ~n1175 & n4438 ) | ( ~n1175 & n4448 ) | ( n4438 & n4448 ) ;
  assign n4450 = ( ~n4420 & n4444 ) | ( ~n4420 & n4449 ) | ( n4444 & n4449 ) ;
  assign n4451 = ( n1175 & n4438 ) | ( n1175 & n4443 ) | ( n4438 & n4443 ) ;
  buffer buf_n4452( .i (n1174), .o (n4452) );
  assign n4453 = ( n4438 & n4448 ) | ( n4438 & n4452 ) | ( n4448 & n4452 ) ;
  assign n4454 = ( ~n4420 & n4451 ) | ( ~n4420 & n4453 ) | ( n4451 & n4453 ) ;
  assign n4455 = ( n1177 & n4450 ) | ( n1177 & ~n4454 ) | ( n4450 & ~n4454 ) ;
  buffer buf_n4456( .i (n4455), .o (n4456) );
  assign n4457 = n2462 & n2515 ;
  assign n4458 = n4390 & ~n4457 ;
  buffer buf_n4396( .i (n4395), .o (n4396) );
  assign n4459 = n1136 & n2513 ;
  assign n4460 = ~n2434 & n4459 ;
  assign n4461 = ( n2462 & n2524 ) | ( n2462 & n4460 ) | ( n2524 & n4460 ) ;
  assign n4462 = n4396 | n4461 ;
  assign n4463 = n4458 | n4462 ;
  assign n4464 = n2524 & n4395 ;
  assign n4465 = ( n2525 & n4390 ) | ( n2525 & n4464 ) | ( n4390 & n4464 ) ;
  assign n4466 = n4383 & ~n4465 ;
  assign n4467 = n4463 & n4466 ;
  buffer buf_n4468( .i (n4467), .o (n4468) );
  assign n4469 = ( n4407 & n4456 ) | ( n4407 & ~n4468 ) | ( n4456 & ~n4468 ) ;
  assign n4470 = ~n4407 & n4456 ;
  assign n4471 = n4456 & ~n4468 ;
  assign n4472 = ( n4469 & n4470 ) | ( n4469 & ~n4471 ) | ( n4470 & ~n4471 ) ;
  buffer buf_n4473( .i (n4472), .o (n4473) );
  assign n4475 = n2768 & ~n4473 ;
  buffer buf_n355( .i (x50), .o (n355) );
  buffer buf_n356( .i (n355), .o (n356) );
  buffer buf_n357( .i (n356), .o (n357) );
  buffer buf_n358( .i (n357), .o (n358) );
  buffer buf_n359( .i (n358), .o (n359) );
  buffer buf_n360( .i (n359), .o (n360) );
  buffer buf_n361( .i (n360), .o (n361) );
  assign n4476 = ~n361 & n3765 ;
  buffer buf_n4477( .i (n4476), .o (n4477) );
  buffer buf_n4478( .i (n4477), .o (n4478) );
  buffer buf_n4479( .i (n4478), .o (n4479) );
  buffer buf_n4480( .i (n4479), .o (n4480) );
  buffer buf_n4481( .i (n4480), .o (n4481) );
  buffer buf_n4482( .i (n4481), .o (n4482) );
  buffer buf_n4483( .i (n4482), .o (n4483) );
  buffer buf_n4484( .i (n4483), .o (n4484) );
  buffer buf_n4485( .i (n655), .o (n4485) );
  assign n4486 = n1128 | n4485 ;
  assign n4487 = n1128 & n1913 ;
  assign n4488 = ( n837 & ~n4486 ) | ( n837 & n4487 ) | ( ~n4486 & n4487 ) ;
  buffer buf_n4489( .i (n699), .o (n4489) );
  buffer buf_n4490( .i (n1127), .o (n4490) );
  assign n4491 = n4489 | n4490 ;
  assign n4492 = n1915 & n4490 ;
  assign n4493 = ( n837 & n4491 ) | ( n837 & ~n4492 ) | ( n4491 & ~n4492 ) ;
  assign n4494 = ~n4488 & n4493 ;
  buffer buf_n4495( .i (n4494), .o (n4495) );
  buffer buf_n4496( .i (n4495), .o (n4496) );
  assign n4497 = n919 & ~n1913 ;
  assign n4498 = n919 | n1915 ;
  assign n4499 = ( n1165 & n4497 ) | ( n1165 & ~n4498 ) | ( n4497 & ~n4498 ) ;
  buffer buf_n4500( .i (n918), .o (n4500) );
  assign n4501 = n4489 & ~n4500 ;
  assign n4502 = n4485 & n4500 ;
  assign n4503 = ( ~n1165 & n4501 ) | ( ~n1165 & n4502 ) | ( n4501 & n4502 ) ;
  assign n4504 = n4499 | n4503 ;
  buffer buf_n4505( .i (n4504), .o (n4505) );
  assign n4506 = ~n1154 & n4485 ;
  assign n4507 = n1154 & ~n1913 ;
  assign n4508 = ( n889 & n4506 ) | ( n889 & n4507 ) | ( n4506 & n4507 ) ;
  buffer buf_n4509( .i (n1153), .o (n4509) );
  assign n4510 = n4489 & ~n4509 ;
  assign n4511 = ~n1915 & n4509 ;
  buffer buf_n4512( .i (n888), .o (n4512) );
  assign n4513 = ( n4510 & n4511 ) | ( n4510 & ~n4512 ) | ( n4511 & ~n4512 ) ;
  assign n4514 = n4508 | n4513 ;
  buffer buf_n4515( .i (n4514), .o (n4515) );
  assign n4516 = ( n4495 & n4505 ) | ( n4495 & n4515 ) | ( n4505 & n4515 ) ;
  assign n4517 = ( ~n4495 & n4505 ) | ( ~n4495 & n4515 ) | ( n4505 & n4515 ) ;
  assign n4518 = ( n4496 & ~n4516 ) | ( n4496 & n4517 ) | ( ~n4516 & n4517 ) ;
  buffer buf_n4519( .i (n4518), .o (n4519) );
  buffer buf_n4520( .i (n4519), .o (n4520) );
  assign n4521 = n800 & n948 ;
  buffer buf_n4522( .i (n4521), .o (n4522) );
  assign n4523 = ( n688 & n695 ) | ( n688 & n4522 ) | ( n695 & n4522 ) ;
  assign n4524 = n800 | n948 ;
  buffer buf_n4525( .i (n4524), .o (n4525) );
  assign n4526 = ( n688 & n695 ) | ( n688 & n4525 ) | ( n695 & n4525 ) ;
  assign n4527 = ~n4523 & n4526 ;
  buffer buf_n4528( .i (n4527), .o (n4528) );
  assign n4529 = ( ~n1880 & n1891 ) | ( ~n1880 & n4528 ) | ( n1891 & n4528 ) ;
  assign n4530 = ( n1880 & n1891 ) | ( n1880 & n4528 ) | ( n1891 & n4528 ) ;
  assign n4531 = ( n1881 & n4529 ) | ( n1881 & ~n4530 ) | ( n4529 & ~n4530 ) ;
  buffer buf_n4532( .i (n4531), .o (n4532) );
  buffer buf_n658( .i (n657), .o (n658) );
  buffer buf_n702( .i (n701), .o (n702) );
  assign n4533 = n658 | n702 ;
  assign n4534 = ( n658 & n702 ) | ( n658 & n753 ) | ( n702 & n753 ) ;
  assign n4535 = ( n1145 & n4533 ) | ( n1145 & ~n4534 ) | ( n4533 & ~n4534 ) ;
  buffer buf_n689( .i (n688), .o (n689) );
  buffer buf_n690( .i (n689), .o (n690) );
  assign n4536 = n690 | n1922 ;
  assign n4537 = ( n690 & ~n1145 ) | ( n690 & n1922 ) | ( ~n1145 & n1922 ) ;
  assign n4538 = ( n4535 & ~n4536 ) | ( n4535 & n4537 ) | ( ~n4536 & n4537 ) ;
  buffer buf_n4539( .i (n4538), .o (n4539) );
  buffer buf_n4540( .i (n4539), .o (n4540) );
  assign n4541 = ( n4519 & n4532 ) | ( n4519 & n4540 ) | ( n4532 & n4540 ) ;
  assign n4542 = ( ~n4519 & n4532 ) | ( ~n4519 & n4540 ) | ( n4532 & n4540 ) ;
  assign n4543 = ( n4520 & ~n4541 ) | ( n4520 & n4542 ) | ( ~n4541 & n4542 ) ;
  buffer buf_n4544( .i (n4543), .o (n4544) );
  buffer buf_n4545( .i (n4544), .o (n4545) );
  buffer buf_n4546( .i (n4545), .o (n4546) );
  assign n4547 = n2677 | n4546 ;
  assign n4548 = ~n4484 & n4547 ;
  buffer buf_n4549( .i (n4548), .o (n4549) );
  buffer buf_n4550( .i (n4549), .o (n4550) );
  buffer buf_n4551( .i (n4550), .o (n4551) );
  buffer buf_n4552( .i (n4551), .o (n4552) );
  buffer buf_n4553( .i (n4552), .o (n4553) );
  assign n4554 = ~n4475 & n4553 ;
  buffer buf_n4555( .i (n4554), .o (n4555) );
  buffer buf_n343( .i (x48), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  buffer buf_n346( .i (n345), .o (n346) );
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  buffer buf_n349( .i (n348), .o (n349) );
  assign n4556 = n349 | n1512 ;
  buffer buf_n4557( .i (n4556), .o (n4557) );
  assign n4558 = n1531 & n4557 ;
  buffer buf_n4559( .i (n4558), .o (n4559) );
  buffer buf_n4560( .i (n4559), .o (n4560) );
  buffer buf_n4561( .i (n4560), .o (n4561) );
  buffer buf_n4562( .i (n4561), .o (n4562) );
  buffer buf_n4563( .i (n4562), .o (n4563) );
  buffer buf_n4564( .i (n4563), .o (n4564) );
  buffer buf_n4565( .i (n4564), .o (n4565) );
  buffer buf_n4566( .i (n4565), .o (n4566) );
  buffer buf_n4567( .i (n4566), .o (n4567) );
  buffer buf_n4568( .i (n4567), .o (n4568) );
  buffer buf_n4569( .i (n4568), .o (n4569) );
  assign n4570 = n689 & n708 ;
  buffer buf_n696( .i (n695), .o (n696) );
  buffer buf_n4571( .i (n2041), .o (n4571) );
  assign n4572 = n696 & ~n4571 ;
  assign n4573 = ( n1010 & n4570 ) | ( n1010 & n4572 ) | ( n4570 & n4572 ) ;
  assign n4574 = n702 | n4571 ;
  assign n4575 = ~n658 & n4571 ;
  assign n4576 = ( n1010 & n4574 ) | ( n1010 & ~n4575 ) | ( n4574 & ~n4575 ) ;
  assign n4577 = ~n4573 & n4576 ;
  buffer buf_n4578( .i (n4577), .o (n4578) );
  buffer buf_n4579( .i (n4578), .o (n4579) );
  buffer buf_n4580( .i (n4579), .o (n4580) );
  buffer buf_n631( .i (n630), .o (n631) );
  assign n4581 = n631 & ~n689 ;
  assign n4582 = n631 | n696 ;
  assign n4583 = ( n1093 & n4581 ) | ( n1093 & ~n4582 ) | ( n4581 & ~n4582 ) ;
  assign n4584 = ~n631 & n702 ;
  assign n4585 = n631 & n658 ;
  buffer buf_n4586( .i (n1092), .o (n4586) );
  assign n4587 = ( n4584 & n4585 ) | ( n4584 & ~n4586 ) | ( n4585 & ~n4586 ) ;
  assign n4588 = n4583 | n4587 ;
  buffer buf_n4589( .i (n4588), .o (n4589) );
  buffer buf_n4590( .i (n4589), .o (n4590) );
  buffer buf_n4591( .i (n686), .o (n4591) );
  assign n4592 = n735 & n4591 ;
  buffer buf_n4593( .i (n693), .o (n4593) );
  assign n4594 = ~n735 & n4593 ;
  assign n4595 = ( n997 & n4592 ) | ( n997 & n4594 ) | ( n4592 & n4594 ) ;
  buffer buf_n4596( .i (n734), .o (n4596) );
  assign n4597 = n4489 | n4596 ;
  assign n4598 = ~n4485 & n4596 ;
  assign n4599 = ( n997 & n4597 ) | ( n997 & ~n4598 ) | ( n4597 & ~n4598 ) ;
  assign n4600 = ~n4595 & n4599 ;
  buffer buf_n4601( .i (n4600), .o (n4601) );
  assign n4602 = n655 & ~n1029 ;
  assign n4603 = ~n686 & n1029 ;
  assign n4604 = ( n724 & n4602 ) | ( n724 & n4603 ) | ( n4602 & n4603 ) ;
  assign n4605 = n699 & ~n1029 ;
  buffer buf_n4606( .i (n1028), .o (n4606) );
  assign n4607 = ~n693 & n4606 ;
  assign n4608 = ( ~n724 & n4605 ) | ( ~n724 & n4607 ) | ( n4605 & n4607 ) ;
  assign n4609 = n4604 | n4608 ;
  buffer buf_n4610( .i (n4609), .o (n4610) );
  buffer buf_n4611( .i (n4610), .o (n4611) );
  assign n4612 = ~n4601 & n4611 ;
  assign n4613 = n4601 & ~n4611 ;
  assign n4614 = n4612 | n4613 ;
  buffer buf_n4615( .i (n4614), .o (n4615) );
  assign n4616 = ( n4579 & n4590 ) | ( n4579 & n4615 ) | ( n4590 & n4615 ) ;
  assign n4617 = ( ~n4579 & n4590 ) | ( ~n4579 & n4615 ) | ( n4590 & n4615 ) ;
  assign n4618 = ( n4580 & ~n4616 ) | ( n4580 & n4617 ) | ( ~n4616 & n4617 ) ;
  buffer buf_n4619( .i (n4618), .o (n4619) );
  buffer buf_n2021( .i (n2020), .o (n2021) );
  buffer buf_n2022( .i (n2021), .o (n2022) );
  buffer buf_n2023( .i (n2022), .o (n2023) );
  assign n4620 = n639 & ~n4591 ;
  assign n4621 = n639 | n4593 ;
  assign n4622 = ( n1042 & n4620 ) | ( n1042 & ~n4621 ) | ( n4620 & ~n4621 ) ;
  buffer buf_n4623( .i (n699), .o (n4623) );
  assign n4624 = ~n639 & n4623 ;
  buffer buf_n4625( .i (n638), .o (n4625) );
  buffer buf_n4626( .i (n655), .o (n4626) );
  assign n4627 = n4625 & n4626 ;
  assign n4628 = ( ~n1042 & n4624 ) | ( ~n1042 & n4627 ) | ( n4624 & n4627 ) ;
  assign n4629 = n4622 | n4628 ;
  buffer buf_n4630( .i (n4629), .o (n4630) );
  buffer buf_n4631( .i (n4630), .o (n4631) );
  assign n4632 = n620 & ~n4591 ;
  assign n4633 = n620 | n4593 ;
  assign n4634 = ( n1083 & n4632 ) | ( n1083 & ~n4633 ) | ( n4632 & ~n4633 ) ;
  buffer buf_n4635( .i (n619), .o (n4635) );
  assign n4636 = n4623 & ~n4635 ;
  assign n4637 = n4626 & n4635 ;
  assign n4638 = ( ~n1083 & n4636 ) | ( ~n1083 & n4637 ) | ( n4636 & n4637 ) ;
  assign n4639 = n4634 | n4638 ;
  buffer buf_n4640( .i (n4639), .o (n4640) );
  assign n4641 = n716 & ~n4591 ;
  assign n4642 = n716 | n4593 ;
  assign n4643 = ( n1021 & n4641 ) | ( n1021 & ~n4642 ) | ( n4641 & ~n4642 ) ;
  buffer buf_n4644( .i (n715), .o (n4644) );
  assign n4645 = n4623 & ~n4644 ;
  assign n4646 = n4626 & n4644 ;
  assign n4647 = ( ~n1021 & n4645 ) | ( ~n1021 & n4646 ) | ( n4645 & n4646 ) ;
  assign n4648 = n4643 | n4647 ;
  buffer buf_n4649( .i (n4648), .o (n4649) );
  assign n4650 = ( ~n4630 & n4640 ) | ( ~n4630 & n4649 ) | ( n4640 & n4649 ) ;
  assign n4651 = ( n4630 & n4640 ) | ( n4630 & n4649 ) | ( n4640 & n4649 ) ;
  assign n4652 = ( n4631 & n4650 ) | ( n4631 & ~n4651 ) | ( n4650 & ~n4651 ) ;
  buffer buf_n4653( .i (n4652), .o (n4653) );
  assign n4654 = n649 & n689 ;
  assign n4655 = ~n649 & n696 ;
  assign n4656 = ( n1059 & n4654 ) | ( n1059 & n4655 ) | ( n4654 & n4655 ) ;
  buffer buf_n4657( .i (n701), .o (n4657) );
  assign n4658 = n649 | n4657 ;
  buffer buf_n4659( .i (n1998), .o (n4659) );
  buffer buf_n4660( .i (n657), .o (n4660) );
  assign n4661 = n4659 & ~n4660 ;
  assign n4662 = ( n1059 & n4658 ) | ( n1059 & ~n4661 ) | ( n4658 & ~n4661 ) ;
  assign n4663 = ~n4656 & n4662 ;
  buffer buf_n4664( .i (n4663), .o (n4664) );
  buffer buf_n4665( .i (n4664), .o (n4665) );
  assign n4666 = ( ~n2022 & n4653 ) | ( ~n2022 & n4665 ) | ( n4653 & n4665 ) ;
  assign n4667 = ( n2022 & n4653 ) | ( n2022 & n4665 ) | ( n4653 & n4665 ) ;
  assign n4668 = ( n2023 & n4666 ) | ( n2023 & ~n4667 ) | ( n4666 & ~n4667 ) ;
  buffer buf_n4669( .i (n4668), .o (n4669) );
  assign n4670 = ( ~n2675 & n4619 ) | ( ~n2675 & n4669 ) | ( n4619 & n4669 ) ;
  assign n4671 = ( n2675 & n4619 ) | ( n2675 & n4669 ) | ( n4619 & n4669 ) ;
  assign n4672 = n4670 & ~n4671 ;
  buffer buf_n4673( .i (n4672), .o (n4673) );
  buffer buf_n4674( .i (n4673), .o (n4674) );
  buffer buf_n4675( .i (n4674), .o (n4675) );
  assign n4676 = ~n2112 & n2155 ;
  buffer buf_n4677( .i (n4676), .o (n4677) );
  buffer buf_n2084( .i (n2083), .o (n2084) );
  buffer buf_n1305( .i (x156), .o (n1305) );
  buffer buf_n1306( .i (n1305), .o (n1306) );
  buffer buf_n1307( .i (n1306), .o (n1307) );
  buffer buf_n1308( .i (n1307), .o (n1308) );
  buffer buf_n1309( .i (n1308), .o (n1309) );
  assign n4678 = n998 & n1309 ;
  assign n4679 = n2122 & n4678 ;
  buffer buf_n4680( .i (n4679), .o (n4680) );
  buffer buf_n1310( .i (n1309), .o (n1310) );
  assign n4682 = n999 | n1310 ;
  assign n4683 = n2123 | n4682 ;
  assign n4684 = ~n4680 & n4683 ;
  buffer buf_n4685( .i (n4684), .o (n4685) );
  assign n4687 = n2084 & ~n4685 ;
  buffer buf_n4681( .i (n4680), .o (n4681) );
  buffer buf_n1311( .i (n1310), .o (n1311) );
  buffer buf_n1312( .i (n1311), .o (n1312) );
  assign n4688 = ( n1001 & n1312 ) | ( n1001 & n2124 ) | ( n1312 & n2124 ) ;
  assign n4689 = ~n4681 & n4688 ;
  assign n4690 = ~n2084 & n4689 ;
  assign n4691 = ( ~n4677 & n4687 ) | ( ~n4677 & n4690 ) | ( n4687 & n4690 ) ;
  buffer buf_n4686( .i (n4685), .o (n4686) );
  assign n4692 = n2087 | n4686 ;
  assign n4693 = n2086 & n4685 ;
  assign n4694 = ( n1036 & n2076 ) | ( n1036 & n2125 ) | ( n2076 & n2125 ) ;
  assign n4695 = ( n2086 & n4685 ) | ( n2086 & n4694 ) | ( n4685 & n4694 ) ;
  assign n4696 = ( ~n4677 & n4693 ) | ( ~n4677 & n4695 ) | ( n4693 & n4695 ) ;
  assign n4697 = ( n4691 & n4692 ) | ( n4691 & ~n4696 ) | ( n4692 & ~n4696 ) ;
  buffer buf_n4698( .i (n4697), .o (n4698) );
  assign n4699 = ~n2279 & n4698 ;
  buffer buf_n2624( .i (n2623), .o (n2624) );
  assign n4700 = n2624 & ~n4698 ;
  assign n4701 = ~n2161 & n2623 ;
  assign n4702 = ( n2279 & ~n4698 ) | ( n2279 & n4701 ) | ( ~n4698 & n4701 ) ;
  assign n4703 = ( n4699 & ~n4700 ) | ( n4699 & n4702 ) | ( ~n4700 & n4702 ) ;
  buffer buf_n4704( .i (n4703), .o (n4704) );
  buffer buf_n2314( .i (n2313), .o (n2314) );
  buffer buf_n2191( .i (n2190), .o (n2191) );
  assign n4705 = ( n2191 & ~n2268 ) | ( n2191 & n2604 ) | ( ~n2268 & n2604 ) ;
  buffer buf_n4706( .i (n4705), .o (n4706) );
  buffer buf_n2266( .i (n2265), .o (n2266) );
  assign n4707 = ( n1086 & ~n1094 ) | ( n1086 & n2206 ) | ( ~n1094 & n2206 ) ;
  assign n4708 = ( n1086 & ~n2186 ) | ( n1086 & n2206 ) | ( ~n2186 & n2206 ) ;
  assign n4709 = ( ~n2266 & n4707 ) | ( ~n2266 & n4708 ) | ( n4707 & n4708 ) ;
  buffer buf_n4710( .i (n4709), .o (n4710) );
  assign n4711 = ( n2284 & ~n2626 ) | ( n2284 & n4710 ) | ( ~n2626 & n4710 ) ;
  assign n4712 = ~n2188 & n2259 ;
  buffer buf_n4713( .i (n4712), .o (n4713) );
  assign n4714 = ( n2284 & n4710 ) | ( n2284 & n4713 ) | ( n4710 & n4713 ) ;
  assign n4715 = ( n4706 & n4711 ) | ( n4706 & n4714 ) | ( n4711 & n4714 ) ;
  buffer buf_n4716( .i (n2283), .o (n4716) );
  assign n4717 = ( n2626 & ~n4710 ) | ( n2626 & n4716 ) | ( ~n4710 & n4716 ) ;
  assign n4718 = ( n4710 & n4713 ) | ( n4710 & ~n4716 ) | ( n4713 & ~n4716 ) ;
  assign n4719 = ( n4706 & ~n4717 ) | ( n4706 & n4718 ) | ( ~n4717 & n4718 ) ;
  assign n4720 = ( n2286 & ~n4715 ) | ( n2286 & n4719 ) | ( ~n4715 & n4719 ) ;
  buffer buf_n4721( .i (n4720), .o (n4721) );
  buffer buf_n2614( .i (n2613), .o (n2614) );
  buffer buf_n2615( .i (n2614), .o (n2615) );
  buffer buf_n2620( .i (n2619), .o (n2620) );
  assign n4722 = ( n2105 & ~n2157 ) | ( n2105 & n2620 ) | ( ~n2157 & n2620 ) ;
  buffer buf_n2109( .i (n2108), .o (n2109) );
  buffer buf_n2110( .i (n2109), .o (n2110) );
  assign n4723 = ~n2110 & n2150 ;
  buffer buf_n4724( .i (n4723), .o (n4724) );
  buffer buf_n4725( .i (n4724), .o (n4725) );
  assign n4726 = ( ~n2615 & n4722 ) | ( ~n2615 & n4725 ) | ( n4722 & n4725 ) ;
  buffer buf_n4727( .i (n4726), .o (n4727) );
  assign n4728 = ( n2313 & n4721 ) | ( n2313 & n4727 ) | ( n4721 & n4727 ) ;
  assign n4729 = ( ~n2313 & n4721 ) | ( ~n2313 & n4727 ) | ( n4721 & n4727 ) ;
  assign n4730 = ( n2314 & ~n4728 ) | ( n2314 & n4729 ) | ( ~n4728 & n4729 ) ;
  buffer buf_n4731( .i (n4730), .o (n4731) );
  assign n4732 = n4704 | n4731 ;
  assign n4733 = ( ~n2764 & n4704 ) | ( ~n2764 & n4731 ) | ( n4704 & n4731 ) ;
  assign n4734 = ( n4675 & n4732 ) | ( n4675 & ~n4733 ) | ( n4732 & ~n4733 ) ;
  buffer buf_n4735( .i (n4734), .o (n4735) );
  buffer buf_n4736( .i (n4735), .o (n4736) );
  assign n4737 = n4569 | n4736 ;
  buffer buf_n4738( .i (n4737), .o (n4738) );
  buffer buf_n4739( .i (n4738), .o (n4739) );
  buffer buf_n266( .i (x37), .o (n266) );
  assign n4740 = ~n266 & n1523 ;
  buffer buf_n4741( .i (n4740), .o (n4741) );
  buffer buf_n4742( .i (n4741), .o (n4742) );
  buffer buf_n4743( .i (n4742), .o (n4743) );
  buffer buf_n4744( .i (n4743), .o (n4744) );
  buffer buf_n4745( .i (n4744), .o (n4745) );
  buffer buf_n4746( .i (n4745), .o (n4746) );
  buffer buf_n4747( .i (n4746), .o (n4747) );
  buffer buf_n4748( .i (n4747), .o (n4748) );
  buffer buf_n4749( .i (n4748), .o (n4749) );
  buffer buf_n4750( .i (n4749), .o (n4750) );
  buffer buf_n4751( .i (n4750), .o (n4751) );
  buffer buf_n4752( .i (n4751), .o (n4752) );
  buffer buf_n4753( .i (n4752), .o (n4753) );
  buffer buf_n4754( .i (n4753), .o (n4754) );
  buffer buf_n4755( .i (n4754), .o (n4755) );
  buffer buf_n4756( .i (n4755), .o (n4756) );
  buffer buf_n4757( .i (n4756), .o (n4757) );
  buffer buf_n4758( .i (n4757), .o (n4758) );
  assign n4759 = n4735 | n4758 ;
  assign n4760 = n2831 & n4759 ;
  buffer buf_n4761( .i (n4760), .o (n4761) );
  buffer buf_n47( .i (x3), .o (n47) );
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  assign n4762 = n49 | n4035 ;
  buffer buf_n155( .i (x22), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  buffer buf_n157( .i (n156), .o (n157) );
  assign n4763 = ~n157 & n4035 ;
  assign n4764 = ( n4037 & ~n4762 ) | ( n4037 & n4763 ) | ( ~n4762 & n4763 ) ;
  buffer buf_n4765( .i (n4764), .o (n4765) );
  buffer buf_n4766( .i (n4765), .o (n4766) );
  buffer buf_n4767( .i (n4766), .o (n4767) );
  buffer buf_n4768( .i (n4767), .o (n4768) );
  buffer buf_n4769( .i (n4768), .o (n4769) );
  buffer buf_n4770( .i (n4769), .o (n4770) );
  buffer buf_n4771( .i (n4770), .o (n4771) );
  buffer buf_n4772( .i (n4771), .o (n4772) );
  buffer buf_n4773( .i (n4772), .o (n4773) );
  buffer buf_n4774( .i (n4773), .o (n4774) );
  buffer buf_n4775( .i (n4774), .o (n4775) );
  buffer buf_n4776( .i (n4775), .o (n4776) );
  buffer buf_n4777( .i (n4776), .o (n4777) );
  buffer buf_n4778( .i (n4777), .o (n4778) );
  buffer buf_n4779( .i (n4778), .o (n4779) );
  buffer buf_n4780( .i (n4779), .o (n4780) );
  buffer buf_n4781( .i (n4780), .o (n4781) );
  buffer buf_n255( .i (x36), .o (n255) );
  buffer buf_n256( .i (n255), .o (n256) );
  buffer buf_n257( .i (n256), .o (n257) );
  buffer buf_n258( .i (n257), .o (n258) );
  buffer buf_n259( .i (n258), .o (n259) );
  buffer buf_n260( .i (n259), .o (n260) );
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  assign n4782 = ~n264 & n1532 ;
  buffer buf_n4783( .i (n4782), .o (n4783) );
  buffer buf_n4784( .i (n4783), .o (n4784) );
  assign n4785 = n2674 & ~n4783 ;
  assign n4786 = ( n4544 & n4784 ) | ( n4544 & ~n4785 ) | ( n4784 & ~n4785 ) ;
  buffer buf_n4787( .i (n4786), .o (n4787) );
  buffer buf_n4788( .i (n4787), .o (n4788) );
  buffer buf_n4789( .i (n4788), .o (n4789) );
  buffer buf_n4790( .i (n4789), .o (n4790) );
  buffer buf_n4791( .i (n4790), .o (n4791) );
  buffer buf_n4792( .i (n4791), .o (n4792) );
  buffer buf_n4793( .i (n4792), .o (n4793) );
  assign n4794 = n2767 | n4792 ;
  assign n4795 = ( n4473 & n4793 ) | ( n4473 & n4794 ) | ( n4793 & n4794 ) ;
  assign n4796 = n2821 & ~n4780 ;
  assign n4797 = ( n4781 & n4795 ) | ( n4781 & ~n4796 ) | ( n4795 & ~n4796 ) ;
  assign n4798 = n4761 | n4797 ;
  assign n4799 = n2965 & ~n4758 ;
  assign n4800 = ~n4736 & n4799 ;
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  assign n4801 = n161 & n4115 ;
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n52( .i (n51), .o (n52) );
  buffer buf_n53( .i (n52), .o (n53) );
  assign n4802 = n53 & ~n4115 ;
  buffer buf_n4803( .i (n1491), .o (n4803) );
  assign n4804 = ( n4801 & n4802 ) | ( n4801 & n4803 ) | ( n4802 & n4803 ) ;
  buffer buf_n4805( .i (n4804), .o (n4805) );
  buffer buf_n4806( .i (n4805), .o (n4806) );
  buffer buf_n4807( .i (n4806), .o (n4807) );
  buffer buf_n4808( .i (n4807), .o (n4808) );
  buffer buf_n4809( .i (n4808), .o (n4809) );
  buffer buf_n4810( .i (n4809), .o (n4810) );
  buffer buf_n4811( .i (n4810), .o (n4811) );
  buffer buf_n4812( .i (n4811), .o (n4812) );
  assign n4813 = n2942 & ~n4810 ;
  buffer buf_n4814( .i (n4813), .o (n4814) );
  assign n4815 = n264 & n1532 ;
  buffer buf_n4816( .i (n4815), .o (n4816) );
  buffer buf_n4817( .i (n4816), .o (n4817) );
  buffer buf_n4818( .i (n4817), .o (n4818) );
  assign n4819 = n2674 & ~n4816 ;
  buffer buf_n4820( .i (n4819), .o (n4820) );
  assign n4821 = ( n4545 & ~n4818 ) | ( n4545 & n4820 ) | ( ~n4818 & n4820 ) ;
  buffer buf_n4822( .i (n4821), .o (n4822) );
  buffer buf_n4823( .i (n4822), .o (n4823) );
  assign n4824 = ( ~n4812 & n4814 ) | ( ~n4812 & n4823 ) | ( n4814 & n4823 ) ;
  buffer buf_n4825( .i (n4824), .o (n4825) );
  buffer buf_n4826( .i (n4825), .o (n4826) );
  buffer buf_n4827( .i (n4826), .o (n4827) );
  assign n4828 = n2761 | n4818 ;
  buffer buf_n4829( .i (n2760), .o (n4829) );
  assign n4830 = n4820 & ~n4829 ;
  assign n4831 = ( n4546 & ~n4828 ) | ( n4546 & n4830 ) | ( ~n4828 & n4830 ) ;
  buffer buf_n4832( .i (n4831), .o (n4832) );
  assign n4833 = ( ~n4812 & n4814 ) | ( ~n4812 & n4832 ) | ( n4814 & n4832 ) ;
  buffer buf_n4834( .i (n4833), .o (n4834) );
  buffer buf_n4835( .i (n4834), .o (n4835) );
  buffer buf_n4836( .i (n4835), .o (n4836) );
  assign n4837 = ( n4473 & n4827 ) | ( n4473 & n4836 ) | ( n4827 & n4836 ) ;
  assign n4838 = ~n4800 & n4837 ;
  buffer buf_n4839( .i (n4838), .o (n4839) );
  assign n4840 = n3240 & ~n4758 ;
  assign n4841 = ~n4736 & n4840 ;
  buffer buf_n4842( .i (n4841), .o (n4842) );
  buffer buf_n4474( .i (n4473), .o (n4474) );
  buffer buf_n566( .i (x78), .o (n566) );
  assign n4843 = n566 & n1314 ;
  buffer buf_n4844( .i (n4843), .o (n4844) );
  buffer buf_n4845( .i (n4844), .o (n4845) );
  buffer buf_n4846( .i (n4845), .o (n4846) );
  buffer buf_n564( .i (x77), .o (n564) );
  assign n4847 = n564 & ~n1314 ;
  buffer buf_n4848( .i (n4847), .o (n4848) );
  buffer buf_n4849( .i (n4848), .o (n4849) );
  buffer buf_n4850( .i (n4849), .o (n4850) );
  assign n4851 = ( n3245 & n4846 ) | ( n3245 & n4850 ) | ( n4846 & n4850 ) ;
  buffer buf_n4852( .i (n4851), .o (n4852) );
  buffer buf_n4853( .i (n4852), .o (n4853) );
  buffer buf_n4854( .i (n4853), .o (n4854) );
  buffer buf_n4855( .i (n4854), .o (n4855) );
  buffer buf_n4856( .i (n4855), .o (n4856) );
  buffer buf_n4857( .i (n4856), .o (n4857) );
  buffer buf_n4858( .i (n4857), .o (n4858) );
  buffer buf_n4859( .i (n4858), .o (n4859) );
  buffer buf_n4860( .i (n4859), .o (n4860) );
  buffer buf_n4861( .i (n4860), .o (n4861) );
  buffer buf_n4862( .i (n4861), .o (n4862) );
  assign n4863 = n3218 | n4860 ;
  buffer buf_n4864( .i (n4863), .o (n4864) );
  assign n4865 = ( ~n4823 & n4862 ) | ( ~n4823 & n4864 ) | ( n4862 & n4864 ) ;
  buffer buf_n4866( .i (n4865), .o (n4866) );
  buffer buf_n4867( .i (n4866), .o (n4867) );
  buffer buf_n4868( .i (n4867), .o (n4868) );
  buffer buf_n4869( .i (n4868), .o (n4869) );
  assign n4870 = ( ~n4832 & n4862 ) | ( ~n4832 & n4864 ) | ( n4862 & n4864 ) ;
  buffer buf_n4871( .i (n4870), .o (n4871) );
  buffer buf_n4872( .i (n4871), .o (n4872) );
  buffer buf_n4873( .i (n4872), .o (n4873) );
  buffer buf_n4874( .i (n4873), .o (n4874) );
  assign n4875 = ( ~n4474 & n4869 ) | ( ~n4474 & n4874 ) | ( n4869 & n4874 ) ;
  assign n4876 = n4842 | n4875 ;
  assign n4877 = n3302 & ~n4758 ;
  assign n4878 = ~n4736 & n4877 ;
  buffer buf_n4879( .i (n4878), .o (n4879) );
  assign n4880 = n566 & n1324 ;
  buffer buf_n4881( .i (n4880), .o (n4881) );
  buffer buf_n4882( .i (n4881), .o (n4882) );
  assign n4883 = n564 & ~n1324 ;
  buffer buf_n4884( .i (n4883), .o (n4884) );
  buffer buf_n4885( .i (n4884), .o (n4885) );
  assign n4886 = ( n3307 & n4882 ) | ( n3307 & n4885 ) | ( n4882 & n4885 ) ;
  buffer buf_n4887( .i (n4886), .o (n4887) );
  buffer buf_n4888( .i (n4887), .o (n4888) );
  buffer buf_n4889( .i (n4888), .o (n4889) );
  buffer buf_n4890( .i (n4889), .o (n4890) );
  buffer buf_n4891( .i (n4890), .o (n4891) );
  buffer buf_n4892( .i (n4891), .o (n4892) );
  buffer buf_n4893( .i (n4892), .o (n4893) );
  buffer buf_n4894( .i (n4893), .o (n4894) );
  buffer buf_n4895( .i (n4894), .o (n4895) );
  buffer buf_n4896( .i (n4895), .o (n4896) );
  buffer buf_n4897( .i (n4896), .o (n4897) );
  buffer buf_n4898( .i (n4897), .o (n4898) );
  assign n4899 = n3279 | n4896 ;
  buffer buf_n4900( .i (n4899), .o (n4900) );
  assign n4901 = ( ~n4823 & n4898 ) | ( ~n4823 & n4900 ) | ( n4898 & n4900 ) ;
  buffer buf_n4902( .i (n4901), .o (n4902) );
  buffer buf_n4903( .i (n4902), .o (n4903) );
  buffer buf_n4904( .i (n4903), .o (n4904) );
  buffer buf_n4905( .i (n4904), .o (n4905) );
  assign n4906 = ( ~n4832 & n4898 ) | ( ~n4832 & n4900 ) | ( n4898 & n4900 ) ;
  buffer buf_n4907( .i (n4906), .o (n4907) );
  buffer buf_n4908( .i (n4907), .o (n4908) );
  buffer buf_n4909( .i (n4908), .o (n4909) );
  buffer buf_n4910( .i (n4909), .o (n4910) );
  assign n4911 = ( ~n4474 & n4905 ) | ( ~n4474 & n4910 ) | ( n4905 & n4910 ) ;
  assign n4912 = n4879 | n4911 ;
  assign y0 = n509 ;
  assign y1 = n772 ;
  assign y2 = n1372 ;
  assign y3 = ~n1202 ;
  assign y4 = ~n915 ;
  assign y5 = ~n975 ;
  assign y6 = n1552 ;
  assign y7 = ~n1227 ;
  assign y8 = ~n1202 ;
  assign y9 = ~n1202 ;
  assign y10 = ~n884 ;
  assign y11 = ~n945 ;
  assign y12 = n1574 ;
  assign y13 = ~n683 ;
  assign y14 = ~n1252 ;
  assign y15 = ~n1303 ;
  assign y16 = ~n1278 ;
  assign y17 = n1597 ;
  assign y18 = n1620 ;
  assign y19 = ~n1643 ;
  assign y20 = ~n1667 ;
  assign y21 = n478 ;
  assign y22 = n509 ;
  assign y23 = n25 ;
  assign y24 = n1227 ;
  assign y25 = n797 ;
  assign y26 = ~n1227 ;
  assign y27 = ~n1709 ;
  assign y28 = ~n1690 ;
  assign y29 = n25 ;
  assign y30 = n25 ;
  assign y31 = n25 ;
  assign y32 = n4913 ;
  assign y33 = n797 ;
  assign y34 = ~n797 ;
  assign y35 = ~n1731 ;
  assign y36 = ~n1755 ;
  assign y37 = ~n1755 ;
  assign y38 = ~n1774 ;
  assign y39 = n1798 ;
  assign y40 = n1821 ;
  assign y41 = n1846 ;
  assign y42 = n1871 ;
  assign y43 = n1960 ;
  assign y44 = n2069 ;
  assign y45 = n2329 ;
  assign y46 = n2535 ;
  assign y47 = n2535 ;
  assign y48 = n2329 ;
  assign y49 = ~n2567 ;
  assign y50 = n2602 ;
  assign y51 = n2641 ;
  assign y52 = n2665 ;
  assign y53 = n2641 ;
  assign y54 = n2665 ;
  assign y55 = n2717 ;
  assign y56 = n2740 ;
  assign y57 = n2781 ;
  assign y58 = n2802 ;
  assign y59 = ~n2853 ;
  assign y60 = n2876 ;
  assign y61 = n2897 ;
  assign y62 = n2935 ;
  assign y63 = ~n2985 ;
  assign y64 = n3016 ;
  assign y65 = n3038 ;
  assign y66 = n3060 ;
  assign y67 = n3080 ;
  assign y68 = ~n3115 ;
  assign y69 = n3157 ;
  assign y70 = ~n3201 ;
  assign y71 = n3206 ;
  assign y72 = n3266 ;
  assign y73 = n3329 ;
  assign y74 = ~n3353 ;
  assign y75 = ~n3369 ;
  assign y76 = ~n3384 ;
  assign y77 = ~n3401 ;
  assign y78 = ~n3425 ;
  assign y79 = ~n3438 ;
  assign y80 = ~n3450 ;
  assign y81 = ~n3465 ;
  assign y82 = n3488 ;
  assign y83 = n3510 ;
  assign y84 = n3539 ;
  assign y85 = n3564 ;
  assign y86 = n3587 ;
  assign y87 = n3611 ;
  assign y88 = n3642 ;
  assign y89 = n3665 ;
  assign y90 = n3700 ;
  assign y91 = n3707 ;
  assign y92 = ~n3740 ;
  assign y93 = n3763 ;
  assign y94 = ~n3789 ;
  assign y95 = ~n3812 ;
  assign y96 = n3830 ;
  assign y97 = ~n3869 ;
  assign y98 = n3891 ;
  assign y99 = n3913 ;
  assign y100 = n3951 ;
  assign y101 = n3983 ;
  assign y102 = n4008 ;
  assign y103 = ~n4032 ;
  assign y104 = n4058 ;
  assign y105 = n4084 ;
  assign y106 = ~n4112 ;
  assign y107 = n4133 ;
  assign y108 = n4164 ;
  assign y109 = n4193 ;
  assign y110 = n4220 ;
  assign y111 = n4246 ;
  assign y112 = n4273 ;
  assign y113 = n4297 ;
  assign y114 = n4322 ;
  assign y115 = n4347 ;
  assign y116 = n4375 ;
  assign y117 = n4555 ;
  assign y118 = n4739 ;
  assign y119 = ~n4798 ;
  assign y120 = ~n4839 ;
  assign y121 = ~n4876 ;
  assign y122 = ~n4912 ;
endmodule
