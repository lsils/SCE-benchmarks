module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n46 , n47 , n48 , n49 , n50 , n51 , n53 , n54 , n55 , n56 , n57 , n58 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 ;
  buffer buf_n19( .i (x2), .o (n19) );
  buffer buf_n46( .i (x5), .o (n46) );
  assign n67 = n19 & n46 ;
  buffer buf_n68( .i (n67), .o (n68) );
  buffer buf_n69( .i (n68), .o (n69) );
  buffer buf_n70( .i (n69), .o (n70) );
  buffer buf_n71( .i (n70), .o (n71) );
  buffer buf_n20( .i (n19), .o (n20) );
  buffer buf_n53( .i (x6), .o (n53) );
  buffer buf_n54( .i (n53), .o (n54) );
  assign n75 = n20 & n54 ;
  buffer buf_n76( .i (n75), .o (n76) );
  buffer buf_n27( .i (x3), .o (n27) );
  buffer buf_n28( .i (n27), .o (n28) );
  buffer buf_n60( .i (x7), .o (n60) );
  buffer buf_n61( .i (n60), .o (n61) );
  assign n80 = n28 | n61 ;
  buffer buf_n81( .i (n80), .o (n81) );
  assign n83 = n76 | n81 ;
  buffer buf_n84( .i (n83), .o (n84) );
  assign n85 = n71 & n84 ;
  buffer buf_n11( .i (x1), .o (n11) );
  buffer buf_n12( .i (n11), .o (n12) );
  buffer buf_n13( .i (n12), .o (n13) );
  buffer buf_n14( .i (n13), .o (n14) );
  buffer buf_n15( .i (n14), .o (n15) );
  buffer buf_n16( .i (n15), .o (n16) );
  buffer buf_n47( .i (n46), .o (n47) );
  assign n86 = n28 & n47 ;
  buffer buf_n87( .i (n86), .o (n87) );
  buffer buf_n88( .i (n87), .o (n88) );
  buffer buf_n55( .i (n54), .o (n55) );
  buffer buf_n56( .i (n55), .o (n56) );
  buffer buf_n62( .i (n61), .o (n62) );
  buffer buf_n63( .i (n62), .o (n63) );
  assign n92 = n56 & n63 ;
  assign n93 = n88 & n92 ;
  assign n94 = n16 | n93 ;
  assign n95 = n85 | n94 ;
  buffer buf_n57( .i (n56), .o (n57) );
  buffer buf_n58( .i (n57), .o (n58) );
  assign n96 = n58 & n84 ;
  buffer buf_n48( .i (n47), .o (n48) );
  buffer buf_n49( .i (n48), .o (n49) );
  buffer buf_n50( .i (n49), .o (n50) );
  buffer buf_n51( .i (n50), .o (n51) );
  buffer buf_n21( .i (n20), .o (n21) );
  buffer buf_n22( .i (n21), .o (n22) );
  assign n97 = n22 & n63 ;
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n29( .i (n28), .o (n29) );
  buffer buf_n30( .i (n29), .o (n30) );
  buffer buf_n31( .i (n30), .o (n31) );
  assign n100 = n31 | n50 ;
  assign n101 = ( n51 & n98 ) | ( n51 & n100 ) | ( n98 & n100 ) ;
  assign n102 = n96 | n101 ;
  assign n103 = n95 & n102 ;
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n2( .i (x0), .o (n2) );
  buffer buf_n3( .i (n2), .o (n3) );
  buffer buf_n4( .i (n3), .o (n4) );
  buffer buf_n5( .i (n4), .o (n5) );
  buffer buf_n6( .i (n5), .o (n6) );
  buffer buf_n7( .i (n6), .o (n7) );
  buffer buf_n38( .i (x4), .o (n38) );
  buffer buf_n39( .i (n38), .o (n39) );
  buffer buf_n40( .i (n39), .o (n40) );
  buffer buf_n41( .i (n40), .o (n41) );
  buffer buf_n42( .i (n41), .o (n42) );
  buffer buf_n43( .i (n42), .o (n43) );
  assign n105 = n7 & n43 ;
  buffer buf_n106( .i (n105), .o (n106) );
  buffer buf_n107( .i (n106), .o (n107) );
  buffer buf_n108( .i (n107), .o (n108) );
  assign n109 = n104 & n108 ;
  buffer buf_n110( .i (n109), .o (n110) );
  buffer buf_n111( .i (n110), .o (n111) );
  buffer buf_n112( .i (n111), .o (n112) );
  assign n113 = ~n104 & n108 ;
  buffer buf_n114( .i (n113), .o (n114) );
  buffer buf_n115( .i (n114), .o (n115) );
  buffer buf_n64( .i (n63), .o (n64) );
  assign n116 = n40 & n55 ;
  buffer buf_n117( .i (n116), .o (n117) );
  assign n118 = n64 & n117 ;
  assign n119 = ~n3 & n20 ;
  buffer buf_n120( .i (n119), .o (n120) );
  assign n124 = n11 & n53 ;
  buffer buf_n125( .i (n124), .o (n125) );
  assign n130 = n40 | n125 ;
  assign n131 = n120 & n130 ;
  assign n132 = ~n11 & n19 ;
  buffer buf_n133( .i (n132), .o (n133) );
  assign n138 = n38 | n53 ;
  buffer buf_n139( .i (n138), .o (n139) );
  assign n143 = n133 & ~n139 ;
  assign n144 = ( ~n2 & n19 ) | ( ~n2 & n53 ) | ( n19 & n53 ) ;
  buffer buf_n145( .i (n144), .o (n145) );
  assign n147 = n55 & ~n145 ;
  assign n148 = ( n5 & n143 ) | ( n5 & n147 ) | ( n143 & n147 ) ;
  assign n149 = n131 | n148 ;
  assign n150 = ~n118 & n149 ;
  buffer buf_n151( .i (n150), .o (n151) );
  assign n153 = n14 & ~n30 ;
  buffer buf_n154( .i (n153), .o (n154) );
  assign n155 = n41 & ~n49 ;
  buffer buf_n156( .i (n155), .o (n156) );
  assign n157 = n154 & n156 ;
  buffer buf_n158( .i (n157), .o (n158) );
  assign n159 = n151 & n158 ;
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n77( .i (n76), .o (n77) );
  buffer buf_n78( .i (n77), .o (n78) );
  assign n162 = n28 & n61 ;
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  assign n174 = n78 | n165 ;
  buffer buf_n175( .i (n174), .o (n175) );
  assign n176 = n106 & n175 ;
  buffer buf_n23( .i (n22), .o (n23) );
  buffer buf_n24( .i (n23), .o (n24) );
  buffer buf_n25( .i (n24), .o (n25) );
  assign n177 = n2 & n46 ;
  buffer buf_n178( .i (n177), .o (n178) );
  buffer buf_n179( .i (n178), .o (n179) );
  buffer buf_n180( .i (n179), .o (n180) );
  assign n185 = ~n15 & n180 ;
  assign n186 = n12 & n39 ;
  buffer buf_n187( .i (n186), .o (n187) );
  buffer buf_n188( .i (n187), .o (n188) );
  assign n190 = n4 | n48 ;
  buffer buf_n191( .i (n190), .o (n191) );
  assign n193 = n188 & ~n191 ;
  assign n194 = n185 | n193 ;
  assign n195 = ~n25 & n194 ;
  buffer buf_n189( .i (n188), .o (n189) );
  assign n196 = n4 & n68 ;
  buffer buf_n197( .i (n196), .o (n197) );
  buffer buf_n198( .i (n197), .o (n198) );
  assign n199 = n49 | n56 ;
  assign n200 = n188 & ~n199 ;
  assign n201 = ( n189 & n198 ) | ( n189 & n200 ) | ( n198 & n200 ) ;
  assign n202 = n87 & n120 ;
  buffer buf_n203( .i (n202), .o (n203) );
  assign n204 = n13 & n62 ;
  buffer buf_n205( .i (n204), .o (n205) );
  assign n207 = ~n42 & n205 ;
  assign n208 = n203 & n207 ;
  assign n209 = n201 | n208 ;
  assign n210 = n195 | n209 ;
  assign n211 = ~n176 & n210 ;
  assign n212 = n160 | n211 ;
  buffer buf_n213( .i (n212), .o (n213) );
  buffer buf_n214( .i (n213), .o (n214) );
  buffer buf_n82( .i (n81), .o (n82) );
  assign n215 = ~n82 & n197 ;
  assign n216 = ~n55 & n178 ;
  buffer buf_n217( .i (n216), .o (n217) );
  assign n220 = n42 | n217 ;
  assign n221 = n215 | n220 ;
  buffer buf_n146( .i (n145), .o (n146) );
  assign n226 = n63 | n146 ;
  buffer buf_n227( .i (n226), .o (n227) );
  assign n228 = n22 | n30 ;
  assign n229 = n15 & n228 ;
  assign n230 = n227 & n229 ;
  assign n231 = n221 & ~n230 ;
  buffer buf_n232( .i (n231), .o (n232) );
  assign n233 = ~n5 & n41 ;
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  buffer buf_n236( .i (n235), .o (n236) );
  buffer buf_n44( .i (n43), .o (n44) );
  assign n222 = n22 | n56 ;
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  assign n237 = n44 & ~n224 ;
  buffer buf_n181( .i (n180), .o (n181) );
  buffer buf_n182( .i (n181), .o (n182) );
  assign n238 = n182 | n235 ;
  assign n239 = ( n236 & ~n237 ) | ( n236 & n238 ) | ( ~n237 & n238 ) ;
  assign n240 = ~n232 & n239 ;
  buffer buf_n241( .i (n240), .o (n241) );
  buffer buf_n242( .i (n241), .o (n242) );
  assign n243 = n114 | n242 ;
  assign n244 = ( n115 & ~n214 ) | ( n115 & n243 ) | ( ~n214 & n243 ) ;
  buffer buf_n8( .i (n7), .o (n8) );
  buffer buf_n79( .i (n78), .o (n79) );
  assign n245 = n8 & n79 ;
  assign n246 = n14 & n49 ;
  buffer buf_n247( .i (n246), .o (n247) );
  buffer buf_n248( .i (n247), .o (n248) );
  assign n253 = ~n223 & n247 ;
  buffer buf_n249( .i (n54), .o (n249) );
  buffer buf_n250( .i (n249), .o (n250) );
  assign n251 = ~n30 & n250 ;
  buffer buf_n252( .i (n251), .o (n252) );
  assign n254 = n234 & ~n252 ;
  assign n255 = ( n248 & n253 ) | ( n248 & ~n254 ) | ( n253 & ~n254 ) ;
  assign n256 = n245 | n255 ;
  assign n257 = n42 & n82 ;
  buffer buf_n258( .i (n257), .o (n258) );
  assign n259 = n7 & n223 ;
  assign n260 = ~n258 & n259 ;
  assign n261 = ~n41 & n250 ;
  buffer buf_n262( .i (n261), .o (n262) );
  assign n264 = n24 & n262 ;
  buffer buf_n265( .i (n48), .o (n265) );
  assign n266 = n14 | n265 ;
  buffer buf_n267( .i (n266), .o (n267) );
  assign n268 = ~n165 & n267 ;
  assign n269 = ~n264 & n268 ;
  assign n270 = ~n260 & n269 ;
  assign n271 = n256 & n270 ;
  buffer buf_n152( .i (n151), .o (n152) );
  buffer buf_n65( .i (n64), .o (n65) );
  buffer buf_n66( .i (n65), .o (n66) );
  buffer buf_n192( .i (n191), .o (n192) );
  assign n272 = ~n181 & n192 ;
  assign n273 = n66 & ~n272 ;
  buffer buf_n263( .i (n262), .o (n263) );
  assign n274 = n16 | n156 ;
  assign n275 = n263 | n274 ;
  buffer buf_n126( .i (n125), .o (n126) );
  buffer buf_n127( .i (n126), .o (n127) );
  buffer buf_n128( .i (n127), .o (n128) );
  assign n276 = n128 | n154 ;
  buffer buf_n277( .i (n276), .o (n277) );
  assign n278 = ( n273 & n275 ) | ( n273 & ~n277 ) | ( n275 & ~n277 ) ;
  assign n279 = n152 & n278 ;
  assign n280 = n271 | n279 ;
  buffer buf_n281( .i (n280), .o (n281) );
  buffer buf_n121( .i (n120), .o (n121) );
  buffer buf_n122( .i (n121), .o (n122) );
  buffer buf_n123( .i (n122), .o (n123) );
  assign n282 = n66 | n123 ;
  assign n283 = ~n24 & n43 ;
  assign n284 = n128 & n192 ;
  assign n285 = ~n283 & n284 ;
  assign n286 = n282 & n285 ;
  buffer buf_n287( .i (n286), .o (n287) );
  buffer buf_n288( .i (n287), .o (n288) );
  buffer buf_n289( .i (n288), .o (n289) );
  assign n290 = ~n281 & n289 ;
  buffer buf_n183( .i (n182), .o (n183) );
  buffer buf_n184( .i (n183), .o (n184) );
  buffer buf_n9( .i (n8), .o (n9) );
  buffer buf_n140( .i (n139), .o (n140) );
  assign n291 = n140 & n163 ;
  assign n292 = ( n23 & n117 ) | ( n23 & n291 ) | ( n117 & n291 ) ;
  buffer buf_n293( .i (n292), .o (n293) );
  buffer buf_n294( .i (n293), .o (n294) );
  assign n295 = n9 & n294 ;
  assign n296 = n184 | n295 ;
  assign n297 = ~n104 & n296 ;
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  assign n298 = ~n219 & n248 ;
  assign n299 = n43 & ~n203 ;
  buffer buf_n300( .i (n299), .o (n300) );
  assign n301 = ~n298 & n300 ;
  assign n302 = n232 & ~n301 ;
  buffer buf_n134( .i (n133), .o (n134) );
  buffer buf_n135( .i (n134), .o (n135) );
  buffer buf_n136( .i (n135), .o (n136) );
  assign n303 = n58 & n136 ;
  buffer buf_n304( .i (n303), .o (n304) );
  assign n305 = n7 & n16 ;
  assign n306 = ~n224 & n305 ;
  assign n307 = n304 | n306 ;
  buffer buf_n166( .i (n165), .o (n166) );
  assign n308 = n44 & n166 ;
  buffer buf_n309( .i (n308), .o (n309) );
  assign n310 = n307 & n309 ;
  assign n311 = n302 | n310 ;
  assign n312 = n297 | n311 ;
  assign n313 = n213 | n312 ;
  assign n314 = n290 | n313 ;
  buffer buf_n99( .i (n98), .o (n99) );
  assign n315 = n31 & n57 ;
  buffer buf_n316( .i (n315), .o (n316) );
  assign n317 = n99 & n316 ;
  buffer buf_n318( .i (n317), .o (n318) );
  buffer buf_n225( .i (n224), .o (n225) );
  assign n319 = n175 & n225 ;
  buffer buf_n167( .i (n166), .o (n167) );
  assign n320 = n167 | n225 ;
  assign n321 = ( n318 & ~n319 ) | ( n318 & n320 ) | ( ~n319 & n320 ) ;
  buffer buf_n322( .i (n321), .o (n322) );
  buffer buf_n323( .i (n322), .o (n323) );
  assign n324 = n114 & n323 ;
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n32( .i (n31), .o (n32) );
  assign n325 = n250 & ~n265 ;
  buffer buf_n326( .i (n325), .o (n326) );
  assign n327 = n32 & n326 ;
  buffer buf_n328( .i (n13), .o (n328) );
  buffer buf_n329( .i (n21), .o (n329) );
  assign n330 = n328 & ~n329 ;
  buffer buf_n331( .i (n330), .o (n331) );
  buffer buf_n332( .i (n331), .o (n332) );
  buffer buf_n141( .i (n140), .o (n141) );
  buffer buf_n142( .i (n141), .o (n142) );
  assign n333 = ~n142 & n331 ;
  assign n334 = ( n327 & n332 ) | ( n327 & n333 ) | ( n332 & n333 ) ;
  buffer buf_n137( .i (n136), .o (n137) );
  assign n335 = n32 & ~n262 ;
  assign n336 = n98 & n262 ;
  assign n337 = ( n137 & ~n335 ) | ( n137 & n336 ) | ( ~n335 & n336 ) ;
  assign n338 = n334 | n337 ;
  buffer buf_n89( .i (n88), .o (n89) );
  buffer buf_n90( .i (n89), .o (n90) );
  assign n339 = n44 | n90 ;
  assign n340 = ~n9 & n339 ;
  assign n341 = n338 & n340 ;
  buffer buf_n342( .i (n6), .o (n342) );
  buffer buf_n343( .i (n40), .o (n343) );
  buffer buf_n344( .i (n343), .o (n344) );
  buffer buf_n345( .i (n344), .o (n345) );
  assign n346 = n342 & ~n345 ;
  buffer buf_n347( .i (n346), .o (n347) );
  buffer buf_n348( .i (n347), .o (n348) );
  assign n349 = n247 | n252 ;
  assign n350 = n25 & n349 ;
  assign n351 = ~n65 & n326 ;
  buffer buf_n352( .i (n351), .o (n352) );
  assign n353 = n65 & n267 ;
  buffer buf_n354( .i (n353), .o (n354) );
  assign n355 = ( n350 & n352 ) | ( n350 & ~n354 ) | ( n352 & ~n354 ) ;
  assign n356 = n348 & n355 ;
  assign n357 = n341 | n356 ;
  assign n358 = n161 | n357 ;
  assign n359 = n281 | n358 ;
  assign n360 = n324 | n359 ;
  buffer buf_n72( .i (n71), .o (n72) );
  buffer buf_n73( .i (n72), .o (n73) );
  buffer buf_n74( .i (n73), .o (n74) );
  assign n375 = n65 & n342 ;
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n129( .i (n128), .o (n129) );
  assign n385 = ~n99 & n129 ;
  buffer buf_n386( .i (n385), .o (n386) );
  assign n387 = ( n74 & n377 ) | ( n74 & n386 ) | ( n377 & n386 ) ;
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n33( .i (n32), .o (n33) );
  buffer buf_n34( .i (n33), .o (n34) );
  buffer buf_n35( .i (n34), .o (n35) );
  buffer buf_n36( .i (n35), .o (n36) );
  buffer buf_n378( .i (n377), .o (n378) );
  assign n389 = ( n74 & ~n377 ) | ( n74 & n386 ) | ( ~n377 & n386 ) ;
  assign n390 = ( ~n36 & n378 ) | ( ~n36 & n389 ) | ( n378 & n389 ) ;
  assign n391 = ~n388 & n390 ;
  assign n361 = ~n58 & n71 ;
  assign n362 = n129 | n361 ;
  buffer buf_n363( .i (n362), .o (n363) );
  buffer buf_n364( .i (n363), .o (n364) );
  assign n367 = ~n51 & n78 ;
  assign n368 = ( n66 & n248 ) | ( n66 & n367 ) | ( n248 & n367 ) ;
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  assign n392 = n364 & ~n370 ;
  buffer buf_n393( .i (n392), .o (n393) );
  assign n379 = n33 & n44 ;
  assign n380 = ~n376 & n379 ;
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n394( .i (n363), .o (n394) );
  assign n395 = ( ~n370 & n381 ) | ( ~n370 & n394 ) | ( n381 & n394 ) ;
  buffer buf_n396( .i (n395), .o (n396) );
  assign n397 = ( n391 & ~n393 ) | ( n391 & n396 ) | ( ~n393 & n396 ) ;
  buffer buf_n365( .i (n364), .o (n365) );
  buffer buf_n366( .i (n365), .o (n366) );
  assign n371 = n167 & n347 ;
  buffer buf_n372( .i (n371), .o (n372) );
  assign n373 = ( ~n364 & n370 ) | ( ~n364 & n372 ) | ( n370 & n372 ) ;
  buffer buf_n374( .i (n373), .o (n374) );
  assign n382 = n36 & ~n381 ;
  assign n383 = ( n364 & n370 ) | ( n364 & n372 ) | ( n370 & n372 ) ;
  assign n384 = n382 & ~n383 ;
  assign n398 = ( n366 & n374 ) | ( n366 & n384 ) | ( n374 & n384 ) ;
  assign n399 = n397 | n398 ;
  buffer buf_n17( .i (n16), .o (n17) );
  buffer buf_n402( .i (n64), .o (n402) );
  assign n403 = n89 & n402 ;
  assign n400 = n76 & ~n163 ;
  buffer buf_n401( .i (n400), .o (n401) );
  assign n404 = ~n89 & n401 ;
  assign n405 = ( ~n17 & n403 ) | ( ~n17 & n404 ) | ( n403 & n404 ) ;
  buffer buf_n406( .i (n405), .o (n406) );
  buffer buf_n91( .i (n90), .o (n91) );
  assign n408 = ( ~n64 & n77 ) | ( ~n64 & n88 ) | ( n77 & n88 ) ;
  buffer buf_n409( .i (n408), .o (n409) );
  assign n410 = ~n79 & n409 ;
  buffer buf_n206( .i (n205), .o (n206) );
  assign n407 = n206 & ~n401 ;
  assign n411 = n407 | n409 ;
  assign n412 = ( ~n91 & n410 ) | ( ~n91 & n411 ) | ( n410 & n411 ) ;
  assign n413 = n406 | n412 ;
  buffer buf_n414( .i (n413), .o (n414) );
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  buffer buf_n417( .i (n416), .o (n417) );
  assign n418 = n99 | n316 ;
  buffer buf_n419( .i (n418), .o (n419) );
  assign n420 = ~n318 & n419 ;
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n168( .i (n167), .o (n168) );
  buffer buf_n169( .i (n168), .o (n169) );
  buffer buf_n170( .i (n169), .o (n170) );
  buffer buf_n171( .i (n170), .o (n171) );
  buffer buf_n172( .i (n171), .o (n172) );
  buffer buf_n173( .i (n172), .o (n173) );
  assign y0 = n112 ;
  assign y1 = n244 ;
  assign y2 = n314 ;
  assign y3 = n360 ;
  assign y4 = n399 ;
  assign y5 = n417 ;
  assign y6 = n424 ;
  assign y7 = n173 ;
endmodule
