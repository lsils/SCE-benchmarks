module buffer( i , o );
  input i ;
  output o ;
endmodule
module inverter( i , o );
  input i ;
  output o ;
endmodule
module top( G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G5 , G6 , G7 , G8 , G9 , G1324 , G1325 , G1326 , G1327 , G1328 , G1329 , G1330 , G1331 , G1332 , G1333 , G1334 , G1335 , G1336 , G1337 , G1338 , G1339 , G1340 , G1341 , G1342 , G1343 , G1344 , G1345 , G1346 , G1347 , G1348 , G1349 , G1350 , G1351 , G1352 , G1353 , G1354 , G1355 );
  input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G5 , G6 , G7 , G8 , G9 ;
  output G1324 , G1325 , G1326 , G1327 , G1328 , G1329 , G1330 , G1331 , G1332 , G1333 , G1334 , G1335 , G1336 , G1337 , G1338 , G1339 , G1340 , G1341 , G1342 , G1343 , G1344 , G1345 , G1346 , G1347 , G1348 , G1349 , G1350 , G1351 , G1352 , G1353 , G1354 , G1355 ;
  wire n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 ;
  assign n42 = G33 & G41 ;
  buffer buf_n43( .i (n42), .o (n43) );
  assign n44 = G17 | G19 ;
  assign n45 = G17 & G19 ;
  assign n46 = n44 & ~n45 ;
  buffer buf_n47( .i (n46), .o (n47) );
  assign n48 = ~G18 & G20 ;
  assign n49 = G18 & ~G20 ;
  assign n50 = n48 | n49 ;
  buffer buf_n51( .i (n50), .o (n51) );
  assign n52 = ~n47 & n51 ;
  assign n53 = n47 & ~n51 ;
  assign n54 = n52 | n53 ;
  buffer buf_n55( .i (n54), .o (n55) );
  assign n57 = ~n43 & n55 ;
  assign n58 = n43 & ~n55 ;
  assign n59 = n57 | n58 ;
  buffer buf_n60( .i (n59), .o (n60) );
  assign n61 = G22 | G23 ;
  assign n62 = G22 & G23 ;
  assign n63 = n61 & ~n62 ;
  buffer buf_n64( .i (n63), .o (n64) );
  assign n65 = G21 & ~G24 ;
  assign n66 = ~G21 & G24 ;
  assign n67 = n65 | n66 ;
  buffer buf_n68( .i (n67), .o (n68) );
  assign n69 = ~n64 & n68 ;
  assign n70 = n64 & ~n68 ;
  assign n71 = n69 | n70 ;
  buffer buf_n72( .i (n71), .o (n72) );
  assign n74 = G13 | G5 ;
  assign n75 = G13 & G5 ;
  assign n76 = n74 & ~n75 ;
  buffer buf_n77( .i (n76), .o (n77) );
  assign n78 = G1 & ~G9 ;
  assign n79 = ~G1 & G9 ;
  assign n80 = n78 | n79 ;
  buffer buf_n81( .i (n80), .o (n81) );
  assign n82 = n77 | n81 ;
  assign n83 = n77 & n81 ;
  assign n84 = n82 & ~n83 ;
  buffer buf_n85( .i (n84), .o (n85) );
  assign n86 = n72 & n85 ;
  assign n87 = n72 | n85 ;
  assign n88 = ~n86 & n87 ;
  buffer buf_n89( .i (n88), .o (n89) );
  assign n90 = ~n60 & n89 ;
  assign n91 = n60 & ~n89 ;
  assign n92 = n90 | n91 ;
  buffer buf_n93( .i (n92), .o (n93) );
  buffer buf_n94( .i (n93), .o (n94) );
  buffer buf_n95( .i (n94), .o (n95) );
  buffer buf_n96( .i (n95), .o (n96) );
  buffer buf_n97( .i (n96), .o (n97) );
  buffer buf_n98( .i (n97), .o (n98) );
  buffer buf_n99( .i (n98), .o (n99) );
  buffer buf_n100( .i (n99), .o (n100) );
  buffer buf_n101( .i (n100), .o (n101) );
  buffer buf_n102( .i (n101), .o (n102) );
  buffer buf_n103( .i (n102), .o (n103) );
  buffer buf_n104( .i (n103), .o (n104) );
  buffer buf_n105( .i (n104), .o (n105) );
  assign n106 = G3 | G4 ;
  assign n107 = G3 & G4 ;
  assign n108 = n106 & ~n107 ;
  buffer buf_n109( .i (n108), .o (n109) );
  assign n110 = G1 & ~G2 ;
  assign n111 = ~G1 & G2 ;
  assign n112 = n110 | n111 ;
  buffer buf_n113( .i (n112), .o (n113) );
  assign n114 = ~n109 & n113 ;
  assign n115 = n109 & ~n113 ;
  assign n116 = n114 | n115 ;
  buffer buf_n117( .i (n116), .o (n117) );
  assign n118 = G39 & G41 ;
  buffer buf_n119( .i (n118), .o (n119) );
  assign n120 = n117 & ~n119 ;
  assign n121 = ~n117 & n119 ;
  assign n122 = n120 | n121 ;
  buffer buf_n123( .i (n122), .o (n123) );
  assign n124 = G10 | G12 ;
  assign n125 = G10 & G12 ;
  assign n126 = n124 & ~n125 ;
  buffer buf_n127( .i (n126), .o (n127) );
  assign n128 = ~G11 & G9 ;
  assign n129 = G11 & ~G9 ;
  assign n130 = n128 | n129 ;
  buffer buf_n131( .i (n130), .o (n131) );
  assign n132 = ~n127 & n131 ;
  assign n133 = n127 & ~n131 ;
  assign n134 = n132 | n133 ;
  buffer buf_n135( .i (n134), .o (n135) );
  assign n136 = G19 | G23 ;
  assign n137 = G19 & G23 ;
  assign n138 = n136 & ~n137 ;
  buffer buf_n139( .i (n138), .o (n139) );
  assign n140 = G27 & ~G31 ;
  assign n141 = ~G27 & G31 ;
  assign n142 = n140 | n141 ;
  buffer buf_n143( .i (n142), .o (n143) );
  assign n144 = n139 | n143 ;
  assign n145 = n139 & n143 ;
  assign n146 = n144 & ~n145 ;
  buffer buf_n147( .i (n146), .o (n147) );
  assign n148 = n135 & n147 ;
  assign n149 = n135 | n147 ;
  assign n150 = ~n148 & n149 ;
  buffer buf_n151( .i (n150), .o (n151) );
  assign n152 = ~n123 & n151 ;
  assign n153 = n123 & ~n151 ;
  assign n154 = n152 | n153 ;
  buffer buf_n155( .i (n154), .o (n155) );
  buffer buf_n156( .i (n155), .o (n156) );
  assign n167 = G7 | G8 ;
  assign n168 = G7 & G8 ;
  assign n169 = n167 & ~n168 ;
  buffer buf_n170( .i (n169), .o (n170) );
  assign n171 = ~G5 & G6 ;
  assign n172 = G5 & ~G6 ;
  assign n173 = n171 | n172 ;
  buffer buf_n174( .i (n173), .o (n174) );
  assign n175 = ~n170 & n174 ;
  assign n176 = n170 & ~n174 ;
  assign n177 = n175 | n176 ;
  buffer buf_n178( .i (n177), .o (n178) );
  assign n179 = G40 & G41 ;
  buffer buf_n180( .i (n179), .o (n180) );
  assign n181 = n178 & ~n180 ;
  assign n182 = ~n178 & n180 ;
  assign n183 = n181 | n182 ;
  buffer buf_n184( .i (n183), .o (n184) );
  assign n185 = G14 | G16 ;
  assign n186 = G14 & G16 ;
  assign n187 = n185 & ~n186 ;
  buffer buf_n188( .i (n187), .o (n188) );
  assign n189 = G13 & ~G15 ;
  assign n190 = ~G13 & G15 ;
  assign n191 = n189 | n190 ;
  buffer buf_n192( .i (n191), .o (n192) );
  assign n193 = ~n188 & n192 ;
  assign n194 = n188 & ~n192 ;
  assign n195 = n193 | n194 ;
  buffer buf_n196( .i (n195), .o (n196) );
  assign n197 = G20 | G24 ;
  assign n198 = G20 & G24 ;
  assign n199 = n197 & ~n198 ;
  buffer buf_n200( .i (n199), .o (n200) );
  assign n201 = ~G28 & G32 ;
  assign n202 = G28 & ~G32 ;
  assign n203 = n201 | n202 ;
  buffer buf_n204( .i (n203), .o (n204) );
  assign n205 = n200 | n204 ;
  assign n206 = n200 & n204 ;
  assign n207 = n205 & ~n206 ;
  buffer buf_n208( .i (n207), .o (n208) );
  assign n209 = n196 & n208 ;
  assign n210 = n196 | n208 ;
  assign n211 = ~n209 & n210 ;
  buffer buf_n212( .i (n211), .o (n212) );
  assign n213 = ~n184 & n212 ;
  assign n214 = n184 & ~n212 ;
  assign n215 = n213 | n214 ;
  buffer buf_n216( .i (n215), .o (n216) );
  buffer buf_n217( .i (n216), .o (n217) );
  assign n228 = n156 & ~n217 ;
  buffer buf_n229( .i (n228), .o (n229) );
  buffer buf_n230( .i (n229), .o (n230) );
  buffer buf_n231( .i (n230), .o (n231) );
  buffer buf_n232( .i (n231), .o (n232) );
  buffer buf_n233( .i (n232), .o (n233) );
  buffer buf_n234( .i (n233), .o (n234) );
  buffer buf_n235( .i (n234), .o (n235) );
  assign n236 = G37 & G41 ;
  buffer buf_n237( .i (n236), .o (n237) );
  assign n238 = n117 & ~n237 ;
  assign n239 = ~n117 & n237 ;
  assign n240 = n238 | n239 ;
  buffer buf_n241( .i (n240), .o (n241) );
  assign n242 = G21 & ~G25 ;
  assign n243 = ~G21 & G25 ;
  assign n244 = n242 | n243 ;
  buffer buf_n245( .i (n244), .o (n245) );
  assign n246 = G17 | G29 ;
  assign n247 = G17 & G29 ;
  assign n248 = n246 & ~n247 ;
  buffer buf_n249( .i (n248), .o (n249) );
  assign n250 = n245 | n249 ;
  assign n251 = n245 & n249 ;
  assign n252 = n250 & ~n251 ;
  buffer buf_n253( .i (n252), .o (n253) );
  assign n254 = n178 & n253 ;
  assign n255 = n178 | n253 ;
  assign n256 = ~n254 & n255 ;
  buffer buf_n257( .i (n256), .o (n257) );
  assign n258 = ~n241 & n257 ;
  assign n259 = n241 & ~n257 ;
  assign n260 = n258 | n259 ;
  buffer buf_n261( .i (n260), .o (n261) );
  buffer buf_n262( .i (n261), .o (n262) );
  assign n273 = G38 & G41 ;
  buffer buf_n274( .i (n273), .o (n274) );
  assign n275 = n135 & ~n274 ;
  assign n276 = ~n135 & n274 ;
  assign n277 = n275 | n276 ;
  buffer buf_n278( .i (n277), .o (n278) );
  assign n279 = ~G18 & G26 ;
  assign n280 = G18 & ~G26 ;
  assign n281 = n279 | n280 ;
  buffer buf_n282( .i (n281), .o (n282) );
  assign n283 = G22 | G30 ;
  assign n284 = G22 & G30 ;
  assign n285 = n283 & ~n284 ;
  buffer buf_n286( .i (n285), .o (n286) );
  assign n287 = n282 | n286 ;
  assign n288 = n282 & n286 ;
  assign n289 = n287 & ~n288 ;
  buffer buf_n290( .i (n289), .o (n290) );
  assign n291 = n196 & n290 ;
  assign n292 = n196 | n290 ;
  assign n293 = ~n291 & n292 ;
  buffer buf_n294( .i (n293), .o (n294) );
  assign n295 = ~n278 & n294 ;
  assign n296 = n278 & ~n294 ;
  assign n297 = n295 | n296 ;
  buffer buf_n298( .i (n297), .o (n298) );
  buffer buf_n299( .i (n298), .o (n299) );
  assign n310 = n262 & ~n299 ;
  buffer buf_n311( .i (n310), .o (n311) );
  buffer buf_n312( .i (n311), .o (n312) );
  buffer buf_n313( .i (n312), .o (n313) );
  buffer buf_n314( .i (n313), .o (n314) );
  buffer buf_n315( .i (n314), .o (n315) );
  assign n316 = G34 & G41 ;
  buffer buf_n317( .i (n316), .o (n317) );
  assign n318 = G29 | G30 ;
  assign n319 = G29 & G30 ;
  assign n320 = n318 & ~n319 ;
  buffer buf_n321( .i (n320), .o (n321) );
  assign n322 = ~G31 & G32 ;
  assign n323 = G31 & ~G32 ;
  assign n324 = n322 | n323 ;
  buffer buf_n325( .i (n324), .o (n325) );
  assign n326 = ~n321 & n325 ;
  assign n327 = n321 & ~n325 ;
  assign n328 = n326 | n327 ;
  buffer buf_n329( .i (n328), .o (n329) );
  assign n331 = ~n317 & n329 ;
  assign n332 = n317 & ~n329 ;
  assign n333 = n331 | n332 ;
  buffer buf_n334( .i (n333), .o (n334) );
  assign n335 = G25 | G28 ;
  assign n336 = G25 & G28 ;
  assign n337 = n335 & ~n336 ;
  buffer buf_n338( .i (n337), .o (n338) );
  assign n339 = G26 & ~G27 ;
  assign n340 = ~G26 & G27 ;
  assign n341 = n339 | n340 ;
  buffer buf_n342( .i (n341), .o (n342) );
  assign n343 = ~n338 & n342 ;
  assign n344 = n338 & ~n342 ;
  assign n345 = n343 | n344 ;
  buffer buf_n346( .i (n345), .o (n346) );
  assign n348 = G14 | G2 ;
  assign n349 = G14 & G2 ;
  assign n350 = n348 & ~n349 ;
  buffer buf_n351( .i (n350), .o (n351) );
  assign n352 = G10 & ~G6 ;
  assign n353 = ~G10 & G6 ;
  assign n354 = n352 | n353 ;
  buffer buf_n355( .i (n354), .o (n355) );
  assign n356 = n351 | n355 ;
  assign n357 = n351 & n355 ;
  assign n358 = n356 & ~n357 ;
  buffer buf_n359( .i (n358), .o (n359) );
  assign n360 = n346 & n359 ;
  assign n361 = n346 | n359 ;
  assign n362 = ~n360 & n361 ;
  buffer buf_n363( .i (n362), .o (n363) );
  assign n364 = ~n334 & n363 ;
  assign n365 = n334 & ~n363 ;
  assign n366 = n364 | n365 ;
  buffer buf_n367( .i (n366), .o (n367) );
  assign n380 = ~n93 & n367 ;
  buffer buf_n381( .i (n380), .o (n381) );
  buffer buf_n56( .i (n55), .o (n56) );
  assign n390 = G35 & G41 ;
  buffer buf_n391( .i (n390), .o (n391) );
  assign n392 = n56 & ~n391 ;
  assign n393 = ~n56 & n391 ;
  assign n394 = n392 | n393 ;
  buffer buf_n395( .i (n394), .o (n395) );
  buffer buf_n347( .i (n346), .o (n347) );
  assign n396 = G11 & ~G15 ;
  assign n397 = ~G11 & G15 ;
  assign n398 = n396 | n397 ;
  buffer buf_n399( .i (n398), .o (n399) );
  assign n400 = G3 | G7 ;
  assign n401 = G3 & G7 ;
  assign n402 = n400 & ~n401 ;
  buffer buf_n403( .i (n402), .o (n403) );
  assign n404 = n399 | n403 ;
  assign n405 = n399 & n403 ;
  assign n406 = n404 & ~n405 ;
  buffer buf_n407( .i (n406), .o (n407) );
  assign n408 = n347 & n407 ;
  assign n409 = n347 | n407 ;
  assign n410 = ~n408 & n409 ;
  buffer buf_n411( .i (n410), .o (n411) );
  assign n412 = ~n395 & n411 ;
  assign n413 = n395 & ~n411 ;
  assign n414 = n412 | n413 ;
  buffer buf_n415( .i (n414), .o (n415) );
  buffer buf_n416( .i (n415), .o (n416) );
  assign n427 = n381 & ~n416 ;
  buffer buf_n428( .i (n427), .o (n428) );
  assign n434 = n93 & ~n367 ;
  buffer buf_n435( .i (n434), .o (n435) );
  assign n444 = ~n416 & n435 ;
  buffer buf_n445( .i (n444), .o (n445) );
  assign n451 = n428 | n445 ;
  buffer buf_n73( .i (n72), .o (n73) );
  assign n452 = G36 & G41 ;
  buffer buf_n453( .i (n452), .o (n453) );
  assign n454 = n73 & ~n453 ;
  assign n455 = ~n73 & n453 ;
  assign n456 = n454 | n455 ;
  buffer buf_n457( .i (n456), .o (n457) );
  buffer buf_n330( .i (n329), .o (n330) );
  assign n458 = G12 & ~G4 ;
  assign n459 = ~G12 & G4 ;
  assign n460 = n458 | n459 ;
  buffer buf_n461( .i (n460), .o (n461) );
  assign n462 = G16 | G8 ;
  assign n463 = G16 & G8 ;
  assign n464 = n462 & ~n463 ;
  buffer buf_n465( .i (n464), .o (n465) );
  assign n466 = n461 | n465 ;
  assign n467 = n461 & n465 ;
  assign n468 = n466 & ~n467 ;
  buffer buf_n469( .i (n468), .o (n469) );
  assign n470 = n330 & n469 ;
  assign n471 = n330 | n469 ;
  assign n472 = ~n470 & n471 ;
  buffer buf_n473( .i (n472), .o (n473) );
  assign n474 = ~n457 & n473 ;
  assign n475 = n457 & ~n473 ;
  assign n476 = n474 | n475 ;
  buffer buf_n477( .i (n476), .o (n477) );
  buffer buf_n478( .i (n477), .o (n478) );
  buffer buf_n479( .i (n478), .o (n479) );
  buffer buf_n480( .i (n479), .o (n480) );
  buffer buf_n481( .i (n480), .o (n481) );
  assign n489 = n451 & ~n481 ;
  assign n490 = n416 & ~n478 ;
  buffer buf_n491( .i (n490), .o (n491) );
  buffer buf_n417( .i (n416), .o (n417) );
  assign n496 = ~n417 & n479 ;
  assign n497 = n491 | n496 ;
  buffer buf_n368( .i (n367), .o (n368) );
  buffer buf_n369( .i (n368), .o (n369) );
  buffer buf_n370( .i (n369), .o (n370) );
  buffer buf_n371( .i (n370), .o (n371) );
  assign n498 = n97 | n371 ;
  assign n499 = n497 & ~n498 ;
  assign n500 = n489 | n499 ;
  buffer buf_n501( .i (n500), .o (n501) );
  assign n504 = n315 & n501 ;
  buffer buf_n505( .i (n504), .o (n505) );
  assign n506 = n235 & n505 ;
  buffer buf_n507( .i (n506), .o (n507) );
  assign n508 = n105 & n507 ;
  buffer buf_n509( .i (n508), .o (n509) );
  assign n510 = G1 & ~n509 ;
  assign n511 = ~G1 & n509 ;
  assign n512 = ~n510 & ~n511 ;
  buffer buf_n372( .i (n371), .o (n372) );
  buffer buf_n373( .i (n372), .o (n373) );
  buffer buf_n374( .i (n373), .o (n374) );
  buffer buf_n375( .i (n374), .o (n375) );
  buffer buf_n376( .i (n375), .o (n376) );
  buffer buf_n377( .i (n376), .o (n377) );
  buffer buf_n378( .i (n377), .o (n378) );
  buffer buf_n379( .i (n378), .o (n379) );
  assign n513 = n379 & n507 ;
  buffer buf_n514( .i (n513), .o (n514) );
  assign n515 = G2 & ~n514 ;
  assign n516 = ~G2 & n514 ;
  assign n517 = ~n515 & ~n516 ;
  buffer buf_n418( .i (n417), .o (n418) );
  buffer buf_n419( .i (n418), .o (n419) );
  buffer buf_n420( .i (n419), .o (n420) );
  buffer buf_n421( .i (n420), .o (n421) );
  buffer buf_n422( .i (n421), .o (n422) );
  buffer buf_n423( .i (n422), .o (n423) );
  buffer buf_n424( .i (n423), .o (n424) );
  buffer buf_n425( .i (n424), .o (n425) );
  buffer buf_n426( .i (n425), .o (n426) );
  assign n518 = n426 & n507 ;
  buffer buf_n519( .i (n518), .o (n519) );
  assign n520 = G3 & ~n519 ;
  assign n521 = ~G3 & n519 ;
  assign n522 = ~n520 & ~n521 ;
  buffer buf_n482( .i (n481), .o (n482) );
  buffer buf_n483( .i (n482), .o (n483) );
  buffer buf_n484( .i (n483), .o (n484) );
  buffer buf_n485( .i (n484), .o (n485) );
  buffer buf_n486( .i (n485), .o (n486) );
  buffer buf_n487( .i (n486), .o (n487) );
  buffer buf_n488( .i (n487), .o (n488) );
  assign n523 = n488 & n507 ;
  buffer buf_n524( .i (n523), .o (n524) );
  assign n525 = G4 & ~n524 ;
  assign n526 = ~G4 & n524 ;
  assign n527 = ~n525 & ~n526 ;
  assign n528 = ~n156 & n217 ;
  buffer buf_n529( .i (n528), .o (n529) );
  buffer buf_n530( .i (n529), .o (n530) );
  buffer buf_n531( .i (n530), .o (n531) );
  buffer buf_n532( .i (n531), .o (n532) );
  buffer buf_n533( .i (n532), .o (n533) );
  buffer buf_n534( .i (n533), .o (n534) );
  buffer buf_n535( .i (n534), .o (n535) );
  assign n536 = n505 & n535 ;
  buffer buf_n537( .i (n536), .o (n537) );
  assign n538 = n105 & n537 ;
  buffer buf_n539( .i (n538), .o (n539) );
  assign n540 = G5 & ~n539 ;
  assign n541 = ~G5 & n539 ;
  assign n542 = ~n540 & ~n541 ;
  assign n543 = n379 & n537 ;
  buffer buf_n544( .i (n543), .o (n544) );
  assign n545 = G6 & ~n544 ;
  assign n546 = ~G6 & n544 ;
  assign n547 = ~n545 & ~n546 ;
  assign n548 = n426 & n537 ;
  buffer buf_n549( .i (n548), .o (n549) );
  assign n550 = G7 & ~n549 ;
  assign n551 = ~G7 & n549 ;
  assign n552 = ~n550 & ~n551 ;
  assign n553 = n488 & n537 ;
  buffer buf_n554( .i (n553), .o (n554) );
  assign n555 = G8 & ~n554 ;
  assign n556 = ~G8 & n554 ;
  assign n557 = ~n555 & ~n556 ;
  assign n558 = ~n262 & n299 ;
  buffer buf_n559( .i (n558), .o (n559) );
  buffer buf_n560( .i (n559), .o (n560) );
  buffer buf_n561( .i (n560), .o (n561) );
  buffer buf_n562( .i (n561), .o (n562) );
  buffer buf_n563( .i (n562), .o (n563) );
  buffer buf_n564( .i (n563), .o (n564) );
  buffer buf_n565( .i (n564), .o (n565) );
  buffer buf_n502( .i (n501), .o (n502) );
  assign n566 = n234 & n502 ;
  assign n567 = n565 & n566 ;
  buffer buf_n568( .i (n567), .o (n568) );
  assign n569 = n105 & n568 ;
  buffer buf_n570( .i (n569), .o (n570) );
  assign n571 = G9 & ~n570 ;
  assign n572 = ~G9 & n570 ;
  assign n573 = ~n571 & ~n572 ;
  assign n574 = n379 & n568 ;
  buffer buf_n575( .i (n574), .o (n575) );
  assign n576 = G10 & ~n575 ;
  assign n577 = ~G10 & n575 ;
  assign n578 = ~n576 & ~n577 ;
  assign n579 = n426 & n568 ;
  buffer buf_n580( .i (n579), .o (n580) );
  assign n581 = G11 & ~n580 ;
  assign n582 = ~G11 & n580 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = n488 & n568 ;
  buffer buf_n585( .i (n584), .o (n585) );
  assign n586 = G12 & ~n585 ;
  assign n587 = ~G12 & n585 ;
  assign n588 = ~n586 & ~n587 ;
  buffer buf_n503( .i (n502), .o (n503) );
  assign n589 = n534 & n564 ;
  assign n590 = n503 & n589 ;
  buffer buf_n591( .i (n590), .o (n591) );
  assign n592 = n105 & n591 ;
  buffer buf_n593( .i (n592), .o (n593) );
  assign n594 = G13 | n593 ;
  assign n595 = G13 & n593 ;
  assign n596 = ~n594 | n595 ;
  assign n597 = n379 & n591 ;
  buffer buf_n598( .i (n597), .o (n598) );
  assign n599 = G14 | n598 ;
  assign n600 = G14 & n598 ;
  assign n601 = ~n599 | n600 ;
  assign n602 = n426 & n591 ;
  buffer buf_n603( .i (n602), .o (n603) );
  assign n604 = G15 & ~n603 ;
  assign n605 = ~G15 & n603 ;
  assign n606 = ~n604 & ~n605 ;
  assign n607 = n488 & n591 ;
  buffer buf_n608( .i (n607), .o (n608) );
  assign n609 = G16 | n608 ;
  assign n610 = G16 & n608 ;
  assign n611 = ~n609 | n610 ;
  buffer buf_n263( .i (n262), .o (n263) );
  buffer buf_n264( .i (n263), .o (n264) );
  buffer buf_n265( .i (n264), .o (n265) );
  buffer buf_n266( .i (n265), .o (n266) );
  buffer buf_n267( .i (n266), .o (n267) );
  buffer buf_n268( .i (n267), .o (n268) );
  buffer buf_n269( .i (n268), .o (n269) );
  buffer buf_n270( .i (n269), .o (n270) );
  buffer buf_n271( .i (n270), .o (n271) );
  buffer buf_n272( .i (n271), .o (n272) );
  buffer buf_n436( .i (n435), .o (n436) );
  buffer buf_n437( .i (n436), .o (n437) );
  buffer buf_n438( .i (n437), .o (n438) );
  buffer buf_n439( .i (n438), .o (n439) );
  buffer buf_n440( .i (n439), .o (n440) );
  buffer buf_n441( .i (n440), .o (n441) );
  buffer buf_n442( .i (n441), .o (n442) );
  buffer buf_n443( .i (n442), .o (n443) );
  buffer buf_n492( .i (n491), .o (n492) );
  buffer buf_n493( .i (n492), .o (n493) );
  buffer buf_n494( .i (n493), .o (n494) );
  buffer buf_n495( .i (n494), .o (n495) );
  assign n612 = n311 | n559 ;
  buffer buf_n157( .i (n156), .o (n157) );
  buffer buf_n158( .i (n157), .o (n158) );
  buffer buf_n218( .i (n217), .o (n218) );
  buffer buf_n219( .i (n218), .o (n219) );
  assign n613 = n158 | n219 ;
  assign n614 = n612 & ~n613 ;
  assign n615 = n229 | n529 ;
  buffer buf_n300( .i (n299), .o (n300) );
  buffer buf_n301( .i (n300), .o (n301) );
  assign n616 = n264 | n301 ;
  assign n617 = n615 & ~n616 ;
  assign n618 = n614 | n617 ;
  buffer buf_n619( .i (n618), .o (n619) );
  assign n622 = n495 & n619 ;
  buffer buf_n623( .i (n622), .o (n623) );
  assign n624 = n443 & n623 ;
  buffer buf_n625( .i (n624), .o (n625) );
  assign n626 = n272 & n625 ;
  buffer buf_n627( .i (n626), .o (n627) );
  assign n628 = G17 & ~n627 ;
  assign n629 = ~G17 & n627 ;
  assign n630 = ~n628 & ~n629 ;
  buffer buf_n302( .i (n301), .o (n302) );
  buffer buf_n303( .i (n302), .o (n303) );
  buffer buf_n304( .i (n303), .o (n304) );
  buffer buf_n305( .i (n304), .o (n305) );
  buffer buf_n306( .i (n305), .o (n306) );
  buffer buf_n307( .i (n306), .o (n307) );
  buffer buf_n308( .i (n307), .o (n308) );
  buffer buf_n309( .i (n308), .o (n309) );
  assign n631 = n309 & n625 ;
  buffer buf_n632( .i (n631), .o (n632) );
  assign n633 = G18 & ~n632 ;
  assign n634 = ~G18 & n632 ;
  assign n635 = ~n633 & ~n634 ;
  buffer buf_n159( .i (n158), .o (n159) );
  buffer buf_n160( .i (n159), .o (n160) );
  buffer buf_n161( .i (n160), .o (n161) );
  buffer buf_n162( .i (n161), .o (n162) );
  buffer buf_n163( .i (n162), .o (n163) );
  buffer buf_n164( .i (n163), .o (n164) );
  buffer buf_n165( .i (n164), .o (n165) );
  buffer buf_n166( .i (n165), .o (n166) );
  assign n636 = n166 & n625 ;
  buffer buf_n637( .i (n636), .o (n637) );
  assign n638 = G19 & ~n637 ;
  assign n639 = ~G19 & n637 ;
  assign n640 = ~n638 & ~n639 ;
  buffer buf_n220( .i (n219), .o (n220) );
  buffer buf_n221( .i (n220), .o (n221) );
  buffer buf_n222( .i (n221), .o (n222) );
  buffer buf_n223( .i (n222), .o (n223) );
  buffer buf_n224( .i (n223), .o (n224) );
  buffer buf_n225( .i (n224), .o (n225) );
  buffer buf_n226( .i (n225), .o (n226) );
  buffer buf_n227( .i (n226), .o (n227) );
  assign n641 = n227 & n625 ;
  buffer buf_n642( .i (n641), .o (n642) );
  assign n643 = G20 & ~n642 ;
  assign n644 = ~G20 & n642 ;
  assign n645 = ~n643 & ~n644 ;
  buffer buf_n620( .i (n619), .o (n620) );
  buffer buf_n621( .i (n620), .o (n621) );
  buffer buf_n446( .i (n445), .o (n446) );
  buffer buf_n447( .i (n446), .o (n447) );
  buffer buf_n448( .i (n447), .o (n448) );
  buffer buf_n449( .i (n448), .o (n449) );
  buffer buf_n450( .i (n449), .o (n450) );
  assign n646 = n450 & n485 ;
  assign n647 = n621 & n646 ;
  buffer buf_n648( .i (n647), .o (n648) );
  assign n649 = n272 & n648 ;
  buffer buf_n650( .i (n649), .o (n650) );
  assign n651 = G21 & ~n650 ;
  assign n652 = ~G21 & n650 ;
  assign n653 = ~n651 & ~n652 ;
  assign n654 = n309 & n648 ;
  buffer buf_n655( .i (n654), .o (n655) );
  assign n656 = G22 & ~n655 ;
  assign n657 = ~G22 & n655 ;
  assign n658 = ~n656 & ~n657 ;
  assign n659 = n166 & n648 ;
  buffer buf_n660( .i (n659), .o (n660) );
  assign n661 = G23 & ~n660 ;
  assign n662 = ~G23 & n660 ;
  assign n663 = ~n661 & ~n662 ;
  assign n664 = n227 & n648 ;
  buffer buf_n665( .i (n664), .o (n665) );
  assign n666 = G24 & ~n665 ;
  assign n667 = ~G24 & n665 ;
  assign n668 = ~n666 & ~n667 ;
  buffer buf_n382( .i (n381), .o (n382) );
  buffer buf_n383( .i (n382), .o (n383) );
  buffer buf_n384( .i (n383), .o (n384) );
  buffer buf_n385( .i (n384), .o (n385) );
  buffer buf_n386( .i (n385), .o (n386) );
  buffer buf_n387( .i (n386), .o (n387) );
  buffer buf_n388( .i (n387), .o (n388) );
  buffer buf_n389( .i (n388), .o (n389) );
  assign n669 = n389 & n623 ;
  buffer buf_n670( .i (n669), .o (n670) );
  assign n671 = n272 & n670 ;
  buffer buf_n672( .i (n671), .o (n672) );
  assign n673 = G25 & ~n672 ;
  assign n674 = ~G25 & n672 ;
  assign n675 = ~n673 & ~n674 ;
  assign n676 = n309 & n670 ;
  buffer buf_n677( .i (n676), .o (n677) );
  assign n678 = G26 & ~n677 ;
  assign n679 = ~G26 & n677 ;
  assign n680 = ~n678 & ~n679 ;
  assign n681 = n166 & n670 ;
  buffer buf_n682( .i (n681), .o (n682) );
  assign n683 = G27 & ~n682 ;
  assign n684 = ~G27 & n682 ;
  assign n685 = ~n683 & ~n684 ;
  assign n686 = n227 & n670 ;
  buffer buf_n687( .i (n686), .o (n687) );
  assign n688 = G28 & ~n687 ;
  assign n689 = ~G28 & n687 ;
  assign n690 = ~n688 & ~n689 ;
  buffer buf_n429( .i (n428), .o (n429) );
  buffer buf_n430( .i (n429), .o (n430) );
  buffer buf_n431( .i (n430), .o (n431) );
  buffer buf_n432( .i (n431), .o (n432) );
  buffer buf_n433( .i (n432), .o (n433) );
  assign n691 = n433 & n485 ;
  assign n692 = n621 & n691 ;
  buffer buf_n693( .i (n692), .o (n693) );
  assign n694 = n272 & n693 ;
  buffer buf_n695( .i (n694), .o (n695) );
  assign n696 = G29 | n695 ;
  assign n697 = G29 & n695 ;
  assign n698 = ~n696 | n697 ;
  assign n699 = n309 & n693 ;
  buffer buf_n700( .i (n699), .o (n700) );
  assign n701 = G30 & ~n700 ;
  assign n702 = ~G30 & n700 ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = n166 & n693 ;
  buffer buf_n705( .i (n704), .o (n705) );
  assign n706 = G31 & ~n705 ;
  assign n707 = ~G31 & n705 ;
  assign n708 = ~n706 & ~n707 ;
  assign n709 = n227 & n693 ;
  buffer buf_n710( .i (n709), .o (n710) );
  assign n711 = G32 | n710 ;
  assign n712 = G32 & n710 ;
  assign n713 = ~n711 | n712 ;
  assign G1324 = n512 ;
  assign G1325 = n517 ;
  assign G1326 = n522 ;
  assign G1327 = n527 ;
  assign G1328 = n542 ;
  assign G1329 = n547 ;
  assign G1330 = n552 ;
  assign G1331 = n557 ;
  assign G1332 = n573 ;
  assign G1333 = n578 ;
  assign G1334 = n583 ;
  assign G1335 = n588 ;
  assign G1336 = n596 ;
  assign G1337 = n601 ;
  assign G1338 = n606 ;
  assign G1339 = n611 ;
  assign G1340 = n630 ;
  assign G1341 = n635 ;
  assign G1342 = n640 ;
  assign G1343 = n645 ;
  assign G1344 = n653 ;
  assign G1345 = n658 ;
  assign G1346 = n663 ;
  assign G1347 = n668 ;
  assign G1348 = n675 ;
  assign G1349 = n680 ;
  assign G1350 = n685 ;
  assign G1351 = n690 ;
  assign G1352 = n698 ;
  assign G1353 = n703 ;
  assign G1354 = n708 ;
  assign G1355 = n713 ;
endmodule
